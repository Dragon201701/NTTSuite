
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed May 19 22:44:15 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [9:0] adra;
  input [9:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_5_tr0, modExp_while_C_24_tr0, VEC_LOOP_1_COMP_LOOP_C_1_tr0,
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24_tr0, VEC_LOOP_1_COMP_LOOP_C_40_tr0,
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0, VEC_LOOP_1_COMP_LOOP_C_80_tr0,
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0, VEC_LOOP_1_COMP_LOOP_C_120_tr0,
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0, VEC_LOOP_1_COMP_LOOP_C_160_tr0,
      VEC_LOOP_C_0_tr0, VEC_LOOP_2_COMP_LOOP_C_1_tr0, VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24_tr0,
      VEC_LOOP_2_COMP_LOOP_C_40_tr0, VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0,
      VEC_LOOP_2_COMP_LOOP_C_80_tr0, VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0,
      VEC_LOOP_2_COMP_LOOP_C_120_tr0, VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0,
      VEC_LOOP_2_COMP_LOOP_C_160_tr0, VEC_LOOP_C_1_tr0, STAGE_LOOP_C_6_tr0
);
  input clk;
  input rst;
  output [9:0] fsm_output;
  reg [9:0] fsm_output;
  input STAGE_LOOP_C_5_tr0;
  input modExp_while_C_24_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_1_tr0;
  input VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_40_tr0;
  input VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_80_tr0;
  input VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_120_tr0;
  input VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0;
  input VEC_LOOP_1_COMP_LOOP_C_160_tr0;
  input VEC_LOOP_C_0_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_1_tr0;
  input VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_40_tr0;
  input VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_80_tr0;
  input VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_120_tr0;
  input VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0;
  input VEC_LOOP_2_COMP_LOOP_C_160_tr0;
  input VEC_LOOP_C_1_tr0;
  input STAGE_LOOP_C_6_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 10'd0,
    STAGE_LOOP_C_0 = 10'd1,
    STAGE_LOOP_C_1 = 10'd2,
    STAGE_LOOP_C_2 = 10'd3,
    STAGE_LOOP_C_3 = 10'd4,
    STAGE_LOOP_C_4 = 10'd5,
    STAGE_LOOP_C_5 = 10'd6,
    modExp_while_C_0 = 10'd7,
    modExp_while_C_1 = 10'd8,
    modExp_while_C_2 = 10'd9,
    modExp_while_C_3 = 10'd10,
    modExp_while_C_4 = 10'd11,
    modExp_while_C_5 = 10'd12,
    modExp_while_C_6 = 10'd13,
    modExp_while_C_7 = 10'd14,
    modExp_while_C_8 = 10'd15,
    modExp_while_C_9 = 10'd16,
    modExp_while_C_10 = 10'd17,
    modExp_while_C_11 = 10'd18,
    modExp_while_C_12 = 10'd19,
    modExp_while_C_13 = 10'd20,
    modExp_while_C_14 = 10'd21,
    modExp_while_C_15 = 10'd22,
    modExp_while_C_16 = 10'd23,
    modExp_while_C_17 = 10'd24,
    modExp_while_C_18 = 10'd25,
    modExp_while_C_19 = 10'd26,
    modExp_while_C_20 = 10'd27,
    modExp_while_C_21 = 10'd28,
    modExp_while_C_22 = 10'd29,
    modExp_while_C_23 = 10'd30,
    modExp_while_C_24 = 10'd31,
    VEC_LOOP_1_COMP_LOOP_C_0 = 10'd32,
    VEC_LOOP_1_COMP_LOOP_C_1 = 10'd33,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0 = 10'd34,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1 = 10'd35,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2 = 10'd36,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3 = 10'd37,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4 = 10'd38,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5 = 10'd39,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6 = 10'd40,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7 = 10'd41,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8 = 10'd42,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9 = 10'd43,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10 = 10'd44,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11 = 10'd45,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12 = 10'd46,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13 = 10'd47,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14 = 10'd48,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15 = 10'd49,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16 = 10'd50,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17 = 10'd51,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18 = 10'd52,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19 = 10'd53,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20 = 10'd54,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21 = 10'd55,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22 = 10'd56,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23 = 10'd57,
    VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24 = 10'd58,
    VEC_LOOP_1_COMP_LOOP_C_2 = 10'd59,
    VEC_LOOP_1_COMP_LOOP_C_3 = 10'd60,
    VEC_LOOP_1_COMP_LOOP_C_4 = 10'd61,
    VEC_LOOP_1_COMP_LOOP_C_5 = 10'd62,
    VEC_LOOP_1_COMP_LOOP_C_6 = 10'd63,
    VEC_LOOP_1_COMP_LOOP_C_7 = 10'd64,
    VEC_LOOP_1_COMP_LOOP_C_8 = 10'd65,
    VEC_LOOP_1_COMP_LOOP_C_9 = 10'd66,
    VEC_LOOP_1_COMP_LOOP_C_10 = 10'd67,
    VEC_LOOP_1_COMP_LOOP_C_11 = 10'd68,
    VEC_LOOP_1_COMP_LOOP_C_12 = 10'd69,
    VEC_LOOP_1_COMP_LOOP_C_13 = 10'd70,
    VEC_LOOP_1_COMP_LOOP_C_14 = 10'd71,
    VEC_LOOP_1_COMP_LOOP_C_15 = 10'd72,
    VEC_LOOP_1_COMP_LOOP_C_16 = 10'd73,
    VEC_LOOP_1_COMP_LOOP_C_17 = 10'd74,
    VEC_LOOP_1_COMP_LOOP_C_18 = 10'd75,
    VEC_LOOP_1_COMP_LOOP_C_19 = 10'd76,
    VEC_LOOP_1_COMP_LOOP_C_20 = 10'd77,
    VEC_LOOP_1_COMP_LOOP_C_21 = 10'd78,
    VEC_LOOP_1_COMP_LOOP_C_22 = 10'd79,
    VEC_LOOP_1_COMP_LOOP_C_23 = 10'd80,
    VEC_LOOP_1_COMP_LOOP_C_24 = 10'd81,
    VEC_LOOP_1_COMP_LOOP_C_25 = 10'd82,
    VEC_LOOP_1_COMP_LOOP_C_26 = 10'd83,
    VEC_LOOP_1_COMP_LOOP_C_27 = 10'd84,
    VEC_LOOP_1_COMP_LOOP_C_28 = 10'd85,
    VEC_LOOP_1_COMP_LOOP_C_29 = 10'd86,
    VEC_LOOP_1_COMP_LOOP_C_30 = 10'd87,
    VEC_LOOP_1_COMP_LOOP_C_31 = 10'd88,
    VEC_LOOP_1_COMP_LOOP_C_32 = 10'd89,
    VEC_LOOP_1_COMP_LOOP_C_33 = 10'd90,
    VEC_LOOP_1_COMP_LOOP_C_34 = 10'd91,
    VEC_LOOP_1_COMP_LOOP_C_35 = 10'd92,
    VEC_LOOP_1_COMP_LOOP_C_36 = 10'd93,
    VEC_LOOP_1_COMP_LOOP_C_37 = 10'd94,
    VEC_LOOP_1_COMP_LOOP_C_38 = 10'd95,
    VEC_LOOP_1_COMP_LOOP_C_39 = 10'd96,
    VEC_LOOP_1_COMP_LOOP_C_40 = 10'd97,
    VEC_LOOP_1_COMP_LOOP_C_41 = 10'd98,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0 = 10'd99,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1 = 10'd100,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2 = 10'd101,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3 = 10'd102,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4 = 10'd103,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5 = 10'd104,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6 = 10'd105,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7 = 10'd106,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8 = 10'd107,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9 = 10'd108,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10 = 10'd109,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11 = 10'd110,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12 = 10'd111,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13 = 10'd112,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14 = 10'd113,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15 = 10'd114,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16 = 10'd115,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17 = 10'd116,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18 = 10'd117,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19 = 10'd118,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20 = 10'd119,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21 = 10'd120,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22 = 10'd121,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23 = 10'd122,
    VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24 = 10'd123,
    VEC_LOOP_1_COMP_LOOP_C_42 = 10'd124,
    VEC_LOOP_1_COMP_LOOP_C_43 = 10'd125,
    VEC_LOOP_1_COMP_LOOP_C_44 = 10'd126,
    VEC_LOOP_1_COMP_LOOP_C_45 = 10'd127,
    VEC_LOOP_1_COMP_LOOP_C_46 = 10'd128,
    VEC_LOOP_1_COMP_LOOP_C_47 = 10'd129,
    VEC_LOOP_1_COMP_LOOP_C_48 = 10'd130,
    VEC_LOOP_1_COMP_LOOP_C_49 = 10'd131,
    VEC_LOOP_1_COMP_LOOP_C_50 = 10'd132,
    VEC_LOOP_1_COMP_LOOP_C_51 = 10'd133,
    VEC_LOOP_1_COMP_LOOP_C_52 = 10'd134,
    VEC_LOOP_1_COMP_LOOP_C_53 = 10'd135,
    VEC_LOOP_1_COMP_LOOP_C_54 = 10'd136,
    VEC_LOOP_1_COMP_LOOP_C_55 = 10'd137,
    VEC_LOOP_1_COMP_LOOP_C_56 = 10'd138,
    VEC_LOOP_1_COMP_LOOP_C_57 = 10'd139,
    VEC_LOOP_1_COMP_LOOP_C_58 = 10'd140,
    VEC_LOOP_1_COMP_LOOP_C_59 = 10'd141,
    VEC_LOOP_1_COMP_LOOP_C_60 = 10'd142,
    VEC_LOOP_1_COMP_LOOP_C_61 = 10'd143,
    VEC_LOOP_1_COMP_LOOP_C_62 = 10'd144,
    VEC_LOOP_1_COMP_LOOP_C_63 = 10'd145,
    VEC_LOOP_1_COMP_LOOP_C_64 = 10'd146,
    VEC_LOOP_1_COMP_LOOP_C_65 = 10'd147,
    VEC_LOOP_1_COMP_LOOP_C_66 = 10'd148,
    VEC_LOOP_1_COMP_LOOP_C_67 = 10'd149,
    VEC_LOOP_1_COMP_LOOP_C_68 = 10'd150,
    VEC_LOOP_1_COMP_LOOP_C_69 = 10'd151,
    VEC_LOOP_1_COMP_LOOP_C_70 = 10'd152,
    VEC_LOOP_1_COMP_LOOP_C_71 = 10'd153,
    VEC_LOOP_1_COMP_LOOP_C_72 = 10'd154,
    VEC_LOOP_1_COMP_LOOP_C_73 = 10'd155,
    VEC_LOOP_1_COMP_LOOP_C_74 = 10'd156,
    VEC_LOOP_1_COMP_LOOP_C_75 = 10'd157,
    VEC_LOOP_1_COMP_LOOP_C_76 = 10'd158,
    VEC_LOOP_1_COMP_LOOP_C_77 = 10'd159,
    VEC_LOOP_1_COMP_LOOP_C_78 = 10'd160,
    VEC_LOOP_1_COMP_LOOP_C_79 = 10'd161,
    VEC_LOOP_1_COMP_LOOP_C_80 = 10'd162,
    VEC_LOOP_1_COMP_LOOP_C_81 = 10'd163,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_0 = 10'd164,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_1 = 10'd165,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_2 = 10'd166,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_3 = 10'd167,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_4 = 10'd168,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_5 = 10'd169,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_6 = 10'd170,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_7 = 10'd171,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_8 = 10'd172,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_9 = 10'd173,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_10 = 10'd174,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_11 = 10'd175,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_12 = 10'd176,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_13 = 10'd177,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_14 = 10'd178,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_15 = 10'd179,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_16 = 10'd180,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_17 = 10'd181,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_18 = 10'd182,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_19 = 10'd183,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_20 = 10'd184,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_21 = 10'd185,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_22 = 10'd186,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_23 = 10'd187,
    VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24 = 10'd188,
    VEC_LOOP_1_COMP_LOOP_C_82 = 10'd189,
    VEC_LOOP_1_COMP_LOOP_C_83 = 10'd190,
    VEC_LOOP_1_COMP_LOOP_C_84 = 10'd191,
    VEC_LOOP_1_COMP_LOOP_C_85 = 10'd192,
    VEC_LOOP_1_COMP_LOOP_C_86 = 10'd193,
    VEC_LOOP_1_COMP_LOOP_C_87 = 10'd194,
    VEC_LOOP_1_COMP_LOOP_C_88 = 10'd195,
    VEC_LOOP_1_COMP_LOOP_C_89 = 10'd196,
    VEC_LOOP_1_COMP_LOOP_C_90 = 10'd197,
    VEC_LOOP_1_COMP_LOOP_C_91 = 10'd198,
    VEC_LOOP_1_COMP_LOOP_C_92 = 10'd199,
    VEC_LOOP_1_COMP_LOOP_C_93 = 10'd200,
    VEC_LOOP_1_COMP_LOOP_C_94 = 10'd201,
    VEC_LOOP_1_COMP_LOOP_C_95 = 10'd202,
    VEC_LOOP_1_COMP_LOOP_C_96 = 10'd203,
    VEC_LOOP_1_COMP_LOOP_C_97 = 10'd204,
    VEC_LOOP_1_COMP_LOOP_C_98 = 10'd205,
    VEC_LOOP_1_COMP_LOOP_C_99 = 10'd206,
    VEC_LOOP_1_COMP_LOOP_C_100 = 10'd207,
    VEC_LOOP_1_COMP_LOOP_C_101 = 10'd208,
    VEC_LOOP_1_COMP_LOOP_C_102 = 10'd209,
    VEC_LOOP_1_COMP_LOOP_C_103 = 10'd210,
    VEC_LOOP_1_COMP_LOOP_C_104 = 10'd211,
    VEC_LOOP_1_COMP_LOOP_C_105 = 10'd212,
    VEC_LOOP_1_COMP_LOOP_C_106 = 10'd213,
    VEC_LOOP_1_COMP_LOOP_C_107 = 10'd214,
    VEC_LOOP_1_COMP_LOOP_C_108 = 10'd215,
    VEC_LOOP_1_COMP_LOOP_C_109 = 10'd216,
    VEC_LOOP_1_COMP_LOOP_C_110 = 10'd217,
    VEC_LOOP_1_COMP_LOOP_C_111 = 10'd218,
    VEC_LOOP_1_COMP_LOOP_C_112 = 10'd219,
    VEC_LOOP_1_COMP_LOOP_C_113 = 10'd220,
    VEC_LOOP_1_COMP_LOOP_C_114 = 10'd221,
    VEC_LOOP_1_COMP_LOOP_C_115 = 10'd222,
    VEC_LOOP_1_COMP_LOOP_C_116 = 10'd223,
    VEC_LOOP_1_COMP_LOOP_C_117 = 10'd224,
    VEC_LOOP_1_COMP_LOOP_C_118 = 10'd225,
    VEC_LOOP_1_COMP_LOOP_C_119 = 10'd226,
    VEC_LOOP_1_COMP_LOOP_C_120 = 10'd227,
    VEC_LOOP_1_COMP_LOOP_C_121 = 10'd228,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_0 = 10'd229,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_1 = 10'd230,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_2 = 10'd231,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_3 = 10'd232,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_4 = 10'd233,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_5 = 10'd234,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_6 = 10'd235,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_7 = 10'd236,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_8 = 10'd237,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_9 = 10'd238,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_10 = 10'd239,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_11 = 10'd240,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_12 = 10'd241,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_13 = 10'd242,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_14 = 10'd243,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_15 = 10'd244,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_16 = 10'd245,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_17 = 10'd246,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_18 = 10'd247,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_19 = 10'd248,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_20 = 10'd249,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_21 = 10'd250,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_22 = 10'd251,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_23 = 10'd252,
    VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24 = 10'd253,
    VEC_LOOP_1_COMP_LOOP_C_122 = 10'd254,
    VEC_LOOP_1_COMP_LOOP_C_123 = 10'd255,
    VEC_LOOP_1_COMP_LOOP_C_124 = 10'd256,
    VEC_LOOP_1_COMP_LOOP_C_125 = 10'd257,
    VEC_LOOP_1_COMP_LOOP_C_126 = 10'd258,
    VEC_LOOP_1_COMP_LOOP_C_127 = 10'd259,
    VEC_LOOP_1_COMP_LOOP_C_128 = 10'd260,
    VEC_LOOP_1_COMP_LOOP_C_129 = 10'd261,
    VEC_LOOP_1_COMP_LOOP_C_130 = 10'd262,
    VEC_LOOP_1_COMP_LOOP_C_131 = 10'd263,
    VEC_LOOP_1_COMP_LOOP_C_132 = 10'd264,
    VEC_LOOP_1_COMP_LOOP_C_133 = 10'd265,
    VEC_LOOP_1_COMP_LOOP_C_134 = 10'd266,
    VEC_LOOP_1_COMP_LOOP_C_135 = 10'd267,
    VEC_LOOP_1_COMP_LOOP_C_136 = 10'd268,
    VEC_LOOP_1_COMP_LOOP_C_137 = 10'd269,
    VEC_LOOP_1_COMP_LOOP_C_138 = 10'd270,
    VEC_LOOP_1_COMP_LOOP_C_139 = 10'd271,
    VEC_LOOP_1_COMP_LOOP_C_140 = 10'd272,
    VEC_LOOP_1_COMP_LOOP_C_141 = 10'd273,
    VEC_LOOP_1_COMP_LOOP_C_142 = 10'd274,
    VEC_LOOP_1_COMP_LOOP_C_143 = 10'd275,
    VEC_LOOP_1_COMP_LOOP_C_144 = 10'd276,
    VEC_LOOP_1_COMP_LOOP_C_145 = 10'd277,
    VEC_LOOP_1_COMP_LOOP_C_146 = 10'd278,
    VEC_LOOP_1_COMP_LOOP_C_147 = 10'd279,
    VEC_LOOP_1_COMP_LOOP_C_148 = 10'd280,
    VEC_LOOP_1_COMP_LOOP_C_149 = 10'd281,
    VEC_LOOP_1_COMP_LOOP_C_150 = 10'd282,
    VEC_LOOP_1_COMP_LOOP_C_151 = 10'd283,
    VEC_LOOP_1_COMP_LOOP_C_152 = 10'd284,
    VEC_LOOP_1_COMP_LOOP_C_153 = 10'd285,
    VEC_LOOP_1_COMP_LOOP_C_154 = 10'd286,
    VEC_LOOP_1_COMP_LOOP_C_155 = 10'd287,
    VEC_LOOP_1_COMP_LOOP_C_156 = 10'd288,
    VEC_LOOP_1_COMP_LOOP_C_157 = 10'd289,
    VEC_LOOP_1_COMP_LOOP_C_158 = 10'd290,
    VEC_LOOP_1_COMP_LOOP_C_159 = 10'd291,
    VEC_LOOP_1_COMP_LOOP_C_160 = 10'd292,
    VEC_LOOP_C_0 = 10'd293,
    VEC_LOOP_2_COMP_LOOP_C_0 = 10'd294,
    VEC_LOOP_2_COMP_LOOP_C_1 = 10'd295,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0 = 10'd296,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1 = 10'd297,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2 = 10'd298,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3 = 10'd299,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4 = 10'd300,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5 = 10'd301,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6 = 10'd302,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7 = 10'd303,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8 = 10'd304,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9 = 10'd305,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10 = 10'd306,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11 = 10'd307,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12 = 10'd308,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13 = 10'd309,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14 = 10'd310,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15 = 10'd311,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16 = 10'd312,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17 = 10'd313,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18 = 10'd314,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19 = 10'd315,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20 = 10'd316,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21 = 10'd317,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22 = 10'd318,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23 = 10'd319,
    VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24 = 10'd320,
    VEC_LOOP_2_COMP_LOOP_C_2 = 10'd321,
    VEC_LOOP_2_COMP_LOOP_C_3 = 10'd322,
    VEC_LOOP_2_COMP_LOOP_C_4 = 10'd323,
    VEC_LOOP_2_COMP_LOOP_C_5 = 10'd324,
    VEC_LOOP_2_COMP_LOOP_C_6 = 10'd325,
    VEC_LOOP_2_COMP_LOOP_C_7 = 10'd326,
    VEC_LOOP_2_COMP_LOOP_C_8 = 10'd327,
    VEC_LOOP_2_COMP_LOOP_C_9 = 10'd328,
    VEC_LOOP_2_COMP_LOOP_C_10 = 10'd329,
    VEC_LOOP_2_COMP_LOOP_C_11 = 10'd330,
    VEC_LOOP_2_COMP_LOOP_C_12 = 10'd331,
    VEC_LOOP_2_COMP_LOOP_C_13 = 10'd332,
    VEC_LOOP_2_COMP_LOOP_C_14 = 10'd333,
    VEC_LOOP_2_COMP_LOOP_C_15 = 10'd334,
    VEC_LOOP_2_COMP_LOOP_C_16 = 10'd335,
    VEC_LOOP_2_COMP_LOOP_C_17 = 10'd336,
    VEC_LOOP_2_COMP_LOOP_C_18 = 10'd337,
    VEC_LOOP_2_COMP_LOOP_C_19 = 10'd338,
    VEC_LOOP_2_COMP_LOOP_C_20 = 10'd339,
    VEC_LOOP_2_COMP_LOOP_C_21 = 10'd340,
    VEC_LOOP_2_COMP_LOOP_C_22 = 10'd341,
    VEC_LOOP_2_COMP_LOOP_C_23 = 10'd342,
    VEC_LOOP_2_COMP_LOOP_C_24 = 10'd343,
    VEC_LOOP_2_COMP_LOOP_C_25 = 10'd344,
    VEC_LOOP_2_COMP_LOOP_C_26 = 10'd345,
    VEC_LOOP_2_COMP_LOOP_C_27 = 10'd346,
    VEC_LOOP_2_COMP_LOOP_C_28 = 10'd347,
    VEC_LOOP_2_COMP_LOOP_C_29 = 10'd348,
    VEC_LOOP_2_COMP_LOOP_C_30 = 10'd349,
    VEC_LOOP_2_COMP_LOOP_C_31 = 10'd350,
    VEC_LOOP_2_COMP_LOOP_C_32 = 10'd351,
    VEC_LOOP_2_COMP_LOOP_C_33 = 10'd352,
    VEC_LOOP_2_COMP_LOOP_C_34 = 10'd353,
    VEC_LOOP_2_COMP_LOOP_C_35 = 10'd354,
    VEC_LOOP_2_COMP_LOOP_C_36 = 10'd355,
    VEC_LOOP_2_COMP_LOOP_C_37 = 10'd356,
    VEC_LOOP_2_COMP_LOOP_C_38 = 10'd357,
    VEC_LOOP_2_COMP_LOOP_C_39 = 10'd358,
    VEC_LOOP_2_COMP_LOOP_C_40 = 10'd359,
    VEC_LOOP_2_COMP_LOOP_C_41 = 10'd360,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0 = 10'd361,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1 = 10'd362,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2 = 10'd363,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3 = 10'd364,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4 = 10'd365,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5 = 10'd366,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6 = 10'd367,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7 = 10'd368,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8 = 10'd369,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9 = 10'd370,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10 = 10'd371,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11 = 10'd372,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12 = 10'd373,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13 = 10'd374,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14 = 10'd375,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15 = 10'd376,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16 = 10'd377,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17 = 10'd378,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18 = 10'd379,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19 = 10'd380,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20 = 10'd381,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21 = 10'd382,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22 = 10'd383,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23 = 10'd384,
    VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24 = 10'd385,
    VEC_LOOP_2_COMP_LOOP_C_42 = 10'd386,
    VEC_LOOP_2_COMP_LOOP_C_43 = 10'd387,
    VEC_LOOP_2_COMP_LOOP_C_44 = 10'd388,
    VEC_LOOP_2_COMP_LOOP_C_45 = 10'd389,
    VEC_LOOP_2_COMP_LOOP_C_46 = 10'd390,
    VEC_LOOP_2_COMP_LOOP_C_47 = 10'd391,
    VEC_LOOP_2_COMP_LOOP_C_48 = 10'd392,
    VEC_LOOP_2_COMP_LOOP_C_49 = 10'd393,
    VEC_LOOP_2_COMP_LOOP_C_50 = 10'd394,
    VEC_LOOP_2_COMP_LOOP_C_51 = 10'd395,
    VEC_LOOP_2_COMP_LOOP_C_52 = 10'd396,
    VEC_LOOP_2_COMP_LOOP_C_53 = 10'd397,
    VEC_LOOP_2_COMP_LOOP_C_54 = 10'd398,
    VEC_LOOP_2_COMP_LOOP_C_55 = 10'd399,
    VEC_LOOP_2_COMP_LOOP_C_56 = 10'd400,
    VEC_LOOP_2_COMP_LOOP_C_57 = 10'd401,
    VEC_LOOP_2_COMP_LOOP_C_58 = 10'd402,
    VEC_LOOP_2_COMP_LOOP_C_59 = 10'd403,
    VEC_LOOP_2_COMP_LOOP_C_60 = 10'd404,
    VEC_LOOP_2_COMP_LOOP_C_61 = 10'd405,
    VEC_LOOP_2_COMP_LOOP_C_62 = 10'd406,
    VEC_LOOP_2_COMP_LOOP_C_63 = 10'd407,
    VEC_LOOP_2_COMP_LOOP_C_64 = 10'd408,
    VEC_LOOP_2_COMP_LOOP_C_65 = 10'd409,
    VEC_LOOP_2_COMP_LOOP_C_66 = 10'd410,
    VEC_LOOP_2_COMP_LOOP_C_67 = 10'd411,
    VEC_LOOP_2_COMP_LOOP_C_68 = 10'd412,
    VEC_LOOP_2_COMP_LOOP_C_69 = 10'd413,
    VEC_LOOP_2_COMP_LOOP_C_70 = 10'd414,
    VEC_LOOP_2_COMP_LOOP_C_71 = 10'd415,
    VEC_LOOP_2_COMP_LOOP_C_72 = 10'd416,
    VEC_LOOP_2_COMP_LOOP_C_73 = 10'd417,
    VEC_LOOP_2_COMP_LOOP_C_74 = 10'd418,
    VEC_LOOP_2_COMP_LOOP_C_75 = 10'd419,
    VEC_LOOP_2_COMP_LOOP_C_76 = 10'd420,
    VEC_LOOP_2_COMP_LOOP_C_77 = 10'd421,
    VEC_LOOP_2_COMP_LOOP_C_78 = 10'd422,
    VEC_LOOP_2_COMP_LOOP_C_79 = 10'd423,
    VEC_LOOP_2_COMP_LOOP_C_80 = 10'd424,
    VEC_LOOP_2_COMP_LOOP_C_81 = 10'd425,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_0 = 10'd426,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_1 = 10'd427,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_2 = 10'd428,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_3 = 10'd429,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_4 = 10'd430,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_5 = 10'd431,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_6 = 10'd432,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_7 = 10'd433,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_8 = 10'd434,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_9 = 10'd435,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_10 = 10'd436,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_11 = 10'd437,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_12 = 10'd438,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_13 = 10'd439,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_14 = 10'd440,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_15 = 10'd441,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_16 = 10'd442,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_17 = 10'd443,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_18 = 10'd444,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_19 = 10'd445,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_20 = 10'd446,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_21 = 10'd447,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_22 = 10'd448,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_23 = 10'd449,
    VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24 = 10'd450,
    VEC_LOOP_2_COMP_LOOP_C_82 = 10'd451,
    VEC_LOOP_2_COMP_LOOP_C_83 = 10'd452,
    VEC_LOOP_2_COMP_LOOP_C_84 = 10'd453,
    VEC_LOOP_2_COMP_LOOP_C_85 = 10'd454,
    VEC_LOOP_2_COMP_LOOP_C_86 = 10'd455,
    VEC_LOOP_2_COMP_LOOP_C_87 = 10'd456,
    VEC_LOOP_2_COMP_LOOP_C_88 = 10'd457,
    VEC_LOOP_2_COMP_LOOP_C_89 = 10'd458,
    VEC_LOOP_2_COMP_LOOP_C_90 = 10'd459,
    VEC_LOOP_2_COMP_LOOP_C_91 = 10'd460,
    VEC_LOOP_2_COMP_LOOP_C_92 = 10'd461,
    VEC_LOOP_2_COMP_LOOP_C_93 = 10'd462,
    VEC_LOOP_2_COMP_LOOP_C_94 = 10'd463,
    VEC_LOOP_2_COMP_LOOP_C_95 = 10'd464,
    VEC_LOOP_2_COMP_LOOP_C_96 = 10'd465,
    VEC_LOOP_2_COMP_LOOP_C_97 = 10'd466,
    VEC_LOOP_2_COMP_LOOP_C_98 = 10'd467,
    VEC_LOOP_2_COMP_LOOP_C_99 = 10'd468,
    VEC_LOOP_2_COMP_LOOP_C_100 = 10'd469,
    VEC_LOOP_2_COMP_LOOP_C_101 = 10'd470,
    VEC_LOOP_2_COMP_LOOP_C_102 = 10'd471,
    VEC_LOOP_2_COMP_LOOP_C_103 = 10'd472,
    VEC_LOOP_2_COMP_LOOP_C_104 = 10'd473,
    VEC_LOOP_2_COMP_LOOP_C_105 = 10'd474,
    VEC_LOOP_2_COMP_LOOP_C_106 = 10'd475,
    VEC_LOOP_2_COMP_LOOP_C_107 = 10'd476,
    VEC_LOOP_2_COMP_LOOP_C_108 = 10'd477,
    VEC_LOOP_2_COMP_LOOP_C_109 = 10'd478,
    VEC_LOOP_2_COMP_LOOP_C_110 = 10'd479,
    VEC_LOOP_2_COMP_LOOP_C_111 = 10'd480,
    VEC_LOOP_2_COMP_LOOP_C_112 = 10'd481,
    VEC_LOOP_2_COMP_LOOP_C_113 = 10'd482,
    VEC_LOOP_2_COMP_LOOP_C_114 = 10'd483,
    VEC_LOOP_2_COMP_LOOP_C_115 = 10'd484,
    VEC_LOOP_2_COMP_LOOP_C_116 = 10'd485,
    VEC_LOOP_2_COMP_LOOP_C_117 = 10'd486,
    VEC_LOOP_2_COMP_LOOP_C_118 = 10'd487,
    VEC_LOOP_2_COMP_LOOP_C_119 = 10'd488,
    VEC_LOOP_2_COMP_LOOP_C_120 = 10'd489,
    VEC_LOOP_2_COMP_LOOP_C_121 = 10'd490,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_0 = 10'd491,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_1 = 10'd492,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_2 = 10'd493,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_3 = 10'd494,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_4 = 10'd495,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_5 = 10'd496,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_6 = 10'd497,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_7 = 10'd498,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_8 = 10'd499,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_9 = 10'd500,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_10 = 10'd501,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_11 = 10'd502,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_12 = 10'd503,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_13 = 10'd504,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_14 = 10'd505,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_15 = 10'd506,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_16 = 10'd507,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_17 = 10'd508,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_18 = 10'd509,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_19 = 10'd510,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_20 = 10'd511,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_21 = 10'd512,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_22 = 10'd513,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_23 = 10'd514,
    VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24 = 10'd515,
    VEC_LOOP_2_COMP_LOOP_C_122 = 10'd516,
    VEC_LOOP_2_COMP_LOOP_C_123 = 10'd517,
    VEC_LOOP_2_COMP_LOOP_C_124 = 10'd518,
    VEC_LOOP_2_COMP_LOOP_C_125 = 10'd519,
    VEC_LOOP_2_COMP_LOOP_C_126 = 10'd520,
    VEC_LOOP_2_COMP_LOOP_C_127 = 10'd521,
    VEC_LOOP_2_COMP_LOOP_C_128 = 10'd522,
    VEC_LOOP_2_COMP_LOOP_C_129 = 10'd523,
    VEC_LOOP_2_COMP_LOOP_C_130 = 10'd524,
    VEC_LOOP_2_COMP_LOOP_C_131 = 10'd525,
    VEC_LOOP_2_COMP_LOOP_C_132 = 10'd526,
    VEC_LOOP_2_COMP_LOOP_C_133 = 10'd527,
    VEC_LOOP_2_COMP_LOOP_C_134 = 10'd528,
    VEC_LOOP_2_COMP_LOOP_C_135 = 10'd529,
    VEC_LOOP_2_COMP_LOOP_C_136 = 10'd530,
    VEC_LOOP_2_COMP_LOOP_C_137 = 10'd531,
    VEC_LOOP_2_COMP_LOOP_C_138 = 10'd532,
    VEC_LOOP_2_COMP_LOOP_C_139 = 10'd533,
    VEC_LOOP_2_COMP_LOOP_C_140 = 10'd534,
    VEC_LOOP_2_COMP_LOOP_C_141 = 10'd535,
    VEC_LOOP_2_COMP_LOOP_C_142 = 10'd536,
    VEC_LOOP_2_COMP_LOOP_C_143 = 10'd537,
    VEC_LOOP_2_COMP_LOOP_C_144 = 10'd538,
    VEC_LOOP_2_COMP_LOOP_C_145 = 10'd539,
    VEC_LOOP_2_COMP_LOOP_C_146 = 10'd540,
    VEC_LOOP_2_COMP_LOOP_C_147 = 10'd541,
    VEC_LOOP_2_COMP_LOOP_C_148 = 10'd542,
    VEC_LOOP_2_COMP_LOOP_C_149 = 10'd543,
    VEC_LOOP_2_COMP_LOOP_C_150 = 10'd544,
    VEC_LOOP_2_COMP_LOOP_C_151 = 10'd545,
    VEC_LOOP_2_COMP_LOOP_C_152 = 10'd546,
    VEC_LOOP_2_COMP_LOOP_C_153 = 10'd547,
    VEC_LOOP_2_COMP_LOOP_C_154 = 10'd548,
    VEC_LOOP_2_COMP_LOOP_C_155 = 10'd549,
    VEC_LOOP_2_COMP_LOOP_C_156 = 10'd550,
    VEC_LOOP_2_COMP_LOOP_C_157 = 10'd551,
    VEC_LOOP_2_COMP_LOOP_C_158 = 10'd552,
    VEC_LOOP_2_COMP_LOOP_C_159 = 10'd553,
    VEC_LOOP_2_COMP_LOOP_C_160 = 10'd554,
    VEC_LOOP_C_1 = 10'd555,
    STAGE_LOOP_C_6 = 10'd556,
    main_C_1 = 10'd557;

  reg [9:0] state_var;
  reg [9:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 10'b0000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 10'b0000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 10'b0000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 10'b0000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 10'b0000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 10'b0000000110;
        if ( STAGE_LOOP_C_5_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 10'b0000000111;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 10'b0000001000;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 10'b0000001001;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 10'b0000001010;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 10'b0000001011;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 10'b0000001100;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 10'b0000001101;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 10'b0000001110;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 10'b0000001111;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 10'b0000010000;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 10'b0000010001;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 10'b0000010010;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 10'b0000010011;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 10'b0000010100;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 10'b0000010101;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 10'b0000010110;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 10'b0000010111;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 10'b0000011000;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 10'b0000011001;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 10'b0000011010;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 10'b0000011011;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 10'b0000011100;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 10'b0000011101;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 10'b0000011110;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 10'b0000011111;
        if ( modExp_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_0 : begin
        fsm_output = 10'b0000100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_C_1 : begin
        fsm_output = 10'b0000100001;
        if ( VEC_LOOP_1_COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 10'b0000100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 10'b0000100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 10'b0000100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 10'b0000100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 10'b0000100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 10'b0000100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 10'b0000101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 10'b0000101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 10'b0000101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 10'b0000101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 10'b0000101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 10'b0000101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 10'b0000101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 10'b0000101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 10'b0000110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 10'b0000110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 10'b0000110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 10'b0000110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 10'b0000110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 10'b0000110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 10'b0000110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 10'b0000110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 10'b0000111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 10'b0000111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 10'b0000111010;
        if ( VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_2 : begin
        fsm_output = 10'b0000111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_C_3 : begin
        fsm_output = 10'b0000111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_C_4 : begin
        fsm_output = 10'b0000111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_C_5 : begin
        fsm_output = 10'b0000111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_C_6 : begin
        fsm_output = 10'b0000111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_C_7 : begin
        fsm_output = 10'b0001000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_C_8 : begin
        fsm_output = 10'b0001000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_C_9 : begin
        fsm_output = 10'b0001000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_C_10 : begin
        fsm_output = 10'b0001000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_C_11 : begin
        fsm_output = 10'b0001000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_C_12 : begin
        fsm_output = 10'b0001000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_C_13 : begin
        fsm_output = 10'b0001000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_C_14 : begin
        fsm_output = 10'b0001000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_C_15 : begin
        fsm_output = 10'b0001001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_C_16 : begin
        fsm_output = 10'b0001001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_C_17 : begin
        fsm_output = 10'b0001001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_C_18 : begin
        fsm_output = 10'b0001001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_C_19 : begin
        fsm_output = 10'b0001001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_C_20 : begin
        fsm_output = 10'b0001001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_C_21 : begin
        fsm_output = 10'b0001001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_C_22 : begin
        fsm_output = 10'b0001001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_C_23 : begin
        fsm_output = 10'b0001010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_C_24 : begin
        fsm_output = 10'b0001010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_25;
      end
      VEC_LOOP_1_COMP_LOOP_C_25 : begin
        fsm_output = 10'b0001010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_26;
      end
      VEC_LOOP_1_COMP_LOOP_C_26 : begin
        fsm_output = 10'b0001010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_27;
      end
      VEC_LOOP_1_COMP_LOOP_C_27 : begin
        fsm_output = 10'b0001010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_28;
      end
      VEC_LOOP_1_COMP_LOOP_C_28 : begin
        fsm_output = 10'b0001010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_29;
      end
      VEC_LOOP_1_COMP_LOOP_C_29 : begin
        fsm_output = 10'b0001010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_30;
      end
      VEC_LOOP_1_COMP_LOOP_C_30 : begin
        fsm_output = 10'b0001010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_31;
      end
      VEC_LOOP_1_COMP_LOOP_C_31 : begin
        fsm_output = 10'b0001011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_32;
      end
      VEC_LOOP_1_COMP_LOOP_C_32 : begin
        fsm_output = 10'b0001011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_33;
      end
      VEC_LOOP_1_COMP_LOOP_C_33 : begin
        fsm_output = 10'b0001011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_34;
      end
      VEC_LOOP_1_COMP_LOOP_C_34 : begin
        fsm_output = 10'b0001011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_35;
      end
      VEC_LOOP_1_COMP_LOOP_C_35 : begin
        fsm_output = 10'b0001011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_36;
      end
      VEC_LOOP_1_COMP_LOOP_C_36 : begin
        fsm_output = 10'b0001011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_37;
      end
      VEC_LOOP_1_COMP_LOOP_C_37 : begin
        fsm_output = 10'b0001011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_38;
      end
      VEC_LOOP_1_COMP_LOOP_C_38 : begin
        fsm_output = 10'b0001011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_39;
      end
      VEC_LOOP_1_COMP_LOOP_C_39 : begin
        fsm_output = 10'b0001100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_40;
      end
      VEC_LOOP_1_COMP_LOOP_C_40 : begin
        fsm_output = 10'b0001100001;
        if ( VEC_LOOP_1_COMP_LOOP_C_40_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_41;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_41 : begin
        fsm_output = 10'b0001100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 10'b0001100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 10'b0001100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 10'b0001100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 10'b0001100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 10'b0001100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 10'b0001101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 10'b0001101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 10'b0001101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 10'b0001101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 10'b0001101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 10'b0001101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 10'b0001101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 10'b0001101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 10'b0001110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 10'b0001110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 10'b0001110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 10'b0001110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 10'b0001110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 10'b0001110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 10'b0001110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 10'b0001110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 10'b0001111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 10'b0001111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 10'b0001111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 10'b0001111011;
        if ( VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_42;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_42 : begin
        fsm_output = 10'b0001111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_43;
      end
      VEC_LOOP_1_COMP_LOOP_C_43 : begin
        fsm_output = 10'b0001111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_44;
      end
      VEC_LOOP_1_COMP_LOOP_C_44 : begin
        fsm_output = 10'b0001111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_45;
      end
      VEC_LOOP_1_COMP_LOOP_C_45 : begin
        fsm_output = 10'b0001111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_46;
      end
      VEC_LOOP_1_COMP_LOOP_C_46 : begin
        fsm_output = 10'b0010000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_47;
      end
      VEC_LOOP_1_COMP_LOOP_C_47 : begin
        fsm_output = 10'b0010000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_48;
      end
      VEC_LOOP_1_COMP_LOOP_C_48 : begin
        fsm_output = 10'b0010000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_49;
      end
      VEC_LOOP_1_COMP_LOOP_C_49 : begin
        fsm_output = 10'b0010000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_50;
      end
      VEC_LOOP_1_COMP_LOOP_C_50 : begin
        fsm_output = 10'b0010000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_51;
      end
      VEC_LOOP_1_COMP_LOOP_C_51 : begin
        fsm_output = 10'b0010000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_52;
      end
      VEC_LOOP_1_COMP_LOOP_C_52 : begin
        fsm_output = 10'b0010000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_53;
      end
      VEC_LOOP_1_COMP_LOOP_C_53 : begin
        fsm_output = 10'b0010000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_54;
      end
      VEC_LOOP_1_COMP_LOOP_C_54 : begin
        fsm_output = 10'b0010001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_55;
      end
      VEC_LOOP_1_COMP_LOOP_C_55 : begin
        fsm_output = 10'b0010001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_56;
      end
      VEC_LOOP_1_COMP_LOOP_C_56 : begin
        fsm_output = 10'b0010001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_57;
      end
      VEC_LOOP_1_COMP_LOOP_C_57 : begin
        fsm_output = 10'b0010001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_58;
      end
      VEC_LOOP_1_COMP_LOOP_C_58 : begin
        fsm_output = 10'b0010001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_59;
      end
      VEC_LOOP_1_COMP_LOOP_C_59 : begin
        fsm_output = 10'b0010001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_60;
      end
      VEC_LOOP_1_COMP_LOOP_C_60 : begin
        fsm_output = 10'b0010001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_61;
      end
      VEC_LOOP_1_COMP_LOOP_C_61 : begin
        fsm_output = 10'b0010001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_62;
      end
      VEC_LOOP_1_COMP_LOOP_C_62 : begin
        fsm_output = 10'b0010010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_63;
      end
      VEC_LOOP_1_COMP_LOOP_C_63 : begin
        fsm_output = 10'b0010010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_64;
      end
      VEC_LOOP_1_COMP_LOOP_C_64 : begin
        fsm_output = 10'b0010010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_65;
      end
      VEC_LOOP_1_COMP_LOOP_C_65 : begin
        fsm_output = 10'b0010010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_66;
      end
      VEC_LOOP_1_COMP_LOOP_C_66 : begin
        fsm_output = 10'b0010010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_67;
      end
      VEC_LOOP_1_COMP_LOOP_C_67 : begin
        fsm_output = 10'b0010010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_68;
      end
      VEC_LOOP_1_COMP_LOOP_C_68 : begin
        fsm_output = 10'b0010010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_69;
      end
      VEC_LOOP_1_COMP_LOOP_C_69 : begin
        fsm_output = 10'b0010010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_70;
      end
      VEC_LOOP_1_COMP_LOOP_C_70 : begin
        fsm_output = 10'b0010011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_71;
      end
      VEC_LOOP_1_COMP_LOOP_C_71 : begin
        fsm_output = 10'b0010011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_72;
      end
      VEC_LOOP_1_COMP_LOOP_C_72 : begin
        fsm_output = 10'b0010011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_73;
      end
      VEC_LOOP_1_COMP_LOOP_C_73 : begin
        fsm_output = 10'b0010011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_74;
      end
      VEC_LOOP_1_COMP_LOOP_C_74 : begin
        fsm_output = 10'b0010011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_75;
      end
      VEC_LOOP_1_COMP_LOOP_C_75 : begin
        fsm_output = 10'b0010011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_76;
      end
      VEC_LOOP_1_COMP_LOOP_C_76 : begin
        fsm_output = 10'b0010011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_77;
      end
      VEC_LOOP_1_COMP_LOOP_C_77 : begin
        fsm_output = 10'b0010011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_78;
      end
      VEC_LOOP_1_COMP_LOOP_C_78 : begin
        fsm_output = 10'b0010100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_79;
      end
      VEC_LOOP_1_COMP_LOOP_C_79 : begin
        fsm_output = 10'b0010100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_80;
      end
      VEC_LOOP_1_COMP_LOOP_C_80 : begin
        fsm_output = 10'b0010100010;
        if ( VEC_LOOP_1_COMP_LOOP_C_80_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_81;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_81 : begin
        fsm_output = 10'b0010100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_0;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 10'b0010100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 10'b0010100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 10'b0010100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 10'b0010100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 10'b0010101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 10'b0010101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 10'b0010101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 10'b0010101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 10'b0010101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 10'b0010101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 10'b0010101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 10'b0010101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 10'b0010110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 10'b0010110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 10'b0010110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 10'b0010110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 10'b0010110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 10'b0010110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 10'b0010110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 10'b0010110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 10'b0010111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 10'b0010111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 10'b0010111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 10'b0010111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 10'b0010111100;
        if ( VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_82;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_82 : begin
        fsm_output = 10'b0010111101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_83;
      end
      VEC_LOOP_1_COMP_LOOP_C_83 : begin
        fsm_output = 10'b0010111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_84;
      end
      VEC_LOOP_1_COMP_LOOP_C_84 : begin
        fsm_output = 10'b0010111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_85;
      end
      VEC_LOOP_1_COMP_LOOP_C_85 : begin
        fsm_output = 10'b0011000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_86;
      end
      VEC_LOOP_1_COMP_LOOP_C_86 : begin
        fsm_output = 10'b0011000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_87;
      end
      VEC_LOOP_1_COMP_LOOP_C_87 : begin
        fsm_output = 10'b0011000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_88;
      end
      VEC_LOOP_1_COMP_LOOP_C_88 : begin
        fsm_output = 10'b0011000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_89;
      end
      VEC_LOOP_1_COMP_LOOP_C_89 : begin
        fsm_output = 10'b0011000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_90;
      end
      VEC_LOOP_1_COMP_LOOP_C_90 : begin
        fsm_output = 10'b0011000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_91;
      end
      VEC_LOOP_1_COMP_LOOP_C_91 : begin
        fsm_output = 10'b0011000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_92;
      end
      VEC_LOOP_1_COMP_LOOP_C_92 : begin
        fsm_output = 10'b0011000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_93;
      end
      VEC_LOOP_1_COMP_LOOP_C_93 : begin
        fsm_output = 10'b0011001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_94;
      end
      VEC_LOOP_1_COMP_LOOP_C_94 : begin
        fsm_output = 10'b0011001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_95;
      end
      VEC_LOOP_1_COMP_LOOP_C_95 : begin
        fsm_output = 10'b0011001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_96;
      end
      VEC_LOOP_1_COMP_LOOP_C_96 : begin
        fsm_output = 10'b0011001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_97;
      end
      VEC_LOOP_1_COMP_LOOP_C_97 : begin
        fsm_output = 10'b0011001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_98;
      end
      VEC_LOOP_1_COMP_LOOP_C_98 : begin
        fsm_output = 10'b0011001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_99;
      end
      VEC_LOOP_1_COMP_LOOP_C_99 : begin
        fsm_output = 10'b0011001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_100;
      end
      VEC_LOOP_1_COMP_LOOP_C_100 : begin
        fsm_output = 10'b0011001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_101;
      end
      VEC_LOOP_1_COMP_LOOP_C_101 : begin
        fsm_output = 10'b0011010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_102;
      end
      VEC_LOOP_1_COMP_LOOP_C_102 : begin
        fsm_output = 10'b0011010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_103;
      end
      VEC_LOOP_1_COMP_LOOP_C_103 : begin
        fsm_output = 10'b0011010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_104;
      end
      VEC_LOOP_1_COMP_LOOP_C_104 : begin
        fsm_output = 10'b0011010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_105;
      end
      VEC_LOOP_1_COMP_LOOP_C_105 : begin
        fsm_output = 10'b0011010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_106;
      end
      VEC_LOOP_1_COMP_LOOP_C_106 : begin
        fsm_output = 10'b0011010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_107;
      end
      VEC_LOOP_1_COMP_LOOP_C_107 : begin
        fsm_output = 10'b0011010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_108;
      end
      VEC_LOOP_1_COMP_LOOP_C_108 : begin
        fsm_output = 10'b0011010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_109;
      end
      VEC_LOOP_1_COMP_LOOP_C_109 : begin
        fsm_output = 10'b0011011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_110;
      end
      VEC_LOOP_1_COMP_LOOP_C_110 : begin
        fsm_output = 10'b0011011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_111;
      end
      VEC_LOOP_1_COMP_LOOP_C_111 : begin
        fsm_output = 10'b0011011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_112;
      end
      VEC_LOOP_1_COMP_LOOP_C_112 : begin
        fsm_output = 10'b0011011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_113;
      end
      VEC_LOOP_1_COMP_LOOP_C_113 : begin
        fsm_output = 10'b0011011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_114;
      end
      VEC_LOOP_1_COMP_LOOP_C_114 : begin
        fsm_output = 10'b0011011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_115;
      end
      VEC_LOOP_1_COMP_LOOP_C_115 : begin
        fsm_output = 10'b0011011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_116;
      end
      VEC_LOOP_1_COMP_LOOP_C_116 : begin
        fsm_output = 10'b0011011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_117;
      end
      VEC_LOOP_1_COMP_LOOP_C_117 : begin
        fsm_output = 10'b0011100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_118;
      end
      VEC_LOOP_1_COMP_LOOP_C_118 : begin
        fsm_output = 10'b0011100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_119;
      end
      VEC_LOOP_1_COMP_LOOP_C_119 : begin
        fsm_output = 10'b0011100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_120;
      end
      VEC_LOOP_1_COMP_LOOP_C_120 : begin
        fsm_output = 10'b0011100011;
        if ( VEC_LOOP_1_COMP_LOOP_C_120_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_121;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_121 : begin
        fsm_output = 10'b0011100100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_0;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 10'b0011100101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_1;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 10'b0011100110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_2;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 10'b0011100111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_3;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 10'b0011101000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_4;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 10'b0011101001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_5;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 10'b0011101010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_6;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 10'b0011101011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_7;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 10'b0011101100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_8;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 10'b0011101101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_9;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 10'b0011101110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_10;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 10'b0011101111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_11;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 10'b0011110000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_12;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 10'b0011110001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_13;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 10'b0011110010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_14;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 10'b0011110011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_15;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 10'b0011110100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_16;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 10'b0011110101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_17;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 10'b0011110110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_18;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 10'b0011110111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_19;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 10'b0011111000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_20;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 10'b0011111001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_21;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 10'b0011111010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_22;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 10'b0011111011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_23;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 10'b0011111100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24;
      end
      VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 10'b0011111101;
        if ( VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_122;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_1_COMP_LOOP_C_122 : begin
        fsm_output = 10'b0011111110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_123;
      end
      VEC_LOOP_1_COMP_LOOP_C_123 : begin
        fsm_output = 10'b0011111111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_124;
      end
      VEC_LOOP_1_COMP_LOOP_C_124 : begin
        fsm_output = 10'b0100000000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_125;
      end
      VEC_LOOP_1_COMP_LOOP_C_125 : begin
        fsm_output = 10'b0100000001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_126;
      end
      VEC_LOOP_1_COMP_LOOP_C_126 : begin
        fsm_output = 10'b0100000010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_127;
      end
      VEC_LOOP_1_COMP_LOOP_C_127 : begin
        fsm_output = 10'b0100000011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_128;
      end
      VEC_LOOP_1_COMP_LOOP_C_128 : begin
        fsm_output = 10'b0100000100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_129;
      end
      VEC_LOOP_1_COMP_LOOP_C_129 : begin
        fsm_output = 10'b0100000101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_130;
      end
      VEC_LOOP_1_COMP_LOOP_C_130 : begin
        fsm_output = 10'b0100000110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_131;
      end
      VEC_LOOP_1_COMP_LOOP_C_131 : begin
        fsm_output = 10'b0100000111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_132;
      end
      VEC_LOOP_1_COMP_LOOP_C_132 : begin
        fsm_output = 10'b0100001000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_133;
      end
      VEC_LOOP_1_COMP_LOOP_C_133 : begin
        fsm_output = 10'b0100001001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_134;
      end
      VEC_LOOP_1_COMP_LOOP_C_134 : begin
        fsm_output = 10'b0100001010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_135;
      end
      VEC_LOOP_1_COMP_LOOP_C_135 : begin
        fsm_output = 10'b0100001011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_136;
      end
      VEC_LOOP_1_COMP_LOOP_C_136 : begin
        fsm_output = 10'b0100001100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_137;
      end
      VEC_LOOP_1_COMP_LOOP_C_137 : begin
        fsm_output = 10'b0100001101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_138;
      end
      VEC_LOOP_1_COMP_LOOP_C_138 : begin
        fsm_output = 10'b0100001110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_139;
      end
      VEC_LOOP_1_COMP_LOOP_C_139 : begin
        fsm_output = 10'b0100001111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_140;
      end
      VEC_LOOP_1_COMP_LOOP_C_140 : begin
        fsm_output = 10'b0100010000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_141;
      end
      VEC_LOOP_1_COMP_LOOP_C_141 : begin
        fsm_output = 10'b0100010001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_142;
      end
      VEC_LOOP_1_COMP_LOOP_C_142 : begin
        fsm_output = 10'b0100010010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_143;
      end
      VEC_LOOP_1_COMP_LOOP_C_143 : begin
        fsm_output = 10'b0100010011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_144;
      end
      VEC_LOOP_1_COMP_LOOP_C_144 : begin
        fsm_output = 10'b0100010100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_145;
      end
      VEC_LOOP_1_COMP_LOOP_C_145 : begin
        fsm_output = 10'b0100010101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_146;
      end
      VEC_LOOP_1_COMP_LOOP_C_146 : begin
        fsm_output = 10'b0100010110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_147;
      end
      VEC_LOOP_1_COMP_LOOP_C_147 : begin
        fsm_output = 10'b0100010111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_148;
      end
      VEC_LOOP_1_COMP_LOOP_C_148 : begin
        fsm_output = 10'b0100011000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_149;
      end
      VEC_LOOP_1_COMP_LOOP_C_149 : begin
        fsm_output = 10'b0100011001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_150;
      end
      VEC_LOOP_1_COMP_LOOP_C_150 : begin
        fsm_output = 10'b0100011010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_151;
      end
      VEC_LOOP_1_COMP_LOOP_C_151 : begin
        fsm_output = 10'b0100011011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_152;
      end
      VEC_LOOP_1_COMP_LOOP_C_152 : begin
        fsm_output = 10'b0100011100;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_153;
      end
      VEC_LOOP_1_COMP_LOOP_C_153 : begin
        fsm_output = 10'b0100011101;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_154;
      end
      VEC_LOOP_1_COMP_LOOP_C_154 : begin
        fsm_output = 10'b0100011110;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_155;
      end
      VEC_LOOP_1_COMP_LOOP_C_155 : begin
        fsm_output = 10'b0100011111;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_156;
      end
      VEC_LOOP_1_COMP_LOOP_C_156 : begin
        fsm_output = 10'b0100100000;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_157;
      end
      VEC_LOOP_1_COMP_LOOP_C_157 : begin
        fsm_output = 10'b0100100001;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_158;
      end
      VEC_LOOP_1_COMP_LOOP_C_158 : begin
        fsm_output = 10'b0100100010;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_159;
      end
      VEC_LOOP_1_COMP_LOOP_C_159 : begin
        fsm_output = 10'b0100100011;
        state_var_NS = VEC_LOOP_1_COMP_LOOP_C_160;
      end
      VEC_LOOP_1_COMP_LOOP_C_160 : begin
        fsm_output = 10'b0100100100;
        if ( VEC_LOOP_1_COMP_LOOP_C_160_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 10'b0100100101;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_6;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_0 : begin
        fsm_output = 10'b0100100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_C_1 : begin
        fsm_output = 10'b0100100111;
        if ( VEC_LOOP_2_COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 10'b0100101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 10'b0100101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 10'b0100101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 10'b0100101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 10'b0100101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 10'b0100101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 10'b0100101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 10'b0100101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 10'b0100110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 10'b0100110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 10'b0100110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 10'b0100110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 10'b0100110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 10'b0100110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 10'b0100110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 10'b0100110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 10'b0100111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 10'b0100111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 10'b0100111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 10'b0100111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 10'b0100111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 10'b0100111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 10'b0100111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 10'b0100111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 10'b0101000000;
        if ( VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_2 : begin
        fsm_output = 10'b0101000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_C_3 : begin
        fsm_output = 10'b0101000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_C_4 : begin
        fsm_output = 10'b0101000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_C_5 : begin
        fsm_output = 10'b0101000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_C_6 : begin
        fsm_output = 10'b0101000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_C_7 : begin
        fsm_output = 10'b0101000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_C_8 : begin
        fsm_output = 10'b0101000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_C_9 : begin
        fsm_output = 10'b0101001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_C_10 : begin
        fsm_output = 10'b0101001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_C_11 : begin
        fsm_output = 10'b0101001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_C_12 : begin
        fsm_output = 10'b0101001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_C_13 : begin
        fsm_output = 10'b0101001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_C_14 : begin
        fsm_output = 10'b0101001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_C_15 : begin
        fsm_output = 10'b0101001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_C_16 : begin
        fsm_output = 10'b0101001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_C_17 : begin
        fsm_output = 10'b0101010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_C_18 : begin
        fsm_output = 10'b0101010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_C_19 : begin
        fsm_output = 10'b0101010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_C_20 : begin
        fsm_output = 10'b0101010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_C_21 : begin
        fsm_output = 10'b0101010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_C_22 : begin
        fsm_output = 10'b0101010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_C_23 : begin
        fsm_output = 10'b0101010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_C_24 : begin
        fsm_output = 10'b0101010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_25;
      end
      VEC_LOOP_2_COMP_LOOP_C_25 : begin
        fsm_output = 10'b0101011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_26;
      end
      VEC_LOOP_2_COMP_LOOP_C_26 : begin
        fsm_output = 10'b0101011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_27;
      end
      VEC_LOOP_2_COMP_LOOP_C_27 : begin
        fsm_output = 10'b0101011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_28;
      end
      VEC_LOOP_2_COMP_LOOP_C_28 : begin
        fsm_output = 10'b0101011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_29;
      end
      VEC_LOOP_2_COMP_LOOP_C_29 : begin
        fsm_output = 10'b0101011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_30;
      end
      VEC_LOOP_2_COMP_LOOP_C_30 : begin
        fsm_output = 10'b0101011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_31;
      end
      VEC_LOOP_2_COMP_LOOP_C_31 : begin
        fsm_output = 10'b0101011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_32;
      end
      VEC_LOOP_2_COMP_LOOP_C_32 : begin
        fsm_output = 10'b0101011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_33;
      end
      VEC_LOOP_2_COMP_LOOP_C_33 : begin
        fsm_output = 10'b0101100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_34;
      end
      VEC_LOOP_2_COMP_LOOP_C_34 : begin
        fsm_output = 10'b0101100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_35;
      end
      VEC_LOOP_2_COMP_LOOP_C_35 : begin
        fsm_output = 10'b0101100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_36;
      end
      VEC_LOOP_2_COMP_LOOP_C_36 : begin
        fsm_output = 10'b0101100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_37;
      end
      VEC_LOOP_2_COMP_LOOP_C_37 : begin
        fsm_output = 10'b0101100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_38;
      end
      VEC_LOOP_2_COMP_LOOP_C_38 : begin
        fsm_output = 10'b0101100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_39;
      end
      VEC_LOOP_2_COMP_LOOP_C_39 : begin
        fsm_output = 10'b0101100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_40;
      end
      VEC_LOOP_2_COMP_LOOP_C_40 : begin
        fsm_output = 10'b0101100111;
        if ( VEC_LOOP_2_COMP_LOOP_C_40_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_41;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_41 : begin
        fsm_output = 10'b0101101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 10'b0101101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 10'b0101101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 10'b0101101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 10'b0101101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 10'b0101101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 10'b0101101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 10'b0101101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 10'b0101110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 10'b0101110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 10'b0101110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 10'b0101110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 10'b0101110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 10'b0101110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 10'b0101110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 10'b0101110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 10'b0101111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 10'b0101111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 10'b0101111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 10'b0101111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 10'b0101111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 10'b0101111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 10'b0101111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 10'b0101111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 10'b0110000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 10'b0110000001;
        if ( VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_42;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_42 : begin
        fsm_output = 10'b0110000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_43;
      end
      VEC_LOOP_2_COMP_LOOP_C_43 : begin
        fsm_output = 10'b0110000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_44;
      end
      VEC_LOOP_2_COMP_LOOP_C_44 : begin
        fsm_output = 10'b0110000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_45;
      end
      VEC_LOOP_2_COMP_LOOP_C_45 : begin
        fsm_output = 10'b0110000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_46;
      end
      VEC_LOOP_2_COMP_LOOP_C_46 : begin
        fsm_output = 10'b0110000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_47;
      end
      VEC_LOOP_2_COMP_LOOP_C_47 : begin
        fsm_output = 10'b0110000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_48;
      end
      VEC_LOOP_2_COMP_LOOP_C_48 : begin
        fsm_output = 10'b0110001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_49;
      end
      VEC_LOOP_2_COMP_LOOP_C_49 : begin
        fsm_output = 10'b0110001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_50;
      end
      VEC_LOOP_2_COMP_LOOP_C_50 : begin
        fsm_output = 10'b0110001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_51;
      end
      VEC_LOOP_2_COMP_LOOP_C_51 : begin
        fsm_output = 10'b0110001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_52;
      end
      VEC_LOOP_2_COMP_LOOP_C_52 : begin
        fsm_output = 10'b0110001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_53;
      end
      VEC_LOOP_2_COMP_LOOP_C_53 : begin
        fsm_output = 10'b0110001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_54;
      end
      VEC_LOOP_2_COMP_LOOP_C_54 : begin
        fsm_output = 10'b0110001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_55;
      end
      VEC_LOOP_2_COMP_LOOP_C_55 : begin
        fsm_output = 10'b0110001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_56;
      end
      VEC_LOOP_2_COMP_LOOP_C_56 : begin
        fsm_output = 10'b0110010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_57;
      end
      VEC_LOOP_2_COMP_LOOP_C_57 : begin
        fsm_output = 10'b0110010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_58;
      end
      VEC_LOOP_2_COMP_LOOP_C_58 : begin
        fsm_output = 10'b0110010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_59;
      end
      VEC_LOOP_2_COMP_LOOP_C_59 : begin
        fsm_output = 10'b0110010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_60;
      end
      VEC_LOOP_2_COMP_LOOP_C_60 : begin
        fsm_output = 10'b0110010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_61;
      end
      VEC_LOOP_2_COMP_LOOP_C_61 : begin
        fsm_output = 10'b0110010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_62;
      end
      VEC_LOOP_2_COMP_LOOP_C_62 : begin
        fsm_output = 10'b0110010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_63;
      end
      VEC_LOOP_2_COMP_LOOP_C_63 : begin
        fsm_output = 10'b0110010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_64;
      end
      VEC_LOOP_2_COMP_LOOP_C_64 : begin
        fsm_output = 10'b0110011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_65;
      end
      VEC_LOOP_2_COMP_LOOP_C_65 : begin
        fsm_output = 10'b0110011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_66;
      end
      VEC_LOOP_2_COMP_LOOP_C_66 : begin
        fsm_output = 10'b0110011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_67;
      end
      VEC_LOOP_2_COMP_LOOP_C_67 : begin
        fsm_output = 10'b0110011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_68;
      end
      VEC_LOOP_2_COMP_LOOP_C_68 : begin
        fsm_output = 10'b0110011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_69;
      end
      VEC_LOOP_2_COMP_LOOP_C_69 : begin
        fsm_output = 10'b0110011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_70;
      end
      VEC_LOOP_2_COMP_LOOP_C_70 : begin
        fsm_output = 10'b0110011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_71;
      end
      VEC_LOOP_2_COMP_LOOP_C_71 : begin
        fsm_output = 10'b0110011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_72;
      end
      VEC_LOOP_2_COMP_LOOP_C_72 : begin
        fsm_output = 10'b0110100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_73;
      end
      VEC_LOOP_2_COMP_LOOP_C_73 : begin
        fsm_output = 10'b0110100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_74;
      end
      VEC_LOOP_2_COMP_LOOP_C_74 : begin
        fsm_output = 10'b0110100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_75;
      end
      VEC_LOOP_2_COMP_LOOP_C_75 : begin
        fsm_output = 10'b0110100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_76;
      end
      VEC_LOOP_2_COMP_LOOP_C_76 : begin
        fsm_output = 10'b0110100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_77;
      end
      VEC_LOOP_2_COMP_LOOP_C_77 : begin
        fsm_output = 10'b0110100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_78;
      end
      VEC_LOOP_2_COMP_LOOP_C_78 : begin
        fsm_output = 10'b0110100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_79;
      end
      VEC_LOOP_2_COMP_LOOP_C_79 : begin
        fsm_output = 10'b0110100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_80;
      end
      VEC_LOOP_2_COMP_LOOP_C_80 : begin
        fsm_output = 10'b0110101000;
        if ( VEC_LOOP_2_COMP_LOOP_C_80_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_81;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_81 : begin
        fsm_output = 10'b0110101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_0;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 10'b0110101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 10'b0110101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 10'b0110101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 10'b0110101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 10'b0110101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 10'b0110101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 10'b0110110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 10'b0110110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 10'b0110110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 10'b0110110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 10'b0110110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 10'b0110110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 10'b0110110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 10'b0110110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 10'b0110111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 10'b0110111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 10'b0110111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 10'b0110111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 10'b0110111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 10'b0110111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 10'b0110111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 10'b0110111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 10'b0111000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 10'b0111000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 10'b0111000010;
        if ( VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_82;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_82 : begin
        fsm_output = 10'b0111000011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_83;
      end
      VEC_LOOP_2_COMP_LOOP_C_83 : begin
        fsm_output = 10'b0111000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_84;
      end
      VEC_LOOP_2_COMP_LOOP_C_84 : begin
        fsm_output = 10'b0111000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_85;
      end
      VEC_LOOP_2_COMP_LOOP_C_85 : begin
        fsm_output = 10'b0111000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_86;
      end
      VEC_LOOP_2_COMP_LOOP_C_86 : begin
        fsm_output = 10'b0111000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_87;
      end
      VEC_LOOP_2_COMP_LOOP_C_87 : begin
        fsm_output = 10'b0111001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_88;
      end
      VEC_LOOP_2_COMP_LOOP_C_88 : begin
        fsm_output = 10'b0111001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_89;
      end
      VEC_LOOP_2_COMP_LOOP_C_89 : begin
        fsm_output = 10'b0111001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_90;
      end
      VEC_LOOP_2_COMP_LOOP_C_90 : begin
        fsm_output = 10'b0111001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_91;
      end
      VEC_LOOP_2_COMP_LOOP_C_91 : begin
        fsm_output = 10'b0111001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_92;
      end
      VEC_LOOP_2_COMP_LOOP_C_92 : begin
        fsm_output = 10'b0111001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_93;
      end
      VEC_LOOP_2_COMP_LOOP_C_93 : begin
        fsm_output = 10'b0111001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_94;
      end
      VEC_LOOP_2_COMP_LOOP_C_94 : begin
        fsm_output = 10'b0111001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_95;
      end
      VEC_LOOP_2_COMP_LOOP_C_95 : begin
        fsm_output = 10'b0111010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_96;
      end
      VEC_LOOP_2_COMP_LOOP_C_96 : begin
        fsm_output = 10'b0111010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_97;
      end
      VEC_LOOP_2_COMP_LOOP_C_97 : begin
        fsm_output = 10'b0111010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_98;
      end
      VEC_LOOP_2_COMP_LOOP_C_98 : begin
        fsm_output = 10'b0111010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_99;
      end
      VEC_LOOP_2_COMP_LOOP_C_99 : begin
        fsm_output = 10'b0111010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_100;
      end
      VEC_LOOP_2_COMP_LOOP_C_100 : begin
        fsm_output = 10'b0111010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_101;
      end
      VEC_LOOP_2_COMP_LOOP_C_101 : begin
        fsm_output = 10'b0111010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_102;
      end
      VEC_LOOP_2_COMP_LOOP_C_102 : begin
        fsm_output = 10'b0111010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_103;
      end
      VEC_LOOP_2_COMP_LOOP_C_103 : begin
        fsm_output = 10'b0111011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_104;
      end
      VEC_LOOP_2_COMP_LOOP_C_104 : begin
        fsm_output = 10'b0111011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_105;
      end
      VEC_LOOP_2_COMP_LOOP_C_105 : begin
        fsm_output = 10'b0111011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_106;
      end
      VEC_LOOP_2_COMP_LOOP_C_106 : begin
        fsm_output = 10'b0111011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_107;
      end
      VEC_LOOP_2_COMP_LOOP_C_107 : begin
        fsm_output = 10'b0111011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_108;
      end
      VEC_LOOP_2_COMP_LOOP_C_108 : begin
        fsm_output = 10'b0111011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_109;
      end
      VEC_LOOP_2_COMP_LOOP_C_109 : begin
        fsm_output = 10'b0111011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_110;
      end
      VEC_LOOP_2_COMP_LOOP_C_110 : begin
        fsm_output = 10'b0111011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_111;
      end
      VEC_LOOP_2_COMP_LOOP_C_111 : begin
        fsm_output = 10'b0111100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_112;
      end
      VEC_LOOP_2_COMP_LOOP_C_112 : begin
        fsm_output = 10'b0111100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_113;
      end
      VEC_LOOP_2_COMP_LOOP_C_113 : begin
        fsm_output = 10'b0111100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_114;
      end
      VEC_LOOP_2_COMP_LOOP_C_114 : begin
        fsm_output = 10'b0111100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_115;
      end
      VEC_LOOP_2_COMP_LOOP_C_115 : begin
        fsm_output = 10'b0111100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_116;
      end
      VEC_LOOP_2_COMP_LOOP_C_116 : begin
        fsm_output = 10'b0111100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_117;
      end
      VEC_LOOP_2_COMP_LOOP_C_117 : begin
        fsm_output = 10'b0111100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_118;
      end
      VEC_LOOP_2_COMP_LOOP_C_118 : begin
        fsm_output = 10'b0111100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_119;
      end
      VEC_LOOP_2_COMP_LOOP_C_119 : begin
        fsm_output = 10'b0111101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_120;
      end
      VEC_LOOP_2_COMP_LOOP_C_120 : begin
        fsm_output = 10'b0111101001;
        if ( VEC_LOOP_2_COMP_LOOP_C_120_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_121;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_121 : begin
        fsm_output = 10'b0111101010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_0;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 10'b0111101011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_1;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 10'b0111101100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_2;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 10'b0111101101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_3;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 10'b0111101110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_4;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 10'b0111101111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_5;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 10'b0111110000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_6;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 10'b0111110001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_7;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 10'b0111110010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_8;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 10'b0111110011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_9;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 10'b0111110100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_10;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 10'b0111110101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_11;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 10'b0111110110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_12;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 10'b0111110111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_13;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 10'b0111111000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_14;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 10'b0111111001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_15;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 10'b0111111010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_16;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 10'b0111111011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_17;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 10'b0111111100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_18;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 10'b0111111101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_19;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 10'b0111111110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_20;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 10'b0111111111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_21;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 10'b1000000000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_22;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 10'b1000000001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_23;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 10'b1000000010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24;
      end
      VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 10'b1000000011;
        if ( VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0 ) begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_122;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      VEC_LOOP_2_COMP_LOOP_C_122 : begin
        fsm_output = 10'b1000000100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_123;
      end
      VEC_LOOP_2_COMP_LOOP_C_123 : begin
        fsm_output = 10'b1000000101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_124;
      end
      VEC_LOOP_2_COMP_LOOP_C_124 : begin
        fsm_output = 10'b1000000110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_125;
      end
      VEC_LOOP_2_COMP_LOOP_C_125 : begin
        fsm_output = 10'b1000000111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_126;
      end
      VEC_LOOP_2_COMP_LOOP_C_126 : begin
        fsm_output = 10'b1000001000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_127;
      end
      VEC_LOOP_2_COMP_LOOP_C_127 : begin
        fsm_output = 10'b1000001001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_128;
      end
      VEC_LOOP_2_COMP_LOOP_C_128 : begin
        fsm_output = 10'b1000001010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_129;
      end
      VEC_LOOP_2_COMP_LOOP_C_129 : begin
        fsm_output = 10'b1000001011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_130;
      end
      VEC_LOOP_2_COMP_LOOP_C_130 : begin
        fsm_output = 10'b1000001100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_131;
      end
      VEC_LOOP_2_COMP_LOOP_C_131 : begin
        fsm_output = 10'b1000001101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_132;
      end
      VEC_LOOP_2_COMP_LOOP_C_132 : begin
        fsm_output = 10'b1000001110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_133;
      end
      VEC_LOOP_2_COMP_LOOP_C_133 : begin
        fsm_output = 10'b1000001111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_134;
      end
      VEC_LOOP_2_COMP_LOOP_C_134 : begin
        fsm_output = 10'b1000010000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_135;
      end
      VEC_LOOP_2_COMP_LOOP_C_135 : begin
        fsm_output = 10'b1000010001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_136;
      end
      VEC_LOOP_2_COMP_LOOP_C_136 : begin
        fsm_output = 10'b1000010010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_137;
      end
      VEC_LOOP_2_COMP_LOOP_C_137 : begin
        fsm_output = 10'b1000010011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_138;
      end
      VEC_LOOP_2_COMP_LOOP_C_138 : begin
        fsm_output = 10'b1000010100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_139;
      end
      VEC_LOOP_2_COMP_LOOP_C_139 : begin
        fsm_output = 10'b1000010101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_140;
      end
      VEC_LOOP_2_COMP_LOOP_C_140 : begin
        fsm_output = 10'b1000010110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_141;
      end
      VEC_LOOP_2_COMP_LOOP_C_141 : begin
        fsm_output = 10'b1000010111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_142;
      end
      VEC_LOOP_2_COMP_LOOP_C_142 : begin
        fsm_output = 10'b1000011000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_143;
      end
      VEC_LOOP_2_COMP_LOOP_C_143 : begin
        fsm_output = 10'b1000011001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_144;
      end
      VEC_LOOP_2_COMP_LOOP_C_144 : begin
        fsm_output = 10'b1000011010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_145;
      end
      VEC_LOOP_2_COMP_LOOP_C_145 : begin
        fsm_output = 10'b1000011011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_146;
      end
      VEC_LOOP_2_COMP_LOOP_C_146 : begin
        fsm_output = 10'b1000011100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_147;
      end
      VEC_LOOP_2_COMP_LOOP_C_147 : begin
        fsm_output = 10'b1000011101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_148;
      end
      VEC_LOOP_2_COMP_LOOP_C_148 : begin
        fsm_output = 10'b1000011110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_149;
      end
      VEC_LOOP_2_COMP_LOOP_C_149 : begin
        fsm_output = 10'b1000011111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_150;
      end
      VEC_LOOP_2_COMP_LOOP_C_150 : begin
        fsm_output = 10'b1000100000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_151;
      end
      VEC_LOOP_2_COMP_LOOP_C_151 : begin
        fsm_output = 10'b1000100001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_152;
      end
      VEC_LOOP_2_COMP_LOOP_C_152 : begin
        fsm_output = 10'b1000100010;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_153;
      end
      VEC_LOOP_2_COMP_LOOP_C_153 : begin
        fsm_output = 10'b1000100011;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_154;
      end
      VEC_LOOP_2_COMP_LOOP_C_154 : begin
        fsm_output = 10'b1000100100;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_155;
      end
      VEC_LOOP_2_COMP_LOOP_C_155 : begin
        fsm_output = 10'b1000100101;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_156;
      end
      VEC_LOOP_2_COMP_LOOP_C_156 : begin
        fsm_output = 10'b1000100110;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_157;
      end
      VEC_LOOP_2_COMP_LOOP_C_157 : begin
        fsm_output = 10'b1000100111;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_158;
      end
      VEC_LOOP_2_COMP_LOOP_C_158 : begin
        fsm_output = 10'b1000101000;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_159;
      end
      VEC_LOOP_2_COMP_LOOP_C_159 : begin
        fsm_output = 10'b1000101001;
        state_var_NS = VEC_LOOP_2_COMP_LOOP_C_160;
      end
      VEC_LOOP_2_COMP_LOOP_C_160 : begin
        fsm_output = 10'b1000101010;
        if ( VEC_LOOP_2_COMP_LOOP_C_160_tr0 ) begin
          state_var_NS = VEC_LOOP_C_1;
        end
        else begin
          state_var_NS = VEC_LOOP_2_COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_1 : begin
        fsm_output = 10'b1000101011;
        if ( VEC_LOOP_C_1_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_6;
        end
        else begin
          state_var_NS = VEC_LOOP_1_COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 10'b1000101100;
        if ( STAGE_LOOP_C_6_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 10'b1000101101;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 10'b0000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [9:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [9:0] fsm_output;
  wire or_tmp_29;
  wire or_tmp_31;
  wire or_tmp_51;
  wire or_tmp_61;
  wire or_tmp_71;
  wire or_tmp_72;
  wire mux_tmp_72;
  wire or_tmp_77;
  wire or_tmp_79;
  wire mux_tmp_84;
  wire mux_tmp_86;
  wire mux_tmp_92;
  wire and_dcpl_13;
  wire nor_tmp_34;
  wire not_tmp_77;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire and_dcpl_43;
  wire and_dcpl_44;
  wire and_dcpl_45;
  wire and_dcpl_46;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire nor_tmp_40;
  wire not_tmp_91;
  wire mux_tmp_162;
  wire or_tmp_148;
  wire and_dcpl_60;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_76;
  wire and_dcpl_82;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire not_tmp_108;
  wire or_tmp_264;
  wire or_tmp_278;
  wire or_tmp_321;
  wire or_tmp_334;
  wire or_tmp_374;
  wire or_tmp_387;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire mux_tmp_317;
  wire mux_tmp_318;
  wire or_tmp_404;
  wire mux_tmp_319;
  wire nor_tmp_63;
  wire nor_tmp_64;
  wire or_tmp_415;
  wire mux_tmp_325;
  wire mux_tmp_329;
  wire mux_tmp_335;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire mux_tmp_340;
  wire or_tmp_416;
  wire mux_tmp_345;
  wire mux_tmp_350;
  wire mux_tmp_373;
  wire or_tmp_421;
  wire or_tmp_423;
  wire or_tmp_426;
  wire mux_tmp_375;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_382;
  wire or_tmp_436;
  wire or_tmp_437;
  wire or_tmp_438;
  wire mux_tmp_393;
  wire not_tmp_170;
  wire mux_tmp_398;
  wire and_dcpl_105;
  wire and_dcpl_107;
  wire not_tmp_173;
  wire or_tmp_449;
  wire or_tmp_451;
  wire or_tmp_455;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire mux_tmp_431;
  wire and_tmp_6;
  wire or_tmp_470;
  wire nand_tmp_42;
  wire and_dcpl_111;
  wire and_dcpl_117;
  wire or_tmp_476;
  wire and_tmp_7;
  wire and_dcpl_119;
  wire and_dcpl_123;
  wire or_tmp_483;
  wire mux_tmp_440;
  wire or_tmp_484;
  wire and_tmp_8;
  wire mux_tmp_448;
  wire mux_tmp_455;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_134;
  wire mux_tmp_504;
  wire and_dcpl_138;
  wire nor_tmp_81;
  wire mux_tmp_506;
  wire nor_tmp_83;
  wire mux_tmp_509;
  wire or_tmp_539;
  wire nor_tmp_86;
  wire mux_tmp_522;
  wire or_tmp_548;
  wire mux_tmp_530;
  wire not_tmp_231;
  wire or_tmp_562;
  wire mux_tmp_537;
  wire or_tmp_567;
  wire mux_tmp_546;
  wire mux_tmp_549;
  wire or_tmp_573;
  wire and_dcpl_147;
  wire mux_tmp_579;
  wire and_dcpl_154;
  wire not_tmp_260;
  wire or_tmp_621;
  wire or_tmp_623;
  wire mux_tmp_588;
  wire mux_tmp_589;
  wire mux_tmp_594;
  wire mux_tmp_599;
  wire or_tmp_635;
  wire or_tmp_637;
  wire nor_tmp_103;
  wire mux_tmp_624;
  wire or_tmp_654;
  wire or_tmp_656;
  wire mux_tmp_637;
  wire or_tmp_670;
  wire mux_tmp_668;
  wire mux_tmp_711;
  wire mux_tmp_722;
  wire or_tmp_716;
  wire mux_tmp_723;
  wire and_tmp_14;
  wire and_dcpl_175;
  wire not_tmp_321;
  wire or_tmp_760;
  wire mux_tmp_760;
  wire or_tmp_762;
  wire or_tmp_769;
  wire mux_tmp_763;
  wire mux_tmp_771;
  wire and_dcpl_176;
  wire not_tmp_324;
  wire and_dcpl_179;
  wire mux_tmp_787;
  reg exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva;
  reg VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  reg [11:0] VEC_LOOP_j_1_12_0_sva_11_0;
  reg VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_5_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [10:0] COMP_LOOP_acc_11_psp_1_sva;
  wire [11:0] nl_COMP_LOOP_acc_11_psp_1_sva;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [6:0] COMP_LOOP_k_9_2_1_sva_6_0;
  reg [63:0] tmp_10_lpi_4_dfm;
  reg [11:0] reg_VEC_LOOP_1_acc_1_psp_ftd_1;
  wire and_160_m1c;
  wire and_163_m1c;
  wire and_141_m1c;
  wire nor_359_m1c;
  wire nand_95_cse;
  wire or_304_cse;
  wire nor_269_cse;
  wire or_315_cse;
  wire and_270_cse;
  reg reg_vec_rsc_triosy_0_3_obj_ld_cse;
  wire nor_70_cse;
  wire and_256_cse;
  wire or_590_cse;
  wire and_300_cse;
  wire or_94_cse;
  wire and_205_cse;
  wire or_814_cse;
  wire or_913_cse;
  wire nor_236_cse;
  wire or_596_cse;
  wire or_369_cse;
  wire nor_268_cse;
  wire or_370_cse;
  wire nor_241_cse;
  wire and_303_cse;
  wire or_756_cse;
  wire nand_119_cse;
  wire or_55_cse;
  wire or_826_cse;
  wire or_899_cse;
  wire and_213_cse;
  wire nor_330_cse;
  wire or_154_cse;
  wire or_54_cse;
  wire nor_312_cse;
  wire mux_190_cse;
  wire mux_189_cse;
  wire mux_186_cse;
  wire mux_561_cse;
  wire mux_560_cse;
  wire mux_749_cse;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire mux_258_cse;
  wire mux_748_cse;
  wire mux_745_cse;
  reg [9:0] COMP_LOOP_acc_psp_1_sva;
  wire [63:0] modExp_base_1_sva_mx1;
  wire modExp_while_and_3;
  wire modExp_while_and_5;
  wire mux_423_itm;
  wire mux_433_itm;
  wire mux_801_itm;
  wire and_dcpl_196;
  wire or_tmp_841;
  wire mux_tmp_824;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_204;
  wire and_dcpl_208;
  wire and_dcpl_215;
  wire and_dcpl_221;
  wire [9:0] z_out_1;
  wire [10:0] nl_z_out_1;
  wire and_dcpl_230;
  wire and_dcpl_242;
  wire and_dcpl_244;
  wire [11:0] z_out_2;
  wire and_dcpl_253;
  wire [11:0] z_out_3;
  wire [12:0] nl_z_out_3;
  wire or_tmp_858;
  wire mux_tmp_833;
  wire and_dcpl_283;
  wire and_dcpl_288;
  wire and_dcpl_292;
  wire and_dcpl_302;
  wire and_dcpl_310;
  wire [64:0] z_out_5;
  wire [65:0] nl_z_out_5;
  wire and_dcpl_314;
  wire and_dcpl_315;
  wire and_dcpl_316;
  wire and_dcpl_319;
  wire not_tmp_415;
  wire mux_tmp_843;
  wire mux_tmp_844;
  wire mux_tmp_845;
  wire mux_tmp_849;
  wire and_dcpl_321;
  wire and_dcpl_323;
  wire and_dcpl_325;
  wire and_dcpl_326;
  wire and_dcpl_327;
  wire and_dcpl_331;
  wire and_dcpl_333;
  wire and_dcpl_334;
  wire and_dcpl_338;
  wire and_dcpl_339;
  wire and_dcpl_342;
  wire and_dcpl_343;
  wire and_dcpl_345;
  wire and_dcpl_346;
  wire and_dcpl_349;
  wire and_dcpl_351;
  wire and_dcpl_352;
  wire and_dcpl_354;
  wire and_dcpl_356;
  wire and_dcpl_357;
  wire and_dcpl_361;
  wire and_dcpl_367;
  wire [63:0] z_out_6;
  wire [64:0] nl_z_out_6;
  wire mux_tmp_860;
  wire or_tmp_890;
  wire mux_tmp_866;
  wire [63:0] z_out_7;
  wire [127:0] nl_z_out_7;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg modExp_exp_1_3_1_sva;
  reg modExp_exp_1_2_1_sva;
  reg modExp_exp_1_1_1_sva;
  reg modExp_exp_1_0_1_sva_1;
  reg [63:0] modExp_base_1_sva;
  reg [63:0] VEC_LOOP_1_COMP_LOOP_1_acc_8_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_1_12_0_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire COMP_LOOP_or_1_cse;
  wire COMP_LOOP_or_3_cse;
  wire or_254_cse;
  wire or_614_cse;
  wire or_611_cse;
  wire mux_680_cse;
  wire nor_332_cse;
  wire STAGE_LOOP_or_ssc;
  wire and_365_cse;
  wire and_392_cse;
  wire mux_165_cse;
  wire mux_163_cse;
  wire or_tmp_911;
  wire mux_tmp_877;
  wire or_tmp_917;
  wire or_tmp_923;
  wire mux_tmp_886;
  wire or_tmp_942;
  wire mux_tmp_907;
  wire mux_tmp_910;
  wire or_tmp_948;
  wire or_tmp_949;
  wire or_tmp_952;
  wire mux_tmp_915;
  wire or_tmp_953;
  wire mux_tmp_916;
  wire mux_tmp_919;
  wire mux_tmp_921;
  wire or_tmp_960;
  wire [64:0] operator_64_false_mux1h_2_rgt;
  wire or_tmp_971;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire and_524_cse;
  wire or_1038_cse;
  wire or_1047_cse;
  wire or_462_cse;
  wire mux_894_cse;
  wire mux_860_itm;
  wire mux_866_itm;
  wire operator_64_false_1_or_2_itm;
  wire COMP_LOOP_or_27_itm;
  wire STAGE_LOOP_nor_itm;
  wire STAGE_LOOP_nor_53_itm;
  wire STAGE_LOOP_or_1_itm;
  wire STAGE_LOOP_or_2_itm;
  wire mux_826_cse;

  wire[0:0] mux_188_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] or_237_nl;
  wire[0:0] or_236_nl;
  wire[0:0] mux_185_nl;
  wire[0:0] mux_184_nl;
  wire[0:0] or_231_nl;
  wire[0:0] or_228_nl;
  wire[0:0] nand_12_nl;
  wire[0:0] or_234_nl;
  wire[0:0] and_275_nl;
  wire[0:0] nor_260_nl;
  wire[0:0] modulo_result_or_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] or_452_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nor_237_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] or_446_nl;
  wire[0:0] or_443_nl;
  wire[0:0] nor_239_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] or_439_nl;
  wire[0:0] or_436_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] or_477_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] or_474_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] or_469_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] nor_228_nl;
  wire[63:0] mux1h_nl;
  wire[0:0] or_994_nl;
  wire[0:0] mux_672_nl;
  wire[0:0] nor_178_nl;
  wire[0:0] mux_671_nl;
  wire[0:0] mux_670_nl;
  wire[0:0] or_709_nl;
  wire[0:0] and_225_nl;
  wire[0:0] mux_669_nl;
  wire[0:0] mux_667_nl;
  wire[0:0] or_705_nl;
  wire[0:0] or_703_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] mux_664_nl;
  wire[0:0] mux_661_nl;
  wire[0:0] mux_660_nl;
  wire[0:0] mux_659_nl;
  wire[0:0] mux_658_nl;
  wire[0:0] or_702_nl;
  wire[0:0] mux_657_nl;
  wire[0:0] mux_656_nl;
  wire[0:0] or_701_nl;
  wire[0:0] mux_650_nl;
  wire[0:0] mux_649_nl;
  wire[0:0] or_699_nl;
  wire[0:0] mux_648_nl;
  wire[0:0] mux_647_nl;
  wire[0:0] mux_639_nl;
  wire[0:0] mux_638_nl;
  wire[0:0] or_695_nl;
  wire[0:0] mux_628_nl;
  wire[0:0] mux_627_nl;
  wire[0:0] mux_626_nl;
  wire[0:0] mux_625_nl;
  wire[0:0] modExp_while_if_and_1_nl;
  wire[0:0] modExp_while_if_and_2_nl;
  wire[0:0] and_126_nl;
  wire[0:0] mux_463_nl;
  wire[0:0] mux_462_nl;
  wire[0:0] mux_461_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] nor_222_nl;
  wire[0:0] mux_459_nl;
  wire[0:0] mux_458_nl;
  wire[0:0] mux_457_nl;
  wire[0:0] or_533_nl;
  wire[0:0] mux_456_nl;
  wire[0:0] nor_223_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] nor_224_nl;
  wire[0:0] mux_453_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] nor_225_nl;
  wire[0:0] or_527_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] or_526_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] or_524_nl;
  wire[0:0] or_523_nl;
  wire[0:0] or_522_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] or_520_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] or_519_nl;
  wire[0:0] or_1035_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] or_1037_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] or_1036_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] and_525_nl;
  wire[0:0] or_1032_nl;
  wire[0:0] or_1028_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] or_1018_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] or_1011_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] or_1063_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] nand_nl;
  wire[0:0] or_1061_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] or_1059_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] or_1055_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] nand_145_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] or_1054_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] or_1052_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] or_1051_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] or_1042_nl;
  wire[0:0] mux_911_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] or_1041_nl;
  wire[0:0] or_992_nl;
  wire[0:0] mux_478_nl;
  wire[0:0] nand_117_nl;
  wire[0:0] or_912_nl;
  wire[0:0] mux_477_nl;
  wire[0:0] mux_476_nl;
  wire[0:0] or_548_nl;
  wire[0:0] nand_85_nl;
  wire[0:0] or_546_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] or_1069_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] or_1067_nl;
  wire[0:0] nand_143_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] mux_500_nl;
  wire[0:0] or_897_nl;
  wire[0:0] mux_499_nl;
  wire[0:0] or_563_nl;
  wire[0:0] or_562_nl;
  wire[0:0] mux_498_nl;
  wire[0:0] nor_216_nl;
  wire[0:0] and_144_nl;
  wire[0:0] r_or_nl;
  wire[0:0] r_or_1_nl;
  wire[0:0] mux_529_nl;
  wire[0:0] mux_528_nl;
  wire[0:0] mux_527_nl;
  wire[0:0] mux_526_nl;
  wire[0:0] and_240_nl;
  wire[0:0] mux_525_nl;
  wire[0:0] mux_524_nl;
  wire[0:0] mux_523_nl;
  wire[0:0] mux_521_nl;
  wire[0:0] mux_520_nl;
  wire[0:0] mux_519_nl;
  wire[0:0] nor_209_nl;
  wire[0:0] and_149_nl;
  wire[0:0] mux_518_nl;
  wire[0:0] mux_517_nl;
  wire[0:0] mux_516_nl;
  wire[0:0] mux_515_nl;
  wire[0:0] or_581_nl;
  wire[0:0] mux_514_nl;
  wire[0:0] or_579_nl;
  wire[0:0] mux_513_nl;
  wire[0:0] or_577_nl;
  wire[0:0] mux_512_nl;
  wire[0:0] and_148_nl;
  wire[0:0] mux_511_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] mux_507_nl;
  wire[0:0] nor_325_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] mux_563_nl;
  wire[0:0] and_235_nl;
  wire[0:0] mux_562_nl;
  wire[0:0] nor_203_nl;
  wire[0:0] nor_204_nl;
  wire[0:0] nor_205_nl;
  wire[0:0] mux_559_nl;
  wire[0:0] or_607_nl;
  wire[0:0] or_606_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] mux_568_nl;
  wire[0:0] and_234_nl;
  wire[0:0] mux_567_nl;
  wire[0:0] nor_200_nl;
  wire[0:0] nor_201_nl;
  wire[0:0] nor_202_nl;
  wire[0:0] mux_564_nl;
  wire[0:0] or_618_nl;
  wire[0:0] or_617_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] mux_573_nl;
  wire[0:0] and_233_nl;
  wire[0:0] mux_572_nl;
  wire[0:0] nor_197_nl;
  wire[0:0] nor_198_nl;
  wire[0:0] nor_199_nl;
  wire[0:0] mux_569_nl;
  wire[0:0] or_629_nl;
  wire[0:0] or_628_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] mux_578_nl;
  wire[0:0] and_230_nl;
  wire[0:0] mux_577_nl;
  wire[0:0] and_231_nl;
  wire[0:0] and_232_nl;
  wire[0:0] nor_196_nl;
  wire[0:0] mux_574_nl;
  wire[0:0] or_636_nl;
  wire[0:0] or_635_nl;
  wire[0:0] mux_557_nl;
  wire[0:0] mux_556_nl;
  wire[0:0] mux_555_nl;
  wire[0:0] mux_554_nl;
  wire[0:0] mux_553_nl;
  wire[0:0] mux_552_nl;
  wire[0:0] mux_551_nl;
  wire[0:0] mux_550_nl;
  wire[0:0] mux_548_nl;
  wire[0:0] mux_547_nl;
  wire[0:0] mux_545_nl;
  wire[0:0] mux_544_nl;
  wire[0:0] mux_543_nl;
  wire[0:0] mux_542_nl;
  wire[0:0] mux_541_nl;
  wire[0:0] mux_540_nl;
  wire[0:0] mux_539_nl;
  wire[0:0] or_603_nl;
  wire[0:0] or_601_nl;
  wire[0:0] mux_538_nl;
  wire[0:0] mux_536_nl;
  wire[0:0] or_598_nl;
  wire[0:0] or_1002_nl;
  wire[0:0] mux_535_nl;
  wire[0:0] or_594_nl;
  wire[0:0] mux_534_nl;
  wire[0:0] or_593_nl;
  wire[0:0] or_592_nl;
  wire[0:0] or_591_nl;
  wire[0:0] COMP_LOOP_mux1h_15_nl;
  wire[8:0] acc_nl;
  wire[9:0] nl_acc_nl;
  wire[6:0] operator_64_false_1_mux_3_nl;
  wire[0:0] operator_64_false_1_or_5_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] and_531_nl;
  wire[6:0] operator_64_false_1_mux_4_nl;
  wire[0:0] COMP_LOOP_and_11_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] mux_616_nl;
  wire[0:0] nor_184_nl;
  wire[0:0] nor_185_nl;
  wire[0:0] mux_615_nl;
  wire[0:0] mux_614_nl;
  wire[0:0] mux_613_nl;
  wire[0:0] mux_612_nl;
  wire[0:0] mux_611_nl;
  wire[0:0] mux_610_nl;
  wire[0:0] mux_609_nl;
  wire[0:0] mux_608_nl;
  wire[0:0] or_673_nl;
  wire[0:0] mux_607_nl;
  wire[0:0] mux_606_nl;
  wire[0:0] mux_605_nl;
  wire[0:0] mux_604_nl;
  wire[0:0] mux_603_nl;
  wire[0:0] or_671_nl;
  wire[0:0] mux_602_nl;
  wire[0:0] mux_601_nl;
  wire[0:0] mux_600_nl;
  wire[0:0] mux_597_nl;
  wire[0:0] mux_596_nl;
  wire[0:0] mux_595_nl;
  wire[0:0] or_665_nl;
  wire[0:0] mux_593_nl;
  wire[0:0] or_71_nl;
  wire[0:0] mux_592_nl;
  wire[0:0] mux_591_nl;
  wire[0:0] or_662_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] mux_590_nl;
  wire[0:0] or_661_nl;
  wire[0:0] nor_186_nl;
  wire[0:0] mux_587_nl;
  wire[0:0] or_656_nl;
  wire[0:0] or_655_nl;
  wire[9:0] VEC_LOOP_1_COMP_LOOP_1_acc_11_nl;
  wire[10:0] nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl;
  wire[0:0] and_221_nl;
  wire[0:0] nor_174_nl;
  wire[63:0] VEC_LOOP_1_COMP_LOOP_1_acc_8_nl;
  wire[64:0] nl_VEC_LOOP_1_COMP_LOOP_1_acc_8_nl;
  wire[0:0] mux_682_nl;
  wire[0:0] nor_173_nl;
  wire[0:0] mux_681_nl;
  wire[0:0] or_721_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] mux_679_nl;
  wire[0:0] and_222_nl;
  wire[0:0] mux_678_nl;
  wire[0:0] nor_175_nl;
  wire[0:0] and_223_nl;
  wire[0:0] and_224_nl;
  wire[0:0] mux_677_nl;
  wire[0:0] nor_176_nl;
  wire[0:0] nor_177_nl;
  wire[0:0] mux_709_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] and_297_nl;
  wire[0:0] mux_702_nl;
  wire[0:0] mux_701_nl;
  wire[0:0] mux_700_nl;
  wire[0:0] mux_699_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] or_93_nl;
  wire[10:0] COMP_LOOP_mux_42_nl;
  wire[0:0] mux_721_nl;
  wire[0:0] mux_720_nl;
  wire[0:0] mux_719_nl;
  wire[0:0] mux_718_nl;
  wire[0:0] mux_717_nl;
  wire[0:0] mux_716_nl;
  wire[0:0] or_758_nl;
  wire[0:0] mux_715_nl;
  wire[0:0] mux_714_nl;
  wire[0:0] mux_713_nl;
  wire[0:0] or_757_nl;
  wire[0:0] mux_712_nl;
  wire[0:0] and_217_nl;
  wire[0:0] mux_731_nl;
  wire[0:0] nor_171_nl;
  wire[0:0] mux_730_nl;
  wire[0:0] or_763_nl;
  wire[0:0] or_762_nl;
  wire[0:0] or_761_nl;
  wire[0:0] mux_729_nl;
  wire[0:0] mux_728_nl;
  wire[0:0] mux_727_nl;
  wire[0:0] mux_726_nl;
  wire[0:0] mux_725_nl;
  wire[0:0] mux_724_nl;
  wire[0:0] or_787_nl;
  wire[0:0] mux_747_nl;
  wire[0:0] mux_746_nl;
  wire[0:0] or_786_nl;
  wire[0:0] or_785_nl;
  wire[0:0] or_780_nl;
  wire[0:0] COMP_LOOP_mux_39_nl;
  wire[0:0] mux_751_nl;
  wire[0:0] mux_750_nl;
  wire[0:0] or_890_nl;
  wire[0:0] mux_732_nl;
  wire[0:0] and_212_nl;
  wire[0:0] nor_170_nl;
  wire[0:0] mux_752_nl;
  wire[0:0] and_210_nl;
  wire[0:0] nor_165_nl;
  wire[0:0] COMP_LOOP_mux1h_27_nl;
  wire[0:0] mux_782_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] mux_780_nl;
  wire[0:0] mux_779_nl;
  wire[0:0] mux_778_nl;
  wire[0:0] mux_777_nl;
  wire[0:0] mux_776_nl;
  wire[0:0] mux_775_nl;
  wire[0:0] mux_774_nl;
  wire[0:0] mux_773_nl;
  wire[0:0] mux_772_nl;
  wire[0:0] mux_769_nl;
  wire[0:0] mux_768_nl;
  wire[0:0] or_824_nl;
  wire[0:0] or_820_nl;
  wire[0:0] mux_767_nl;
  wire[0:0] mux_766_nl;
  wire[0:0] mux_765_nl;
  wire[0:0] mux_764_nl;
  wire[0:0] mux_762_nl;
  wire[0:0] mux_761_nl;
  wire[0:0] or_810_nl;
  wire[0:0] COMP_LOOP_mux1h_44_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] or_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] or_989_nl;
  wire[0:0] or_990_nl;
  wire[0:0] or_991_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] or_852_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] or_851_nl;
  wire[0:0] or_850_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] nor_142_nl;
  wire[0:0] nor_143_nl;
  wire[0:0] or_91_nl;
  wire[0:0] or_103_nl;
  wire[0:0] or_102_nl;
  wire[0:0] mux_158_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] or_901_nl;
  wire[0:0] nand_100_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] nor_310_nl;
  wire[0:0] nor_311_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] or_467_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] or_465_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] or_475_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] nor_232_nl;
  wire[0:0] nor_233_nl;
  wire[0:0] nand_40_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] nand_39_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] or_909_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] nand_87_nl;
  wire[0:0] or_498_nl;
  wire[0:0] or_496_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] or_910_nl;
  wire[0:0] or_911_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] or_491_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] or_503_nl;
  wire[0:0] or_501_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] or_508_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] or_507_nl;
  wire[0:0] or_505_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] nor_227_nl;
  wire[0:0] and_253_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] or_531_nl;
  wire[0:0] mux_673_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] mux_503_nl;
  wire[0:0] or_571_nl;
  wire[0:0] or_570_nl;
  wire[0:0] mux_505_nl;
  wire[0:0] or_572_nl;
  wire[0:0] and_306_nl;
  wire[0:0] mux_508_nl;
  wire[0:0] nor_211_nl;
  wire[0:0] or_587_nl;
  wire[0:0] nor_208_nl;
  wire[0:0] and_239_nl;
  wire[0:0] mux_532_nl;
  wire[0:0] mux_531_nl;
  wire[0:0] or_588_nl;
  wire[0:0] or_600_nl;
  wire[0:0] nor_nl;
  wire[0:0] mux_585_nl;
  wire[0:0] mux_584_nl;
  wire[0:0] nor_189_nl;
  wire[0:0] nor_190_nl;
  wire[0:0] mux_583_nl;
  wire[0:0] nor_191_nl;
  wire[0:0] nor_192_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] and_229_nl;
  wire[0:0] mux_581_nl;
  wire[0:0] nor_193_nl;
  wire[0:0] nor_194_nl;
  wire[0:0] nor_195_nl;
  wire[0:0] mux_580_nl;
  wire[0:0] or_643_nl;
  wire[0:0] or_642_nl;
  wire[0:0] or_659_nl;
  wire[0:0] mux_598_nl;
  wire[0:0] or_669_nl;
  wire[0:0] mux_623_nl;
  wire[0:0] or_73_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] or_694_nl;
  wire[0:0] mux_636_nl;
  wire[0:0] or_708_nl;
  wire[0:0] mux_758_nl;
  wire[0:0] mux_757_nl;
  wire[0:0] nor_158_nl;
  wire[0:0] mux_756_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] or_797_nl;
  wire[0:0] nor_159_nl;
  wire[0:0] and_208_nl;
  wire[0:0] mux_755_nl;
  wire[0:0] nor_160_nl;
  wire[0:0] mux_754_nl;
  wire[0:0] nor_161_nl;
  wire[0:0] and_209_nl;
  wire[0:0] mux_753_nl;
  wire[0:0] nor_162_nl;
  wire[0:0] nor_163_nl;
  wire[0:0] nor_164_nl;
  wire[0:0] or_801_nl;
  wire[0:0] and_292_nl;
  wire[0:0] nor_150_nl;
  wire[0:0] nor_151_nl;
  wire[0:0] mux_785_nl;
  wire[0:0] or_832_nl;
  wire[0:0] mux_784_nl;
  wire[0:0] or_831_nl;
  wire[0:0] or_27_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] nor_132_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] mux_790_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] or_843_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] mux_496_nl;
  wire[0:0] nor_217_nl;
  wire[0:0] mux_495_nl;
  wire[0:0] or_9_nl;
  wire[0:0] or_556_nl;
  wire[0:0] mux_502_nl;
  wire[0:0] mux_501_nl;
  wire[0:0] or_914_nl;
  wire[0:0] or_915_nl;
  wire[0:0] or_916_nl;
  wire[0:0] or_184_nl;
  wire[0:0] or_180_nl;
  wire[0:0] and_61_nl;
  wire[0:0] and_63_nl;
  wire[0:0] mux_167_nl;
  wire[0:0] nor_307_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] or_186_nl;
  wire[0:0] mux_164_nl;
  wire[0:0] nor_308_nl;
  wire[0:0] nor_309_nl;
  wire[0:0] and_65_nl;
  wire[0:0] mux_170_nl;
  wire[0:0] and_283_nl;
  wire[0:0] mux_169_nl;
  wire[0:0] nor_304_nl;
  wire[0:0] nor_305_nl;
  wire[0:0] nor_306_nl;
  wire[0:0] mux_168_nl;
  wire[0:0] or_190_nl;
  wire[0:0] or_189_nl;
  wire[0:0] and_70_nl;
  wire[0:0] mux_173_nl;
  wire[0:0] and_282_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] nor_301_nl;
  wire[0:0] nor_302_nl;
  wire[0:0] nor_303_nl;
  wire[0:0] and_77_nl;
  wire[0:0] mux_176_nl;
  wire[0:0] nor_299_nl;
  wire[0:0] mux_175_nl;
  wire[0:0] or_209_nl;
  wire[0:0] or_208_nl;
  wire[0:0] nor_300_nl;
  wire[0:0] mux_174_nl;
  wire[0:0] or_205_nl;
  wire[0:0] or_204_nl;
  wire[0:0] nor_292_nl;
  wire[0:0] nor_293_nl;
  wire[0:0] mux_183_nl;
  wire[0:0] nand_11_nl;
  wire[0:0] mux_182_nl;
  wire[0:0] nor_294_nl;
  wire[0:0] mux_181_nl;
  wire[0:0] or_224_nl;
  wire[0:0] or_223_nl;
  wire[0:0] mux_180_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] nor_296_nl;
  wire[0:0] or_217_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] nand_10_nl;
  wire[0:0] mux_178_nl;
  wire[0:0] nor_297_nl;
  wire[0:0] nor_298_nl;
  wire[0:0] mux_177_nl;
  wire[0:0] or_213_nl;
  wire[0:0] or_211_nl;
  wire[0:0] mux_207_nl;
  wire[0:0] nor_282_nl;
  wire[0:0] mux_206_nl;
  wire[0:0] mux_205_nl;
  wire[0:0] or_267_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] or_266_nl;
  wire[0:0] or_264_nl;
  wire[0:0] or_263_nl;
  wire[0:0] or_261_nl;
  wire[0:0] mux_203_nl;
  wire[0:0] mux_202_nl;
  wire[0:0] or_260_nl;
  wire[0:0] mux_201_nl;
  wire[0:0] or_259_nl;
  wire[0:0] or_258_nl;
  wire[0:0] or_257_nl;
  wire[0:0] or_256_nl;
  wire[0:0] nor_283_nl;
  wire[0:0] mux_200_nl;
  wire[0:0] or_253_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] and_280_nl;
  wire[0:0] mux_198_nl;
  wire[0:0] and_281_nl;
  wire[0:0] mux_197_nl;
  wire[0:0] nor_284_nl;
  wire[0:0] nor_285_nl;
  wire[0:0] mux_196_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] mux_194_nl;
  wire[0:0] mux_193_nl;
  wire[0:0] nor_286_nl;
  wire[0:0] nor_287_nl;
  wire[0:0] nor_288_nl;
  wire[0:0] or_246_nl;
  wire[0:0] nor_289_nl;
  wire[0:0] nor_290_nl;
  wire[0:0] nor_291_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] or_242_nl;
  wire[0:0] nor_274_nl;
  wire[0:0] nor_275_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] and_279_nl;
  wire[0:0] mux_213_nl;
  wire[0:0] nor_277_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] nor_278_nl;
  wire[0:0] nor_279_nl;
  wire[0:0] or_275_nl;
  wire[0:0] mux_211_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] nor_280_nl;
  wire[0:0] nor_281_nl;
  wire[0:0] mux_209_nl;
  wire[0:0] or_271_nl;
  wire[0:0] or_269_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] nor_267_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] or_324_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] or_322_nl;
  wire[0:0] or_320_nl;
  wire[0:0] or_318_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] nand_22_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] or_314_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] or_313_nl;
  wire[0:0] or_311_nl;
  wire[0:0] and_276_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] nor_270_nl;
  wire[0:0] nor_271_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_277_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] or_308_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] or_307_nl;
  wire[0:0] or_306_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] or_299_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] or_303_nl;
  wire[0:0] or_302_nl;
  wire[0:0] or_301_nl;
  wire[0:0] or_300_nl;
  wire[0:0] and_278_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] nor_272_nl;
  wire[0:0] nor_273_nl;
  wire[0:0] and_274_nl;
  wire[0:0] nor_261_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] nand_24_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] nor_262_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] or_338_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] nor_263_nl;
  wire[0:0] nor_264_nl;
  wire[0:0] or_332_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] nor_265_nl;
  wire[0:0] nor_266_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] or_328_nl;
  wire[0:0] or_326_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] nor_255_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] or_379_nl;
  wire[0:0] or_377_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] or_375_nl;
  wire[0:0] nor_54_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] or_373_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] or_372_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] or_371_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] or_367_nl;
  wire[0:0] and_271_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] nor_256_nl;
  wire[0:0] nor_257_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] and_272_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] or_364_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] or_363_nl;
  wire[0:0] or_362_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] or_356_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] or_360_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] or_358_nl;
  wire[0:0] nor_51_nl;
  wire[0:0] or_357_nl;
  wire[0:0] and_273_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] nor_258_nl;
  wire[0:0] nor_259_nl;
  wire[0:0] and_267_nl;
  wire[0:0] nor_248_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nand_32_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] and_269_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] nor_250_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] nor_251_nl;
  wire[0:0] nor_252_nl;
  wire[0:0] or_387_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] nand_30_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] nor_253_nl;
  wire[0:0] nor_254_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] nand_112_nl;
  wire[0:0] or_381_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] nor_240_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] or_431_nl;
  wire[0:0] or_429_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] or_427_nl;
  wire[0:0] and_261_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] or_425_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] or_424_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] nand_38_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] and_263_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] nor_243_nl;
  wire[0:0] nor_244_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] and_264_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] or_417_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] or_416_nl;
  wire[0:0] nand_91_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] or_409_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] nand_92_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] or_411_nl;
  wire[0:0] and_265_nl;
  wire[0:0] or_410_nl;
  wire[0:0] and_266_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] nor_245_nl;
  wire[0:0] nor_246_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] and_522_nl;
  wire[0:0] mux_827_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] or_999_nl;
  wire[0:0] or_1000_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] or_997_nl;
  wire[0:0] or_998_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] or_938_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] nand_140_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] or_945_nl;
  wire[0:0] or_993_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] or_942_nl;
  wire[0:0] or_940_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] or_951_nl;
  wire[0:0] or_950_nl;
  wire[0:0] or_959_nl;
  wire[0:0] or_957_nl;
  wire[0:0] nand_125_nl;
  wire[0:0] or_956_nl;
  wire[0:0] or_965_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] or_966_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] nand_126_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] or_963_nl;
  wire[0:0] or_961_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] or_970_nl;
  wire[0:0] or_968_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] or_973_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] or_972_nl;
  wire[0:0] or_976_nl;
  wire[0:0] or_975_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] or_1007_nl;
  wire[0:0] or_1005_nl;
  wire[0:0] nand_147_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] or_1053_nl;
  wire[1:0] operator_64_false_1_operator_64_false_1_or_1_nl;
  wire[1:0] operator_64_false_1_mux_5_nl;
  wire[0:0] operator_64_false_1_mux1h_9_nl;
  wire[0:0] operator_64_false_1_mux1h_10_nl;
  wire[0:0] operator_64_false_1_mux1h_11_nl;
  wire[0:0] operator_64_false_1_mux1h_12_nl;
  wire[0:0] operator_64_false_1_mux1h_13_nl;
  wire[0:0] operator_64_false_1_mux1h_14_nl;
  wire[0:0] operator_64_false_1_mux1h_15_nl;
  wire[0:0] operator_64_false_1_mux1h_16_nl;
  wire[6:0] operator_64_false_1_operator_64_false_1_mux_1_nl;
  wire[0:0] operator_64_false_1_or_6_nl;
  wire[12:0] acc_2_nl;
  wire[13:0] nl_acc_2_nl;
  wire[2:0] COMP_LOOP_mux1h_83_nl;
  wire[8:0] COMP_LOOP_mux1h_84_nl;
  wire[0:0] COMP_LOOP_or_34_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_or_3_nl;
  wire[1:0] COMP_LOOP_mux_41_nl;
  wire[11:0] COMP_LOOP_mux1h_85_nl;
  wire[0:0] and_532_nl;
  wire[0:0] COMP_LOOP_or_35_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_5_nl;
  wire[63:0] COMP_LOOP_mux1h_86_nl;
  wire[63:0] COMP_LOOP_or_36_nl;
  wire[63:0] COMP_LOOP_mux1h_87_nl;
  wire[0:0] COMP_LOOP_or_37_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_or_1_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_103_nl;
  wire[0:0] STAGE_LOOP_mux_55_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_104_nl;
  wire[0:0] STAGE_LOOP_mux_56_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_105_nl;
  wire[0:0] STAGE_LOOP_mux_57_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_106_nl;
  wire[0:0] STAGE_LOOP_mux_58_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_107_nl;
  wire[0:0] STAGE_LOOP_mux_59_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_108_nl;
  wire[0:0] STAGE_LOOP_mux_60_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_109_nl;
  wire[0:0] STAGE_LOOP_mux_61_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_110_nl;
  wire[0:0] STAGE_LOOP_mux_62_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_111_nl;
  wire[0:0] STAGE_LOOP_mux_63_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_112_nl;
  wire[0:0] STAGE_LOOP_mux_64_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_113_nl;
  wire[0:0] STAGE_LOOP_mux_65_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_114_nl;
  wire[0:0] STAGE_LOOP_mux_66_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_115_nl;
  wire[0:0] STAGE_LOOP_mux_67_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_116_nl;
  wire[0:0] STAGE_LOOP_mux_68_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_117_nl;
  wire[0:0] STAGE_LOOP_mux_69_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_118_nl;
  wire[0:0] STAGE_LOOP_mux_70_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_119_nl;
  wire[0:0] STAGE_LOOP_mux_71_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_120_nl;
  wire[0:0] STAGE_LOOP_mux_72_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_121_nl;
  wire[0:0] STAGE_LOOP_mux_73_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_122_nl;
  wire[0:0] STAGE_LOOP_mux_74_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_123_nl;
  wire[0:0] STAGE_LOOP_mux_75_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_124_nl;
  wire[0:0] STAGE_LOOP_mux_76_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_125_nl;
  wire[0:0] STAGE_LOOP_mux_77_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_126_nl;
  wire[0:0] STAGE_LOOP_mux_78_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_127_nl;
  wire[0:0] STAGE_LOOP_mux_79_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_128_nl;
  wire[0:0] STAGE_LOOP_mux_80_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_129_nl;
  wire[0:0] STAGE_LOOP_mux_81_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_130_nl;
  wire[0:0] STAGE_LOOP_mux_82_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_131_nl;
  wire[0:0] STAGE_LOOP_mux_83_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_132_nl;
  wire[0:0] STAGE_LOOP_mux_84_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_133_nl;
  wire[0:0] STAGE_LOOP_mux_85_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_134_nl;
  wire[0:0] STAGE_LOOP_mux_86_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_135_nl;
  wire[0:0] STAGE_LOOP_mux_87_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_136_nl;
  wire[0:0] STAGE_LOOP_mux_88_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_137_nl;
  wire[0:0] STAGE_LOOP_mux_89_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_138_nl;
  wire[0:0] STAGE_LOOP_mux_90_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_139_nl;
  wire[0:0] STAGE_LOOP_mux_91_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_140_nl;
  wire[0:0] STAGE_LOOP_mux_92_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_141_nl;
  wire[0:0] STAGE_LOOP_mux_93_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_142_nl;
  wire[0:0] STAGE_LOOP_mux_94_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_143_nl;
  wire[0:0] STAGE_LOOP_mux_95_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_144_nl;
  wire[0:0] STAGE_LOOP_mux_96_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_145_nl;
  wire[0:0] STAGE_LOOP_mux_97_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_146_nl;
  wire[0:0] STAGE_LOOP_mux_98_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_147_nl;
  wire[0:0] STAGE_LOOP_mux_99_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_148_nl;
  wire[0:0] STAGE_LOOP_mux_100_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_149_nl;
  wire[0:0] STAGE_LOOP_mux_101_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_150_nl;
  wire[0:0] STAGE_LOOP_mux_102_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_151_nl;
  wire[0:0] STAGE_LOOP_mux_103_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_152_nl;
  wire[0:0] STAGE_LOOP_mux_104_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_153_nl;
  wire[0:0] STAGE_LOOP_mux_105_nl;
  wire[1:0] STAGE_LOOP_and_4_nl;
  wire[1:0] STAGE_LOOP_mux1h_6_nl;
  wire[0:0] STAGE_LOOP_nor_106_nl;
  wire[8:0] STAGE_LOOP_mux1h_7_nl;
  wire[7:0] COMP_LOOP_acc_61_nl;
  wire[8:0] nl_COMP_LOOP_acc_61_nl;
  wire[8:0] COMP_LOOP_acc_62_nl;
  wire[9:0] nl_COMP_LOOP_acc_62_nl;
  wire[0:0] STAGE_LOOP_or_10_nl;
  wire[0:0] STAGE_LOOP_or_11_nl;
  wire[0:0] STAGE_LOOP_mux1h_8_nl;
  wire[0:0] STAGE_LOOP_or_12_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_154_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_155_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_156_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_157_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_158_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_159_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_160_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_161_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_162_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_163_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_164_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_165_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_166_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_167_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_168_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_169_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_170_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_171_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_172_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_173_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_174_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_175_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_176_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_177_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_178_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_179_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_180_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_181_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_182_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_183_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_184_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_185_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_186_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_187_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_188_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_189_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_190_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_191_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_192_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_193_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_194_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_195_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_196_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_197_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_198_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_199_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_200_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_201_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_202_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_203_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_204_nl;
  wire[0:0] STAGE_LOOP_STAGE_LOOP_and_205_nl;
  wire[1:0] STAGE_LOOP_and_5_nl;
  wire[1:0] STAGE_LOOP_mux1h_9_nl;
  wire[0:0] STAGE_LOOP_nor_107_nl;
  wire[9:0] STAGE_LOOP_mux1h_10_nl;
  wire[0:0] STAGE_LOOP_or_13_nl;
  wire[0:0] STAGE_LOOP_or_14_nl;
  wire[63:0] modExp_while_if_mux1h_1_nl;
  wire[0:0] and_533_nl;
  wire[0:0] modExp_while_if_modExp_while_if_nand_1_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] or_1078_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] or_1080_nl;
  wire[0:0] and_534_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] and_535_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] and_536_nl;
  wire[63:0] modExp_while_if_modExp_while_if_mux1h_1_nl;
  wire[0:0] modExp_while_if_modExp_while_if_nor_1_nl;
  wire[0:0] modExp_while_if_and_6_nl;
  wire[0:0] modExp_while_if_and_7_nl;
  wire[0:0] modExp_while_if_and_8_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_5_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_5_tr0 = ~ (z_out_5[64]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0 = ~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_40_tr0 = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_80_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_80_tr0 = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_120_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_120_tr0 = ~
      VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_6[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0 = ~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_40_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_40_tr0 = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_80_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_80_tr0 = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_120_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_120_tr0 = ~
      VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0
      = ~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0 = z_out_6[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_6_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_6_tr0 = ~ (z_out_5[2]);
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_3_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_5_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_5_tr0[0:0]),
      .modExp_while_C_24_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_1_COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_1_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_C_24_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_1_COMP_LOOP_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_40_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_2_modExp_1_while_C_24_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_C_80_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_80_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_3_modExp_1_while_C_24_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_C_120_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_C_120_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_1_COMP_LOOP_4_modExp_1_while_C_24_tr0[0:0]),
      .VEC_LOOP_1_COMP_LOOP_C_160_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_1_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_1_modExp_1_while_C_24_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_2_COMP_LOOP_C_40_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_40_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_2_modExp_1_while_C_24_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_80_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_80_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_3_modExp_1_while_C_24_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_120_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_C_120_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_2_COMP_LOOP_4_modExp_1_while_C_24_tr0[0:0]),
      .VEC_LOOP_2_COMP_LOOP_C_160_tr0(exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva),
      .VEC_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_1_tr0[0:0]),
      .STAGE_LOOP_C_6_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_6_tr0[0:0])
    );
  assign mux_187_nl = MUX_s_1_2_2(or_304_cse, or_369_cse, fsm_output[1]);
  assign or_237_nl = (~ (fsm_output[1])) | (~ (fsm_output[8])) | (fsm_output[9])
      | (fsm_output[7]);
  assign mux_188_nl = MUX_s_1_2_2(mux_187_nl, or_237_nl, fsm_output[2]);
  assign or_236_nl = (fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[9])
      | (~ (fsm_output[7]));
  assign mux_189_cse = MUX_s_1_2_2(mux_188_nl, or_236_nl, fsm_output[3]);
  assign or_231_nl = (fsm_output[9:7]!=3'b010);
  assign mux_184_nl = MUX_s_1_2_2(or_369_cse, or_231_nl, fsm_output[1]);
  assign mux_185_nl = MUX_s_1_2_2(mux_184_nl, nand_95_cse, fsm_output[2]);
  assign or_228_nl = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[9]))
      | (fsm_output[7]);
  assign mux_186_cse = MUX_s_1_2_2(mux_185_nl, or_228_nl, fsm_output[3]);
  assign nand_12_nl = ~((fsm_output[6]) & (~ mux_189_cse));
  assign or_234_nl = (fsm_output[6]) | mux_186_cse;
  assign mux_190_cse = MUX_s_1_2_2(nand_12_nl, or_234_nl, fsm_output[0]);
  assign nand_95_cse = ~((fsm_output[1]) & (fsm_output[7]) & (fsm_output[8]) & (~
      (fsm_output[9])));
  assign or_304_cse = (fsm_output[9:7]!=3'b000);
  assign nor_269_cse = ~((fsm_output[9:7]!=3'b001));
  assign or_315_cse = (fsm_output[2]) | (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])) |
      (fsm_output[1]) | (~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign nor_268_cse = ~((VEC_LOOP_j_1_12_0_sva_11_0[1]) | (fsm_output[9:7]!=3'b000));
  assign and_275_nl = (fsm_output[6]) & (~ mux_189_cse);
  assign nor_260_nl = ~((fsm_output[6]) | mux_186_cse);
  assign mux_258_cse = MUX_s_1_2_2(and_275_nl, nor_260_nl, fsm_output[0]);
  assign and_270_cse = VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm & (COMP_LOOP_acc_11_psp_1_sva[0]);
  assign or_369_cse = (fsm_output[9:7]!=3'b001);
  assign or_370_cse = (~ (VEC_LOOP_j_1_12_0_sva_11_0[1])) | (fsm_output[9:7]!=3'b000);
  assign nor_241_cse = ~((~ (VEC_LOOP_j_1_12_0_sva_11_0[1])) | (fsm_output[9:7]!=3'b000));
  assign nor_70_cse = ~((fsm_output[8]) | (~ (fsm_output[2])));
  assign and_256_cse = (fsm_output[3:2]==2'b11);
  assign nor_236_cse = ~((fsm_output[3:2]!=2'b00));
  assign or_154_cse = (fsm_output[7:6]!=2'b00);
  assign or_709_nl = (~ (fsm_output[2])) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_670_nl = MUX_s_1_2_2(or_tmp_670, or_709_nl, fsm_output[7]);
  assign mux_671_nl = MUX_s_1_2_2(mux_670_nl, mux_tmp_668, fsm_output[1]);
  assign nor_178_nl = ~((fsm_output[8]) | mux_671_nl);
  assign or_705_nl = (fsm_output[2]) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign or_703_nl = (fsm_output[2]) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_667_nl = MUX_s_1_2_2(or_705_nl, or_703_nl, fsm_output[7]);
  assign mux_669_nl = MUX_s_1_2_2(mux_tmp_668, mux_667_nl, fsm_output[1]);
  assign and_225_nl = (fsm_output[8]) & (~ mux_669_nl);
  assign mux_672_nl = MUX_s_1_2_2(nor_178_nl, and_225_nl, fsm_output[3]);
  assign or_702_nl = (~ (fsm_output[2])) | (fsm_output[4]);
  assign mux_658_nl = MUX_s_1_2_2((~ nor_tmp_103), or_702_nl, fsm_output[1]);
  assign mux_659_nl = MUX_s_1_2_2(or_tmp_654, mux_658_nl, fsm_output[3]);
  assign mux_656_nl = MUX_s_1_2_2((~ or_tmp_61), (fsm_output[4]), fsm_output[1]);
  assign or_701_nl = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[1])
      | (fsm_output[2]) | (fsm_output[4]);
  assign mux_657_nl = MUX_s_1_2_2(mux_656_nl, or_701_nl, fsm_output[3]);
  assign mux_660_nl = MUX_s_1_2_2(mux_659_nl, mux_657_nl, fsm_output[8]);
  assign mux_661_nl = MUX_s_1_2_2(mux_660_nl, mux_tmp_624, fsm_output[7]);
  assign or_699_nl = (fsm_output[3]) | (~(VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      | (fsm_output[2:1]!=2'b11))) | (fsm_output[4]);
  assign mux_648_nl = MUX_s_1_2_2((fsm_output[4]), or_tmp_656, fsm_output[3]);
  assign mux_649_nl = MUX_s_1_2_2(or_699_nl, mux_648_nl, fsm_output[8]);
  assign mux_650_nl = MUX_s_1_2_2(mux_tmp_637, mux_649_nl, fsm_output[7]);
  assign mux_664_nl = MUX_s_1_2_2(mux_661_nl, mux_650_nl, fsm_output[6]);
  assign or_695_nl = (fsm_output[4:1]!=4'b0000);
  assign mux_638_nl = MUX_s_1_2_2(or_695_nl, or_756_cse, fsm_output[8]);
  assign mux_639_nl = MUX_s_1_2_2(mux_638_nl, mux_tmp_637, fsm_output[7]);
  assign mux_625_nl = MUX_s_1_2_2((~ nor_tmp_103), or_tmp_61, fsm_output[1]);
  assign mux_626_nl = MUX_s_1_2_2(or_tmp_51, mux_625_nl, fsm_output[3]);
  assign mux_627_nl = MUX_s_1_2_2(mux_626_nl, or_756_cse, fsm_output[8]);
  assign mux_628_nl = MUX_s_1_2_2(mux_627_nl, mux_tmp_624, fsm_output[7]);
  assign mux_647_nl = MUX_s_1_2_2(mux_639_nl, mux_628_nl, fsm_output[6]);
  assign mux_950_nl = MUX_s_1_2_2(mux_664_nl, mux_647_nl, fsm_output[0]);
  assign or_994_nl = and_dcpl_104 | (mux_672_nl & and_dcpl_109 & (fsm_output[5])
      & (~((not_tmp_260 & (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)) |
      (mux_950_nl & (~ (fsm_output[9])))))) | (~ mux_423_itm);
  assign modExp_while_if_and_1_nl = modExp_while_and_3 & not_tmp_260;
  assign modExp_while_if_and_2_nl = modExp_while_and_5 & not_tmp_260;
  assign mux1h_nl = MUX1HOT_v_64_5_2(z_out_7, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      modulo_result_rem_cmp_z, z_out_6, (z_out_5[63:0]), {or_994_nl , and_dcpl_138
      , modExp_while_if_and_1_nl , modExp_while_if_and_2_nl , and_dcpl_108});
  assign and_126_nl = and_dcpl_33 & and_dcpl_102;
  assign or_533_nl = (fsm_output[1]) | (~ (fsm_output[7]));
  assign mux_457_nl = MUX_s_1_2_2(or_533_nl, or_tmp_484, fsm_output[8]);
  assign mux_458_nl = MUX_s_1_2_2(mux_457_nl, (~ and_dcpl_86), fsm_output[2]);
  assign mux_459_nl = MUX_s_1_2_2(or_826_cse, mux_458_nl, fsm_output[3]);
  assign nor_222_nl = ~((fsm_output[6]) | mux_459_nl);
  assign nor_223_nl = ~((fsm_output[3]) | mux_tmp_455);
  assign nor_224_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[1]))
      | (fsm_output[7]));
  assign mux_453_nl = MUX_s_1_2_2(and_dcpl_66, and_tmp_6, fsm_output[2]);
  assign mux_454_nl = MUX_s_1_2_2(nor_224_nl, mux_453_nl, fsm_output[3]);
  assign mux_456_nl = MUX_s_1_2_2(nor_223_nl, mux_454_nl, fsm_output[6]);
  assign mux_460_nl = MUX_s_1_2_2(nor_222_nl, mux_456_nl, fsm_output[0]);
  assign nor_225_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | and_dcpl_65);
  assign or_527_nl = (fsm_output[2]) | (~ and_tmp_8);
  assign mux_450_nl = MUX_s_1_2_2(nor_225_nl, or_527_nl, fsm_output[3]);
  assign mux_451_nl = MUX_s_1_2_2(mux_tmp_448, mux_450_nl, fsm_output[6]);
  assign mux_449_nl = MUX_s_1_2_2(mux_tmp_448, mux_tmp_440, fsm_output[6]);
  assign mux_452_nl = MUX_s_1_2_2(mux_451_nl, mux_449_nl, fsm_output[0]);
  assign mux_461_nl = MUX_s_1_2_2(mux_460_nl, mux_452_nl, fsm_output[4]);
  assign mux_443_nl = MUX_s_1_2_2(or_tmp_470, or_826_cse, fsm_output[2]);
  assign or_524_nl = (fsm_output[2]) | (fsm_output[8]) | (fsm_output[7]);
  assign mux_444_nl = MUX_s_1_2_2(mux_443_nl, or_524_nl, fsm_output[3]);
  assign or_526_nl = (fsm_output[6]) | mux_444_nl;
  assign or_523_nl = (fsm_output[6]) | or_tmp_476;
  assign mux_445_nl = MUX_s_1_2_2(or_526_nl, or_523_nl, fsm_output[0]);
  assign mux_446_nl = MUX_s_1_2_2(or_814_cse, mux_445_nl, fsm_output[4]);
  assign mux_462_nl = MUX_s_1_2_2(mux_461_nl, mux_446_nl, fsm_output[9]);
  assign or_519_nl = (fsm_output[8]) | and_dcpl_65;
  assign mux_441_nl = MUX_s_1_2_2(or_519_nl, and_tmp_8, fsm_output[2]);
  assign or_520_nl = (fsm_output[3]) | (~ mux_441_nl);
  assign mux_442_nl = MUX_s_1_2_2(or_520_nl, mux_tmp_440, or_913_cse);
  assign or_522_nl = (fsm_output[9]) | (~((fsm_output[4]) | mux_442_nl));
  assign mux_463_nl = MUX_s_1_2_2(mux_462_nl, or_522_nl, fsm_output[5]);
  assign operator_64_false_mux1h_2_rgt = MUX1HOT_v_65_3_2(z_out_5, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
      ({1'b0 , mux1h_nl}), {and_126_nl , and_dcpl_123 , (~ mux_463_nl)});
  assign and_524_cse = (fsm_output[1:0]==2'b11);
  assign or_1038_cse = (fsm_output[5]) | (~ (fsm_output[9]));
  assign or_1035_nl = (fsm_output[5]) | (fsm_output[9]);
  assign mux_894_cse = MUX_s_1_2_2(or_1035_nl, or_55_cse, fsm_output[4]);
  assign or_1047_cse = (~ (fsm_output[4])) | (fsm_output[5]) | (fsm_output[9]);
  assign and_141_m1c = and_dcpl_48 & nor_236_cse & and_dcpl_130;
  assign modExp_result_and_rgt = (~ modExp_while_and_5) & and_141_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_5 & and_141_m1c;
  assign or_590_cse = (fsm_output[1:0]!=2'b00);
  assign or_913_cse = (~ (fsm_output[0])) | (fsm_output[6]);
  assign or_596_cse = (~ (fsm_output[6])) | (fsm_output[0]);
  assign nand_119_cse = ~((fsm_output[3:2]==2'b11));
  assign or_614_cse = (~ (fsm_output[2])) | (fsm_output[3]) | (fsm_output[8]);
  assign mux_561_cse = MUX_s_1_2_2(or_tmp_573, or_614_cse, fsm_output[7]);
  assign or_611_cse = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign mux_560_cse = MUX_s_1_2_2(or_611_cse, or_tmp_573, fsm_output[7]);
  assign and_300_cse = (fsm_output[2:1]==2'b11);
  assign nor_330_cse = ~((~ (fsm_output[8])) | (fsm_output[3]) | (fsm_output[0])
      | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]));
  assign and_221_nl = (fsm_output[8]) & (fsm_output[3]);
  assign nor_174_nl = ~((fsm_output[8]) | (fsm_output[3]));
  assign mux_680_cse = MUX_s_1_2_2(and_221_nl, nor_174_nl, fsm_output[1]);
  assign COMP_LOOP_or_1_cse = (and_dcpl_33 & and_dcpl_41) | (and_dcpl_47 & (fsm_output[8])
      & and_dcpl_76 & and_dcpl_41);
  assign or_94_cse = (fsm_output[2:1]!=2'b00);
  assign or_756_cse = (fsm_output[4:3]!=2'b00);
  assign and_213_cse = (fsm_output[5:4]==2'b11);
  assign or_787_nl = (~ (fsm_output[0])) | (fsm_output[6]) | (fsm_output[9]) | (~
      (fsm_output[8])) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[5]);
  assign mux_749_cse = MUX_s_1_2_2(or_tmp_451, or_787_nl, fsm_output[7]);
  assign or_786_nl = (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[5]);
  assign or_785_nl = (fsm_output[9:8]!=2'b00) | not_tmp_173;
  assign mux_746_nl = MUX_s_1_2_2(or_786_nl, or_785_nl, fsm_output[6]);
  assign mux_747_nl = MUX_s_1_2_2(or_tmp_449, mux_746_nl, fsm_output[0]);
  assign mux_748_cse = MUX_s_1_2_2(mux_747_nl, or_tmp_451, fsm_output[7]);
  assign or_780_nl = (~ (fsm_output[6])) | (fsm_output[9]) | (fsm_output[8]) | not_tmp_173;
  assign mux_745_cse = MUX_s_1_2_2(or_tmp_449, or_780_nl, fsm_output[0]);
  assign and_205_cse = (fsm_output[7:6]==2'b11);
  assign or_814_cse = (fsm_output[8:6]!=3'b000);
  assign or_826_cse = (fsm_output[8:7]!=2'b00);
  assign COMP_LOOP_or_3_cse = (and_dcpl_49 & and_dcpl_45) | (and_dcpl_38 & and_dcpl_60)
      | (and_dcpl_66 & and_256_cse & and_dcpl_45) | (and_dcpl_73 & and_256_cse &
      and_dcpl_60) | (and_dcpl_31 & (fsm_output[8]) & nor_236_cse & and_dcpl_82)
      | (and_dcpl_87 & and_dcpl_29) | (and_dcpl_87 & and_dcpl_82) | (and_dcpl_32
      & and_dcpl_76 & and_dcpl_28 & (fsm_output[9]) & (~ (fsm_output[5])));
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      (tmp_10_lpi_4_dfm[63:1]), and_dcpl_134);
  assign modExp_base_1_sva_mx1 = MUX_v_64_2_2(modulo_result_rem_cmp_z, z_out_6, modulo_result_rem_cmp_z[63]);
  assign modExp_while_and_3 = (~ (modulo_result_rem_cmp_z[63])) & VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  assign modExp_while_and_5 = (modulo_result_rem_cmp_z[63]) & VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  assign nor_332_cse = ~((fsm_output[4:3]!=2'b00));
  assign or_tmp_29 = nor_332_cse | (fsm_output[9]) | (~ (fsm_output[5]));
  assign and_303_cse = (fsm_output[4:3]==2'b11);
  assign or_tmp_31 = and_303_cse | (fsm_output[9]) | (~ (fsm_output[5]));
  assign or_55_cse = (fsm_output[9]) | (~ (fsm_output[5]));
  assign or_54_cse = (~ (fsm_output[4])) | (fsm_output[9]) | (~ (fsm_output[5]));
  assign or_tmp_51 = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4]);
  assign or_tmp_61 = (fsm_output[2]) | (~ (fsm_output[4]));
  assign or_tmp_71 = (~((fsm_output[8:7]!=2'b01))) | (fsm_output[9]);
  assign or_tmp_72 = (fsm_output[9:8]!=2'b01);
  assign or_91_nl = (fsm_output[9:8]!=2'b00);
  assign mux_tmp_72 = MUX_s_1_2_2(or_91_nl, or_tmp_72, fsm_output[7]);
  assign or_tmp_77 = (fsm_output[9:7]!=3'b011);
  assign or_tmp_79 = (fsm_output[9:8]!=2'b10);
  assign mux_tmp_84 = MUX_s_1_2_2(or_tmp_79, or_tmp_72, fsm_output[7]);
  assign mux_tmp_86 = MUX_s_1_2_2(or_tmp_79, (fsm_output[9]), fsm_output[7]);
  assign or_103_nl = (fsm_output[8]) | (~ (fsm_output[1])) | (fsm_output[2]);
  assign or_102_nl = (~ (fsm_output[8])) | (fsm_output[1]) | (fsm_output[2]);
  assign mux_tmp_92 = MUX_s_1_2_2(or_103_nl, or_102_nl, fsm_output[3]);
  assign and_dcpl_13 = ~((fsm_output[9]) | (fsm_output[5]));
  assign nor_tmp_34 = (fsm_output[5]) & (fsm_output[9]);
  assign nor_312_cse = ~((fsm_output[8:6]!=3'b000));
  assign or_901_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[8]);
  assign mux_157_nl = MUX_s_1_2_2(or_901_nl, nor_312_cse, fsm_output[9]);
  assign nand_100_nl = ~((fsm_output[9]) & (((fsm_output[2]) & (fsm_output[3]) &
      (fsm_output[5])) | (fsm_output[8:6]!=3'b000)));
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, nand_100_nl, or_590_cse);
  assign nand_101_nl = ~((fsm_output[9]) & ((fsm_output[8:5]!=4'b0000)));
  assign not_tmp_77 = MUX_s_1_2_2(mux_158_nl, nand_101_nl, fsm_output[4]);
  assign and_dcpl_28 = ~((fsm_output[6]) | (fsm_output[0]) | (fsm_output[4]));
  assign and_dcpl_29 = and_dcpl_28 & and_dcpl_13;
  assign and_dcpl_31 = ~((fsm_output[7]) | (fsm_output[1]));
  assign and_dcpl_32 = and_dcpl_31 & (~ (fsm_output[8]));
  assign and_dcpl_33 = and_dcpl_32 & nor_236_cse;
  assign and_dcpl_38 = and_dcpl_32 & and_256_cse;
  assign and_dcpl_40 = (~ (fsm_output[9])) & (fsm_output[5]);
  assign and_dcpl_41 = and_dcpl_28 & and_dcpl_40;
  assign and_dcpl_43 = (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_dcpl_44 = and_dcpl_43 & (fsm_output[4]);
  assign and_dcpl_45 = and_dcpl_44 & and_dcpl_40;
  assign and_dcpl_46 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_47 = (~ (fsm_output[7])) & (fsm_output[1]);
  assign and_dcpl_48 = and_dcpl_47 & (~ (fsm_output[8]));
  assign and_dcpl_49 = and_dcpl_48 & and_dcpl_46;
  assign and_dcpl_51 = (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_dcpl_52 = and_dcpl_51 & (fsm_output[4]);
  assign nor_tmp_40 = (fsm_output[8]) & (fsm_output[1]);
  assign nor_310_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[1]));
  assign nor_311_nl = ~((fsm_output[2]) | (~ nor_tmp_40));
  assign not_tmp_91 = MUX_s_1_2_2(nor_310_nl, nor_311_nl, fsm_output[3]);
  assign mux_tmp_162 = MUX_s_1_2_2(or_596_cse, or_913_cse, fsm_output[7]);
  assign or_tmp_148 = (fsm_output[9]) | (~ (fsm_output[7])) | (fsm_output[0]) | (~
      (fsm_output[6]));
  assign and_dcpl_60 = and_dcpl_52 & and_dcpl_40;
  assign and_dcpl_65 = (fsm_output[7]) & (~ (fsm_output[1]));
  assign and_dcpl_66 = and_dcpl_65 & (~ (fsm_output[8]));
  assign and_dcpl_72 = (fsm_output[7]) & (fsm_output[1]);
  assign and_dcpl_73 = and_dcpl_72 & (~ (fsm_output[8]));
  assign and_dcpl_76 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_82 = (fsm_output[6]) & (fsm_output[0]) & (~ (fsm_output[4])) &
      and_dcpl_13;
  assign and_dcpl_86 = and_dcpl_72 & (fsm_output[8]);
  assign and_dcpl_87 = and_dcpl_86 & nor_236_cse;
  assign not_tmp_108 = ~((fsm_output[2]) & (fsm_output[9]));
  assign or_tmp_264 = (fsm_output[2]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b01) |
      (fsm_output[1]) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[9:7]!=3'b011);
  assign or_tmp_278 = (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b01) | (~ (fsm_output[1]))
      | (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign or_tmp_321 = (fsm_output[2]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b10) |
      (fsm_output[1]) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[9:7]!=3'b011);
  assign or_tmp_334 = (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b10) | (~ (fsm_output[1]))
      | (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign or_tmp_374 = (fsm_output[2]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b11) |
      (fsm_output[1]) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[9:7]!=3'b011);
  assign or_tmp_387 = (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b11) | (~ (fsm_output[1]))
      | (fsm_output[7]) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign and_dcpl_101 = and_dcpl_43 & (~ (fsm_output[4]));
  assign and_dcpl_102 = and_dcpl_101 & and_dcpl_13;
  assign and_dcpl_103 = and_dcpl_48 & and_dcpl_76;
  assign and_dcpl_104 = and_dcpl_103 & and_dcpl_102;
  assign mux_tmp_317 = MUX_s_1_2_2((~ or_756_cse), and_303_cse, fsm_output[2]);
  assign mux_tmp_318 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[3]);
  assign or_tmp_404 = (fsm_output[4:3]!=2'b10);
  assign mux_tmp_319 = MUX_s_1_2_2((~ or_tmp_404), mux_tmp_318, fsm_output[2]);
  assign nor_tmp_63 = (fsm_output[4:2]==3'b111);
  assign or_899_cse = (fsm_output[3:2]!=2'b00);
  assign nor_tmp_64 = or_899_cse & (fsm_output[4]);
  assign or_tmp_415 = ~(nand_119_cse & (fsm_output[4]));
  assign mux_324_nl = MUX_s_1_2_2(nor_tmp_64, or_tmp_415, fsm_output[5]);
  assign mux_323_nl = MUX_s_1_2_2((~ mux_tmp_317), nor_tmp_64, fsm_output[5]);
  assign mux_tmp_325 = MUX_s_1_2_2((~ mux_324_nl), mux_323_nl, fsm_output[8]);
  assign mux_327_nl = MUX_s_1_2_2(and_303_cse, or_tmp_415, fsm_output[5]);
  assign mux_326_nl = MUX_s_1_2_2((~ nor_tmp_63), and_303_cse, fsm_output[5]);
  assign mux_328_nl = MUX_s_1_2_2((~ mux_327_nl), mux_326_nl, fsm_output[8]);
  assign mux_tmp_329 = MUX_s_1_2_2(mux_328_nl, mux_tmp_325, fsm_output[1]);
  assign mux_tmp_335 = MUX_s_1_2_2((fsm_output[3]), (fsm_output[4]), fsm_output[2]);
  assign mux_336_nl = MUX_s_1_2_2(mux_tmp_335, or_tmp_415, fsm_output[5]);
  assign mux_334_nl = MUX_s_1_2_2((~ mux_tmp_317), and_303_cse, fsm_output[5]);
  assign mux_tmp_337 = MUX_s_1_2_2((~ mux_336_nl), mux_334_nl, fsm_output[8]);
  assign mux_332_nl = MUX_s_1_2_2((~ nor_tmp_64), (fsm_output[4]), fsm_output[5]);
  assign mux_330_nl = MUX_s_1_2_2(mux_tmp_318, (fsm_output[3]), fsm_output[2]);
  assign mux_331_nl = MUX_s_1_2_2((~ mux_330_nl), nor_tmp_64, fsm_output[5]);
  assign mux_333_nl = MUX_s_1_2_2(mux_332_nl, mux_331_nl, fsm_output[8]);
  assign mux_tmp_338 = MUX_s_1_2_2(mux_tmp_337, mux_333_nl, fsm_output[1]);
  assign mux_tmp_340 = MUX_s_1_2_2((~ and_303_cse), nor_tmp_64, fsm_output[5]);
  assign or_tmp_416 = (fsm_output[4:3]!=2'b01);
  assign mux_tmp_345 = MUX_s_1_2_2(mux_tmp_318, or_tmp_416, fsm_output[2]);
  assign mux_tmp_350 = MUX_s_1_2_2(and_303_cse, mux_tmp_345, fsm_output[5]);
  assign mux_tmp_373 = MUX_s_1_2_2((~ (fsm_output[5])), (fsm_output[5]), fsm_output[4]);
  assign or_tmp_421 = (~((~ (fsm_output[8])) | (fsm_output[2]))) | (fsm_output[9])
      | mux_tmp_373;
  assign or_tmp_423 = (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[5]));
  assign or_tmp_426 = (~ (fsm_output[2])) | (fsm_output[9]) | mux_tmp_373;
  assign mux_374_nl = MUX_s_1_2_2(or_55_cse, or_tmp_423, fsm_output[2]);
  assign mux_tmp_375 = MUX_s_1_2_2(or_tmp_426, mux_374_nl, fsm_output[8]);
  assign or_462_cse = (fsm_output[2]) | (fsm_output[9]) | (fsm_output[4]) | (~ (fsm_output[5]));
  assign mux_376_nl = MUX_s_1_2_2(or_462_cse, or_55_cse, fsm_output[8]);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, mux_tmp_375, fsm_output[1]);
  assign mux_tmp_378 = MUX_s_1_2_2(mux_377_nl, or_tmp_421, fsm_output[3]);
  assign or_467_nl = (fsm_output[2]) | (fsm_output[9]) | (~ (fsm_output[5]));
  assign mux_tmp_379 = MUX_s_1_2_2(or_tmp_426, or_467_nl, fsm_output[8]);
  assign mux_tmp_380 = MUX_s_1_2_2(or_tmp_426, or_55_cse, fsm_output[8]);
  assign mux_381_nl = MUX_s_1_2_2(mux_tmp_380, mux_tmp_379, fsm_output[1]);
  assign or_465_nl = (~((fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[2])))
      | (fsm_output[9]) | mux_tmp_373;
  assign mux_tmp_382 = MUX_s_1_2_2(mux_381_nl, or_465_nl, fsm_output[3]);
  assign or_tmp_436 = (fsm_output[9]) | (~ (fsm_output[4]));
  assign or_tmp_437 = (fsm_output[5:4]!=2'b01);
  assign or_tmp_438 = (fsm_output[5:4]!=2'b10);
  assign mux_tmp_393 = MUX_s_1_2_2((~ (fsm_output[4])), or_tmp_438, fsm_output[9]);
  assign not_tmp_170 = ~((fsm_output[5:4]==2'b11));
  assign mux_396_nl = MUX_s_1_2_2(not_tmp_170, or_tmp_438, fsm_output[9]);
  assign mux_397_nl = MUX_s_1_2_2(mux_396_nl, mux_tmp_393, fsm_output[2]);
  assign or_475_nl = (fsm_output[9]) | not_tmp_170;
  assign mux_395_nl = MUX_s_1_2_2(or_tmp_423, or_475_nl, fsm_output[2]);
  assign mux_tmp_398 = MUX_s_1_2_2(mux_397_nl, mux_395_nl, fsm_output[8]);
  assign and_dcpl_105 = ~((fsm_output[7]) | (fsm_output[2]));
  assign nor_232_nl = ~((fsm_output[8]) | (~ (fsm_output[1])));
  assign nor_233_nl = ~((~ (fsm_output[8])) | (fsm_output[1]));
  assign mux_416_nl = MUX_s_1_2_2(nor_232_nl, nor_233_nl, fsm_output[3]);
  assign and_dcpl_107 = mux_416_nl & and_dcpl_105 & and_dcpl_41;
  assign not_tmp_173 = ~((fsm_output[5:3]==3'b111));
  assign or_tmp_449 = (fsm_output[6]) | (fsm_output[9]) | (fsm_output[8]) | not_tmp_173;
  assign or_tmp_451 = (fsm_output[0]) | (~ (fsm_output[6])) | (fsm_output[9]) | (~
      (fsm_output[8])) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[5]);
  assign nand_40_nl = ~((fsm_output[2]) & (~ mux_748_cse));
  assign nand_39_nl = ~((fsm_output[7]) & (~ mux_745_cse));
  assign mux_419_nl = MUX_s_1_2_2(mux_749_cse, nand_39_nl, fsm_output[2]);
  assign mux_423_itm = MUX_s_1_2_2(nand_40_nl, mux_419_nl, fsm_output[1]);
  assign or_tmp_455 = (~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[9]) | (~
      (fsm_output[0])) | (fsm_output[6]);
  assign nand_87_nl = ~((fsm_output[4]) & (fsm_output[9]) & (fsm_output[0]) & (~
      (fsm_output[6])));
  assign or_498_nl = (fsm_output[4]) | (fsm_output[9]) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign mux_427_nl = MUX_s_1_2_2(nand_87_nl, or_498_nl, fsm_output[3]);
  assign mux_428_nl = MUX_s_1_2_2(mux_427_nl, or_tmp_455, fsm_output[7]);
  assign or_496_nl = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[4])
      | (fsm_output[9]) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign mux_429_nl = MUX_s_1_2_2(mux_428_nl, or_496_nl, fsm_output[1]);
  assign or_909_nl = (fsm_output[2]) | mux_429_nl;
  assign or_910_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[4]))
      | (fsm_output[9]) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign or_911_nl = (fsm_output[7]) | (~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[9])
      | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_425_nl = MUX_s_1_2_2(or_910_nl, or_911_nl, fsm_output[1]);
  assign or_491_nl = (~ (fsm_output[3])) | (fsm_output[4]) | (fsm_output[9]) | (fsm_output[0])
      | (~ (fsm_output[6]));
  assign mux_424_nl = MUX_s_1_2_2(or_491_nl, or_tmp_455, fsm_output[7]);
  assign nand_113_nl = ~((fsm_output[1]) & (~ mux_424_nl));
  assign mux_426_nl = MUX_s_1_2_2(mux_425_nl, nand_113_nl, fsm_output[2]);
  assign mux_430_nl = MUX_s_1_2_2(or_909_nl, mux_426_nl, fsm_output[8]);
  assign and_dcpl_108 = ~(mux_430_nl | (fsm_output[5]));
  assign and_dcpl_109 = ~((fsm_output[4]) | (fsm_output[9]));
  assign and_dcpl_110 = and_dcpl_109 & (fsm_output[5]);
  assign mux_tmp_431 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[1]);
  assign and_tmp_6 = (fsm_output[8]) & mux_tmp_431;
  assign or_tmp_470 = (fsm_output[8]) | (~ (fsm_output[1])) | (fsm_output[7]);
  assign or_503_nl = (fsm_output[8]) | (fsm_output[1]) | (~ (fsm_output[7]));
  assign mux_432_nl = MUX_s_1_2_2(or_tmp_470, or_503_nl, fsm_output[2]);
  assign or_501_nl = (fsm_output[2]) | (~ and_tmp_6);
  assign mux_433_itm = MUX_s_1_2_2(mux_432_nl, or_501_nl, fsm_output[3]);
  assign nand_tmp_42 = ~((fsm_output[6]) & (~ mux_433_itm));
  assign or_507_nl = (~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[1]) | (~
      (fsm_output[7]));
  assign or_505_nl = (fsm_output[2]) | (~ and_dcpl_86);
  assign mux_434_nl = MUX_s_1_2_2(or_507_nl, or_505_nl, fsm_output[3]);
  assign or_508_nl = (fsm_output[6]) | mux_434_nl;
  assign mux_435_nl = MUX_s_1_2_2(or_508_nl, nand_tmp_42, fsm_output[0]);
  assign and_dcpl_111 = (~ mux_435_nl) & and_dcpl_110;
  assign and_dcpl_117 = (~((~((fsm_output[1]) ^ (fsm_output[2]))) | (fsm_output[7])
      | (fsm_output[8]) | (fsm_output[3]))) & (~ (fsm_output[6])) & (~ (fsm_output[4]))
      & and_dcpl_13;
  assign or_tmp_476 = and_256_cse | (fsm_output[8:7]!=2'b00);
  assign and_tmp_7 = (fsm_output[9]) & ((fsm_output[4]) | (fsm_output[6]) | or_tmp_476);
  assign and_dcpl_119 = (~ (fsm_output[8])) & (fsm_output[2]);
  assign nor_227_nl = ~((fsm_output[0]) | (fsm_output[3]));
  assign and_253_nl = (fsm_output[0]) & (fsm_output[3]);
  assign mux_438_nl = MUX_s_1_2_2(nor_227_nl, and_253_nl, fsm_output[4]);
  assign and_dcpl_123 = mux_438_nl & and_dcpl_47 & and_dcpl_119 & (~ (fsm_output[6]))
      & and_dcpl_13;
  assign or_tmp_483 = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[1]) | (~
      (fsm_output[7]));
  assign mux_439_nl = MUX_s_1_2_2(or_tmp_470, (fsm_output[8]), fsm_output[2]);
  assign mux_tmp_440 = MUX_s_1_2_2((~ mux_439_nl), or_tmp_483, fsm_output[3]);
  assign or_tmp_484 = (~ (fsm_output[1])) | (fsm_output[7]);
  assign and_tmp_8 = (fsm_output[8]) & or_tmp_484;
  assign mux_447_nl = MUX_s_1_2_2(or_tmp_470, and_tmp_8, fsm_output[2]);
  assign mux_tmp_448 = MUX_s_1_2_2((~ mux_447_nl), or_tmp_483, fsm_output[3]);
  assign or_531_nl = (fsm_output[8]) | (fsm_output[1]) | (fsm_output[7]);
  assign mux_tmp_455 = MUX_s_1_2_2(or_826_cse, or_531_nl, fsm_output[2]);
  assign nor_362_nl = ~((~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[3]) |
      (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]));
  assign nor_363_nl = ~((fsm_output[9]) | (~((fsm_output[1]) & (fsm_output[3]) &
      (fsm_output[4]) & (fsm_output[6]) & (fsm_output[7]))));
  assign mux_673_nl = MUX_s_1_2_2(nor_362_nl, nor_363_nl, fsm_output[5]);
  assign and_dcpl_129 = mux_673_nl & and_dcpl_119 & (~ (fsm_output[0]));
  assign and_dcpl_130 = and_dcpl_44 & and_dcpl_13;
  assign and_dcpl_134 = and_dcpl_48 & and_256_cse & and_dcpl_130;
  assign or_571_nl = (fsm_output[8]) | (~ mux_tmp_431);
  assign or_570_nl = (~ (fsm_output[8])) | (~ (fsm_output[1])) | (fsm_output[7]);
  assign mux_503_nl = MUX_s_1_2_2(or_571_nl, or_570_nl, fsm_output[2]);
  assign mux_tmp_504 = MUX_s_1_2_2(mux_503_nl, or_tmp_483, fsm_output[3]);
  assign or_572_nl = (fsm_output[6]) | mux_tmp_504;
  assign mux_505_nl = MUX_s_1_2_2(nand_tmp_42, or_572_nl, fsm_output[0]);
  assign and_dcpl_138 = (~ mux_505_nl) & and_dcpl_110;
  assign nor_tmp_81 = (fsm_output[5:3]==3'b111);
  assign and_306_nl = (fsm_output[3]) & (fsm_output[5]);
  assign mux_tmp_506 = MUX_s_1_2_2(and_306_nl, nor_tmp_81, fsm_output[2]);
  assign nor_tmp_83 = or_899_cse & (fsm_output[5:4]==2'b11);
  assign nor_211_nl = ~((fsm_output[5:4]!=2'b00));
  assign mux_508_nl = MUX_s_1_2_2(nor_211_nl, and_213_cse, fsm_output[3]);
  assign mux_tmp_509 = MUX_s_1_2_2(mux_508_nl, nor_tmp_81, fsm_output[2]);
  assign or_tmp_539 = ~(nand_119_cse & and_213_cse);
  assign nor_tmp_86 = or_tmp_416 & (fsm_output[5]);
  assign mux_tmp_522 = MUX_s_1_2_2(nor_tmp_81, nor_tmp_86, fsm_output[2]);
  assign or_tmp_548 = ~((fsm_output[8]) & (fsm_output[2]) & (~ (fsm_output[3])) &
      (fsm_output[4]));
  assign or_587_nl = (fsm_output[8]) | (fsm_output[2]) | (fsm_output[3]) | (~ (fsm_output[4]));
  assign mux_tmp_530 = MUX_s_1_2_2(or_587_nl, or_tmp_548, fsm_output[1]);
  assign nor_208_nl = ~((fsm_output[7:6]!=2'b10) | mux_tmp_530);
  assign or_588_nl = (fsm_output[8]) | (~ (fsm_output[2])) | (~ (fsm_output[3]))
      | (fsm_output[4]);
  assign mux_531_nl = MUX_s_1_2_2(or_tmp_548, or_588_nl, fsm_output[1]);
  assign mux_532_nl = MUX_s_1_2_2(mux_531_nl, mux_tmp_530, fsm_output[7]);
  assign and_239_nl = (fsm_output[6]) & (~ mux_532_nl);
  assign not_tmp_231 = MUX_s_1_2_2(nor_208_nl, and_239_nl, fsm_output[0]);
  assign or_tmp_562 = (((fsm_output[2]) | (~ (fsm_output[7]))) & (fsm_output[3]))
      | (fsm_output[4]);
  assign or_600_nl = (fsm_output[4:2]!=3'b000);
  assign mux_tmp_537 = MUX_s_1_2_2(or_600_nl, or_tmp_562, fsm_output[8]);
  assign or_tmp_567 = (~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[3]))))
      | (fsm_output[4]);
  assign mux_tmp_546 = MUX_s_1_2_2((~ or_756_cse), or_756_cse, fsm_output[7]);
  assign mux_tmp_549 = MUX_s_1_2_2(mux_tmp_546, or_tmp_567, fsm_output[8]);
  assign or_tmp_573 = (fsm_output[2]) | (~((fsm_output[3]) & (fsm_output[8])));
  assign and_dcpl_147 = and_dcpl_101 & and_dcpl_40;
  assign nor_nl = ~((fsm_output[1]) | (fsm_output[8]));
  assign mux_tmp_579 = MUX_s_1_2_2(nor_nl, nor_tmp_40, fsm_output[2]);
  assign and_dcpl_154 = mux_tmp_579 & (~ (fsm_output[7])) & (~ (fsm_output[3]));
  assign nor_189_nl = ~((fsm_output[6]) | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (~ (fsm_output[5])) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[3]));
  assign nor_190_nl = ~((fsm_output[6]) | (~ (fsm_output[2])) | (~ (fsm_output[4]))
      | (~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[3])));
  assign mux_584_nl = MUX_s_1_2_2(nor_189_nl, nor_190_nl, fsm_output[7]);
  assign nor_191_nl = ~((fsm_output[6]) | (~ (fsm_output[2])) | (fsm_output[4]) |
      (~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[3])));
  assign nor_192_nl = ~((~ (fsm_output[6])) | (fsm_output[2]) | (fsm_output[4]) |
      (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[3]));
  assign mux_583_nl = MUX_s_1_2_2(nor_191_nl, nor_192_nl, fsm_output[7]);
  assign mux_585_nl = MUX_s_1_2_2(mux_584_nl, mux_583_nl, fsm_output[1]);
  assign nor_193_nl = ~((fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[3]));
  assign nor_194_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[4])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[3])));
  assign mux_581_nl = MUX_s_1_2_2(nor_193_nl, nor_194_nl, fsm_output[6]);
  assign and_229_nl = (fsm_output[7]) & mux_581_nl;
  assign or_643_nl = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[3]);
  assign or_642_nl = (fsm_output[2]) | (~ (fsm_output[4])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[3]));
  assign mux_580_nl = MUX_s_1_2_2(or_643_nl, or_642_nl, fsm_output[6]);
  assign nor_195_nl = ~((fsm_output[7]) | mux_580_nl);
  assign mux_582_nl = MUX_s_1_2_2(and_229_nl, nor_195_nl, fsm_output[1]);
  assign not_tmp_260 = MUX_s_1_2_2(mux_585_nl, mux_582_nl, fsm_output[0]);
  assign or_tmp_621 = (~ (fsm_output[2])) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign or_tmp_623 = (fsm_output[4]) | (~ (fsm_output[8]));
  assign or_659_nl = (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_tmp_588 = MUX_s_1_2_2(or_tmp_623, or_659_nl, fsm_output[2]);
  assign mux_tmp_589 = MUX_s_1_2_2(mux_tmp_588, or_tmp_621, fsm_output[1]);
  assign mux_tmp_594 = MUX_s_1_2_2((fsm_output[4]), or_tmp_623, fsm_output[2]);
  assign mux_598_nl = MUX_s_1_2_2((fsm_output[4]), or_tmp_623, or_94_cse);
  assign or_669_nl = (~((fsm_output[2:1]!=2'b00))) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign mux_tmp_599 = MUX_s_1_2_2(mux_598_nl, or_669_nl, fsm_output[3]);
  assign or_tmp_635 = (fsm_output[4]) | (fsm_output[8]);
  assign or_tmp_637 = (fsm_output[2]) | (~ (fsm_output[4])) | (fsm_output[8]);
  assign nor_tmp_103 = (fsm_output[2]) & (fsm_output[4]);
  assign or_73_nl = (fsm_output[2]) | (fsm_output[4]);
  assign mux_623_nl = MUX_s_1_2_2(or_73_nl, (~ nor_tmp_103), fsm_output[3]);
  assign mux_54_nl = MUX_s_1_2_2((fsm_output[4]), or_tmp_51, fsm_output[3]);
  assign mux_tmp_624 = MUX_s_1_2_2(mux_623_nl, mux_54_nl, fsm_output[8]);
  assign or_tmp_654 = (~(VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm | (~ (fsm_output[1]))))
      | (fsm_output[2]) | (fsm_output[4]);
  assign or_tmp_656 = (((~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[1]))
      & (fsm_output[2])) | (fsm_output[4]);
  assign or_694_nl = (fsm_output[3]) | or_tmp_656;
  assign mux_636_nl = MUX_s_1_2_2((fsm_output[4]), or_tmp_654, fsm_output[3]);
  assign mux_tmp_637 = MUX_s_1_2_2(or_694_nl, mux_636_nl, fsm_output[8]);
  assign or_tmp_670 = (~ (fsm_output[2])) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign or_708_nl = (fsm_output[2]) | (fsm_output[0]) | (fsm_output[6]);
  assign mux_tmp_668 = MUX_s_1_2_2(or_708_nl, or_tmp_670, fsm_output[7]);
  assign mux_tmp_711 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign mux_tmp_722 = MUX_s_1_2_2((fsm_output[4]), (fsm_output[7]), fsm_output[5]);
  assign or_tmp_716 = (~ (fsm_output[4])) | (fsm_output[7]);
  assign mux_tmp_723 = MUX_s_1_2_2((~ or_tmp_716), (fsm_output[7]), fsm_output[5]);
  assign and_tmp_14 = (fsm_output[5]) & or_tmp_716;
  assign and_dcpl_175 = and_dcpl_154 & and_dcpl_147;
  assign nand_74_nl = ~((fsm_output[6]) & (fsm_output[1]) & (fsm_output[7]) & (fsm_output[8])
      & (~ (fsm_output[2])));
  assign or_797_nl = (fsm_output[6]) | (fsm_output[1]) | (~ (fsm_output[7])) | (~
      (fsm_output[8])) | (fsm_output[2]);
  assign mux_756_nl = MUX_s_1_2_2(nand_74_nl, or_797_nl, fsm_output[0]);
  assign nor_158_nl = ~((fsm_output[4]) | mux_756_nl);
  assign nor_159_nl = ~((fsm_output[4]) | (fsm_output[0]) | (fsm_output[6]) | (~
      (fsm_output[1])) | (fsm_output[7]) | (fsm_output[8]) | (fsm_output[2]));
  assign mux_757_nl = MUX_s_1_2_2(nor_158_nl, nor_159_nl, fsm_output[5]);
  assign nor_160_nl = ~((fsm_output[0]) | (fsm_output[6]) | (fsm_output[1]) | (fsm_output[7])
      | (~ (fsm_output[8])) | (fsm_output[2]));
  assign nor_161_nl = ~((fsm_output[6]) | (fsm_output[1]) | (~ (fsm_output[7])) |
      (fsm_output[8]) | (~ (fsm_output[2])));
  assign nor_162_nl = ~((~ (fsm_output[7])) | (fsm_output[8]) | (~ (fsm_output[2])));
  assign nor_163_nl = ~((fsm_output[7]) | (fsm_output[8]) | (fsm_output[2]));
  assign mux_753_nl = MUX_s_1_2_2(nor_162_nl, nor_163_nl, fsm_output[1]);
  assign and_209_nl = (fsm_output[6]) & mux_753_nl;
  assign mux_754_nl = MUX_s_1_2_2(nor_161_nl, and_209_nl, fsm_output[0]);
  assign mux_755_nl = MUX_s_1_2_2(nor_160_nl, mux_754_nl, fsm_output[4]);
  assign and_208_nl = (fsm_output[5]) & mux_755_nl;
  assign mux_758_nl = MUX_s_1_2_2(mux_757_nl, and_208_nl, fsm_output[3]);
  assign nor_164_nl = ~((fsm_output[8:0]!=9'b000000011));
  assign not_tmp_321 = MUX_s_1_2_2(mux_758_nl, nor_164_nl, fsm_output[9]);
  assign or_tmp_760 = (~((~ (fsm_output[8])) | (fsm_output[4]))) | (fsm_output[9])
      | (~ (fsm_output[5]));
  assign or_801_nl = (~((fsm_output[8]) | (~ (fsm_output[4])))) | (fsm_output[9])
      | (~ (fsm_output[5]));
  assign mux_tmp_760 = MUX_s_1_2_2(or_tmp_760, or_801_nl, fsm_output[3]);
  assign or_tmp_762 = (~((fsm_output[7]) | (fsm_output[8]) | (~ (fsm_output[4]))))
      | (fsm_output[9]) | (~ (fsm_output[5]));
  assign or_tmp_769 = (~((~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[4])))
      | (fsm_output[9]) | (~ (fsm_output[5]));
  assign mux_tmp_763 = MUX_s_1_2_2(or_1038_cse, or_55_cse, fsm_output[4]);
  assign and_292_nl = (fsm_output[8:7]==2'b11);
  assign mux_tmp_771 = MUX_s_1_2_2(or_54_cse, mux_894_cse, and_292_nl);
  assign and_dcpl_176 = ~((fsm_output[0]) | (fsm_output[9]));
  assign nor_150_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[3]) |
      (~ (fsm_output[8])) | (fsm_output[1]));
  assign nor_151_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (fsm_output[8]) | (~ (fsm_output[1])));
  assign not_tmp_324 = MUX_s_1_2_2(nor_150_nl, nor_151_nl, fsm_output[5]);
  assign or_831_nl = (fsm_output[2]) | (fsm_output[8]) | (~ and_dcpl_72);
  assign mux_784_nl = MUX_s_1_2_2(or_831_nl, or_tmp_483, fsm_output[3]);
  assign or_832_nl = (fsm_output[6]) | mux_784_nl;
  assign mux_785_nl = MUX_s_1_2_2(nand_tmp_42, or_832_nl, fsm_output[0]);
  assign and_dcpl_179 = (~ mux_785_nl) & and_dcpl_110;
  assign or_27_nl = (~ (fsm_output[6])) | (fsm_output[3]);
  assign mux_tmp_787 = MUX_s_1_2_2(mux_894_cse, or_54_cse, or_27_nl);
  assign mux_796_nl = MUX_s_1_2_2(or_1038_cse, or_55_cse, or_756_cse);
  assign mux_797_nl = MUX_s_1_2_2(mux_796_nl, or_tmp_29, fsm_output[6]);
  assign mux_798_nl = MUX_s_1_2_2(mux_797_nl, or_tmp_31, and_524_cse);
  assign mux_799_nl = MUX_s_1_2_2(mux_798_nl, or_tmp_29, fsm_output[7]);
  assign nor_132_nl = ~((~ (fsm_output[7])) | (fsm_output[0]) | (fsm_output[1]) |
      (~ (fsm_output[6])));
  assign mux_795_nl = MUX_s_1_2_2(or_tmp_31, or_tmp_29, nor_132_nl);
  assign mux_800_nl = MUX_s_1_2_2(mux_799_nl, mux_795_nl, fsm_output[2]);
  assign mux_792_nl = MUX_s_1_2_2(mux_tmp_787, or_tmp_29, or_590_cse);
  assign mux_39_nl = MUX_s_1_2_2(mux_894_cse, or_54_cse, fsm_output[3]);
  assign or_843_nl = (~((~((fsm_output[6]) | (~ (fsm_output[3])))) | (fsm_output[4])))
      | (fsm_output[9]) | (~ (fsm_output[5]));
  assign mux_790_nl = MUX_s_1_2_2(mux_39_nl, or_843_nl, fsm_output[1]);
  assign mux_788_nl = MUX_s_1_2_2(mux_tmp_787, or_tmp_29, fsm_output[1]);
  assign mux_791_nl = MUX_s_1_2_2(mux_790_nl, mux_788_nl, fsm_output[0]);
  assign mux_793_nl = MUX_s_1_2_2(mux_792_nl, mux_791_nl, fsm_output[7]);
  assign mux_794_nl = MUX_s_1_2_2(mux_793_nl, or_tmp_29, fsm_output[2]);
  assign mux_801_itm = MUX_s_1_2_2(mux_800_nl, mux_794_nl, fsm_output[8]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_38 & and_dcpl_28 & nor_tmp_34;
  assign VEC_LOOP_j_1_12_0_sva_11_0_mx0c1 = and_dcpl_49 & and_dcpl_101 & nor_tmp_34;
  assign or_9_nl = (fsm_output[8]) | (fsm_output[3]) | (fsm_output[7]) | (fsm_output[6]);
  assign or_556_nl = (fsm_output[6]) | (fsm_output[3]) | mux_tmp_455;
  assign mux_495_nl = MUX_s_1_2_2(or_9_nl, or_556_nl, fsm_output[0]);
  assign nor_217_nl = ~((fsm_output[4]) | mux_495_nl);
  assign mux_496_nl = MUX_s_1_2_2(nor_217_nl, or_814_cse, fsm_output[9]);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(mux_496_nl, and_tmp_7, fsm_output[5]);
  assign or_914_nl = (fsm_output[0]) | (~ (fsm_output[6])) | (fsm_output[3]) | (fsm_output[2])
      | (~ (fsm_output[8])) | (fsm_output[1]);
  assign or_915_nl = (~ (fsm_output[0])) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[1]));
  assign mux_501_nl = MUX_s_1_2_2(or_914_nl, or_915_nl, fsm_output[4]);
  assign or_916_nl = (~ (fsm_output[4])) | (fsm_output[0]) | (fsm_output[6]) | (~
      (fsm_output[3])) | (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[1]));
  assign mux_502_nl = MUX_s_1_2_2(mux_501_nl, or_916_nl, fsm_output[5]);
  assign nor_359_m1c = ~(mux_502_nl | (fsm_output[7]) | (fsm_output[9]));
  assign and_160_m1c = and_dcpl_73 & nor_236_cse & and_dcpl_147;
  assign and_163_m1c = and_dcpl_65 & (fsm_output[8]) & and_dcpl_46 & and_dcpl_147;
  assign or_184_nl = (~ (fsm_output[9])) | (fsm_output[7]) | (~ (fsm_output[0]))
      | (fsm_output[6]);
  assign mux_165_cse = MUX_s_1_2_2(or_184_nl, or_tmp_148, fsm_output[8]);
  assign or_180_nl = (fsm_output[9]) | (fsm_output[7]) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_163_cse = MUX_s_1_2_2(or_tmp_148, or_180_nl, fsm_output[8]);
  assign and_61_nl = not_tmp_91 & (~ (fsm_output[7])) & and_dcpl_52 & and_dcpl_13;
  assign or_186_nl = (fsm_output[9:8]!=2'b00) | mux_tmp_162;
  assign mux_166_nl = MUX_s_1_2_2(or_186_nl, mux_165_cse, fsm_output[3]);
  assign nor_307_nl = ~((fsm_output[2]) | mux_166_nl);
  assign nor_308_nl = ~((fsm_output[3]) | mux_163_cse);
  assign nor_309_nl = ~((fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[9]) |
      mux_tmp_162);
  assign mux_164_nl = MUX_s_1_2_2(nor_308_nl, nor_309_nl, fsm_output[2]);
  assign mux_167_nl = MUX_s_1_2_2(nor_307_nl, mux_164_nl, fsm_output[1]);
  assign and_63_nl = mux_167_nl & (fsm_output[5:4]==2'b10);
  assign nor_304_nl = ~((fsm_output[3]) | (fsm_output[9]) | (fsm_output[7]));
  assign nor_305_nl = ~((~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[7])));
  assign mux_169_nl = MUX_s_1_2_2(nor_304_nl, nor_305_nl, fsm_output[8]);
  assign and_283_nl = (~((fsm_output[6:4]!=3'b110))) & mux_169_nl;
  assign or_190_nl = (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_189_nl = (~ (fsm_output[9])) | (fsm_output[7]);
  assign mux_168_nl = MUX_s_1_2_2(or_190_nl, or_189_nl, fsm_output[3]);
  assign nor_306_nl = ~((~ (fsm_output[4])) | (fsm_output[5]) | (fsm_output[6]) |
      (fsm_output[8]) | mux_168_nl);
  assign mux_170_nl = MUX_s_1_2_2(and_283_nl, nor_306_nl, fsm_output[2]);
  assign and_65_nl = mux_170_nl & (fsm_output[1:0]==2'b01);
  assign nor_301_nl = ~((~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[1])));
  assign nor_302_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[1]));
  assign mux_172_nl = MUX_s_1_2_2(nor_301_nl, nor_302_nl, fsm_output[3]);
  assign and_282_nl = (fsm_output[4]) & (fsm_output[6]) & mux_172_nl;
  assign nor_303_nl = ~((fsm_output[4]) | (fsm_output[6]) | mux_tmp_92);
  assign mux_173_nl = MUX_s_1_2_2(and_282_nl, nor_303_nl, fsm_output[5]);
  assign and_70_nl = mux_173_nl & (fsm_output[7]) & (~ (fsm_output[0])) & (~ (fsm_output[9]));
  assign or_209_nl = (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[7]);
  assign or_208_nl = (fsm_output[2]) | (~((fsm_output[8:7]==2'b11)));
  assign mux_175_nl = MUX_s_1_2_2(or_209_nl, or_208_nl, fsm_output[3]);
  assign nor_299_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | mux_175_nl);
  assign or_205_nl = (fsm_output[8:7]!=2'b01);
  assign or_204_nl = (fsm_output[8:7]!=2'b10);
  assign mux_174_nl = MUX_s_1_2_2(or_205_nl, or_204_nl, fsm_output[2]);
  assign nor_300_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[3]) |
      mux_174_nl);
  assign mux_176_nl = MUX_s_1_2_2(nor_299_nl, nor_300_nl, fsm_output[5]);
  assign and_77_nl = mux_176_nl & (fsm_output[1]) & (fsm_output[0]) & (~ (fsm_output[9]));
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_10_7_2(z_out_1, (z_out_6[12:3]), COMP_LOOP_acc_psp_1_sva,
      (COMP_LOOP_acc_10_cse_12_1_1_sva[11:2]), (COMP_LOOP_acc_1_cse_5_sva[11:2]),
      (COMP_LOOP_acc_11_psp_1_sva[10:1]), (COMP_LOOP_acc_1_cse_2_sva[11:2]), {COMP_LOOP_or_1_cse
      , COMP_LOOP_or_3_cse , and_61_nl , and_63_nl , and_65_nl , and_70_nl , and_77_nl});
  assign vec_rsc_0_0_i_da_d_pff = modExp_base_1_sva_mx1;
  assign nor_292_nl = ~((~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | mux_190_cse);
  assign or_224_nl = (VEC_LOOP_j_1_12_0_sva_11_0[1]) | (fsm_output[9:7]!=3'b000);
  assign or_223_nl = (COMP_LOOP_acc_11_psp_1_sva[0]) | (fsm_output[9:7]!=3'b001);
  assign mux_181_nl = MUX_s_1_2_2(or_224_nl, or_223_nl, fsm_output[1]);
  assign nor_294_nl = ~((~ (fsm_output[2])) | (VEC_LOOP_j_1_12_0_sva_11_0[0]) | mux_181_nl);
  assign nor_295_nl = ~((~ (fsm_output[1])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b00)
      | (fsm_output[9:7]!=3'b010));
  assign nor_296_nl = ~((fsm_output[1]) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) | (COMP_LOOP_acc_11_psp_1_sva[0])
      | (fsm_output[9:7]!=3'b011));
  assign mux_180_nl = MUX_s_1_2_2(nor_295_nl, nor_296_nl, fsm_output[2]);
  assign mux_182_nl = MUX_s_1_2_2(nor_294_nl, mux_180_nl, fsm_output[3]);
  assign nand_11_nl = ~((fsm_output[6]) & mux_182_nl);
  assign nor_297_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b00) | (fsm_output[9:7]!=3'b001));
  assign nor_298_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00) | (fsm_output[9:7]!=3'b010));
  assign mux_178_nl = MUX_s_1_2_2(nor_297_nl, nor_298_nl, fsm_output[1]);
  assign nand_10_nl = ~((fsm_output[2]) & mux_178_nl);
  assign or_213_nl = (~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00)
      | (fsm_output[9:7]!=3'b011);
  assign or_211_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b00) |
      (fsm_output[9:7]!=3'b100);
  assign mux_177_nl = MUX_s_1_2_2(or_213_nl, or_211_nl, fsm_output[2]);
  assign mux_179_nl = MUX_s_1_2_2(nand_10_nl, mux_177_nl, fsm_output[3]);
  assign or_217_nl = (fsm_output[6]) | mux_179_nl;
  assign mux_183_nl = MUX_s_1_2_2(nand_11_nl, or_217_nl, fsm_output[0]);
  assign nor_293_nl = ~((fsm_output[5]) | mux_183_nl);
  assign vec_rsc_0_0_i_wea_d_pff = MUX_s_1_2_2(nor_292_nl, nor_293_nl, fsm_output[4]);
  assign or_254_cse = (z_out_6[2:1]!=2'b00) | (~ (fsm_output[7])) | (~ (fsm_output[2]))
      | (fsm_output[9]);
  assign or_266_nl = (fsm_output[1]) | (fsm_output[7]) | (z_out_6[2:1]!=2'b00) |
      not_tmp_108;
  assign or_264_nl = (~ (fsm_output[1])) | (~ (fsm_output[7])) | (fsm_output[2])
      | (fsm_output[9]);
  assign mux_204_nl = MUX_s_1_2_2(or_266_nl, or_264_nl, fsm_output[8]);
  assign or_267_nl = (fsm_output[3]) | mux_204_nl;
  assign or_263_nl = (fsm_output[3]) | (fsm_output[8]) | (fsm_output[1]) | (fsm_output[7])
      | (z_out_6[2:1]!=2'b00) | not_tmp_108;
  assign or_261_nl = (z_out_6[2:1]!=2'b00);
  assign mux_205_nl = MUX_s_1_2_2(or_267_nl, or_263_nl, or_261_nl);
  assign or_259_nl = (VEC_LOOP_j_1_12_0_sva_11_0[1]) | (fsm_output[7]) | (fsm_output[2])
      | (fsm_output[9]);
  assign or_258_nl = (COMP_LOOP_acc_11_psp_1_sva[0]) | (~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_201_nl = MUX_s_1_2_2(or_259_nl, or_258_nl, fsm_output[1]);
  assign or_260_nl = (VEC_LOOP_j_1_12_0_sva_11_0[0]) | mux_201_nl;
  assign or_257_nl = (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b00) | (~ (fsm_output[1]))
      | (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign mux_202_nl = MUX_s_1_2_2(or_260_nl, or_257_nl, fsm_output[8]);
  assign or_256_nl = (~ (fsm_output[8])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) |
      (fsm_output[1]) | (COMP_LOOP_acc_11_psp_1_sva[0]) | (~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_203_nl = MUX_s_1_2_2(mux_202_nl, or_256_nl, fsm_output[3]);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, mux_203_nl, fsm_output[5]);
  assign nor_282_nl = ~((fsm_output[0]) | mux_206_nl);
  assign or_253_nl = (z_out_6[2:1]!=2'b00) | (fsm_output[7]) | (fsm_output[2]) |
      (fsm_output[9]);
  assign mux_200_nl = MUX_s_1_2_2(or_254_cse, or_253_nl, fsm_output[1]);
  assign nor_283_nl = ~((~((fsm_output[0]) & (fsm_output[5]) & (fsm_output[3]) &
      (~ (fsm_output[8])))) | mux_200_nl);
  assign mux_207_nl = MUX_s_1_2_2(nor_282_nl, nor_283_nl, fsm_output[4]);
  assign nor_284_nl = ~((z_out_6[2:1]!=2'b00) | (fsm_output[7]) | (fsm_output[2])
      | (fsm_output[9]));
  assign nor_285_nl = ~((z_out_6[2:1]!=2'b00) | (~ (fsm_output[7])) | (fsm_output[2])
      | (fsm_output[9]));
  assign mux_197_nl = MUX_s_1_2_2(nor_284_nl, nor_285_nl, fsm_output[1]);
  assign and_281_nl = (~((fsm_output[3]) | (~ (fsm_output[8])))) & mux_197_nl;
  assign nor_286_nl = ~((~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (fsm_output[7])
      | (fsm_output[2]) | (fsm_output[9]));
  assign nor_287_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[9]));
  assign mux_193_nl = MUX_s_1_2_2(nor_286_nl, nor_287_nl, fsm_output[1]);
  assign nor_288_nl = ~((~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00)
      | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[7]))
      | (fsm_output[2]) | (fsm_output[9]));
  assign or_246_nl = (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b00);
  assign mux_194_nl = MUX_s_1_2_2(mux_193_nl, nor_288_nl, or_246_nl);
  assign nor_289_nl = ~((~ (fsm_output[1])) | (~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00) | (fsm_output[7]) | (~ (fsm_output[2]))
      | (fsm_output[9]));
  assign mux_195_nl = MUX_s_1_2_2(mux_194_nl, nor_289_nl, fsm_output[8]);
  assign nor_290_nl = ~((~ (fsm_output[8])) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b00)
      | (fsm_output[1]) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~
      (fsm_output[7])) | (fsm_output[2]) | (fsm_output[9]));
  assign mux_196_nl = MUX_s_1_2_2(mux_195_nl, nor_290_nl, fsm_output[3]);
  assign mux_198_nl = MUX_s_1_2_2(and_281_nl, mux_196_nl, fsm_output[5]);
  assign and_280_nl = (fsm_output[0]) & mux_198_nl;
  assign or_242_nl = (z_out_6[2:1]!=2'b00) | (fsm_output[7]) | (~ (fsm_output[2]))
      | (fsm_output[9]);
  assign mux_192_nl = MUX_s_1_2_2(or_242_nl, or_254_cse, fsm_output[1]);
  assign nor_291_nl = ~((fsm_output[0]) | (~ (fsm_output[5])) | (~ (fsm_output[3]))
      | (fsm_output[8]) | mux_192_nl);
  assign mux_199_nl = MUX_s_1_2_2(and_280_nl, nor_291_nl, fsm_output[4]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_207_nl,
      mux_199_nl, fsm_output[6]);
  assign nor_274_nl = ~((~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01)
      | mux_190_cse);
  assign nor_277_nl = ~((COMP_LOOP_acc_11_psp_1_sva[0]) | (fsm_output[9:7]!=3'b001));
  assign mux_213_nl = MUX_s_1_2_2(nor_268_cse, nor_277_nl, fsm_output[1]);
  assign and_279_nl = (fsm_output[2]) & (VEC_LOOP_j_1_12_0_sva_11_0[0]) & mux_213_nl;
  assign nor_278_nl = ~((~ (fsm_output[1])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b01)
      | (fsm_output[9:7]!=3'b010));
  assign nor_279_nl = ~((fsm_output[1]) | (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]))
      | (COMP_LOOP_acc_11_psp_1_sva[0]) | (fsm_output[9:7]!=3'b011));
  assign mux_212_nl = MUX_s_1_2_2(nor_278_nl, nor_279_nl, fsm_output[2]);
  assign mux_214_nl = MUX_s_1_2_2(and_279_nl, mux_212_nl, fsm_output[3]);
  assign nand_17_nl = ~((fsm_output[6]) & mux_214_nl);
  assign nor_280_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b01) | (fsm_output[9:7]!=3'b001));
  assign nor_281_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01) | (fsm_output[9:7]!=3'b010));
  assign mux_210_nl = MUX_s_1_2_2(nor_280_nl, nor_281_nl, fsm_output[1]);
  assign nand_15_nl = ~((fsm_output[2]) & mux_210_nl);
  assign or_271_nl = (~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01)
      | (fsm_output[9:7]!=3'b011);
  assign or_269_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b01) |
      (fsm_output[9:7]!=3'b100);
  assign mux_209_nl = MUX_s_1_2_2(or_271_nl, or_269_nl, fsm_output[2]);
  assign mux_211_nl = MUX_s_1_2_2(nand_15_nl, mux_209_nl, fsm_output[3]);
  assign or_275_nl = (fsm_output[6]) | mux_211_nl;
  assign mux_215_nl = MUX_s_1_2_2(nand_17_nl, or_275_nl, fsm_output[0]);
  assign nor_275_nl = ~((fsm_output[5]) | mux_215_nl);
  assign vec_rsc_0_1_i_wea_d_pff = MUX_s_1_2_2(nor_274_nl, nor_275_nl, fsm_output[4]);
  assign or_322_nl = (fsm_output[1]) | (fsm_output[7]) | (z_out_6[2:1]!=2'b01) |
      (fsm_output[9:8]!=2'b10);
  assign mux_240_nl = MUX_s_1_2_2(nand_95_cse, or_322_nl, fsm_output[2]);
  assign or_324_nl = (fsm_output[3]) | mux_240_nl;
  assign or_320_nl = (fsm_output[3]) | (~ (fsm_output[2])) | (fsm_output[1]) | (fsm_output[7])
      | (z_out_6[2:1]!=2'b01) | (fsm_output[9:8]!=2'b10);
  assign or_318_nl = (z_out_6[2:1]!=2'b01);
  assign mux_241_nl = MUX_s_1_2_2(or_324_nl, or_320_nl, or_318_nl);
  assign mux_236_nl = MUX_s_1_2_2(nor_268_cse, nor_269_cse, fsm_output[1]);
  assign nand_22_nl = ~((VEC_LOOP_j_1_12_0_sva_11_0[0]) & mux_236_nl);
  assign mux_237_nl = MUX_s_1_2_2(nand_22_nl, or_tmp_278, fsm_output[2]);
  assign mux_238_nl = MUX_s_1_2_2(mux_237_nl, or_315_cse, fsm_output[3]);
  assign or_313_nl = (~ (VEC_LOOP_j_1_12_0_sva_11_0[0])) | (fsm_output[1]) | (VEC_LOOP_j_1_12_0_sva_11_0[1])
      | (fsm_output[9:7]!=3'b000);
  assign mux_235_nl = MUX_s_1_2_2(or_313_nl, or_tmp_278, fsm_output[2]);
  assign or_314_nl = (fsm_output[3]) | mux_235_nl;
  assign or_311_nl = (~ VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm) | (COMP_LOOP_acc_11_psp_1_sva[0]);
  assign mux_239_nl = MUX_s_1_2_2(mux_238_nl, or_314_nl, or_311_nl);
  assign mux_242_nl = MUX_s_1_2_2(mux_241_nl, mux_239_nl, fsm_output[5]);
  assign nor_267_nl = ~((fsm_output[0]) | mux_242_nl);
  assign nor_270_nl = ~((z_out_6[2:1]!=2'b01) | (~ (fsm_output[1])) | (fsm_output[7])
      | (fsm_output[8]) | (fsm_output[9]));
  assign nor_271_nl = ~((z_out_6[2:1]!=2'b01) | (fsm_output[1]) | (~ (fsm_output[7]))
      | (fsm_output[8]) | (fsm_output[9]));
  assign mux_234_nl = MUX_s_1_2_2(nor_270_nl, nor_271_nl, fsm_output[2]);
  assign and_276_nl = (fsm_output[0]) & (fsm_output[5]) & (fsm_output[3]) & mux_234_nl;
  assign mux_243_nl = MUX_s_1_2_2(nor_267_nl, and_276_nl, fsm_output[4]);
  assign or_307_nl = (z_out_6[2:1]!=2'b01) | (fsm_output[9:7]!=3'b010);
  assign or_306_nl = (z_out_6[2:1]!=2'b01) | (fsm_output[9:7]!=3'b011);
  assign mux_231_nl = MUX_s_1_2_2(or_307_nl, or_306_nl, fsm_output[1]);
  assign or_308_nl = (fsm_output[3:2]!=2'b00) | mux_231_nl;
  assign or_299_nl = (fsm_output[2:1]!=2'b01) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01) | (fsm_output[9:7]!=3'b001);
  assign mux_225_nl = MUX_s_1_2_2(or_299_nl, or_tmp_264, fsm_output[3]);
  assign or_303_nl = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01)
      | (fsm_output[9:7]!=3'b001);
  assign mux_226_nl = MUX_s_1_2_2(or_304_cse, or_303_nl, fsm_output[1]);
  assign or_302_nl = (~ (fsm_output[1])) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01) | (fsm_output[9:7]!=3'b001);
  assign or_301_nl = (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b01);
  assign mux_227_nl = MUX_s_1_2_2(mux_226_nl, or_302_nl, or_301_nl);
  assign or_300_nl = (~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01)
      | (fsm_output[9:7]!=3'b010);
  assign mux_228_nl = MUX_s_1_2_2(mux_227_nl, or_300_nl, fsm_output[2]);
  assign mux_229_nl = MUX_s_1_2_2(mux_228_nl, or_tmp_264, fsm_output[3]);
  assign mux_230_nl = MUX_s_1_2_2(mux_225_nl, mux_229_nl, VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  assign mux_232_nl = MUX_s_1_2_2(or_308_nl, mux_230_nl, fsm_output[5]);
  assign and_277_nl = (fsm_output[0]) & (~ mux_232_nl);
  assign nor_272_nl = ~((z_out_6[2:1]!=2'b01) | (fsm_output[9:7]!=3'b000));
  assign nor_273_nl = ~((z_out_6[2:1]!=2'b01) | (fsm_output[9:7]!=3'b001));
  assign mux_224_nl = MUX_s_1_2_2(nor_272_nl, nor_273_nl, fsm_output[1]);
  assign and_278_nl = (~ (fsm_output[0])) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[2])
      & mux_224_nl;
  assign mux_233_nl = MUX_s_1_2_2(and_277_nl, and_278_nl, fsm_output[4]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_243_nl,
      mux_233_nl, fsm_output[6]);
  assign and_274_nl = (~((~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b10)))
      & mux_258_cse;
  assign or_338_nl = (~ (COMP_LOOP_acc_11_psp_1_sva[0])) | (fsm_output[9:7]!=3'b001);
  assign mux_249_nl = MUX_s_1_2_2(or_370_cse, or_338_nl, fsm_output[1]);
  assign nor_262_nl = ~((~ (fsm_output[2])) | (VEC_LOOP_j_1_12_0_sva_11_0[0]) | mux_249_nl);
  assign nor_263_nl = ~((~ (fsm_output[1])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b10)
      | (fsm_output[9:7]!=3'b010));
  assign nor_264_nl = ~((fsm_output[1]) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) | (~
      (COMP_LOOP_acc_11_psp_1_sva[0])) | (fsm_output[9:7]!=3'b011));
  assign mux_248_nl = MUX_s_1_2_2(nor_263_nl, nor_264_nl, fsm_output[2]);
  assign mux_250_nl = MUX_s_1_2_2(nor_262_nl, mux_248_nl, fsm_output[3]);
  assign nand_24_nl = ~((fsm_output[6]) & mux_250_nl);
  assign nor_265_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b10) | (fsm_output[9:7]!=3'b001));
  assign nor_266_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10) | (fsm_output[9:7]!=3'b010));
  assign mux_246_nl = MUX_s_1_2_2(nor_265_nl, nor_266_nl, fsm_output[1]);
  assign nand_23_nl = ~((fsm_output[2]) & mux_246_nl);
  assign or_328_nl = (~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10)
      | (fsm_output[9:7]!=3'b011);
  assign or_326_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b10) |
      (fsm_output[9:7]!=3'b100);
  assign mux_245_nl = MUX_s_1_2_2(or_328_nl, or_326_nl, fsm_output[2]);
  assign mux_247_nl = MUX_s_1_2_2(nand_23_nl, mux_245_nl, fsm_output[3]);
  assign or_332_nl = (fsm_output[6]) | mux_247_nl;
  assign mux_251_nl = MUX_s_1_2_2(nand_24_nl, or_332_nl, fsm_output[0]);
  assign nor_261_nl = ~((fsm_output[5]) | mux_251_nl);
  assign vec_rsc_0_2_i_wea_d_pff = MUX_s_1_2_2(and_274_nl, nor_261_nl, fsm_output[4]);
  assign or_379_nl = (fsm_output[3]) | (~ (fsm_output[2])) | (fsm_output[1]) | (fsm_output[7])
      | (z_out_6[2:1]!=2'b10) | (fsm_output[9:8]!=2'b10);
  assign or_375_nl = (fsm_output[1]) | (fsm_output[7]) | (z_out_6[2:1]!=2'b10) |
      (fsm_output[9:8]!=2'b10);
  assign mux_276_nl = MUX_s_1_2_2(nand_95_cse, or_375_nl, fsm_output[2]);
  assign or_377_nl = (fsm_output[3]) | mux_276_nl;
  assign nor_54_nl = ~((z_out_6[2:1]!=2'b10));
  assign mux_277_nl = MUX_s_1_2_2(or_379_nl, or_377_nl, nor_54_nl);
  assign or_372_nl = (VEC_LOOP_j_1_12_0_sva_11_0[0]) | (fsm_output[1]) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[1]))
      | (fsm_output[9:7]!=3'b000);
  assign mux_274_nl = MUX_s_1_2_2(or_372_nl, or_tmp_334, fsm_output[2]);
  assign or_373_nl = (fsm_output[3]) | mux_274_nl;
  assign mux_271_nl = MUX_s_1_2_2(or_370_cse, or_369_cse, fsm_output[1]);
  assign or_371_nl = (VEC_LOOP_j_1_12_0_sva_11_0[0]) | mux_271_nl;
  assign mux_272_nl = MUX_s_1_2_2(or_371_nl, or_tmp_334, fsm_output[2]);
  assign or_367_nl = (fsm_output[2]) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]) | (fsm_output[1])
      | (~ (fsm_output[7])) | (~ (fsm_output[8])) | (fsm_output[9]);
  assign mux_273_nl = MUX_s_1_2_2(mux_272_nl, or_367_nl, fsm_output[3]);
  assign mux_275_nl = MUX_s_1_2_2(or_373_nl, mux_273_nl, and_270_cse);
  assign mux_278_nl = MUX_s_1_2_2(mux_277_nl, mux_275_nl, fsm_output[5]);
  assign nor_255_nl = ~((fsm_output[0]) | mux_278_nl);
  assign nor_256_nl = ~((z_out_6[2:1]!=2'b10) | (~ (fsm_output[1])) | (fsm_output[7])
      | (fsm_output[8]) | (fsm_output[9]));
  assign nor_257_nl = ~((z_out_6[2:1]!=2'b10) | (fsm_output[1]) | (~ (fsm_output[7]))
      | (fsm_output[8]) | (fsm_output[9]));
  assign mux_270_nl = MUX_s_1_2_2(nor_256_nl, nor_257_nl, fsm_output[2]);
  assign and_271_nl = (fsm_output[0]) & (fsm_output[5]) & (fsm_output[3]) & mux_270_nl;
  assign mux_279_nl = MUX_s_1_2_2(nor_255_nl, and_271_nl, fsm_output[4]);
  assign or_363_nl = (z_out_6[2:1]!=2'b10) | (fsm_output[9:7]!=3'b010);
  assign or_362_nl = (z_out_6[2:1]!=2'b10) | (fsm_output[9:7]!=3'b011);
  assign mux_267_nl = MUX_s_1_2_2(or_363_nl, or_362_nl, fsm_output[1]);
  assign or_364_nl = (fsm_output[3:2]!=2'b00) | mux_267_nl;
  assign or_356_nl = (fsm_output[2:1]!=2'b01) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10) | (fsm_output[9:7]!=3'b001);
  assign mux_261_nl = MUX_s_1_2_2(or_356_nl, or_tmp_321, fsm_output[3]);
  assign or_360_nl = (~ (fsm_output[1])) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10) | (fsm_output[9:7]!=3'b001);
  assign or_358_nl = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10)
      | (fsm_output[9:7]!=3'b001);
  assign mux_262_nl = MUX_s_1_2_2(or_304_cse, or_358_nl, fsm_output[1]);
  assign nor_51_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b10));
  assign mux_263_nl = MUX_s_1_2_2(or_360_nl, mux_262_nl, nor_51_nl);
  assign or_357_nl = (~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10)
      | (fsm_output[9:7]!=3'b010);
  assign mux_264_nl = MUX_s_1_2_2(mux_263_nl, or_357_nl, fsm_output[2]);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, or_tmp_321, fsm_output[3]);
  assign mux_266_nl = MUX_s_1_2_2(mux_261_nl, mux_265_nl, VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  assign mux_268_nl = MUX_s_1_2_2(or_364_nl, mux_266_nl, fsm_output[5]);
  assign and_272_nl = (fsm_output[0]) & (~ mux_268_nl);
  assign nor_258_nl = ~((z_out_6[2:1]!=2'b10) | (fsm_output[9:7]!=3'b000));
  assign nor_259_nl = ~((z_out_6[2:1]!=2'b10) | (fsm_output[9:7]!=3'b001));
  assign mux_260_nl = MUX_s_1_2_2(nor_258_nl, nor_259_nl, fsm_output[1]);
  assign and_273_nl = (~ (fsm_output[0])) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[2])
      & mux_260_nl;
  assign mux_269_nl = MUX_s_1_2_2(and_272_nl, and_273_nl, fsm_output[4]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_279_nl,
      mux_269_nl, fsm_output[6]);
  assign and_267_nl = (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11)
      & mux_258_cse;
  assign nor_250_nl = ~((~ (COMP_LOOP_acc_11_psp_1_sva[0])) | (fsm_output[9:7]!=3'b001));
  assign mux_285_nl = MUX_s_1_2_2(nor_241_cse, nor_250_nl, fsm_output[1]);
  assign and_269_nl = (fsm_output[2]) & (VEC_LOOP_j_1_12_0_sva_11_0[0]) & mux_285_nl;
  assign nor_251_nl = ~((~ (fsm_output[1])) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b11)
      | (fsm_output[9:7]!=3'b010));
  assign nor_252_nl = ~((fsm_output[1]) | (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]))
      | (~ (COMP_LOOP_acc_11_psp_1_sva[0])) | (fsm_output[9:7]!=3'b011));
  assign mux_284_nl = MUX_s_1_2_2(nor_251_nl, nor_252_nl, fsm_output[2]);
  assign mux_286_nl = MUX_s_1_2_2(and_269_nl, mux_284_nl, fsm_output[3]);
  assign nand_32_nl = ~((fsm_output[6]) & mux_286_nl);
  assign nor_253_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b11) | (fsm_output[9:7]!=3'b001));
  assign nor_254_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b11) | (fsm_output[9:7]!=3'b010));
  assign mux_282_nl = MUX_s_1_2_2(nor_253_nl, nor_254_nl, fsm_output[1]);
  assign nand_30_nl = ~((fsm_output[2]) & mux_282_nl);
  assign nand_112_nl = ~((fsm_output[1]) & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b11)
      & (fsm_output[9:7]==3'b011));
  assign or_381_nl = (fsm_output[1]) | (COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b11) |
      (fsm_output[9:7]!=3'b100);
  assign mux_281_nl = MUX_s_1_2_2(nand_112_nl, or_381_nl, fsm_output[2]);
  assign mux_283_nl = MUX_s_1_2_2(nand_30_nl, mux_281_nl, fsm_output[3]);
  assign or_387_nl = (fsm_output[6]) | mux_283_nl;
  assign mux_287_nl = MUX_s_1_2_2(nand_32_nl, or_387_nl, fsm_output[0]);
  assign nor_248_nl = ~((fsm_output[5]) | mux_287_nl);
  assign vec_rsc_0_3_i_wea_d_pff = MUX_s_1_2_2(and_267_nl, nor_248_nl, fsm_output[4]);
  assign or_431_nl = (fsm_output[3]) | (~ (fsm_output[2])) | (fsm_output[1]) | (fsm_output[7])
      | (z_out_6[2:1]!=2'b11) | (fsm_output[9:8]!=2'b10);
  assign or_427_nl = (fsm_output[1]) | (fsm_output[7]) | (z_out_6[2:1]!=2'b11) |
      (fsm_output[9:8]!=2'b10);
  assign mux_312_nl = MUX_s_1_2_2(nand_95_cse, or_427_nl, fsm_output[2]);
  assign or_429_nl = (fsm_output[3]) | mux_312_nl;
  assign and_261_nl = (z_out_6[2:1]==2'b11);
  assign mux_313_nl = MUX_s_1_2_2(or_431_nl, or_429_nl, and_261_nl);
  assign or_424_nl = (~ (VEC_LOOP_j_1_12_0_sva_11_0[0])) | (fsm_output[1]) | (~ (VEC_LOOP_j_1_12_0_sva_11_0[1]))
      | (fsm_output[9:7]!=3'b000);
  assign mux_310_nl = MUX_s_1_2_2(or_424_nl, or_tmp_387, fsm_output[2]);
  assign or_425_nl = (fsm_output[3]) | mux_310_nl;
  assign mux_307_nl = MUX_s_1_2_2(nor_241_cse, nor_269_cse, fsm_output[1]);
  assign nand_38_nl = ~((VEC_LOOP_j_1_12_0_sva_11_0[0]) & mux_307_nl);
  assign mux_308_nl = MUX_s_1_2_2(nand_38_nl, or_tmp_387, fsm_output[2]);
  assign mux_309_nl = MUX_s_1_2_2(mux_308_nl, or_315_cse, fsm_output[3]);
  assign mux_311_nl = MUX_s_1_2_2(or_425_nl, mux_309_nl, and_270_cse);
  assign mux_314_nl = MUX_s_1_2_2(mux_313_nl, mux_311_nl, fsm_output[5]);
  assign nor_240_nl = ~((fsm_output[0]) | mux_314_nl);
  assign nor_243_nl = ~((z_out_6[2:1]!=2'b11) | (~ (fsm_output[1])) | (fsm_output[7])
      | (fsm_output[8]) | (fsm_output[9]));
  assign nor_244_nl = ~((z_out_6[2:1]!=2'b11) | (fsm_output[1]) | (~ (fsm_output[7]))
      | (fsm_output[8]) | (fsm_output[9]));
  assign mux_306_nl = MUX_s_1_2_2(nor_243_nl, nor_244_nl, fsm_output[2]);
  assign and_263_nl = (fsm_output[0]) & (fsm_output[5]) & (fsm_output[3]) & mux_306_nl;
  assign mux_315_nl = MUX_s_1_2_2(nor_240_nl, and_263_nl, fsm_output[4]);
  assign or_416_nl = (z_out_6[2:1]!=2'b11) | (fsm_output[9:7]!=3'b010);
  assign nand_91_nl = ~((z_out_6[2:1]==2'b11) & (fsm_output[9:7]==3'b011));
  assign mux_303_nl = MUX_s_1_2_2(or_416_nl, nand_91_nl, fsm_output[1]);
  assign or_417_nl = (fsm_output[3:2]!=2'b00) | mux_303_nl;
  assign or_409_nl = (fsm_output[2:1]!=2'b01) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b11) | (fsm_output[9:7]!=3'b001);
  assign mux_297_nl = MUX_s_1_2_2(or_409_nl, or_tmp_374, fsm_output[3]);
  assign nand_92_nl = ~((fsm_output[1]) & VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b11) & (fsm_output[9:7]==3'b001));
  assign or_411_nl = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b11)
      | (fsm_output[9:7]!=3'b001);
  assign mux_298_nl = MUX_s_1_2_2(or_304_cse, or_411_nl, fsm_output[1]);
  assign and_265_nl = (COMP_LOOP_acc_1_cse_5_sva[1:0]==2'b11);
  assign mux_299_nl = MUX_s_1_2_2(nand_92_nl, mux_298_nl, and_265_nl);
  assign or_410_nl = (~ (fsm_output[1])) | (COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b11)
      | (fsm_output[9:7]!=3'b010);
  assign mux_300_nl = MUX_s_1_2_2(mux_299_nl, or_410_nl, fsm_output[2]);
  assign mux_301_nl = MUX_s_1_2_2(mux_300_nl, or_tmp_374, fsm_output[3]);
  assign mux_302_nl = MUX_s_1_2_2(mux_297_nl, mux_301_nl, VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm);
  assign mux_304_nl = MUX_s_1_2_2(or_417_nl, mux_302_nl, fsm_output[5]);
  assign and_264_nl = (fsm_output[0]) & (~ mux_304_nl);
  assign nor_245_nl = ~((z_out_6[2:1]!=2'b11) | (fsm_output[9:7]!=3'b000));
  assign nor_246_nl = ~((z_out_6[2:1]!=2'b11) | (fsm_output[9:7]!=3'b001));
  assign mux_296_nl = MUX_s_1_2_2(nor_245_nl, nor_246_nl, fsm_output[1]);
  assign and_266_nl = (~ (fsm_output[0])) & (fsm_output[5]) & (fsm_output[3]) & (fsm_output[2])
      & mux_296_nl;
  assign mux_305_nl = MUX_s_1_2_2(and_264_nl, and_266_nl, fsm_output[4]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_315_nl,
      mux_305_nl, fsm_output[6]);
  assign nor_394_nl = ~((fsm_output[1]) | (~ (fsm_output[5])) | (~ (fsm_output[3]))
      | (~ (fsm_output[2])) | (fsm_output[8]) | (~ (fsm_output[4])));
  assign nor_395_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[3]) |
      (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[4]));
  assign mux_824_nl = MUX_s_1_2_2(nor_394_nl, nor_395_nl, fsm_output[6]);
  assign and_dcpl_196 = mux_824_nl & (~ (fsm_output[9])) & (fsm_output[7]) & (fsm_output[0]);
  assign or_tmp_841 = (~ (fsm_output[3])) | (fsm_output[2]) | (~ (fsm_output[8]));
  assign mux_tmp_824 = MUX_s_1_2_2(or_614_cse, or_tmp_841, fsm_output[1]);
  assign mux_826_cse = MUX_s_1_2_2(or_tmp_841, or_611_cse, fsm_output[1]);
  assign nor_393_nl = ~((fsm_output[7:6]!=2'b10) | mux_tmp_824);
  assign mux_827_nl = MUX_s_1_2_2(mux_826_cse, mux_tmp_824, fsm_output[7]);
  assign and_522_nl = (fsm_output[6]) & (~ mux_827_nl);
  assign mux_828_nl = MUX_s_1_2_2(nor_393_nl, and_522_nl, fsm_output[0]);
  assign and_dcpl_199 = mux_828_nl & (~ (fsm_output[4])) & (fsm_output[5]) & (~ (fsm_output[9]));
  assign and_dcpl_200 = ~((fsm_output[6]) | (fsm_output[0]));
  assign and_dcpl_204 = (~ (fsm_output[3])) & (fsm_output[5]);
  assign and_dcpl_208 = ~((fsm_output[8]) | (fsm_output[4]) | (fsm_output[2]) | (~
      and_dcpl_204) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[7]) | (~ and_dcpl_200));
  assign and_dcpl_215 = (fsm_output[8]) & (~ (fsm_output[4])) & (fsm_output[2]) &
      and_dcpl_204 & (~ (fsm_output[9])) & (fsm_output[1]) & (~ (fsm_output[7]))
      & and_dcpl_200;
  assign and_dcpl_221 = mux_680_cse & (~ (fsm_output[4])) & (~ (fsm_output[2])) &
      (fsm_output[5]) & (~ (fsm_output[9])) & (~ (fsm_output[7])) & and_dcpl_200;
  assign and_dcpl_230 = ~((fsm_output[2]) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[8])
      | (~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[1]) | (fsm_output[7])
      | (~ and_dcpl_200));
  assign and_365_cse = (fsm_output[2]) & (~ (fsm_output[4])) & (~ (fsm_output[3]))
      & (fsm_output[8]) & (fsm_output[5]) & (~ (fsm_output[9])) & (fsm_output[1])
      & (~ (fsm_output[7])) & and_dcpl_200;
  assign or_999_nl = (~ (fsm_output[1])) | (~ (fsm_output[5])) | (fsm_output[8])
      | (~((fsm_output[4:3]==2'b11)));
  assign or_1000_nl = (fsm_output[1]) | (fsm_output[5]) | (~ (fsm_output[8])) | (fsm_output[3])
      | (fsm_output[4]);
  assign mux_830_nl = MUX_s_1_2_2(or_999_nl, or_1000_nl, fsm_output[6]);
  assign and_dcpl_242 = ~(mux_830_nl | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[7])
      | (~ (fsm_output[0])));
  assign or_997_nl = (~ (fsm_output[7])) | (~ (fsm_output[1])) | (fsm_output[5])
      | (~ (fsm_output[8])) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[2]);
  assign or_998_nl = (fsm_output[7]) | (fsm_output[1]) | (~ (fsm_output[5])) | (fsm_output[8])
      | (~((fsm_output[4:2]==3'b111)));
  assign mux_831_nl = MUX_s_1_2_2(or_997_nl, or_998_nl, fsm_output[6]);
  assign and_dcpl_244 = ~(mux_831_nl | (fsm_output[9]) | (fsm_output[0]));
  assign and_dcpl_253 = nor_332_cse & (~ (fsm_output[2])) & (~ (fsm_output[8])) &
      (fsm_output[5]) & (~ (fsm_output[9])) & (~ (fsm_output[1])) & (~ (fsm_output[7]))
      & and_dcpl_200;
  assign nor_382_nl = ~((fsm_output[7]) | (fsm_output[1]) | (~ (fsm_output[9])) |
      (fsm_output[5]) | (fsm_output[3]) | (fsm_output[4]));
  assign nor_383_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[1])) | (fsm_output[9])
      | not_tmp_173);
  assign mux_833_nl = MUX_s_1_2_2(nor_382_nl, nor_383_nl, fsm_output[6]);
  assign and_392_cse = mux_833_nl & (fsm_output[2]) & (~ (fsm_output[8])) & (~ (fsm_output[0]));
  assign or_tmp_858 = (fsm_output[9]) | (fsm_output[8]) | (fsm_output[2]) | (~ (fsm_output[3]))
      | (fsm_output[4]);
  assign or_938_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
      | (~ (fsm_output[3])) | (fsm_output[4]);
  assign mux_tmp_833 = MUX_s_1_2_2(or_tmp_858, or_938_nl, fsm_output[1]);
  assign or_945_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[2]) | (fsm_output[3])
      | (~ (fsm_output[4]));
  assign mux_837_nl = MUX_s_1_2_2(or_945_nl, or_tmp_858, fsm_output[1]);
  assign mux_838_nl = MUX_s_1_2_2(mux_tmp_833, mux_837_nl, fsm_output[7]);
  assign nand_140_nl = ~((fsm_output[6]) & (~ mux_838_nl));
  assign or_942_nl = (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[2]) | (fsm_output[3])
      | (~ (fsm_output[4]));
  assign or_940_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[2]) | (~
      (fsm_output[3])) | (fsm_output[4]);
  assign mux_835_nl = MUX_s_1_2_2(or_942_nl, or_940_nl, fsm_output[1]);
  assign mux_836_nl = MUX_s_1_2_2(mux_835_nl, mux_tmp_833, fsm_output[7]);
  assign or_993_nl = (fsm_output[6]) | mux_836_nl;
  assign mux_839_nl = MUX_s_1_2_2(nand_140_nl, or_993_nl, fsm_output[0]);
  assign and_dcpl_283 = ~(mux_839_nl | (fsm_output[5]));
  assign and_dcpl_288 = ~((fsm_output[8]) | (fsm_output[5]));
  assign and_dcpl_292 = nor_332_cse & (~ (fsm_output[2])) & and_dcpl_288 & (~ (fsm_output[9]))
      & (~ (fsm_output[1])) & (~ (fsm_output[7])) & (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_dcpl_302 = nor_332_cse & (fsm_output[2]) & and_dcpl_288 & (~ (fsm_output[9]))
      & (fsm_output[1]) & (~ (fsm_output[7])) & and_dcpl_200;
  assign and_dcpl_310 = (~ (fsm_output[4])) & (fsm_output[3]) & (fsm_output[2]) &
      (~ (fsm_output[8])) & (fsm_output[5]) & (fsm_output[9]) & (~ (fsm_output[1]))
      & (~ (fsm_output[7])) & and_dcpl_200;
  assign and_dcpl_314 = (fsm_output[9]) & (~ (fsm_output[1])) & (~ (fsm_output[7]))
      & and_dcpl_200;
  assign and_dcpl_315 = (~ (fsm_output[8])) & (fsm_output[5]);
  assign and_dcpl_316 = (fsm_output[2]) & (~ (fsm_output[4]));
  assign and_dcpl_319 = and_dcpl_316 & (fsm_output[3]) & and_dcpl_315 & and_dcpl_314;
  assign not_tmp_415 = MUX_s_1_2_2((fsm_output[6]), (~ (fsm_output[6])), fsm_output[0]);
  assign or_951_nl = (fsm_output[8]) | (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[0]))
      | (fsm_output[6]);
  assign mux_843_nl = MUX_s_1_2_2(mux_165_cse, or_951_nl, fsm_output[1]);
  assign or_950_nl = (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_415;
  assign mux_tmp_843 = MUX_s_1_2_2(mux_843_nl, or_950_nl, fsm_output[5]);
  assign or_959_nl = (fsm_output[9]) | (fsm_output[0]) | (~ (fsm_output[6]));
  assign or_957_nl = (fsm_output[9]) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_tmp_844 = MUX_s_1_2_2(or_959_nl, or_957_nl, fsm_output[7]);
  assign nand_125_nl = ~((fsm_output[1]) & (fsm_output[8]) & (~ mux_tmp_844));
  assign or_956_nl = (~ (fsm_output[1])) | (fsm_output[8]) | (fsm_output[7]) | (fsm_output[9])
      | not_tmp_415;
  assign mux_tmp_845 = MUX_s_1_2_2(nand_125_nl, or_956_nl, fsm_output[5]);
  assign or_965_nl = (fsm_output[8]) | mux_tmp_844;
  assign mux_tmp_849 = MUX_s_1_2_2(or_965_nl, mux_163_cse, fsm_output[1]);
  assign nand_127_nl = ~((fsm_output[8]) & (~ mux_tmp_844));
  assign mux_856_nl = MUX_s_1_2_2(nand_127_nl, mux_165_cse, fsm_output[1]);
  assign mux_857_nl = MUX_s_1_2_2(mux_856_nl, mux_tmp_849, fsm_output[5]);
  assign mux_858_nl = MUX_s_1_2_2(mux_857_nl, mux_tmp_843, fsm_output[4]);
  assign or_966_nl = (fsm_output[1]) | mux_165_cse;
  assign mux_854_nl = MUX_s_1_2_2(mux_tmp_849, or_966_nl, fsm_output[5]);
  assign mux_855_nl = MUX_s_1_2_2(mux_854_nl, mux_tmp_845, fsm_output[4]);
  assign mux_859_nl = MUX_s_1_2_2(mux_858_nl, mux_855_nl, fsm_output[3]);
  assign nand_126_nl = ~((fsm_output[5]) & (fsm_output[1]) & (fsm_output[8]) & (~
      mux_tmp_844));
  assign or_963_nl = (fsm_output[9:7]!=3'b010) | not_tmp_415;
  assign or_961_nl = (fsm_output[9:7]!=3'b011) | not_tmp_415;
  assign mux_848_nl = MUX_s_1_2_2(or_963_nl, or_961_nl, fsm_output[1]);
  assign mux_851_nl = MUX_s_1_2_2(mux_tmp_849, mux_848_nl, fsm_output[5]);
  assign mux_852_nl = MUX_s_1_2_2(nand_126_nl, mux_851_nl, fsm_output[4]);
  assign mux_847_nl = MUX_s_1_2_2(mux_tmp_845, mux_tmp_843, fsm_output[4]);
  assign mux_853_nl = MUX_s_1_2_2(mux_852_nl, mux_847_nl, fsm_output[3]);
  assign mux_860_itm = MUX_s_1_2_2(mux_859_nl, mux_853_nl, fsm_output[2]);
  assign and_dcpl_321 = (~ (fsm_output[9])) & (fsm_output[1]);
  assign and_dcpl_323 = and_dcpl_321 & (~ (fsm_output[7])) & and_dcpl_43;
  assign and_dcpl_325 = and_dcpl_316 & (~ (fsm_output[3]));
  assign and_dcpl_326 = and_dcpl_325 & (~ (fsm_output[8])) & (~ (fsm_output[5]));
  assign and_dcpl_327 = and_dcpl_326 & and_dcpl_323;
  assign and_dcpl_331 = (fsm_output[4:2]==3'b110) & and_dcpl_315 & and_dcpl_323;
  assign and_dcpl_333 = ~((fsm_output[9]) | (fsm_output[1]));
  assign and_dcpl_334 = and_dcpl_333 & (~ (fsm_output[7]));
  assign and_dcpl_338 = (fsm_output[4:2]==3'b111) & and_dcpl_315;
  assign and_dcpl_339 = and_dcpl_338 & and_dcpl_334 & and_dcpl_51;
  assign and_dcpl_342 = and_dcpl_338 & and_dcpl_333 & (fsm_output[7]) & and_dcpl_43;
  assign and_dcpl_343 = and_dcpl_321 & (fsm_output[7]);
  assign and_dcpl_345 = and_dcpl_338 & and_dcpl_343 & and_dcpl_51;
  assign and_dcpl_346 = (fsm_output[6]) & (fsm_output[0]);
  assign and_dcpl_349 = ~((fsm_output[2]) | (fsm_output[4]));
  assign and_dcpl_351 = and_dcpl_349 & (~ (fsm_output[3])) & (fsm_output[8]) & (~
      (fsm_output[5]));
  assign and_dcpl_352 = and_dcpl_351 & and_dcpl_334 & and_dcpl_346;
  assign and_dcpl_354 = and_dcpl_351 & and_dcpl_343 & and_dcpl_200;
  assign and_dcpl_356 = and_dcpl_351 & and_dcpl_343 & and_dcpl_346;
  assign and_dcpl_357 = and_dcpl_326 & and_dcpl_314;
  assign and_dcpl_361 = and_dcpl_325 & (fsm_output[8]) & (fsm_output[5]) & and_dcpl_334
      & and_dcpl_43;
  assign and_dcpl_367 = and_dcpl_349 & (fsm_output[3]) & and_dcpl_315 & (fsm_output[9])
      & (fsm_output[1]) & (~ (fsm_output[7])) & and_dcpl_43;
  assign or_970_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[9]) | (fsm_output[8])
      | not_tmp_173;
  assign or_968_nl = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[9])
      | (fsm_output[8]) | not_tmp_173;
  assign mux_tmp_860 = MUX_s_1_2_2(or_970_nl, or_968_nl, fsm_output[7]);
  assign or_tmp_890 = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[9]) | (~
      (fsm_output[8])) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[5]);
  assign or_973_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[9]) | (~
      (fsm_output[8])) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[5]);
  assign mux_864_nl = MUX_s_1_2_2(or_tmp_890, or_973_nl, fsm_output[7]);
  assign mux_865_nl = MUX_s_1_2_2(mux_tmp_860, mux_864_nl, fsm_output[6]);
  assign or_972_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[5]);
  assign mux_862_nl = MUX_s_1_2_2(or_972_nl, or_tmp_890, fsm_output[7]);
  assign mux_863_nl = MUX_s_1_2_2(mux_862_nl, mux_tmp_860, fsm_output[6]);
  assign mux_866_itm = MUX_s_1_2_2(mux_865_nl, mux_863_nl, fsm_output[0]);
  assign or_976_nl = (fsm_output[3:1]!=3'b010);
  assign or_975_nl = (fsm_output[3:1]!=3'b101);
  assign mux_tmp_866 = MUX_s_1_2_2(or_976_nl, or_975_nl, fsm_output[8]);
  assign STAGE_LOOP_or_ssc = and_dcpl_339 | and_dcpl_345 | and_dcpl_354 | and_dcpl_357;
  assign or_tmp_911 = (~((fsm_output[5:4]!=2'b10))) | (fsm_output[9]);
  assign or_1007_nl = (~((~ (fsm_output[0])) | (~ (fsm_output[4])) | (fsm_output[5])))
      | (fsm_output[9]);
  assign mux_878_nl = MUX_s_1_2_2(or_tmp_911, or_1007_nl, fsm_output[1]);
  assign or_1005_nl = (~((~(and_524_cse | (fsm_output[4]))) | (fsm_output[5]))) |
      (fsm_output[9]);
  assign mux_tmp_877 = MUX_s_1_2_2(mux_878_nl, or_1005_nl, fsm_output[2]);
  assign or_tmp_917 = (~((~((fsm_output[1:0]!=2'b00))) | (fsm_output[5:4]!=2'b01)))
      | (fsm_output[9]);
  assign or_tmp_923 = (~((fsm_output[5:4]!=2'b01))) | (fsm_output[9]);
  assign mux_tmp_886 = MUX_s_1_2_2((~ (fsm_output[9])), (fsm_output[9]), fsm_output[5]);
  assign or_tmp_942 = ~((fsm_output[3]) & (fsm_output[2]) & (fsm_output[4]) & (fsm_output[5])
      & (~ (fsm_output[9])));
  assign nand_147_nl = ~((fsm_output[3]) & VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm
      & (fsm_output[2]) & (fsm_output[4]) & (fsm_output[5]) & (~ (fsm_output[9])));
  assign mux_tmp_907 = MUX_s_1_2_2(nand_147_nl, or_tmp_942, fsm_output[1]);
  assign or_1044_nl = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[2])
      | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[9]);
  assign mux_tmp_910 = MUX_s_1_2_2(or_1044_nl, or_462_cse, fsm_output[3]);
  assign or_tmp_948 = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[2]))
      | (fsm_output[4]) | (~ (fsm_output[5])) | (fsm_output[9]);
  assign or_tmp_949 = (fsm_output[4]) | (fsm_output[5]) | (fsm_output[9]);
  assign or_tmp_952 = (~ (fsm_output[2])) | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[9]);
  assign mux_916_nl = MUX_s_1_2_2(or_tmp_423, or_tmp_949, fsm_output[2]);
  assign mux_tmp_915 = MUX_s_1_2_2(or_tmp_952, mux_916_nl, VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign or_tmp_953 = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[5]) | (fsm_output[9]);
  assign mux_tmp_916 = MUX_s_1_2_2(or_tmp_953, mux_tmp_915, fsm_output[3]);
  assign mux_tmp_919 = MUX_s_1_2_2(or_tmp_948, or_tmp_953, fsm_output[3]);
  assign or_1053_nl = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[4]) | (~ (fsm_output[5]))
      | (fsm_output[9]);
  assign mux_tmp_921 = MUX_s_1_2_2(mux_tmp_919, or_1053_nl, fsm_output[1]);
  assign or_tmp_960 = (fsm_output[4]) | (fsm_output[5]) | (~ (fsm_output[9]));
  assign or_tmp_971 = (~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[0]) | (fsm_output[3])
      | (fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]);
  assign operator_64_false_1_or_2_itm = and_dcpl_199 | and_dcpl_221;
  assign COMP_LOOP_or_27_itm = and_dcpl_242 | and_dcpl_244;
  assign STAGE_LOOP_nor_itm = ~(and_dcpl_319 | and_dcpl_331 | and_dcpl_339 | and_dcpl_342
      | and_dcpl_345 | and_dcpl_352 | and_dcpl_354 | and_dcpl_356 | and_dcpl_357
      | and_dcpl_361 | and_dcpl_367);
  assign STAGE_LOOP_nor_53_itm = ~(and_dcpl_319 | and_dcpl_327 | and_dcpl_331 | and_dcpl_339
      | and_dcpl_342 | and_dcpl_345 | and_dcpl_352 | and_dcpl_354 | and_dcpl_356
      | and_dcpl_357 | and_dcpl_361 | and_dcpl_367);
  assign STAGE_LOOP_or_1_itm = and_dcpl_331 | and_dcpl_339 | and_dcpl_342 | and_dcpl_345;
  assign STAGE_LOOP_or_2_itm = and_dcpl_352 | and_dcpl_354 | and_dcpl_356 | and_dcpl_357;
  always @(posedge clk) begin
    if ( ~ not_tmp_77 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_33 & and_dcpl_29) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, (z_out_6[3:0]), STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_77 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_3_obj_ld_cse <= 1'b0;
      VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= 1'b0;
      modExp_exp_1_0_1_sva_1 <= 1'b0;
      modExp_exp_1_1_1_sva <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_3_obj_ld_cse <= and_dcpl_32 & and_256_cse & (~ (fsm_output[6]))
          & (~ (fsm_output[0])) & (~ (fsm_output[4])) & (fsm_output[9]) & (fsm_output[5])
          & (~ (z_out_5[2]));
      VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= (COMP_LOOP_mux1h_15_nl &
          (~((~ mux_tmp_504) & and_dcpl_147))) | ((~ mux_433_itm) & and_dcpl_51 &
          (~ (fsm_output[4])) & and_dcpl_40);
      modExp_exp_1_0_1_sva_1 <= (COMP_LOOP_mux_39_nl & (~(mux_732_nl & (~ (fsm_output[7]))
          & (~ (fsm_output[4])) & and_dcpl_40))) | (mux_752_nl & (fsm_output[7])
          & (~ (fsm_output[4])) & and_dcpl_40);
      modExp_exp_1_1_1_sva <= COMP_LOOP_mux1h_27_nl & (~(not_tmp_324 & and_dcpl_105
          & and_dcpl_176));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_44_nl & mux_806_nl;
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_4_2(z_out_7, operator_64_false_acc_mut_63_0,
        VEC_LOOP_1_COMP_LOOP_1_acc_8_itm, (z_out_5[63:0]), {modulo_result_or_nl ,
        mux_372_nl , (~ mux_415_nl) , and_dcpl_108});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_5, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_117);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_117);
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_436_nl, and_tmp_7, fsm_output[5]) ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_908_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_944_nl ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_1_12_0_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_123 | VEC_LOOP_j_1_12_0_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_1_12_0_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out_6[11:0]),
          VEC_LOOP_j_1_12_0_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_2_1_sva_6_0 <= 7'b0000000;
    end
    else if ( ~ mux_949_nl ) begin
      COMP_LOOP_k_9_2_1_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (z_out_5[6:0]), or_992_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_while_and_3 | modExp_while_and_5 | modExp_result_sva_mx0c0 | mux_500_nl)
        & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, z_out_6, {modExp_result_sva_mx0c0 , modExp_result_and_rgt
          , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_529_nl ) begin
      modExp_base_1_sva <= MUX1HOT_v_64_4_2(r_sva, modulo_result_rem_cmp_z, z_out_6,
          modExp_result_sva, {and_144_nl , r_or_nl , r_or_1_nl , and_dcpl_138});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_10_lpi_4_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( MUX_s_1_2_2(mux_557_nl, or_1002_nl, fsm_output[9]) ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_5_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
          {and_dcpl_123 , COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl , COMP_LOOP_or_8_nl
          , COMP_LOOP_or_9_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva <= 1'b0;
    end
    else if ( and_dcpl_104 | and_dcpl_107 | and_dcpl_129 ) begin
      exit_VEC_LOOP_1_COMP_LOOP_1_modExp_1_while_sva <= MUX1HOT_s_1_3_2((~ (z_out_6[63])),
          (~ (z_out_1[8])), (~ (readslicef_10_1_9(VEC_LOOP_1_COMP_LOOP_1_acc_11_nl))),
          {and_dcpl_104 , and_dcpl_107 , and_dcpl_129});
    end
  end
  always @(posedge clk) begin
    if ( (mux_682_nl & and_dcpl_109) | and_dcpl_108 ) begin
      VEC_LOOP_1_COMP_LOOP_1_acc_8_itm <= MUX_v_64_2_2(z_out_7, VEC_LOOP_1_COMP_LOOP_1_acc_8_nl,
          and_dcpl_108);
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_or_1_cse ) begin
      COMP_LOOP_acc_psp_1_sva <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_5_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_709_nl, or_tmp_71, fsm_output[6]) ) begin
      COMP_LOOP_acc_1_cse_5_sva <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_1_sva <= 11'b00000000000;
    end
    else if ( mux_721_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_11_psp_1_sva <= nl_COMP_LOOP_acc_11_psp_1_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( mux_731_nl | (fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_2_1_sva <= 1'b0;
      modExp_exp_1_3_1_sva <= 1'b0;
      modExp_exp_1_4_1_sva <= 1'b0;
      modExp_exp_1_5_1_sva <= 1'b0;
      modExp_exp_1_6_1_sva <= 1'b0;
    end
    else if ( mux_801_itm ) begin
      modExp_exp_1_2_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_1_sva_6_0[0]), modExp_exp_1_3_1_sva,
          (COMP_LOOP_k_9_2_1_sva_6_0[1]), {and_dcpl_175 , not_tmp_321 , and_dcpl_179});
      modExp_exp_1_3_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_1_sva_6_0[1]), modExp_exp_1_4_1_sva,
          (COMP_LOOP_k_9_2_1_sva_6_0[2]), {and_dcpl_175 , not_tmp_321 , and_dcpl_179});
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_1_sva_6_0[2]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_2_1_sva_6_0[3]), {and_dcpl_175 , not_tmp_321 , and_dcpl_179});
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_1_sva_6_0[3]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_2_1_sva_6_0[4]), {and_dcpl_175 , not_tmp_321 , and_dcpl_179});
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_2_1_sva_6_0[4]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_2_1_sva_6_0[5]), {and_dcpl_175 , not_tmp_321 , and_dcpl_179});
    end
  end
  always @(posedge clk) begin
    if ( (not_tmp_324 & and_dcpl_105 & (fsm_output[0]) & (~ (fsm_output[9]))) | and_dcpl_111
        | (mux_807_nl & and_dcpl_176) ) begin
      VEC_LOOP_1_COMP_LOOP_2_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out_2[9]),
          (z_out_1[8]), and_dcpl_111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_3_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_6[12:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_VEC_LOOP_1_acc_1_psp_ftd_1 <= 12'b000000000000;
    end
    else if ( ~((fsm_output[7]) | (fsm_output[1]) | (~ (fsm_output[8])) | (~ (fsm_output[2]))
        | (fsm_output[3]) | (fsm_output[6]) | (~ (fsm_output[0])) | (fsm_output[4])
        | or_55_cse) ) begin
      reg_VEC_LOOP_1_acc_1_psp_ftd_1 <= z_out_6[11:0];
    end
  end
  assign modulo_result_or_nl = and_dcpl_104 | and_dcpl_107 | (~ mux_423_itm) | and_dcpl_111;
  assign or_452_nl = nor_236_cse | (fsm_output[4]);
  assign mux_366_nl = MUX_s_1_2_2(mux_tmp_345, or_452_nl, fsm_output[5]);
  assign mux_364_nl = MUX_s_1_2_2(or_tmp_404, or_tmp_416, fsm_output[2]);
  assign mux_365_nl = MUX_s_1_2_2(and_303_cse, mux_364_nl, fsm_output[5]);
  assign mux_367_nl = MUX_s_1_2_2(mux_366_nl, mux_365_nl, fsm_output[8]);
  assign mux_361_nl = MUX_s_1_2_2(or_tmp_416, (~ mux_tmp_318), fsm_output[2]);
  assign mux_362_nl = MUX_s_1_2_2(mux_tmp_345, mux_361_nl, fsm_output[5]);
  assign mux_363_nl = MUX_s_1_2_2(mux_362_nl, mux_tmp_350, fsm_output[8]);
  assign mux_368_nl = MUX_s_1_2_2(mux_367_nl, mux_363_nl, fsm_output[1]);
  assign mux_369_nl = MUX_s_1_2_2((~ mux_368_nl), mux_tmp_338, fsm_output[6]);
  assign mux_357_nl = MUX_s_1_2_2((~ mux_tmp_319), and_303_cse, fsm_output[5]);
  assign mux_358_nl = MUX_s_1_2_2(mux_tmp_340, mux_357_nl, fsm_output[8]);
  assign mux_359_nl = MUX_s_1_2_2(mux_358_nl, mux_tmp_337, fsm_output[1]);
  assign mux_360_nl = MUX_s_1_2_2(mux_tmp_329, mux_359_nl, fsm_output[6]);
  assign mux_370_nl = MUX_s_1_2_2(mux_369_nl, mux_360_nl, fsm_output[7]);
  assign mux_351_nl = MUX_s_1_2_2(or_tmp_416, (~ or_tmp_404), fsm_output[2]);
  assign mux_352_nl = MUX_s_1_2_2(mux_tmp_345, mux_351_nl, fsm_output[5]);
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, mux_tmp_350, fsm_output[8]);
  assign mux_347_nl = MUX_s_1_2_2((fsm_output[4]), (~ (fsm_output[4])), and_256_cse);
  assign mux_348_nl = MUX_s_1_2_2(or_tmp_416, mux_347_nl, fsm_output[5]);
  assign mux_346_nl = MUX_s_1_2_2(mux_tmp_335, mux_tmp_345, fsm_output[5]);
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, mux_346_nl, fsm_output[8]);
  assign mux_354_nl = MUX_s_1_2_2(mux_353_nl, mux_349_nl, fsm_output[1]);
  assign mux_341_nl = MUX_s_1_2_2((~ or_tmp_404), or_756_cse, fsm_output[2]);
  assign mux_342_nl = MUX_s_1_2_2((~ nor_tmp_64), mux_341_nl, fsm_output[5]);
  assign mux_343_nl = MUX_s_1_2_2(mux_342_nl, mux_tmp_340, fsm_output[8]);
  assign mux_344_nl = MUX_s_1_2_2(mux_tmp_325, mux_343_nl, fsm_output[1]);
  assign mux_355_nl = MUX_s_1_2_2((~ mux_354_nl), mux_344_nl, fsm_output[6]);
  assign mux_339_nl = MUX_s_1_2_2(mux_tmp_338, mux_tmp_329, fsm_output[6]);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, mux_339_nl, fsm_output[7]);
  assign mux_371_nl = MUX_s_1_2_2(mux_370_nl, mux_356_nl, fsm_output[0]);
  assign or_446_nl = (fsm_output[8]) | (fsm_output[5]) | (~((fsm_output[4:2]!=3'b001)));
  assign or_443_nl = (fsm_output[8]) | (fsm_output[5]) | nor_tmp_63;
  assign mux_321_nl = MUX_s_1_2_2(or_446_nl, or_443_nl, fsm_output[1]);
  assign nor_237_nl = ~((fsm_output[7:6]!=2'b00) | mux_321_nl);
  assign or_439_nl = (fsm_output[8]) | (fsm_output[5]) | mux_tmp_319;
  assign or_436_nl = (fsm_output[8]) | (fsm_output[5]) | mux_tmp_317;
  assign mux_320_nl = MUX_s_1_2_2(or_439_nl, or_436_nl, fsm_output[1]);
  assign nor_239_nl = ~((fsm_output[7:6]!=2'b00) | mux_320_nl);
  assign mux_322_nl = MUX_s_1_2_2(nor_237_nl, nor_239_nl, fsm_output[0]);
  assign mux_372_nl = MUX_s_1_2_2(mux_371_nl, mux_322_nl, fsm_output[9]);
  assign mux_409_nl = MUX_s_1_2_2(mux_tmp_393, or_1047_cse, fsm_output[2]);
  assign mux_410_nl = MUX_s_1_2_2(mux_409_nl, or_tmp_436, fsm_output[8]);
  assign mux_406_nl = MUX_s_1_2_2(mux_tmp_373, or_tmp_437, fsm_output[9]);
  assign mux_407_nl = MUX_s_1_2_2(or_1047_cse, mux_406_nl, fsm_output[2]);
  assign mux_408_nl = MUX_s_1_2_2(mux_407_nl, or_tmp_436, fsm_output[8]);
  assign mux_411_nl = MUX_s_1_2_2(mux_410_nl, mux_408_nl, fsm_output[1]);
  assign mux_412_nl = MUX_s_1_2_2(mux_tmp_398, mux_411_nl, fsm_output[3]);
  assign mux_413_nl = MUX_s_1_2_2(mux_412_nl, mux_tmp_382, fsm_output[6]);
  assign or_477_nl = nor_70_cse | (fsm_output[9]) | (~ (fsm_output[5]));
  assign mux_403_nl = MUX_s_1_2_2(or_477_nl, mux_tmp_380, fsm_output[1]);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_nl, or_tmp_421, fsm_output[3]);
  assign mux_405_nl = MUX_s_1_2_2(mux_tmp_378, mux_404_nl, fsm_output[6]);
  assign mux_414_nl = MUX_s_1_2_2(mux_413_nl, mux_405_nl, fsm_output[7]);
  assign or_474_nl = (~ (fsm_output[2])) | (fsm_output[9]) | (~ (fsm_output[4]));
  assign mux_394_nl = MUX_s_1_2_2(mux_tmp_393, or_474_nl, fsm_output[8]);
  assign mux_399_nl = MUX_s_1_2_2(mux_tmp_398, mux_394_nl, fsm_output[1]);
  assign mux_391_nl = MUX_s_1_2_2(or_tmp_436, or_tmp_437, nor_70_cse);
  assign mux_388_nl = MUX_s_1_2_2(or_tmp_438, or_tmp_437, fsm_output[9]);
  assign mux_389_nl = MUX_s_1_2_2(or_1047_cse, mux_388_nl, fsm_output[2]);
  assign mux_390_nl = MUX_s_1_2_2(mux_389_nl, or_tmp_436, fsm_output[8]);
  assign mux_392_nl = MUX_s_1_2_2(mux_391_nl, mux_390_nl, fsm_output[1]);
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, mux_392_nl, fsm_output[3]);
  assign mux_386_nl = MUX_s_1_2_2(mux_tmp_375, mux_tmp_379, fsm_output[1]);
  assign or_469_nl = (fsm_output[9]) | mux_tmp_373;
  assign mux_384_nl = MUX_s_1_2_2(or_469_nl, or_1047_cse, nor_70_cse);
  assign mux_385_nl = MUX_s_1_2_2(or_tmp_421, mux_384_nl, fsm_output[1]);
  assign mux_387_nl = MUX_s_1_2_2(mux_386_nl, mux_385_nl, fsm_output[3]);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, mux_387_nl, fsm_output[6]);
  assign mux_383_nl = MUX_s_1_2_2(mux_tmp_382, mux_tmp_378, fsm_output[6]);
  assign mux_402_nl = MUX_s_1_2_2(mux_401_nl, mux_383_nl, fsm_output[7]);
  assign mux_415_nl = MUX_s_1_2_2(mux_414_nl, mux_402_nl, fsm_output[0]);
  assign operator_64_false_1_mux_3_nl = MUX_v_7_2_2((~ COMP_LOOP_k_9_2_1_sva_6_0),
      (~ (STAGE_LOOP_lshift_psp_sva[9:3])), and_dcpl_196);
  assign nor_456_nl = ~((fsm_output[2]) | (fsm_output[8]));
  assign and_531_nl = (fsm_output[2]) & (fsm_output[8]);
  assign mux_952_nl = MUX_s_1_2_2(nor_456_nl, and_531_nl, fsm_output[1]);
  assign operator_64_false_1_or_5_nl = (~(mux_952_nl & and_dcpl_109 & (~ (fsm_output[3]))
      & (fsm_output[5]) & (~ (fsm_output[7])) & and_dcpl_200)) | and_dcpl_196;
  assign operator_64_false_1_mux_4_nl = MUX_v_7_2_2(7'b0000001, COMP_LOOP_k_9_2_1_sva_6_0,
      and_dcpl_196);
  assign nl_acc_nl = ({1'b1 , operator_64_false_1_mux_3_nl , operator_64_false_1_or_5_nl})
      + conv_u2u_8_9({operator_64_false_1_mux_4_nl , 1'b1});
  assign acc_nl = nl_acc_nl[8:0];
  assign COMP_LOOP_and_11_nl = (~ and_dcpl_134) & and_dcpl_123;
  assign nor_184_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[3]) |
      (fsm_output[2]) | (~ nor_tmp_40));
  assign nor_185_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | (~ (fsm_output[3]))
      | (~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[1]));
  assign mux_616_nl = MUX_s_1_2_2(nor_184_nl, nor_185_nl, fsm_output[5]);
  assign COMP_LOOP_or_11_nl = (and_dcpl_154 & and_dcpl_41) | (mux_616_nl & (fsm_output[7])
      & (fsm_output[0]) & (~ (fsm_output[9])));
  assign mux_610_nl = MUX_s_1_2_2(or_tmp_637, or_tmp_635, fsm_output[3]);
  assign or_673_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (fsm_output[8]);
  assign mux_608_nl = MUX_s_1_2_2(or_tmp_637, or_673_nl, fsm_output[1]);
  assign mux_609_nl = MUX_s_1_2_2(mux_608_nl, or_tmp_635, fsm_output[3]);
  assign mux_611_nl = MUX_s_1_2_2(mux_610_nl, mux_609_nl, fsm_output[0]);
  assign mux_604_nl = MUX_s_1_2_2((fsm_output[4]), (~ (fsm_output[8])), fsm_output[2]);
  assign mux_605_nl = MUX_s_1_2_2(mux_604_nl, or_tmp_623, fsm_output[1]);
  assign or_671_nl = (~ (fsm_output[2])) | (fsm_output[8]);
  assign mux_603_nl = MUX_s_1_2_2(or_tmp_621, or_671_nl, fsm_output[1]);
  assign mux_606_nl = MUX_s_1_2_2(mux_605_nl, mux_603_nl, fsm_output[3]);
  assign mux_607_nl = MUX_s_1_2_2(mux_606_nl, mux_tmp_599, fsm_output[0]);
  assign mux_612_nl = MUX_s_1_2_2((~ mux_611_nl), mux_607_nl, fsm_output[5]);
  assign mux_600_nl = MUX_s_1_2_2(mux_tmp_594, mux_tmp_589, fsm_output[3]);
  assign mux_601_nl = MUX_s_1_2_2(mux_600_nl, mux_tmp_599, fsm_output[0]);
  assign mux_602_nl = MUX_s_1_2_2(nor_330_cse, mux_601_nl, fsm_output[5]);
  assign mux_613_nl = MUX_s_1_2_2(mux_612_nl, mux_602_nl, fsm_output[6]);
  assign or_665_nl = (fsm_output[1]) | mux_tmp_588;
  assign mux_595_nl = MUX_s_1_2_2(mux_tmp_594, or_665_nl, fsm_output[3]);
  assign mux_596_nl = MUX_s_1_2_2(nor_330_cse, mux_595_nl, fsm_output[5]);
  assign or_71_nl = (~ (fsm_output[8])) | (fsm_output[3]) | (~ (fsm_output[1])) |
      (fsm_output[2]) | (fsm_output[4]);
  assign or_662_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[4]) | (fsm_output[8]);
  assign nand_55_nl = ~((fsm_output[1]) & (~ mux_tmp_588));
  assign mux_591_nl = MUX_s_1_2_2(or_662_nl, nand_55_nl, fsm_output[3]);
  assign or_661_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[8]);
  assign mux_590_nl = MUX_s_1_2_2(or_661_nl, mux_tmp_589, fsm_output[3]);
  assign mux_592_nl = MUX_s_1_2_2(mux_591_nl, mux_590_nl, fsm_output[0]);
  assign mux_593_nl = MUX_s_1_2_2(or_71_nl, mux_592_nl, fsm_output[5]);
  assign mux_597_nl = MUX_s_1_2_2(mux_596_nl, mux_593_nl, fsm_output[6]);
  assign mux_614_nl = MUX_s_1_2_2(mux_613_nl, mux_597_nl, fsm_output[7]);
  assign or_656_nl = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[4]) | (fsm_output[8]);
  assign or_655_nl = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[4])
      | (fsm_output[8]);
  assign mux_587_nl = MUX_s_1_2_2(or_656_nl, or_655_nl, fsm_output[0]);
  assign nor_186_nl = ~((fsm_output[7:5]!=3'b000) | mux_587_nl);
  assign mux_615_nl = MUX_s_1_2_2(mux_614_nl, nor_186_nl, fsm_output[9]);
  assign COMP_LOOP_mux1h_15_nl = MUX1HOT_s_1_5_2((operator_66_true_div_cmp_z[0]),
      (tmp_10_lpi_4_dfm[0]), (readslicef_9_1_8(acc_nl)), modExp_exp_1_0_1_sva_1,
      VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm, {COMP_LOOP_and_11_nl , and_dcpl_134
      , COMP_LOOP_or_11_nl , not_tmp_260 , mux_615_nl});
  assign mux_750_nl = MUX_s_1_2_2(mux_749_cse, mux_748_cse, fsm_output[1]);
  assign or_890_nl = (fsm_output[1]) | (~ (fsm_output[7])) | mux_745_cse;
  assign mux_751_nl = MUX_s_1_2_2(mux_750_nl, or_890_nl, fsm_output[2]);
  assign COMP_LOOP_mux_39_nl = MUX_s_1_2_2(modExp_exp_1_1_1_sva, modExp_exp_1_0_1_sva_1,
      mux_751_nl);
  assign and_212_nl = (fsm_output[6]) & (~ mux_tmp_92);
  assign nor_170_nl = ~((fsm_output[6]) | (fsm_output[3]) | (~ mux_tmp_579));
  assign mux_732_nl = MUX_s_1_2_2(and_212_nl, nor_170_nl, fsm_output[0]);
  assign and_210_nl = (fsm_output[6]) & not_tmp_91;
  assign nor_165_nl = ~((fsm_output[6]) | mux_tmp_92);
  assign mux_752_nl = MUX_s_1_2_2(and_210_nl, nor_165_nl, fsm_output[0]);
  assign mux_776_nl = MUX_s_1_2_2(mux_tmp_763, or_54_cse, fsm_output[8]);
  assign mux_775_nl = MUX_s_1_2_2(or_54_cse, mux_894_cse, fsm_output[8]);
  assign mux_777_nl = MUX_s_1_2_2(mux_776_nl, mux_775_nl, fsm_output[7]);
  assign mux_778_nl = MUX_s_1_2_2(mux_777_nl, mux_tmp_771, fsm_output[6]);
  assign mux_779_nl = MUX_s_1_2_2(mux_778_nl, or_tmp_760, fsm_output[3]);
  assign mux_772_nl = MUX_s_1_2_2(mux_tmp_763, or_54_cse, or_826_cse);
  assign mux_773_nl = MUX_s_1_2_2(mux_772_nl, mux_tmp_771, fsm_output[6]);
  assign mux_774_nl = MUX_s_1_2_2(mux_773_nl, or_tmp_769, fsm_output[3]);
  assign mux_780_nl = MUX_s_1_2_2(mux_779_nl, mux_774_nl, fsm_output[0]);
  assign or_824_nl = (~((~(and_205_cse | (fsm_output[8]))) | (fsm_output[4]))) |
      (fsm_output[9]) | (~ (fsm_output[5]));
  assign or_820_nl = (~(and_205_cse | (fsm_output[8]) | (~ (fsm_output[4])))) | (fsm_output[9])
      | (~ (fsm_output[5]));
  assign mux_768_nl = MUX_s_1_2_2(or_824_nl, or_820_nl, fsm_output[3]);
  assign mux_769_nl = MUX_s_1_2_2(mux_768_nl, mux_tmp_760, fsm_output[0]);
  assign mux_781_nl = MUX_s_1_2_2(mux_780_nl, mux_769_nl, fsm_output[2]);
  assign mux_764_nl = MUX_s_1_2_2(mux_tmp_763, or_54_cse, or_814_cse);
  assign mux_762_nl = MUX_s_1_2_2(or_tmp_762, or_tmp_769, fsm_output[6]);
  assign mux_765_nl = MUX_s_1_2_2(mux_764_nl, mux_762_nl, fsm_output[3]);
  assign or_810_nl = (~((~((fsm_output[8:7]!=2'b00))) | (fsm_output[4]))) | (fsm_output[9])
      | (~ (fsm_output[5]));
  assign mux_761_nl = MUX_s_1_2_2(or_810_nl, or_tmp_762, fsm_output[3]);
  assign mux_766_nl = MUX_s_1_2_2(mux_765_nl, mux_761_nl, fsm_output[0]);
  assign mux_767_nl = MUX_s_1_2_2(mux_766_nl, mux_tmp_760, fsm_output[2]);
  assign mux_782_nl = MUX_s_1_2_2(mux_781_nl, mux_767_nl, fsm_output[1]);
  assign COMP_LOOP_mux1h_27_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_2_1_sva_6_0[6]),
      modExp_exp_1_2_1_sva, modExp_exp_1_1_1_sva, (COMP_LOOP_k_9_2_1_sva_6_0[0]),
      {and_dcpl_175 , not_tmp_321 , (~ mux_782_nl) , and_dcpl_179});
  assign COMP_LOOP_mux1h_44_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_2_1_sva_6_0[5]),
      modExp_exp_1_1_1_sva, modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_2_1_sva_6_0[6]),
      {and_dcpl_175 , and_dcpl_107 , (~ mux_801_itm) , and_dcpl_179});
  assign or_nl = (~ (fsm_output[0])) | (fsm_output[6]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[8])) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[5]);
  assign or_989_nl = (fsm_output[9:6]!=4'b0010) | not_tmp_173;
  assign or_990_nl = (fsm_output[9:6]!=4'b0011) | not_tmp_173;
  assign mux_804_nl = MUX_s_1_2_2(or_989_nl, or_990_nl, fsm_output[0]);
  assign mux_805_nl = MUX_s_1_2_2(or_nl, mux_804_nl, fsm_output[2]);
  assign or_852_nl = (fsm_output[9:3]!=7'b0111000);
  assign or_851_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[8]) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[5]);
  assign or_850_nl = (fsm_output[9:7]!=3'b000) | not_tmp_173;
  assign mux_802_nl = MUX_s_1_2_2(or_851_nl, or_850_nl, fsm_output[6]);
  assign mux_803_nl = MUX_s_1_2_2(or_852_nl, mux_802_nl, fsm_output[0]);
  assign or_991_nl = (fsm_output[2]) | mux_803_nl;
  assign mux_806_nl = MUX_s_1_2_2(mux_805_nl, or_991_nl, fsm_output[1]);
  assign nor_228_nl = ~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2])
      | (fsm_output[8]) | (fsm_output[1]) | (fsm_output[7]));
  assign mux_436_nl = MUX_s_1_2_2(nor_228_nl, or_814_cse, fsm_output[9]);
  assign mux_901_nl = MUX_s_1_2_2(or_1038_cse, (fsm_output[9]), fsm_output[4]);
  assign mux_902_nl = MUX_s_1_2_2(mux_901_nl, nor_tmp_34, fsm_output[0]);
  assign mux_903_nl = MUX_s_1_2_2(mux_902_nl, mux_tmp_886, fsm_output[1]);
  assign or_1037_nl = (~ (fsm_output[1])) | (fsm_output[4]);
  assign mux_900_nl = MUX_s_1_2_2(nor_tmp_34, mux_tmp_886, or_1037_nl);
  assign mux_904_nl = MUX_s_1_2_2(mux_903_nl, mux_900_nl, fsm_output[2]);
  assign or_1036_nl = (~(and_524_cse | (fsm_output[5:4]!=2'b10))) | (fsm_output[9]);
  assign mux_899_nl = MUX_s_1_2_2(or_1036_nl, or_tmp_923, fsm_output[2]);
  assign mux_905_nl = MUX_s_1_2_2(mux_904_nl, mux_899_nl, fsm_output[7]);
  assign mux_897_nl = MUX_s_1_2_2(or_tmp_911, or_tmp_917, fsm_output[2]);
  assign mux_898_nl = MUX_s_1_2_2(mux_tmp_877, mux_897_nl, fsm_output[7]);
  assign mux_906_nl = MUX_s_1_2_2(mux_905_nl, mux_898_nl, fsm_output[6]);
  assign mux_895_nl = MUX_s_1_2_2(mux_894_cse, or_tmp_923, fsm_output[0]);
  assign nor_429_nl = ~((fsm_output[6]) | (fsm_output[7]) | (~ (fsm_output[2])) |
      (~ (fsm_output[1])));
  assign mux_896_nl = MUX_s_1_2_2(or_tmp_911, mux_895_nl, nor_429_nl);
  assign mux_907_nl = MUX_s_1_2_2(mux_906_nl, mux_896_nl, fsm_output[8]);
  assign mux_889_nl = MUX_s_1_2_2(nor_tmp_34, mux_tmp_886, fsm_output[4]);
  assign mux_886_nl = MUX_s_1_2_2(nor_tmp_34, or_55_cse, fsm_output[4]);
  assign and_525_nl = ((fsm_output[5:4]!=2'b00)) & (fsm_output[9]);
  assign mux_887_nl = MUX_s_1_2_2(mux_886_nl, and_525_nl, and_524_cse);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, mux_887_nl, fsm_output[2]);
  assign or_1032_nl = (~((~((~((fsm_output[2:0]!=3'b000))) | (fsm_output[4]))) |
      (fsm_output[5]))) | (fsm_output[9]);
  assign mux_891_nl = MUX_s_1_2_2(mux_890_nl, or_1032_nl, fsm_output[7]);
  assign or_1028_nl = (~((~((~((~ (fsm_output[7])) | (fsm_output[2]) | (fsm_output[1])
      | (~ (fsm_output[0])))) | (fsm_output[4]))) | (fsm_output[5]))) | (fsm_output[9]);
  assign mux_892_nl = MUX_s_1_2_2(mux_891_nl, or_1028_nl, fsm_output[6]);
  assign or_1025_nl = (~((~((~((fsm_output[2:0]!=3'b010))) | (fsm_output[4]))) |
      (fsm_output[5]))) | (fsm_output[9]);
  assign or_1021_nl = (~((fsm_output[0]) | (fsm_output[4]) | (~ (fsm_output[5]))))
      | (fsm_output[9]);
  assign mux_882_nl = MUX_s_1_2_2(or_1021_nl, or_tmp_923, fsm_output[1]);
  assign or_1018_nl = (~((~((~((fsm_output[1:0]!=2'b10))) | (fsm_output[4]))) | (fsm_output[5])))
      | (fsm_output[9]);
  assign mux_883_nl = MUX_s_1_2_2(mux_882_nl, or_1018_nl, fsm_output[2]);
  assign mux_884_nl = MUX_s_1_2_2(or_1025_nl, mux_883_nl, fsm_output[7]);
  assign or_1011_nl = (~((~((~((fsm_output[1:0]!=2'b01))) | (fsm_output[4]))) | (fsm_output[5])))
      | (fsm_output[9]);
  assign mux_880_nl = MUX_s_1_2_2(or_tmp_917, or_1011_nl, fsm_output[2]);
  assign mux_881_nl = MUX_s_1_2_2(mux_880_nl, mux_tmp_877, fsm_output[7]);
  assign mux_885_nl = MUX_s_1_2_2(mux_884_nl, mux_881_nl, fsm_output[6]);
  assign mux_893_nl = MUX_s_1_2_2(mux_892_nl, mux_885_nl, fsm_output[8]);
  assign mux_908_nl = MUX_s_1_2_2(mux_907_nl, mux_893_nl, fsm_output[3]);
  assign mux_939_nl = MUX_s_1_2_2(mux_tmp_915, or_tmp_948, fsm_output[3]);
  assign mux_940_nl = MUX_s_1_2_2(or_tmp_942, mux_939_nl, fsm_output[1]);
  assign mux_941_nl = MUX_s_1_2_2(mux_940_nl, mux_tmp_907, fsm_output[7]);
  assign nand_nl = ~(VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & (fsm_output[2])
      & (fsm_output[4]) & (fsm_output[5]) & (~ (fsm_output[9])));
  assign or_1061_nl = (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (fsm_output[2])
      | (fsm_output[4]) | (~ (fsm_output[5])) | (fsm_output[9]);
  assign mux_938_nl = MUX_s_1_2_2(nand_nl, or_1061_nl, fsm_output[3]);
  assign or_1063_nl = (fsm_output[7]) | (fsm_output[1]) | mux_938_nl;
  assign mux_942_nl = MUX_s_1_2_2(mux_941_nl, or_1063_nl, fsm_output[8]);
  assign mux_933_nl = MUX_s_1_2_2((fsm_output[9]), or_1038_cse, fsm_output[4]);
  assign mux_934_nl = MUX_s_1_2_2(mux_933_nl, or_tmp_960, fsm_output[2]);
  assign or_1059_nl = (fsm_output[3]) | mux_934_nl;
  assign mux_930_nl = MUX_s_1_2_2(or_tmp_960, or_tmp_949, fsm_output[2]);
  assign mux_931_nl = MUX_s_1_2_2(or_tmp_952, mux_930_nl, VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign or_1055_nl = (~ (fsm_output[2])) | (~ (fsm_output[4])) | (fsm_output[5])
      | (fsm_output[9]);
  assign mux_932_nl = MUX_s_1_2_2(mux_931_nl, or_1055_nl, fsm_output[3]);
  assign mux_935_nl = MUX_s_1_2_2(or_1059_nl, mux_932_nl, fsm_output[1]);
  assign mux_936_nl = MUX_s_1_2_2(mux_935_nl, mux_tmp_921, fsm_output[7]);
  assign or_1054_nl = (~ (fsm_output[2])) | (fsm_output[4]) | (~ (fsm_output[5]))
      | (fsm_output[9]);
  assign mux_928_nl = MUX_s_1_2_2(or_1054_nl, or_tmp_953, fsm_output[3]);
  assign nand_145_nl = ~((fsm_output[1]) & (~ mux_928_nl));
  assign mux_927_nl = MUX_s_1_2_2(mux_tmp_910, mux_tmp_916, fsm_output[1]);
  assign mux_929_nl = MUX_s_1_2_2(nand_145_nl, mux_927_nl, fsm_output[7]);
  assign mux_937_nl = MUX_s_1_2_2(mux_936_nl, mux_929_nl, fsm_output[8]);
  assign mux_943_nl = MUX_s_1_2_2(mux_942_nl, mux_937_nl, fsm_output[0]);
  assign or_1052_nl = (fsm_output[3]) | (~ (fsm_output[2])) | (fsm_output[4]) | (~
      (fsm_output[5])) | (fsm_output[9]);
  assign mux_922_nl = MUX_s_1_2_2(or_1052_nl, mux_tmp_919, fsm_output[1]);
  assign mux_924_nl = MUX_s_1_2_2(mux_tmp_921, mux_922_nl, fsm_output[7]);
  assign or_1051_nl = (~ (fsm_output[3])) | (fsm_output[2]) | (fsm_output[4]) | (~
      (fsm_output[5])) | (fsm_output[9]);
  assign mux_919_nl = MUX_s_1_2_2(or_1051_nl, mux_tmp_916, fsm_output[1]);
  assign mux_913_nl = MUX_s_1_2_2(or_1047_cse, or_tmp_949, fsm_output[2]);
  assign mux_914_nl = MUX_s_1_2_2(mux_913_nl, or_tmp_948, fsm_output[3]);
  assign mux_915_nl = MUX_s_1_2_2(mux_914_nl, mux_tmp_910, fsm_output[1]);
  assign mux_920_nl = MUX_s_1_2_2(mux_919_nl, mux_915_nl, fsm_output[7]);
  assign mux_925_nl = MUX_s_1_2_2(mux_924_nl, mux_920_nl, fsm_output[8]);
  assign or_1041_nl = (~ (fsm_output[3])) | (~ VEC_LOOP_1_COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm)
      | (fsm_output[2]) | (~ (fsm_output[4])) | (~ (fsm_output[5])) | (fsm_output[9]);
  assign mux_910_nl = MUX_s_1_2_2(or_tmp_942, or_1041_nl, fsm_output[1]);
  assign mux_911_nl = MUX_s_1_2_2(mux_910_nl, mux_tmp_907, fsm_output[7]);
  assign or_1042_nl = (fsm_output[8]) | mux_911_nl;
  assign mux_926_nl = MUX_s_1_2_2(mux_925_nl, or_1042_nl, fsm_output[0]);
  assign mux_944_nl = MUX_s_1_2_2(mux_943_nl, mux_926_nl, fsm_output[6]);
  assign nand_117_nl = ~((fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[4]))
      & (fsm_output[0]) & (fsm_output[3]) & (fsm_output[1]) & (~ (fsm_output[8])));
  assign or_548_nl = (fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[1])) | (fsm_output[8]);
  assign nand_85_nl = ~((fsm_output[0]) & (fsm_output[3]) & (fsm_output[1]) & (~
      (fsm_output[8])));
  assign mux_476_nl = MUX_s_1_2_2(or_548_nl, nand_85_nl, fsm_output[4]);
  assign or_546_nl = (fsm_output[4]) | (~ (fsm_output[0])) | (fsm_output[3]) | (fsm_output[1])
      | (~ (fsm_output[8]));
  assign mux_477_nl = MUX_s_1_2_2(mux_476_nl, or_546_nl, fsm_output[5]);
  assign or_912_nl = (fsm_output[9]) | mux_477_nl;
  assign mux_478_nl = MUX_s_1_2_2(nand_117_nl, or_912_nl, fsm_output[2]);
  assign or_992_nl = mux_478_nl | (fsm_output[7:6]!=2'b00);
  assign or_1069_nl = (~ (fsm_output[2])) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[7]) | (fsm_output[6]);
  assign mux_947_nl = MUX_s_1_2_2(or_1069_nl, or_tmp_971, fsm_output[9]);
  assign or_1067_nl = (fsm_output[2]) | (~ (fsm_output[5])) | (~ (fsm_output[0]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[7]) | (fsm_output[6]);
  assign mux_946_nl = MUX_s_1_2_2(or_tmp_971, or_1067_nl, fsm_output[9]);
  assign mux_948_nl = MUX_s_1_2_2(mux_947_nl, mux_946_nl, fsm_output[1]);
  assign nor_434_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[8])
      | (fsm_output[7]) | (fsm_output[6]));
  assign nor_435_nl = ~((fsm_output[0]) | (~ (fsm_output[3])) | (fsm_output[8]) |
      (~((fsm_output[7:6]==2'b11))));
  assign mux_945_nl = MUX_s_1_2_2(nor_434_nl, nor_435_nl, fsm_output[5]);
  assign nand_143_nl = ~((~((~ (fsm_output[1])) | (fsm_output[9]) | (~ (fsm_output[2]))))
      & mux_945_nl);
  assign mux_949_nl = MUX_s_1_2_2(mux_948_nl, nand_143_nl, fsm_output[4]);
  assign or_563_nl = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]);
  assign or_562_nl = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]);
  assign mux_499_nl = MUX_s_1_2_2(or_563_nl, or_562_nl, and_524_cse);
  assign or_897_nl = (fsm_output[5]) | (fsm_output[3]) | mux_499_nl;
  assign nor_216_nl = ~(and_256_cse | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7])
      | (fsm_output[8]));
  assign mux_498_nl = MUX_s_1_2_2(nor_312_cse, nor_216_nl, fsm_output[5]);
  assign mux_500_nl = MUX_s_1_2_2(or_897_nl, mux_498_nl, fsm_output[9]);
  assign and_144_nl = and_dcpl_103 & and_dcpl_29;
  assign r_or_nl = ((~ (modulo_result_rem_cmp_z[63])) & nor_359_m1c) | (not_tmp_231
      & and_dcpl_40 & (~ (modulo_result_rem_cmp_z[63])));
  assign r_or_1_nl = ((modulo_result_rem_cmp_z[63]) & nor_359_m1c) | (not_tmp_231
      & and_dcpl_40 & (modulo_result_rem_cmp_z[63]));
  assign and_240_nl = (fsm_output[6]) & (~ or_tmp_539);
  assign mux_524_nl = MUX_s_1_2_2(mux_tmp_522, nor_tmp_83, fsm_output[6]);
  assign mux_523_nl = MUX_s_1_2_2((~ or_tmp_539), mux_tmp_522, fsm_output[6]);
  assign mux_525_nl = MUX_s_1_2_2(mux_524_nl, mux_523_nl, fsm_output[0]);
  assign mux_526_nl = MUX_s_1_2_2(and_240_nl, mux_525_nl, fsm_output[7]);
  assign nor_209_nl = ~((fsm_output[5:2]!=4'b1010));
  assign mux_519_nl = MUX_s_1_2_2(nor_209_nl, nor_tmp_81, fsm_output[6]);
  assign and_149_nl = (fsm_output[6]) & mux_tmp_506;
  assign mux_520_nl = MUX_s_1_2_2(mux_519_nl, and_149_nl, fsm_output[0]);
  assign mux_521_nl = MUX_s_1_2_2(mux_520_nl, mux_tmp_509, fsm_output[7]);
  assign mux_527_nl = MUX_s_1_2_2(mux_526_nl, mux_521_nl, fsm_output[8]);
  assign or_581_nl = (fsm_output[5:2]!=4'b1000);
  assign mux_515_nl = MUX_s_1_2_2(or_581_nl, or_tmp_539, fsm_output[6]);
  assign or_579_nl = (fsm_output[5:2]!=4'b0001);
  assign or_577_nl = (fsm_output[3]) | (~ and_213_cse);
  assign mux_513_nl = MUX_s_1_2_2((~ nor_tmp_86), or_577_nl, fsm_output[2]);
  assign mux_514_nl = MUX_s_1_2_2(or_579_nl, mux_513_nl, fsm_output[6]);
  assign mux_516_nl = MUX_s_1_2_2(mux_515_nl, mux_514_nl, fsm_output[0]);
  assign mux_517_nl = MUX_s_1_2_2(mux_516_nl, or_tmp_539, fsm_output[7]);
  assign and_148_nl = (fsm_output[6]) & nor_tmp_83;
  assign mux_510_nl = MUX_s_1_2_2(mux_tmp_506, mux_tmp_509, fsm_output[6]);
  assign mux_507_nl = MUX_s_1_2_2(nor_tmp_83, mux_tmp_506, fsm_output[6]);
  assign mux_511_nl = MUX_s_1_2_2(mux_510_nl, mux_507_nl, fsm_output[0]);
  assign mux_512_nl = MUX_s_1_2_2(and_148_nl, mux_511_nl, fsm_output[7]);
  assign mux_518_nl = MUX_s_1_2_2((~ mux_517_nl), mux_512_nl, fsm_output[8]);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, mux_518_nl, fsm_output[1]);
  assign nor_325_nl = ~((fsm_output[8:2]!=7'b0000000));
  assign mux_529_nl = MUX_s_1_2_2(mux_528_nl, nor_325_nl, fsm_output[9]);
  assign nor_203_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b00) | mux_561_cse);
  assign nor_204_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b00) | mux_560_cse);
  assign mux_562_nl = MUX_s_1_2_2(nor_203_nl, nor_204_nl, fsm_output[1]);
  assign and_235_nl = (fsm_output[6]) & mux_562_nl;
  assign or_607_nl = (fsm_output[7]) | (VEC_LOOP_j_1_12_0_sva_11_0[1:0]!=2'b00) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_606_nl = (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[3]) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b00)
      | (~ (fsm_output[8]));
  assign mux_559_nl = MUX_s_1_2_2(or_607_nl, or_606_nl, fsm_output[1]);
  assign nor_205_nl = ~((fsm_output[6]) | mux_559_nl);
  assign mux_563_nl = MUX_s_1_2_2(and_235_nl, nor_205_nl, fsm_output[0]);
  assign COMP_LOOP_or_6_nl = (mux_563_nl & and_dcpl_110) | ((~((VEC_LOOP_j_1_12_0_sva_11_0[0])
      | (COMP_LOOP_acc_11_psp_1_sva[0]))) & and_160_m1c) | ((~((reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      | (COMP_LOOP_acc_11_psp_1_sva[0]))) & and_163_m1c);
  assign nor_200_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b01) | mux_561_cse);
  assign nor_201_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b01) | mux_560_cse);
  assign mux_567_nl = MUX_s_1_2_2(nor_200_nl, nor_201_nl, fsm_output[1]);
  assign and_234_nl = (fsm_output[6]) & mux_567_nl;
  assign or_618_nl = (fsm_output[7]) | (VEC_LOOP_j_1_12_0_sva_11_0[1:0]!=2'b01) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_617_nl = (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[3]) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]!=2'b01)
      | (~ (fsm_output[8]));
  assign mux_564_nl = MUX_s_1_2_2(or_618_nl, or_617_nl, fsm_output[1]);
  assign nor_202_nl = ~((fsm_output[6]) | mux_564_nl);
  assign mux_568_nl = MUX_s_1_2_2(and_234_nl, nor_202_nl, fsm_output[0]);
  assign COMP_LOOP_or_7_nl = (mux_568_nl & and_dcpl_110) | ((VEC_LOOP_j_1_12_0_sva_11_0[0])
      & (~ (COMP_LOOP_acc_11_psp_1_sva[0])) & and_160_m1c) | ((reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      & (~ (COMP_LOOP_acc_11_psp_1_sva[0])) & and_163_m1c);
  assign nor_197_nl = ~((COMP_LOOP_acc_1_cse_2_sva[1:0]!=2'b10) | mux_561_cse);
  assign nor_198_nl = ~((COMP_LOOP_acc_1_cse_5_sva[1:0]!=2'b10) | mux_560_cse);
  assign mux_572_nl = MUX_s_1_2_2(nor_197_nl, nor_198_nl, fsm_output[1]);
  assign and_233_nl = (fsm_output[6]) & mux_572_nl;
  assign or_629_nl = (fsm_output[7]) | (VEC_LOOP_j_1_12_0_sva_11_0[1:0]!=2'b10) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_628_nl = (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[3]) | (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      | (~((reg_VEC_LOOP_1_acc_1_psp_ftd_1[1]) & (fsm_output[8])));
  assign mux_569_nl = MUX_s_1_2_2(or_629_nl, or_628_nl, fsm_output[1]);
  assign nor_199_nl = ~((fsm_output[6]) | mux_569_nl);
  assign mux_573_nl = MUX_s_1_2_2(and_233_nl, nor_199_nl, fsm_output[0]);
  assign COMP_LOOP_or_8_nl = (mux_573_nl & and_dcpl_110) | ((COMP_LOOP_acc_11_psp_1_sva[0])
      & (~ (VEC_LOOP_j_1_12_0_sva_11_0[0])) & and_160_m1c) | ((COMP_LOOP_acc_11_psp_1_sva[0])
      & (~ (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])) & and_163_m1c);
  assign and_231_nl = (COMP_LOOP_acc_1_cse_2_sva[1:0]==2'b11) & (~ mux_561_cse);
  assign and_232_nl = (COMP_LOOP_acc_1_cse_5_sva[1:0]==2'b11) & (~ mux_560_cse);
  assign mux_577_nl = MUX_s_1_2_2(and_231_nl, and_232_nl, fsm_output[1]);
  assign and_230_nl = (fsm_output[6]) & mux_577_nl;
  assign or_636_nl = (fsm_output[7]) | (VEC_LOOP_j_1_12_0_sva_11_0[1:0]!=2'b11) |
      (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8]);
  assign or_635_nl = (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[3]) | (~((reg_VEC_LOOP_1_acc_1_psp_ftd_1[1:0]==2'b11)
      & (fsm_output[8])));
  assign mux_574_nl = MUX_s_1_2_2(or_636_nl, or_635_nl, fsm_output[1]);
  assign nor_196_nl = ~((fsm_output[6]) | mux_574_nl);
  assign mux_578_nl = MUX_s_1_2_2(and_230_nl, nor_196_nl, fsm_output[0]);
  assign COMP_LOOP_or_9_nl = (mux_578_nl & and_dcpl_110) | ((VEC_LOOP_j_1_12_0_sva_11_0[0])
      & (COMP_LOOP_acc_11_psp_1_sva[0]) & and_160_m1c) | ((reg_VEC_LOOP_1_acc_1_psp_ftd_1[0])
      & (COMP_LOOP_acc_11_psp_1_sva[0]) & and_163_m1c);
  assign mux_551_nl = MUX_s_1_2_2((~ or_756_cse), (fsm_output[4]), fsm_output[7]);
  assign mux_552_nl = MUX_s_1_2_2(mux_551_nl, mux_tmp_546, fsm_output[2]);
  assign mux_553_nl = MUX_s_1_2_2(mux_552_nl, or_tmp_567, fsm_output[8]);
  assign mux_554_nl = MUX_s_1_2_2(mux_553_nl, mux_tmp_549, fsm_output[1]);
  assign mux_545_nl = MUX_s_1_2_2(and_303_cse, or_756_cse, fsm_output[7]);
  assign mux_547_nl = MUX_s_1_2_2(mux_tmp_546, mux_545_nl, fsm_output[2]);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, or_tmp_562, fsm_output[8]);
  assign mux_550_nl = MUX_s_1_2_2(mux_tmp_549, mux_548_nl, fsm_output[1]);
  assign mux_555_nl = MUX_s_1_2_2(mux_554_nl, mux_550_nl, fsm_output[0]);
  assign mux_543_nl = MUX_s_1_2_2(or_tmp_562, (fsm_output[4]), fsm_output[8]);
  assign mux_542_nl = MUX_s_1_2_2(or_756_cse, or_tmp_567, fsm_output[8]);
  assign mux_544_nl = MUX_s_1_2_2(mux_543_nl, mux_542_nl, fsm_output[1]);
  assign mux_556_nl = MUX_s_1_2_2(mux_555_nl, mux_544_nl, fsm_output[6]);
  assign or_603_nl = (~((~ (fsm_output[2])) | (fsm_output[7]))) | (fsm_output[4:3]!=2'b00);
  assign or_601_nl = and_256_cse | (fsm_output[4]);
  assign mux_539_nl = MUX_s_1_2_2(or_603_nl, or_601_nl, fsm_output[8]);
  assign mux_540_nl = MUX_s_1_2_2(mux_539_nl, mux_tmp_537, fsm_output[1]);
  assign or_598_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[4]);
  assign mux_536_nl = MUX_s_1_2_2(or_598_nl, or_756_cse, fsm_output[8]);
  assign mux_538_nl = MUX_s_1_2_2(mux_tmp_537, mux_536_nl, fsm_output[1]);
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, mux_538_nl, or_596_cse);
  assign mux_557_nl = MUX_s_1_2_2(mux_556_nl, (~ mux_541_nl), fsm_output[5]);
  assign or_593_nl = (fsm_output[7]) | and_303_cse;
  assign or_592_nl = (fsm_output[7]) | (fsm_output[4]);
  assign mux_534_nl = MUX_s_1_2_2(or_593_nl, or_592_nl, fsm_output[2]);
  assign or_594_nl = (fsm_output[8]) | mux_534_nl;
  assign or_591_nl = (fsm_output[8]) | (fsm_output[7]) | (fsm_output[4]);
  assign mux_535_nl = MUX_s_1_2_2(or_594_nl, or_591_nl, or_590_cse);
  assign or_1002_nl = (fsm_output[6:5]!=2'b00) | mux_535_nl;
  assign nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl = ({(z_out_5[7:0]) , 2'b00}) + ({1'b1
      , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))}) + 10'b0000000001;
  assign VEC_LOOP_1_COMP_LOOP_1_acc_11_nl = nl_VEC_LOOP_1_COMP_LOOP_1_acc_11_nl[9:0];
  assign nl_VEC_LOOP_1_COMP_LOOP_1_acc_8_nl = tmp_10_lpi_4_dfm - modExp_base_1_sva_mx1;
  assign VEC_LOOP_1_COMP_LOOP_1_acc_8_nl = nl_VEC_LOOP_1_COMP_LOOP_1_acc_8_nl[63:0];
  assign or_721_nl = (fsm_output[0]) | (fsm_output[6]) | (fsm_output[1]) | (fsm_output[8])
      | (~ (fsm_output[3]));
  assign nand_58_nl = ~((fsm_output[0]) & mux_680_cse);
  assign mux_681_nl = MUX_s_1_2_2(or_721_nl, nand_58_nl, fsm_output[5]);
  assign nor_173_nl = ~((fsm_output[2]) | mux_681_nl);
  assign nor_175_nl = ~((fsm_output[6]) | (~((fsm_output[1]) & (fsm_output[8]) &
      (fsm_output[3]))));
  assign and_223_nl = (fsm_output[6]) & (fsm_output[1]) & (fsm_output[8]) & (fsm_output[3]);
  assign mux_678_nl = MUX_s_1_2_2(nor_175_nl, and_223_nl, fsm_output[0]);
  assign and_222_nl = (fsm_output[5]) & mux_678_nl;
  assign nor_176_nl = ~((fsm_output[6]) | (fsm_output[1]) | (fsm_output[8]) | (fsm_output[3]));
  assign nor_177_nl = ~((~ (fsm_output[6])) | (fsm_output[1]) | (fsm_output[8]) |
      (fsm_output[3]));
  assign mux_677_nl = MUX_s_1_2_2(nor_176_nl, nor_177_nl, fsm_output[0]);
  assign and_224_nl = (fsm_output[5]) & mux_677_nl;
  assign mux_679_nl = MUX_s_1_2_2(and_222_nl, and_224_nl, fsm_output[2]);
  assign mux_682_nl = MUX_s_1_2_2(nor_173_nl, mux_679_nl, fsm_output[7]);
  assign mux_87_nl = MUX_s_1_2_2(mux_tmp_86, mux_tmp_84, fsm_output[3]);
  assign mux_85_nl = MUX_s_1_2_2(mux_tmp_84, or_tmp_77, fsm_output[3]);
  assign and_297_nl = or_590_cse & (fsm_output[2]);
  assign mux_88_nl = MUX_s_1_2_2(mux_87_nl, mux_85_nl, and_297_nl);
  assign mux_89_nl = MUX_s_1_2_2(mux_tmp_86, mux_88_nl, fsm_output[4]);
  assign mux_699_nl = MUX_s_1_2_2(or_tmp_77, or_tmp_71, fsm_output[3]);
  assign mux_79_nl = MUX_s_1_2_2(mux_tmp_72, or_tmp_71, fsm_output[3]);
  assign mux_700_nl = MUX_s_1_2_2(mux_699_nl, mux_79_nl, or_94_cse);
  assign or_93_nl = and_300_cse | (fsm_output[3]);
  assign mux_78_nl = MUX_s_1_2_2(mux_tmp_72, or_tmp_71, or_93_nl);
  assign mux_701_nl = MUX_s_1_2_2(mux_700_nl, mux_78_nl, fsm_output[0]);
  assign mux_702_nl = MUX_s_1_2_2(mux_701_nl, or_tmp_71, fsm_output[4]);
  assign mux_709_nl = MUX_s_1_2_2(mux_89_nl, mux_702_nl, fsm_output[5]);
  assign COMP_LOOP_mux_42_nl = MUX_v_11_2_2((VEC_LOOP_j_1_12_0_sva_11_0[11:1]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:1]),
      and_365_cse);
  assign nl_COMP_LOOP_acc_11_psp_1_sva  = COMP_LOOP_mux_42_nl + conv_u2u_8_11({COMP_LOOP_k_9_2_1_sva_6_0
      , 1'b1});
  assign mux_717_nl = MUX_s_1_2_2(or_154_cse, (~ mux_tmp_711), and_300_cse);
  assign mux_718_nl = MUX_s_1_2_2(mux_717_nl, or_154_cse, fsm_output[8]);
  assign or_758_nl = (~ (fsm_output[8])) | (fsm_output[2]);
  assign mux_716_nl = MUX_s_1_2_2((~ or_154_cse), mux_tmp_711, or_758_nl);
  assign mux_719_nl = MUX_s_1_2_2((~ mux_718_nl), mux_716_nl, fsm_output[3]);
  assign mux_720_nl = MUX_s_1_2_2((~ or_154_cse), mux_719_nl, fsm_output[4]);
  assign or_757_nl = (fsm_output[2:0]!=3'b000);
  assign mux_713_nl = MUX_s_1_2_2(mux_tmp_711, and_205_cse, or_757_nl);
  assign and_217_nl = (fsm_output[2:0]==3'b111);
  assign mux_712_nl = MUX_s_1_2_2(mux_tmp_711, and_205_cse, and_217_nl);
  assign mux_714_nl = MUX_s_1_2_2(mux_713_nl, mux_712_nl, fsm_output[8]);
  assign mux_715_nl = MUX_s_1_2_2(mux_714_nl, and_205_cse, or_756_cse);
  assign mux_721_nl = MUX_s_1_2_2(mux_720_nl, mux_715_nl, fsm_output[5]);
  assign or_763_nl = and_213_cse | (fsm_output[7]);
  assign or_762_nl = (fsm_output[5]) | (fsm_output[7]);
  assign or_761_nl = (fsm_output[3:0]!=4'b0000);
  assign mux_730_nl = MUX_s_1_2_2(or_763_nl, or_762_nl, or_761_nl);
  assign nor_171_nl = ~((fsm_output[6]) | mux_730_nl);
  assign mux_726_nl = MUX_s_1_2_2(mux_tmp_723, mux_tmp_722, and_524_cse);
  assign mux_727_nl = MUX_s_1_2_2(and_tmp_14, mux_726_nl, fsm_output[3]);
  assign mux_724_nl = MUX_s_1_2_2(and_tmp_14, mux_tmp_723, and_524_cse);
  assign mux_725_nl = MUX_s_1_2_2(mux_724_nl, mux_tmp_722, fsm_output[3]);
  assign mux_728_nl = MUX_s_1_2_2(mux_727_nl, mux_725_nl, fsm_output[2]);
  assign mux_729_nl = MUX_s_1_2_2(mux_728_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_731_nl = MUX_s_1_2_2(nor_171_nl, mux_729_nl, fsm_output[8]);
  assign nor_142_nl = ~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[2])
      | (~ and_dcpl_86));
  assign nor_143_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[6])) | (~ (fsm_output[3]))
      | (~ (fsm_output[2])) | (fsm_output[8]) | (fsm_output[1]) | (fsm_output[7]));
  assign mux_807_nl = MUX_s_1_2_2(nor_142_nl, nor_143_nl, fsm_output[5]);
  assign operator_64_false_1_mux_5_nl = MUX_v_2_2_2((VEC_LOOP_j_1_12_0_sva_11_0[11:10]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]), and_dcpl_215);
  assign operator_64_false_1_operator_64_false_1_or_1_nl = MUX_v_2_2_2(operator_64_false_1_mux_5_nl,
      2'b11, operator_64_false_1_or_2_itm);
  assign operator_64_false_1_mux1h_9_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_7_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[9]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9]), (~ modExp_exp_1_1_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_10_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_6_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[8]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[8]), (~ modExp_exp_1_7_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_11_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_5_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[7]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[7]), (~ modExp_exp_1_6_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_12_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_4_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[6]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[6]), (~ modExp_exp_1_5_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_13_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_3_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[5]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[5]), (~ modExp_exp_1_4_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_14_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_2_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[4]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[4]), (~ modExp_exp_1_3_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_15_nl = MUX1HOT_s_1_4_2((~ modExp_exp_1_1_1_sva),
      (VEC_LOOP_j_1_12_0_sva_11_0[3]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[3]), (~ modExp_exp_1_2_1_sva),
      {and_dcpl_199 , and_dcpl_208 , and_dcpl_215 , and_dcpl_221});
  assign operator_64_false_1_mux1h_16_nl = MUX1HOT_s_1_3_2((~ modExp_exp_1_0_1_sva_1),
      (VEC_LOOP_j_1_12_0_sva_11_0[2]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[2]), {operator_64_false_1_or_2_itm
      , and_dcpl_208 , and_dcpl_215});
  assign operator_64_false_1_or_6_nl = and_dcpl_208 | and_dcpl_215;
  assign operator_64_false_1_operator_64_false_1_mux_1_nl = MUX_v_7_2_2(7'b0000001,
      COMP_LOOP_k_9_2_1_sva_6_0, operator_64_false_1_or_6_nl);
  assign nl_z_out_1 = ({operator_64_false_1_operator_64_false_1_or_1_nl , operator_64_false_1_mux1h_9_nl
      , operator_64_false_1_mux1h_10_nl , operator_64_false_1_mux1h_11_nl , operator_64_false_1_mux1h_12_nl
      , operator_64_false_1_mux1h_13_nl , operator_64_false_1_mux1h_14_nl , operator_64_false_1_mux1h_15_nl
      , operator_64_false_1_mux1h_16_nl}) + conv_u2u_7_10(operator_64_false_1_operator_64_false_1_mux_1_nl);
  assign z_out_1 = nl_z_out_1[9:0];
  assign COMP_LOOP_mux1h_83_nl = MUX1HOT_v_3_3_2((VEC_LOOP_j_1_12_0_sva_11_0[11:9]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:9]), 3'b001, {and_dcpl_230 , and_365_cse
      , COMP_LOOP_or_27_itm});
  assign COMP_LOOP_mux1h_84_nl = MUX1HOT_v_9_3_2((VEC_LOOP_j_1_12_0_sva_11_0[8:0]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[8:0]), (~ (STAGE_LOOP_lshift_psp_sva[9:1])),
      {and_dcpl_230 , and_365_cse , COMP_LOOP_or_27_itm});
  assign COMP_LOOP_or_34_nl = (~(and_dcpl_230 | and_365_cse)) | and_dcpl_242 | and_dcpl_244;
  assign COMP_LOOP_mux_41_nl = MUX_v_2_2_2(2'b01, 2'b10, and_dcpl_244);
  assign COMP_LOOP_COMP_LOOP_or_3_nl = MUX_v_2_2_2(COMP_LOOP_mux_41_nl, 2'b11, and_365_cse);
  assign nl_acc_2_nl = ({COMP_LOOP_mux1h_83_nl , COMP_LOOP_mux1h_84_nl , COMP_LOOP_or_34_nl})
      + conv_u2u_10_13({COMP_LOOP_k_9_2_1_sva_6_0 , COMP_LOOP_COMP_LOOP_or_3_nl ,
      1'b1});
  assign acc_2_nl = nl_acc_2_nl[12:0];
  assign z_out_2 = readslicef_13_12_1(acc_2_nl);
  assign and_532_nl = nor_332_cse & (fsm_output[2]) & (fsm_output[8]) & (fsm_output[5])
      & (~ (fsm_output[9])) & (fsm_output[1]) & (~ (fsm_output[7])) & and_dcpl_200;
  assign COMP_LOOP_or_35_nl = and_dcpl_244 | and_392_cse;
  assign COMP_LOOP_mux1h_85_nl = MUX1HOT_v_12_3_2(VEC_LOOP_j_1_12_0_sva_11_0, reg_VEC_LOOP_1_acc_1_psp_ftd_1,
      ({2'b00 , STAGE_LOOP_lshift_psp_sva}), {and_dcpl_253 , and_532_nl , COMP_LOOP_or_35_nl});
  assign COMP_LOOP_COMP_LOOP_or_4_nl = and_dcpl_253 | and_392_cse;
  assign nl_z_out_3 = COMP_LOOP_mux1h_85_nl + conv_u2u_9_12({COMP_LOOP_k_9_2_1_sva_6_0
      , COMP_LOOP_COMP_LOOP_or_4_nl , 1'b1});
  assign z_out_3 = nl_z_out_3[11:0];
  assign COMP_LOOP_COMP_LOOP_or_5_nl = (~(and_dcpl_283 | and_dcpl_292 | and_392_cse
      | and_dcpl_310)) | and_dcpl_302;
  assign COMP_LOOP_mux1h_86_nl = MUX1HOT_v_64_5_2(tmp_10_lpi_4_dfm, p_sva, ({57'b000000000000000000000000000000000000000000000000000000000
      , COMP_LOOP_k_9_2_1_sva_6_0}), (~ (operator_66_true_div_cmp_z[63:0])), ({61'b0000000000000000000000000000000000000000000000000000000000000
      , (z_out_6[3:1])}), {and_dcpl_283 , and_dcpl_292 , and_392_cse , and_dcpl_302
      , and_dcpl_310});
  assign COMP_LOOP_or_37_nl = and_392_cse | and_dcpl_302;
  assign COMP_LOOP_mux1h_87_nl = MUX1HOT_v_64_3_2(modExp_base_1_sva_mx1, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      64'b0000000000000000000000000000000000000000000000000000000000000011, {and_dcpl_283
      , COMP_LOOP_or_37_nl , and_dcpl_310});
  assign COMP_LOOP_or_36_nl = MUX_v_64_2_2(COMP_LOOP_mux1h_87_nl, 64'b1111111111111111111111111111111111111111111111111111111111111111,
      and_dcpl_292);
  assign nl_z_out_5 = ({COMP_LOOP_COMP_LOOP_or_5_nl , COMP_LOOP_mux1h_86_nl}) + conv_s2u_64_65(COMP_LOOP_or_36_nl);
  assign z_out_5 = nl_z_out_5[64:0];
  assign STAGE_LOOP_STAGE_LOOP_or_1_nl = ((modulo_result_rem_cmp_z[63]) & STAGE_LOOP_nor_itm)
      | and_dcpl_327;
  assign STAGE_LOOP_mux_55_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[62]), (~ (operator_64_false_acc_mut_63_0[62])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_103_nl = STAGE_LOOP_mux_55_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_56_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[61]), (~ (operator_64_false_acc_mut_63_0[61])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_104_nl = STAGE_LOOP_mux_56_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_57_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[60]), (~ (operator_64_false_acc_mut_63_0[60])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_105_nl = STAGE_LOOP_mux_57_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_58_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[59]), (~ (operator_64_false_acc_mut_63_0[59])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_106_nl = STAGE_LOOP_mux_58_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_59_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[58]), (~ (operator_64_false_acc_mut_63_0[58])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_107_nl = STAGE_LOOP_mux_59_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_60_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[57]), (~ (operator_64_false_acc_mut_63_0[57])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_108_nl = STAGE_LOOP_mux_60_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_61_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[56]), (~ (operator_64_false_acc_mut_63_0[56])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_109_nl = STAGE_LOOP_mux_61_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_62_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[55]), (~ (operator_64_false_acc_mut_63_0[55])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_110_nl = STAGE_LOOP_mux_62_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_63_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[54]), (~ (operator_64_false_acc_mut_63_0[54])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_111_nl = STAGE_LOOP_mux_63_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_64_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[53]), (~ (operator_64_false_acc_mut_63_0[53])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_112_nl = STAGE_LOOP_mux_64_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_65_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[52]), (~ (operator_64_false_acc_mut_63_0[52])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_113_nl = STAGE_LOOP_mux_65_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_66_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[51]), (~ (operator_64_false_acc_mut_63_0[51])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_114_nl = STAGE_LOOP_mux_66_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_67_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[50]), (~ (operator_64_false_acc_mut_63_0[50])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_115_nl = STAGE_LOOP_mux_67_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_68_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[49]), (~ (operator_64_false_acc_mut_63_0[49])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_116_nl = STAGE_LOOP_mux_68_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_69_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[48]), (~ (operator_64_false_acc_mut_63_0[48])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_117_nl = STAGE_LOOP_mux_69_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_70_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[47]), (~ (operator_64_false_acc_mut_63_0[47])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_118_nl = STAGE_LOOP_mux_70_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_71_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[46]), (~ (operator_64_false_acc_mut_63_0[46])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_119_nl = STAGE_LOOP_mux_71_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_72_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[45]), (~ (operator_64_false_acc_mut_63_0[45])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_120_nl = STAGE_LOOP_mux_72_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_73_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[44]), (~ (operator_64_false_acc_mut_63_0[44])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_121_nl = STAGE_LOOP_mux_73_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_74_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[43]), (~ (operator_64_false_acc_mut_63_0[43])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_122_nl = STAGE_LOOP_mux_74_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_75_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[42]), (~ (operator_64_false_acc_mut_63_0[42])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_123_nl = STAGE_LOOP_mux_75_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_76_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[41]), (~ (operator_64_false_acc_mut_63_0[41])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_124_nl = STAGE_LOOP_mux_76_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_77_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[40]), (~ (operator_64_false_acc_mut_63_0[40])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_125_nl = STAGE_LOOP_mux_77_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_78_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[39]), (~ (operator_64_false_acc_mut_63_0[39])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_126_nl = STAGE_LOOP_mux_78_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_79_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[38]), (~ (operator_64_false_acc_mut_63_0[38])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_127_nl = STAGE_LOOP_mux_79_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_80_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[37]), (~ (operator_64_false_acc_mut_63_0[37])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_128_nl = STAGE_LOOP_mux_80_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_81_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[36]), (~ (operator_64_false_acc_mut_63_0[36])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_129_nl = STAGE_LOOP_mux_81_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_82_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[35]), (~ (operator_64_false_acc_mut_63_0[35])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_130_nl = STAGE_LOOP_mux_82_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_83_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[34]), (~ (operator_64_false_acc_mut_63_0[34])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_131_nl = STAGE_LOOP_mux_83_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_84_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[33]), (~ (operator_64_false_acc_mut_63_0[33])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_132_nl = STAGE_LOOP_mux_84_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_85_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[32]), (~ (operator_64_false_acc_mut_63_0[32])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_133_nl = STAGE_LOOP_mux_85_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_86_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[31]), (~ (operator_64_false_acc_mut_63_0[31])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_134_nl = STAGE_LOOP_mux_86_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_87_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[30]), (~ (operator_64_false_acc_mut_63_0[30])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_135_nl = STAGE_LOOP_mux_87_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_88_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[29]), (~ (operator_64_false_acc_mut_63_0[29])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_136_nl = STAGE_LOOP_mux_88_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_89_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[28]), (~ (operator_64_false_acc_mut_63_0[28])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_137_nl = STAGE_LOOP_mux_89_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_90_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[27]), (~ (operator_64_false_acc_mut_63_0[27])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_138_nl = STAGE_LOOP_mux_90_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_91_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[26]), (~ (operator_64_false_acc_mut_63_0[26])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_139_nl = STAGE_LOOP_mux_91_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_92_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[25]), (~ (operator_64_false_acc_mut_63_0[25])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_140_nl = STAGE_LOOP_mux_92_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_93_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[24]), (~ (operator_64_false_acc_mut_63_0[24])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_141_nl = STAGE_LOOP_mux_93_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_94_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[23]), (~ (operator_64_false_acc_mut_63_0[23])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_142_nl = STAGE_LOOP_mux_94_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_95_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[22]), (~ (operator_64_false_acc_mut_63_0[22])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_143_nl = STAGE_LOOP_mux_95_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_96_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[21]), (~ (operator_64_false_acc_mut_63_0[21])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_144_nl = STAGE_LOOP_mux_96_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_97_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[20]), (~ (operator_64_false_acc_mut_63_0[20])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_145_nl = STAGE_LOOP_mux_97_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_98_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[19]), (~ (operator_64_false_acc_mut_63_0[19])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_146_nl = STAGE_LOOP_mux_98_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_99_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[18]), (~ (operator_64_false_acc_mut_63_0[18])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_147_nl = STAGE_LOOP_mux_99_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_100_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[17]), (~ (operator_64_false_acc_mut_63_0[17])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_148_nl = STAGE_LOOP_mux_100_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_101_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[16]), (~ (operator_64_false_acc_mut_63_0[16])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_149_nl = STAGE_LOOP_mux_101_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_102_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[15]), (~ (operator_64_false_acc_mut_63_0[15])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_150_nl = STAGE_LOOP_mux_102_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_103_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[14]), (~ (operator_64_false_acc_mut_63_0[14])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_151_nl = STAGE_LOOP_mux_103_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_104_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[13]), (~ (operator_64_false_acc_mut_63_0[13])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_152_nl = STAGE_LOOP_mux_104_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux_105_nl = MUX_s_1_2_2((modulo_result_rem_cmp_z[12]), (~ (operator_64_false_acc_mut_63_0[12])),
      and_dcpl_327);
  assign STAGE_LOOP_STAGE_LOOP_and_153_nl = STAGE_LOOP_mux_105_nl & STAGE_LOOP_nor_itm;
  assign STAGE_LOOP_mux1h_6_nl = MUX1HOT_v_2_4_2((modulo_result_rem_cmp_z[11:10]),
      (~ (operator_64_false_acc_mut_63_0[11:10])), (VEC_LOOP_j_1_12_0_sva_11_0[11:10]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]), {(~ mux_860_itm) , and_dcpl_327 ,
      and_dcpl_361 , and_dcpl_367});
  assign STAGE_LOOP_nor_106_nl = ~(and_dcpl_319 | and_dcpl_331 | and_dcpl_339 | and_dcpl_342
      | and_dcpl_345 | and_dcpl_352 | and_dcpl_354 | and_dcpl_356 | and_dcpl_357);
  assign STAGE_LOOP_and_4_nl = MUX_v_2_2_2(2'b00, STAGE_LOOP_mux1h_6_nl, STAGE_LOOP_nor_106_nl);
  assign nl_COMP_LOOP_acc_61_nl = (STAGE_LOOP_lshift_psp_sva[9:2]) + conv_u2u_7_8(COMP_LOOP_k_9_2_1_sva_6_0);
  assign COMP_LOOP_acc_61_nl = nl_COMP_LOOP_acc_61_nl[7:0];
  assign nl_COMP_LOOP_acc_62_nl = (STAGE_LOOP_lshift_psp_sva[9:1]) + conv_u2u_8_9({COMP_LOOP_k_9_2_1_sva_6_0
      , 1'b1});
  assign COMP_LOOP_acc_62_nl = nl_COMP_LOOP_acc_62_nl[8:0];
  assign STAGE_LOOP_or_10_nl = and_dcpl_331 | and_dcpl_352;
  assign STAGE_LOOP_or_11_nl = and_dcpl_342 | and_dcpl_356;
  assign STAGE_LOOP_mux1h_7_nl = MUX1HOT_v_9_8_2(({6'b000000 , (STAGE_LOOP_i_3_0_sva[3:1])}),
      (modulo_result_rem_cmp_z[9:1]), (~ (operator_64_false_acc_mut_63_0[9:1])),
      ({COMP_LOOP_acc_61_nl , (STAGE_LOOP_lshift_psp_sva[1])}), (z_out_3[9:1]), COMP_LOOP_acc_62_nl,
      (VEC_LOOP_j_1_12_0_sva_11_0[9:1]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9:1]), {and_dcpl_319
      , (~ mux_860_itm) , and_dcpl_327 , STAGE_LOOP_or_10_nl , STAGE_LOOP_or_ssc
      , STAGE_LOOP_or_11_nl , and_dcpl_361 , and_dcpl_367});
  assign STAGE_LOOP_or_12_nl = and_dcpl_331 | and_dcpl_342 | and_dcpl_352 | and_dcpl_356;
  assign STAGE_LOOP_mux1h_8_nl = MUX1HOT_s_1_7_2((STAGE_LOOP_i_3_0_sva[0]), (modulo_result_rem_cmp_z[0]),
      (~ (operator_64_false_acc_mut_63_0[0])), (STAGE_LOOP_lshift_psp_sva[0]), (z_out_3[0]),
      (VEC_LOOP_j_1_12_0_sva_11_0[0]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[0]), {and_dcpl_319
      , (~ mux_860_itm) , and_dcpl_327 , STAGE_LOOP_or_12_nl , STAGE_LOOP_or_ssc
      , and_dcpl_361 , and_dcpl_367});
  assign STAGE_LOOP_STAGE_LOOP_and_154_nl = (p_sva[63]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_155_nl = (p_sva[62]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_156_nl = (p_sva[61]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_157_nl = (p_sva[60]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_158_nl = (p_sva[59]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_159_nl = (p_sva[58]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_160_nl = (p_sva[57]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_161_nl = (p_sva[56]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_162_nl = (p_sva[55]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_163_nl = (p_sva[54]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_164_nl = (p_sva[53]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_165_nl = (p_sva[52]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_166_nl = (p_sva[51]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_167_nl = (p_sva[50]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_168_nl = (p_sva[49]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_169_nl = (p_sva[48]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_170_nl = (p_sva[47]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_171_nl = (p_sva[46]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_172_nl = (p_sva[45]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_173_nl = (p_sva[44]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_174_nl = (p_sva[43]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_175_nl = (p_sva[42]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_176_nl = (p_sva[41]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_177_nl = (p_sva[40]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_178_nl = (p_sva[39]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_179_nl = (p_sva[38]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_180_nl = (p_sva[37]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_181_nl = (p_sva[36]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_182_nl = (p_sva[35]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_183_nl = (p_sva[34]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_184_nl = (p_sva[33]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_185_nl = (p_sva[32]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_186_nl = (p_sva[31]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_187_nl = (p_sva[30]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_188_nl = (p_sva[29]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_189_nl = (p_sva[28]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_190_nl = (p_sva[27]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_191_nl = (p_sva[26]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_192_nl = (p_sva[25]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_193_nl = (p_sva[24]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_194_nl = (p_sva[23]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_195_nl = (p_sva[22]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_196_nl = (p_sva[21]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_197_nl = (p_sva[20]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_198_nl = (p_sva[19]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_199_nl = (p_sva[18]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_200_nl = (p_sva[17]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_201_nl = (p_sva[16]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_202_nl = (p_sva[15]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_203_nl = (p_sva[14]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_204_nl = (p_sva[13]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_STAGE_LOOP_and_205_nl = (p_sva[12]) & STAGE_LOOP_nor_53_itm;
  assign STAGE_LOOP_mux1h_9_nl = MUX1HOT_v_2_3_2((p_sva[11:10]), (VEC_LOOP_j_1_12_0_sva_11_0[11:10]),
      (reg_VEC_LOOP_1_acc_1_psp_ftd_1[11:10]), {(~ mux_860_itm) , STAGE_LOOP_or_1_itm
      , STAGE_LOOP_or_2_itm});
  assign STAGE_LOOP_nor_107_nl = ~(and_dcpl_319 | and_dcpl_327 | and_dcpl_361 | and_dcpl_367);
  assign STAGE_LOOP_and_5_nl = MUX_v_2_2_2(2'b00, STAGE_LOOP_mux1h_9_nl, STAGE_LOOP_nor_107_nl);
  assign STAGE_LOOP_or_13_nl = and_dcpl_319 | and_dcpl_327;
  assign STAGE_LOOP_or_14_nl = and_dcpl_361 | and_dcpl_367;
  assign STAGE_LOOP_mux1h_10_nl = MUX1HOT_v_10_5_2(10'b0000000001, (p_sva[9:0]),
      (VEC_LOOP_j_1_12_0_sva_11_0[9:0]), (reg_VEC_LOOP_1_acc_1_psp_ftd_1[9:0]), STAGE_LOOP_lshift_psp_sva,
      {STAGE_LOOP_or_13_nl , (~ mux_860_itm) , STAGE_LOOP_or_1_itm , STAGE_LOOP_or_2_itm
      , STAGE_LOOP_or_14_nl});
  assign nl_z_out_6 = ({STAGE_LOOP_STAGE_LOOP_or_1_nl , STAGE_LOOP_STAGE_LOOP_and_103_nl
      , STAGE_LOOP_STAGE_LOOP_and_104_nl , STAGE_LOOP_STAGE_LOOP_and_105_nl , STAGE_LOOP_STAGE_LOOP_and_106_nl
      , STAGE_LOOP_STAGE_LOOP_and_107_nl , STAGE_LOOP_STAGE_LOOP_and_108_nl , STAGE_LOOP_STAGE_LOOP_and_109_nl
      , STAGE_LOOP_STAGE_LOOP_and_110_nl , STAGE_LOOP_STAGE_LOOP_and_111_nl , STAGE_LOOP_STAGE_LOOP_and_112_nl
      , STAGE_LOOP_STAGE_LOOP_and_113_nl , STAGE_LOOP_STAGE_LOOP_and_114_nl , STAGE_LOOP_STAGE_LOOP_and_115_nl
      , STAGE_LOOP_STAGE_LOOP_and_116_nl , STAGE_LOOP_STAGE_LOOP_and_117_nl , STAGE_LOOP_STAGE_LOOP_and_118_nl
      , STAGE_LOOP_STAGE_LOOP_and_119_nl , STAGE_LOOP_STAGE_LOOP_and_120_nl , STAGE_LOOP_STAGE_LOOP_and_121_nl
      , STAGE_LOOP_STAGE_LOOP_and_122_nl , STAGE_LOOP_STAGE_LOOP_and_123_nl , STAGE_LOOP_STAGE_LOOP_and_124_nl
      , STAGE_LOOP_STAGE_LOOP_and_125_nl , STAGE_LOOP_STAGE_LOOP_and_126_nl , STAGE_LOOP_STAGE_LOOP_and_127_nl
      , STAGE_LOOP_STAGE_LOOP_and_128_nl , STAGE_LOOP_STAGE_LOOP_and_129_nl , STAGE_LOOP_STAGE_LOOP_and_130_nl
      , STAGE_LOOP_STAGE_LOOP_and_131_nl , STAGE_LOOP_STAGE_LOOP_and_132_nl , STAGE_LOOP_STAGE_LOOP_and_133_nl
      , STAGE_LOOP_STAGE_LOOP_and_134_nl , STAGE_LOOP_STAGE_LOOP_and_135_nl , STAGE_LOOP_STAGE_LOOP_and_136_nl
      , STAGE_LOOP_STAGE_LOOP_and_137_nl , STAGE_LOOP_STAGE_LOOP_and_138_nl , STAGE_LOOP_STAGE_LOOP_and_139_nl
      , STAGE_LOOP_STAGE_LOOP_and_140_nl , STAGE_LOOP_STAGE_LOOP_and_141_nl , STAGE_LOOP_STAGE_LOOP_and_142_nl
      , STAGE_LOOP_STAGE_LOOP_and_143_nl , STAGE_LOOP_STAGE_LOOP_and_144_nl , STAGE_LOOP_STAGE_LOOP_and_145_nl
      , STAGE_LOOP_STAGE_LOOP_and_146_nl , STAGE_LOOP_STAGE_LOOP_and_147_nl , STAGE_LOOP_STAGE_LOOP_and_148_nl
      , STAGE_LOOP_STAGE_LOOP_and_149_nl , STAGE_LOOP_STAGE_LOOP_and_150_nl , STAGE_LOOP_STAGE_LOOP_and_151_nl
      , STAGE_LOOP_STAGE_LOOP_and_152_nl , STAGE_LOOP_STAGE_LOOP_and_153_nl , STAGE_LOOP_and_4_nl
      , STAGE_LOOP_mux1h_7_nl , STAGE_LOOP_mux1h_8_nl}) + ({STAGE_LOOP_STAGE_LOOP_and_154_nl
      , STAGE_LOOP_STAGE_LOOP_and_155_nl , STAGE_LOOP_STAGE_LOOP_and_156_nl , STAGE_LOOP_STAGE_LOOP_and_157_nl
      , STAGE_LOOP_STAGE_LOOP_and_158_nl , STAGE_LOOP_STAGE_LOOP_and_159_nl , STAGE_LOOP_STAGE_LOOP_and_160_nl
      , STAGE_LOOP_STAGE_LOOP_and_161_nl , STAGE_LOOP_STAGE_LOOP_and_162_nl , STAGE_LOOP_STAGE_LOOP_and_163_nl
      , STAGE_LOOP_STAGE_LOOP_and_164_nl , STAGE_LOOP_STAGE_LOOP_and_165_nl , STAGE_LOOP_STAGE_LOOP_and_166_nl
      , STAGE_LOOP_STAGE_LOOP_and_167_nl , STAGE_LOOP_STAGE_LOOP_and_168_nl , STAGE_LOOP_STAGE_LOOP_and_169_nl
      , STAGE_LOOP_STAGE_LOOP_and_170_nl , STAGE_LOOP_STAGE_LOOP_and_171_nl , STAGE_LOOP_STAGE_LOOP_and_172_nl
      , STAGE_LOOP_STAGE_LOOP_and_173_nl , STAGE_LOOP_STAGE_LOOP_and_174_nl , STAGE_LOOP_STAGE_LOOP_and_175_nl
      , STAGE_LOOP_STAGE_LOOP_and_176_nl , STAGE_LOOP_STAGE_LOOP_and_177_nl , STAGE_LOOP_STAGE_LOOP_and_178_nl
      , STAGE_LOOP_STAGE_LOOP_and_179_nl , STAGE_LOOP_STAGE_LOOP_and_180_nl , STAGE_LOOP_STAGE_LOOP_and_181_nl
      , STAGE_LOOP_STAGE_LOOP_and_182_nl , STAGE_LOOP_STAGE_LOOP_and_183_nl , STAGE_LOOP_STAGE_LOOP_and_184_nl
      , STAGE_LOOP_STAGE_LOOP_and_185_nl , STAGE_LOOP_STAGE_LOOP_and_186_nl , STAGE_LOOP_STAGE_LOOP_and_187_nl
      , STAGE_LOOP_STAGE_LOOP_and_188_nl , STAGE_LOOP_STAGE_LOOP_and_189_nl , STAGE_LOOP_STAGE_LOOP_and_190_nl
      , STAGE_LOOP_STAGE_LOOP_and_191_nl , STAGE_LOOP_STAGE_LOOP_and_192_nl , STAGE_LOOP_STAGE_LOOP_and_193_nl
      , STAGE_LOOP_STAGE_LOOP_and_194_nl , STAGE_LOOP_STAGE_LOOP_and_195_nl , STAGE_LOOP_STAGE_LOOP_and_196_nl
      , STAGE_LOOP_STAGE_LOOP_and_197_nl , STAGE_LOOP_STAGE_LOOP_and_198_nl , STAGE_LOOP_STAGE_LOOP_and_199_nl
      , STAGE_LOOP_STAGE_LOOP_and_200_nl , STAGE_LOOP_STAGE_LOOP_and_201_nl , STAGE_LOOP_STAGE_LOOP_and_202_nl
      , STAGE_LOOP_STAGE_LOOP_and_203_nl , STAGE_LOOP_STAGE_LOOP_and_204_nl , STAGE_LOOP_STAGE_LOOP_and_205_nl
      , STAGE_LOOP_and_5_nl , STAGE_LOOP_mux1h_10_nl});
  assign z_out_6 = nl_z_out_6[63:0];
  assign and_533_nl = nor_332_cse & (fsm_output[2]) & and_dcpl_288 & (~ (fsm_output[9]))
      & (fsm_output[1]) & (~ (fsm_output[7])) & (~ (fsm_output[6])) & (fsm_output[0]);
  assign or_1078_nl = (fsm_output[7]) | mux_826_cse;
  assign nand_149_nl = ~((fsm_output[8]) & (fsm_output[2]) & (fsm_output[3]));
  assign mux_957_nl = MUX_s_1_2_2(nand_149_nl, or_614_cse, fsm_output[1]);
  assign mux_956_nl = MUX_s_1_2_2(mux_tmp_824, mux_957_nl, fsm_output[7]);
  assign mux_954_nl = MUX_s_1_2_2(or_1078_nl, mux_956_nl, fsm_output[6]);
  assign or_1080_nl = (fsm_output[7:6]!=2'b10) | mux_tmp_824;
  assign mux_953_nl = MUX_s_1_2_2(mux_954_nl, or_1080_nl, fsm_output[0]);
  assign modExp_while_if_modExp_while_if_nand_1_nl = ~(mux_866_itm & (mux_953_nl
      | (fsm_output[4]) | (~ (fsm_output[5])) | (fsm_output[9])));
  assign nor_461_nl = ~((fsm_output[7]) | (fsm_output[0]) | (fsm_output[6]) | (fsm_output[8])
      | (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[3])));
  assign nor_462_nl = ~((fsm_output[3:1]!=3'b001));
  assign nor_463_nl = ~((fsm_output[3:1]!=3'b100));
  assign mux_960_nl = MUX_s_1_2_2(nor_462_nl, nor_463_nl, fsm_output[8]);
  assign and_535_nl = (fsm_output[0]) & mux_960_nl;
  assign nor_464_nl = ~((fsm_output[6]) | mux_tmp_866);
  assign and_536_nl = (fsm_output[6]) & (~ mux_tmp_866);
  assign mux_961_nl = MUX_s_1_2_2(nor_464_nl, and_536_nl, fsm_output[0]);
  assign mux_959_nl = MUX_s_1_2_2(and_535_nl, mux_961_nl, fsm_output[7]);
  assign mux_958_nl = MUX_s_1_2_2(nor_461_nl, mux_959_nl, fsm_output[5]);
  assign and_534_nl = mux_958_nl & and_dcpl_109;
  assign modExp_while_if_mux1h_1_nl = MUX1HOT_v_64_3_2(modExp_result_sva, operator_64_false_acc_mut_63_0,
      modExp_base_1_sva, {and_533_nl , modExp_while_if_modExp_while_if_nand_1_nl
      , and_534_nl});
  assign modExp_while_if_modExp_while_if_nor_1_nl = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | mux_866_itm);
  assign modExp_while_if_and_6_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b01)
      & (~ mux_866_itm);
  assign modExp_while_if_and_7_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b10)
      & (~ mux_866_itm);
  assign modExp_while_if_and_8_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b11)
      & (~ mux_866_itm);
  assign modExp_while_if_modExp_while_if_mux1h_1_nl = MUX1HOT_v_64_5_2(modExp_base_1_sva,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
      {mux_866_itm , modExp_while_if_modExp_while_if_nor_1_nl , modExp_while_if_and_6_nl
      , modExp_while_if_and_7_nl , modExp_while_if_and_8_nl});
  assign nl_z_out_7 = modExp_while_if_mux1h_1_nl * modExp_while_if_modExp_while_if_mux1h_1_nl;
  assign z_out_7 = nl_z_out_7[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_5_2;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [4:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    MUX1HOT_v_10_5_2 = result;
  end
  endfunction


  function automatic [9:0] MUX1HOT_v_10_7_2;
    input [9:0] input_6;
    input [9:0] input_5;
    input [9:0] input_4;
    input [9:0] input_3;
    input [9:0] input_2;
    input [9:0] input_1;
    input [9:0] input_0;
    input [6:0] sel;
    reg [9:0] result;
  begin
    result = input_0 & {10{sel[0]}};
    result = result | ( input_1 & {10{sel[1]}});
    result = result | ( input_2 & {10{sel[2]}});
    result = result | ( input_3 & {10{sel[3]}});
    result = result | ( input_4 & {10{sel[4]}});
    result = result | ( input_5 & {10{sel[5]}});
    result = result | ( input_6 & {10{sel[6]}});
    MUX1HOT_v_10_7_2 = result;
  end
  endfunction


  function automatic [11:0] MUX1HOT_v_12_3_2;
    input [11:0] input_2;
    input [11:0] input_1;
    input [11:0] input_0;
    input [2:0] sel;
    reg [11:0] result;
  begin
    result = input_0 & {12{sel[0]}};
    result = result | ( input_1 & {12{sel[1]}});
    result = result | ( input_2 & {12{sel[2]}});
    MUX1HOT_v_12_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_4_2;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [3:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    MUX1HOT_v_64_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_5_2;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [4:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    MUX1HOT_v_64_5_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_3_2;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [2:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    MUX1HOT_v_9_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_8_2;
    input [8:0] input_7;
    input [8:0] input_6;
    input [8:0] input_5;
    input [8:0] input_4;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [7:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    result = result | ( input_4 & {9{sel[4]}});
    result = result | ( input_5 & {9{sel[5]}});
    result = result | ( input_6 & {9{sel[6]}});
    result = result | ( input_7 & {9{sel[7]}});
    MUX1HOT_v_9_8_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] conv_s2u_64_65 ;
    input [63:0]  vector ;
  begin
    conv_s2u_64_65 = {vector[63], vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_7_10 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_10 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_10_13 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_13 = {{3{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [9:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [9:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [9:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [9:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [9:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_10_64_1024_1024_64_1_gen
      vec_rsc_0_0_i (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_10_64_1024_1024_64_1_gen
      vec_rsc_0_1_i (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_10_64_1024_1024_64_1_gen
      vec_rsc_0_2_i (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_10_64_1024_1024_64_1_gen
      vec_rsc_0_3_i (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff)
    );
endmodule



