
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features; 
//       please enable Verilog2001 in the flow!

module mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers
   
    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC
   
    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a, 
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a, 
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v5.v 
module mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_1R1W_RBW_DUAL.v 
// Memory Type:            BLOCK
// Operating Mode:         Simple Dual Port (2-Port)
// Clock Mode:             Dual Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_1R1W_RBW_DUAL
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_1R1W_RBW_DUAL #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( clkr,clkr_en,clkw,clkw_en,d,q,radr,wadr,we);

  input  clkr;
  input  clkr_en;
  input  clkw;
  input  clkw_en;
  input [data_width-1:0] d;
  output [data_width-1:0] q;
  input [addr_width-1:0] radr;
  input [addr_width-1:0] wadr;
  input  we;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramq;
  
  // Port Map
  // readA :: CLOCK clkr ENABLE clkr_en DATA_OUT q ADDRESS radr
  // writeA :: CLOCK clkw ENABLE clkw_en DATA_IN d ADDRESS wadr WRITE_ENABLE we

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] radr_reg;
      reg [data_width-1:0] d_reg;
      reg [addr_width-1:0] wadr_reg;
      reg we_reg;
      
      always @(posedge clkr) begin
        if (clkr_en) begin
          radr_reg <= radr;
        end
      end
      always @(posedge clkw) begin
        if (clkw_en) begin
          d_reg <= d;
          wadr_reg <= wadr;
          we_reg <= we;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clkr) begin
        if (clkr_en) begin
            ramq <= mem[radr_reg];
        end
      end
      always @(posedge clkw) begin
        if (clkw_en) begin
            if (we_reg) begin
              mem[wadr_reg] <= d_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clkr) begin
        if (clkr_en) begin
            ramq <= mem[radr];
        end
      end
      always @(posedge clkw) begin
        if (clkw_en) begin
            if (we) begin
              mem[wadr] <= d;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign q = ramq;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpq;
      
      always @(posedge clkr) begin
        if (clkr_en) begin
          tmpq <= ramq;
        end
      end
      
      assign q = tmpq;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1q;
      
      reg [data_width-1:0] tmp2q;
      
      always @(posedge clkr) begin
        if (clkr_en) begin
          tmp1q <= ramq;
        end
      end
      
      always @(posedge clkr) begin
        if (clkr_en) begin
          tmp2q <= tmp1q;
        end
      end
      
      assign q = tmp2q;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Wed Sep 15 01:51:08 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [3:0] adra;
  input [3:0] adra_d;
  input [31:0] da_d;
  output [31:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen
    (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen (
  clkr_en, clkw_en, q, radr, we, d, wadr, clkr, clkr_en_d, clkw_en_d, d_d, q_d, radr_d,
      wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clkr_en;
  output clkw_en;
  input [31:0] q;
  output [3:0] radr;
  output we;
  output [31:0] d;
  output [3:0] wadr;
  input clkr;
  input clkr_en_d;
  input clkw_en_d;
  input [31:0] d_d;
  output [31:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkr_en = (clkr_en_d);
  assign clkw_en = (clkw_en_d);
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module peaseNTT_core_core_fsm (
  clk, rst, fsm_output, INNER_LOOP1_C_0_tr0, INNER_LOOP2_C_0_tr0, STAGE_LOOP_C_2_tr0,
      INNER_LOOP3_C_0_tr0, INNER_LOOP4_C_0_tr0, INNER_LOOP4_C_0_tr1
);
  input clk;
  input rst;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input INNER_LOOP1_C_0_tr0;
  input INNER_LOOP2_C_0_tr0;
  input STAGE_LOOP_C_2_tr0;
  input INNER_LOOP3_C_0_tr0;
  input INNER_LOOP4_C_0_tr0;
  input INNER_LOOP4_C_0_tr1;


  // FSM State Type Declaration for peaseNTT_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    STAGE_LOOP_C_0 = 4'd1,
    INNER_LOOP1_C_0 = 4'd2,
    STAGE_LOOP_C_1 = 4'd3,
    INNER_LOOP2_C_0 = 4'd4,
    STAGE_LOOP_C_2 = 4'd5,
    STAGE_LOOP1_C_0 = 4'd6,
    INNER_LOOP3_C_0 = 4'd7,
    STAGE_LOOP1_C_1 = 4'd8,
    INNER_LOOP4_C_0 = 4'd9,
    main_C_1 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : peaseNTT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = INNER_LOOP1_C_0;
      end
      INNER_LOOP1_C_0 : begin
        fsm_output = 11'b00000000100;
        if ( INNER_LOOP1_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = INNER_LOOP1_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 11'b00000001000;
        state_var_NS = INNER_LOOP2_C_0;
      end
      INNER_LOOP2_C_0 : begin
        fsm_output = 11'b00000010000;
        if ( INNER_LOOP2_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_2;
        end
        else begin
          state_var_NS = INNER_LOOP2_C_0;
        end
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 11'b00000100000;
        if ( STAGE_LOOP_C_2_tr0 ) begin
          state_var_NS = STAGE_LOOP1_C_0;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      STAGE_LOOP1_C_0 : begin
        fsm_output = 11'b00001000000;
        state_var_NS = INNER_LOOP3_C_0;
      end
      INNER_LOOP3_C_0 : begin
        fsm_output = 11'b00010000000;
        if ( INNER_LOOP3_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP1_C_1;
        end
        else begin
          state_var_NS = INNER_LOOP3_C_0;
        end
      end
      STAGE_LOOP1_C_1 : begin
        fsm_output = 11'b00100000000;
        state_var_NS = INNER_LOOP4_C_0;
      end
      INNER_LOOP4_C_0 : begin
        fsm_output = 11'b01000000000;
        if ( INNER_LOOP4_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else if ( INNER_LOOP4_C_0_tr1 ) begin
          state_var_NS = INNER_LOOP4_C_0;
        end
        else begin
          state_var_NS = STAGE_LOOP1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_core_wait_dp
// ------------------------------------------------------------------


module peaseNTT_core_wait_dp (
  yt_rsc_0_0_cgo_iro, yt_rsc_0_0_i_clkr_en_d, yt_rsc_0_16_cgo_iro, yt_rsc_0_16_i_clkr_en_d,
      yt_rsc_1_0_cgo_iro, yt_rsc_1_0_i_clkr_en_d, yt_rsc_1_16_cgo_iro, yt_rsc_1_16_i_clkr_en_d,
      yt_rsc_2_0_cgo_iro, yt_rsc_2_0_i_clkr_en_d, yt_rsc_2_16_cgo_iro, yt_rsc_2_16_i_clkr_en_d,
      yt_rsc_3_0_cgo_iro, yt_rsc_3_0_i_clkr_en_d, yt_rsc_3_16_cgo_iro, yt_rsc_3_16_i_clkr_en_d,
      yt_rsc_4_0_cgo_iro, yt_rsc_4_0_i_clkr_en_d, yt_rsc_4_16_cgo_iro, yt_rsc_4_16_i_clkr_en_d,
      yt_rsc_5_0_cgo_iro, yt_rsc_5_0_i_clkr_en_d, yt_rsc_5_16_cgo_iro, yt_rsc_5_16_i_clkr_en_d,
      yt_rsc_6_0_cgo_iro, yt_rsc_6_0_i_clkr_en_d, yt_rsc_6_16_cgo_iro, yt_rsc_6_16_i_clkr_en_d,
      yt_rsc_7_0_cgo_iro, yt_rsc_7_0_i_clkr_en_d, yt_rsc_7_16_cgo_iro, yt_rsc_7_16_i_clkr_en_d,
      ensig_cgo_iro, ensig_cgo_iro_17, yt_rsc_0_0_cgo, yt_rsc_0_16_cgo, yt_rsc_1_0_cgo,
      yt_rsc_1_16_cgo, yt_rsc_2_0_cgo, yt_rsc_2_16_cgo, yt_rsc_3_0_cgo, yt_rsc_3_16_cgo,
      yt_rsc_4_0_cgo, yt_rsc_4_16_cgo, yt_rsc_5_0_cgo, yt_rsc_5_16_cgo, yt_rsc_6_0_cgo,
      yt_rsc_6_16_cgo, yt_rsc_7_0_cgo, yt_rsc_7_16_cgo, ensig_cgo, mult_t_mul_cmp_en,
      ensig_cgo_17, mult_z_mul_cmp_1_en
);
  input yt_rsc_0_0_cgo_iro;
  output yt_rsc_0_0_i_clkr_en_d;
  input yt_rsc_0_16_cgo_iro;
  output yt_rsc_0_16_i_clkr_en_d;
  input yt_rsc_1_0_cgo_iro;
  output yt_rsc_1_0_i_clkr_en_d;
  input yt_rsc_1_16_cgo_iro;
  output yt_rsc_1_16_i_clkr_en_d;
  input yt_rsc_2_0_cgo_iro;
  output yt_rsc_2_0_i_clkr_en_d;
  input yt_rsc_2_16_cgo_iro;
  output yt_rsc_2_16_i_clkr_en_d;
  input yt_rsc_3_0_cgo_iro;
  output yt_rsc_3_0_i_clkr_en_d;
  input yt_rsc_3_16_cgo_iro;
  output yt_rsc_3_16_i_clkr_en_d;
  input yt_rsc_4_0_cgo_iro;
  output yt_rsc_4_0_i_clkr_en_d;
  input yt_rsc_4_16_cgo_iro;
  output yt_rsc_4_16_i_clkr_en_d;
  input yt_rsc_5_0_cgo_iro;
  output yt_rsc_5_0_i_clkr_en_d;
  input yt_rsc_5_16_cgo_iro;
  output yt_rsc_5_16_i_clkr_en_d;
  input yt_rsc_6_0_cgo_iro;
  output yt_rsc_6_0_i_clkr_en_d;
  input yt_rsc_6_16_cgo_iro;
  output yt_rsc_6_16_i_clkr_en_d;
  input yt_rsc_7_0_cgo_iro;
  output yt_rsc_7_0_i_clkr_en_d;
  input yt_rsc_7_16_cgo_iro;
  output yt_rsc_7_16_i_clkr_en_d;
  input ensig_cgo_iro;
  input ensig_cgo_iro_17;
  input yt_rsc_0_0_cgo;
  input yt_rsc_0_16_cgo;
  input yt_rsc_1_0_cgo;
  input yt_rsc_1_16_cgo;
  input yt_rsc_2_0_cgo;
  input yt_rsc_2_16_cgo;
  input yt_rsc_3_0_cgo;
  input yt_rsc_3_16_cgo;
  input yt_rsc_4_0_cgo;
  input yt_rsc_4_16_cgo;
  input yt_rsc_5_0_cgo;
  input yt_rsc_5_16_cgo;
  input yt_rsc_6_0_cgo;
  input yt_rsc_6_16_cgo;
  input yt_rsc_7_0_cgo;
  input yt_rsc_7_16_cgo;
  input ensig_cgo;
  output mult_t_mul_cmp_en;
  input ensig_cgo_17;
  output mult_z_mul_cmp_1_en;



  // Interconnect Declarations for Component Instantiations 
  assign yt_rsc_0_0_i_clkr_en_d = yt_rsc_0_0_cgo | yt_rsc_0_0_cgo_iro;
  assign yt_rsc_0_16_i_clkr_en_d = yt_rsc_0_16_cgo | yt_rsc_0_16_cgo_iro;
  assign yt_rsc_1_0_i_clkr_en_d = yt_rsc_1_0_cgo | yt_rsc_1_0_cgo_iro;
  assign yt_rsc_1_16_i_clkr_en_d = yt_rsc_1_16_cgo | yt_rsc_1_16_cgo_iro;
  assign yt_rsc_2_0_i_clkr_en_d = yt_rsc_2_0_cgo | yt_rsc_2_0_cgo_iro;
  assign yt_rsc_2_16_i_clkr_en_d = yt_rsc_2_16_cgo | yt_rsc_2_16_cgo_iro;
  assign yt_rsc_3_0_i_clkr_en_d = yt_rsc_3_0_cgo | yt_rsc_3_0_cgo_iro;
  assign yt_rsc_3_16_i_clkr_en_d = yt_rsc_3_16_cgo | yt_rsc_3_16_cgo_iro;
  assign yt_rsc_4_0_i_clkr_en_d = yt_rsc_4_0_cgo | yt_rsc_4_0_cgo_iro;
  assign yt_rsc_4_16_i_clkr_en_d = yt_rsc_4_16_cgo | yt_rsc_4_16_cgo_iro;
  assign yt_rsc_5_0_i_clkr_en_d = yt_rsc_5_0_cgo | yt_rsc_5_0_cgo_iro;
  assign yt_rsc_5_16_i_clkr_en_d = yt_rsc_5_16_cgo | yt_rsc_5_16_cgo_iro;
  assign yt_rsc_6_0_i_clkr_en_d = yt_rsc_6_0_cgo | yt_rsc_6_0_cgo_iro;
  assign yt_rsc_6_16_i_clkr_en_d = yt_rsc_6_16_cgo | yt_rsc_6_16_cgo_iro;
  assign yt_rsc_7_0_i_clkr_en_d = yt_rsc_7_0_cgo | yt_rsc_7_0_cgo_iro;
  assign yt_rsc_7_16_i_clkr_en_d = yt_rsc_7_16_cgo | yt_rsc_7_16_cgo_iro;
  assign mult_t_mul_cmp_en = ensig_cgo | ensig_cgo_iro;
  assign mult_z_mul_cmp_1_en = ensig_cgo_17 | ensig_cgo_iro_17;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_core
// ------------------------------------------------------------------


module peaseNTT_core (
  clk, rst, xt_rsc_triosy_0_0_lz, xt_rsc_triosy_0_1_lz, xt_rsc_triosy_0_2_lz, xt_rsc_triosy_0_3_lz,
      xt_rsc_triosy_0_4_lz, xt_rsc_triosy_0_5_lz, xt_rsc_triosy_0_6_lz, xt_rsc_triosy_0_7_lz,
      xt_rsc_triosy_0_8_lz, xt_rsc_triosy_0_9_lz, xt_rsc_triosy_0_10_lz, xt_rsc_triosy_0_11_lz,
      xt_rsc_triosy_0_12_lz, xt_rsc_triosy_0_13_lz, xt_rsc_triosy_0_14_lz, xt_rsc_triosy_0_15_lz,
      xt_rsc_triosy_0_16_lz, xt_rsc_triosy_0_17_lz, xt_rsc_triosy_0_18_lz, xt_rsc_triosy_0_19_lz,
      xt_rsc_triosy_0_20_lz, xt_rsc_triosy_0_21_lz, xt_rsc_triosy_0_22_lz, xt_rsc_triosy_0_23_lz,
      xt_rsc_triosy_0_24_lz, xt_rsc_triosy_0_25_lz, xt_rsc_triosy_0_26_lz, xt_rsc_triosy_0_27_lz,
      xt_rsc_triosy_0_28_lz, xt_rsc_triosy_0_29_lz, xt_rsc_triosy_0_30_lz, xt_rsc_triosy_0_31_lz,
      xt_rsc_triosy_1_0_lz, xt_rsc_triosy_1_1_lz, xt_rsc_triosy_1_2_lz, xt_rsc_triosy_1_3_lz,
      xt_rsc_triosy_1_4_lz, xt_rsc_triosy_1_5_lz, xt_rsc_triosy_1_6_lz, xt_rsc_triosy_1_7_lz,
      xt_rsc_triosy_1_8_lz, xt_rsc_triosy_1_9_lz, xt_rsc_triosy_1_10_lz, xt_rsc_triosy_1_11_lz,
      xt_rsc_triosy_1_12_lz, xt_rsc_triosy_1_13_lz, xt_rsc_triosy_1_14_lz, xt_rsc_triosy_1_15_lz,
      xt_rsc_triosy_1_16_lz, xt_rsc_triosy_1_17_lz, xt_rsc_triosy_1_18_lz, xt_rsc_triosy_1_19_lz,
      xt_rsc_triosy_1_20_lz, xt_rsc_triosy_1_21_lz, xt_rsc_triosy_1_22_lz, xt_rsc_triosy_1_23_lz,
      xt_rsc_triosy_1_24_lz, xt_rsc_triosy_1_25_lz, xt_rsc_triosy_1_26_lz, xt_rsc_triosy_1_27_lz,
      xt_rsc_triosy_1_28_lz, xt_rsc_triosy_1_29_lz, xt_rsc_triosy_1_30_lz, xt_rsc_triosy_1_31_lz,
      xt_rsc_triosy_2_0_lz, xt_rsc_triosy_2_1_lz, xt_rsc_triosy_2_2_lz, xt_rsc_triosy_2_3_lz,
      xt_rsc_triosy_2_4_lz, xt_rsc_triosy_2_5_lz, xt_rsc_triosy_2_6_lz, xt_rsc_triosy_2_7_lz,
      xt_rsc_triosy_2_8_lz, xt_rsc_triosy_2_9_lz, xt_rsc_triosy_2_10_lz, xt_rsc_triosy_2_11_lz,
      xt_rsc_triosy_2_12_lz, xt_rsc_triosy_2_13_lz, xt_rsc_triosy_2_14_lz, xt_rsc_triosy_2_15_lz,
      xt_rsc_triosy_2_16_lz, xt_rsc_triosy_2_17_lz, xt_rsc_triosy_2_18_lz, xt_rsc_triosy_2_19_lz,
      xt_rsc_triosy_2_20_lz, xt_rsc_triosy_2_21_lz, xt_rsc_triosy_2_22_lz, xt_rsc_triosy_2_23_lz,
      xt_rsc_triosy_2_24_lz, xt_rsc_triosy_2_25_lz, xt_rsc_triosy_2_26_lz, xt_rsc_triosy_2_27_lz,
      xt_rsc_triosy_2_28_lz, xt_rsc_triosy_2_29_lz, xt_rsc_triosy_2_30_lz, xt_rsc_triosy_2_31_lz,
      xt_rsc_triosy_3_0_lz, xt_rsc_triosy_3_1_lz, xt_rsc_triosy_3_2_lz, xt_rsc_triosy_3_3_lz,
      xt_rsc_triosy_3_4_lz, xt_rsc_triosy_3_5_lz, xt_rsc_triosy_3_6_lz, xt_rsc_triosy_3_7_lz,
      xt_rsc_triosy_3_8_lz, xt_rsc_triosy_3_9_lz, xt_rsc_triosy_3_10_lz, xt_rsc_triosy_3_11_lz,
      xt_rsc_triosy_3_12_lz, xt_rsc_triosy_3_13_lz, xt_rsc_triosy_3_14_lz, xt_rsc_triosy_3_15_lz,
      xt_rsc_triosy_3_16_lz, xt_rsc_triosy_3_17_lz, xt_rsc_triosy_3_18_lz, xt_rsc_triosy_3_19_lz,
      xt_rsc_triosy_3_20_lz, xt_rsc_triosy_3_21_lz, xt_rsc_triosy_3_22_lz, xt_rsc_triosy_3_23_lz,
      xt_rsc_triosy_3_24_lz, xt_rsc_triosy_3_25_lz, xt_rsc_triosy_3_26_lz, xt_rsc_triosy_3_27_lz,
      xt_rsc_triosy_3_28_lz, xt_rsc_triosy_3_29_lz, xt_rsc_triosy_3_30_lz, xt_rsc_triosy_3_31_lz,
      xt_rsc_triosy_4_0_lz, xt_rsc_triosy_4_1_lz, xt_rsc_triosy_4_2_lz, xt_rsc_triosy_4_3_lz,
      xt_rsc_triosy_4_4_lz, xt_rsc_triosy_4_5_lz, xt_rsc_triosy_4_6_lz, xt_rsc_triosy_4_7_lz,
      xt_rsc_triosy_4_8_lz, xt_rsc_triosy_4_9_lz, xt_rsc_triosy_4_10_lz, xt_rsc_triosy_4_11_lz,
      xt_rsc_triosy_4_12_lz, xt_rsc_triosy_4_13_lz, xt_rsc_triosy_4_14_lz, xt_rsc_triosy_4_15_lz,
      xt_rsc_triosy_4_16_lz, xt_rsc_triosy_4_17_lz, xt_rsc_triosy_4_18_lz, xt_rsc_triosy_4_19_lz,
      xt_rsc_triosy_4_20_lz, xt_rsc_triosy_4_21_lz, xt_rsc_triosy_4_22_lz, xt_rsc_triosy_4_23_lz,
      xt_rsc_triosy_4_24_lz, xt_rsc_triosy_4_25_lz, xt_rsc_triosy_4_26_lz, xt_rsc_triosy_4_27_lz,
      xt_rsc_triosy_4_28_lz, xt_rsc_triosy_4_29_lz, xt_rsc_triosy_4_30_lz, xt_rsc_triosy_4_31_lz,
      xt_rsc_triosy_5_0_lz, xt_rsc_triosy_5_1_lz, xt_rsc_triosy_5_2_lz, xt_rsc_triosy_5_3_lz,
      xt_rsc_triosy_5_4_lz, xt_rsc_triosy_5_5_lz, xt_rsc_triosy_5_6_lz, xt_rsc_triosy_5_7_lz,
      xt_rsc_triosy_5_8_lz, xt_rsc_triosy_5_9_lz, xt_rsc_triosy_5_10_lz, xt_rsc_triosy_5_11_lz,
      xt_rsc_triosy_5_12_lz, xt_rsc_triosy_5_13_lz, xt_rsc_triosy_5_14_lz, xt_rsc_triosy_5_15_lz,
      xt_rsc_triosy_5_16_lz, xt_rsc_triosy_5_17_lz, xt_rsc_triosy_5_18_lz, xt_rsc_triosy_5_19_lz,
      xt_rsc_triosy_5_20_lz, xt_rsc_triosy_5_21_lz, xt_rsc_triosy_5_22_lz, xt_rsc_triosy_5_23_lz,
      xt_rsc_triosy_5_24_lz, xt_rsc_triosy_5_25_lz, xt_rsc_triosy_5_26_lz, xt_rsc_triosy_5_27_lz,
      xt_rsc_triosy_5_28_lz, xt_rsc_triosy_5_29_lz, xt_rsc_triosy_5_30_lz, xt_rsc_triosy_5_31_lz,
      xt_rsc_triosy_6_0_lz, xt_rsc_triosy_6_1_lz, xt_rsc_triosy_6_2_lz, xt_rsc_triosy_6_3_lz,
      xt_rsc_triosy_6_4_lz, xt_rsc_triosy_6_5_lz, xt_rsc_triosy_6_6_lz, xt_rsc_triosy_6_7_lz,
      xt_rsc_triosy_6_8_lz, xt_rsc_triosy_6_9_lz, xt_rsc_triosy_6_10_lz, xt_rsc_triosy_6_11_lz,
      xt_rsc_triosy_6_12_lz, xt_rsc_triosy_6_13_lz, xt_rsc_triosy_6_14_lz, xt_rsc_triosy_6_15_lz,
      xt_rsc_triosy_6_16_lz, xt_rsc_triosy_6_17_lz, xt_rsc_triosy_6_18_lz, xt_rsc_triosy_6_19_lz,
      xt_rsc_triosy_6_20_lz, xt_rsc_triosy_6_21_lz, xt_rsc_triosy_6_22_lz, xt_rsc_triosy_6_23_lz,
      xt_rsc_triosy_6_24_lz, xt_rsc_triosy_6_25_lz, xt_rsc_triosy_6_26_lz, xt_rsc_triosy_6_27_lz,
      xt_rsc_triosy_6_28_lz, xt_rsc_triosy_6_29_lz, xt_rsc_triosy_6_30_lz, xt_rsc_triosy_6_31_lz,
      xt_rsc_triosy_7_0_lz, xt_rsc_triosy_7_1_lz, xt_rsc_triosy_7_2_lz, xt_rsc_triosy_7_3_lz,
      xt_rsc_triosy_7_4_lz, xt_rsc_triosy_7_5_lz, xt_rsc_triosy_7_6_lz, xt_rsc_triosy_7_7_lz,
      xt_rsc_triosy_7_8_lz, xt_rsc_triosy_7_9_lz, xt_rsc_triosy_7_10_lz, xt_rsc_triosy_7_11_lz,
      xt_rsc_triosy_7_12_lz, xt_rsc_triosy_7_13_lz, xt_rsc_triosy_7_14_lz, xt_rsc_triosy_7_15_lz,
      xt_rsc_triosy_7_16_lz, xt_rsc_triosy_7_17_lz, xt_rsc_triosy_7_18_lz, xt_rsc_triosy_7_19_lz,
      xt_rsc_triosy_7_20_lz, xt_rsc_triosy_7_21_lz, xt_rsc_triosy_7_22_lz, xt_rsc_triosy_7_23_lz,
      xt_rsc_triosy_7_24_lz, xt_rsc_triosy_7_25_lz, xt_rsc_triosy_7_26_lz, xt_rsc_triosy_7_27_lz,
      xt_rsc_triosy_7_28_lz, xt_rsc_triosy_7_29_lz, xt_rsc_triosy_7_30_lz, xt_rsc_triosy_7_31_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_0_0_lz, twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz, twiddle_rsc_triosy_0_3_lz, twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz, twiddle_rsc_triosy_0_6_lz, twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz, twiddle_rsc_triosy_0_9_lz, twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz, twiddle_rsc_triosy_0_12_lz, twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz, twiddle_rsc_triosy_0_15_lz, twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_triosy_0_1_lz, twiddle_h_rsc_triosy_0_2_lz, twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_triosy_0_4_lz, twiddle_h_rsc_triosy_0_5_lz, twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_triosy_0_7_lz, twiddle_h_rsc_triosy_0_8_lz, twiddle_h_rsc_triosy_0_9_lz,
      twiddle_h_rsc_triosy_0_10_lz, twiddle_h_rsc_triosy_0_11_lz, twiddle_h_rsc_triosy_0_12_lz,
      twiddle_h_rsc_triosy_0_13_lz, twiddle_h_rsc_triosy_0_14_lz, twiddle_h_rsc_triosy_0_15_lz,
      yt_rsc_0_0_i_clkr_en_d, yt_rsc_0_0_i_q_d, yt_rsc_0_1_i_q_d, yt_rsc_0_2_i_q_d,
      yt_rsc_0_3_i_q_d, yt_rsc_0_4_i_q_d, yt_rsc_0_5_i_q_d, yt_rsc_0_6_i_q_d, yt_rsc_0_7_i_q_d,
      yt_rsc_0_8_i_q_d, yt_rsc_0_9_i_q_d, yt_rsc_0_10_i_q_d, yt_rsc_0_11_i_q_d, yt_rsc_0_12_i_q_d,
      yt_rsc_0_13_i_q_d, yt_rsc_0_14_i_q_d, yt_rsc_0_15_i_q_d, yt_rsc_0_16_i_clkr_en_d,
      yt_rsc_0_16_i_q_d, yt_rsc_0_17_i_q_d, yt_rsc_0_18_i_q_d, yt_rsc_0_19_i_q_d,
      yt_rsc_0_20_i_q_d, yt_rsc_0_21_i_q_d, yt_rsc_0_22_i_q_d, yt_rsc_0_23_i_q_d,
      yt_rsc_0_24_i_q_d, yt_rsc_0_25_i_q_d, yt_rsc_0_26_i_q_d, yt_rsc_0_27_i_q_d,
      yt_rsc_0_28_i_q_d, yt_rsc_0_29_i_q_d, yt_rsc_0_30_i_q_d, yt_rsc_0_31_i_q_d,
      yt_rsc_1_0_i_clkr_en_d, yt_rsc_1_0_i_q_d, yt_rsc_1_1_i_q_d, yt_rsc_1_2_i_q_d,
      yt_rsc_1_3_i_q_d, yt_rsc_1_4_i_q_d, yt_rsc_1_5_i_q_d, yt_rsc_1_6_i_q_d, yt_rsc_1_7_i_q_d,
      yt_rsc_1_8_i_q_d, yt_rsc_1_9_i_q_d, yt_rsc_1_10_i_q_d, yt_rsc_1_11_i_q_d, yt_rsc_1_12_i_q_d,
      yt_rsc_1_13_i_q_d, yt_rsc_1_14_i_q_d, yt_rsc_1_15_i_q_d, yt_rsc_1_16_i_clkr_en_d,
      yt_rsc_1_16_i_q_d, yt_rsc_1_17_i_q_d, yt_rsc_1_18_i_q_d, yt_rsc_1_19_i_q_d,
      yt_rsc_1_20_i_q_d, yt_rsc_1_21_i_q_d, yt_rsc_1_22_i_q_d, yt_rsc_1_23_i_q_d,
      yt_rsc_1_24_i_q_d, yt_rsc_1_25_i_q_d, yt_rsc_1_26_i_q_d, yt_rsc_1_27_i_q_d,
      yt_rsc_1_28_i_q_d, yt_rsc_1_29_i_q_d, yt_rsc_1_30_i_q_d, yt_rsc_1_31_i_q_d,
      yt_rsc_2_0_i_clkr_en_d, yt_rsc_2_0_i_q_d, yt_rsc_2_1_i_q_d, yt_rsc_2_2_i_q_d,
      yt_rsc_2_3_i_q_d, yt_rsc_2_4_i_q_d, yt_rsc_2_5_i_q_d, yt_rsc_2_6_i_q_d, yt_rsc_2_7_i_q_d,
      yt_rsc_2_8_i_q_d, yt_rsc_2_9_i_q_d, yt_rsc_2_10_i_q_d, yt_rsc_2_11_i_q_d, yt_rsc_2_12_i_q_d,
      yt_rsc_2_13_i_q_d, yt_rsc_2_14_i_q_d, yt_rsc_2_15_i_q_d, yt_rsc_2_16_i_clkr_en_d,
      yt_rsc_2_16_i_q_d, yt_rsc_2_17_i_q_d, yt_rsc_2_18_i_q_d, yt_rsc_2_19_i_q_d,
      yt_rsc_2_20_i_q_d, yt_rsc_2_21_i_q_d, yt_rsc_2_22_i_q_d, yt_rsc_2_23_i_q_d,
      yt_rsc_2_24_i_q_d, yt_rsc_2_25_i_q_d, yt_rsc_2_26_i_q_d, yt_rsc_2_27_i_q_d,
      yt_rsc_2_28_i_q_d, yt_rsc_2_29_i_q_d, yt_rsc_2_30_i_q_d, yt_rsc_2_31_i_q_d,
      yt_rsc_3_0_i_clkr_en_d, yt_rsc_3_0_i_q_d, yt_rsc_3_1_i_q_d, yt_rsc_3_2_i_q_d,
      yt_rsc_3_3_i_q_d, yt_rsc_3_4_i_q_d, yt_rsc_3_5_i_q_d, yt_rsc_3_6_i_q_d, yt_rsc_3_7_i_q_d,
      yt_rsc_3_8_i_q_d, yt_rsc_3_9_i_q_d, yt_rsc_3_10_i_q_d, yt_rsc_3_11_i_q_d, yt_rsc_3_12_i_q_d,
      yt_rsc_3_13_i_q_d, yt_rsc_3_14_i_q_d, yt_rsc_3_15_i_q_d, yt_rsc_3_16_i_clkr_en_d,
      yt_rsc_3_16_i_q_d, yt_rsc_3_17_i_q_d, yt_rsc_3_18_i_q_d, yt_rsc_3_19_i_q_d,
      yt_rsc_3_20_i_q_d, yt_rsc_3_21_i_q_d, yt_rsc_3_22_i_q_d, yt_rsc_3_23_i_q_d,
      yt_rsc_3_24_i_q_d, yt_rsc_3_25_i_q_d, yt_rsc_3_26_i_q_d, yt_rsc_3_27_i_q_d,
      yt_rsc_3_28_i_q_d, yt_rsc_3_29_i_q_d, yt_rsc_3_30_i_q_d, yt_rsc_3_31_i_q_d,
      yt_rsc_4_0_i_clkr_en_d, yt_rsc_4_0_i_q_d, yt_rsc_4_1_i_q_d, yt_rsc_4_2_i_q_d,
      yt_rsc_4_3_i_q_d, yt_rsc_4_4_i_q_d, yt_rsc_4_5_i_q_d, yt_rsc_4_6_i_q_d, yt_rsc_4_7_i_q_d,
      yt_rsc_4_8_i_q_d, yt_rsc_4_9_i_q_d, yt_rsc_4_10_i_q_d, yt_rsc_4_11_i_q_d, yt_rsc_4_12_i_q_d,
      yt_rsc_4_13_i_q_d, yt_rsc_4_14_i_q_d, yt_rsc_4_15_i_q_d, yt_rsc_4_16_i_clkr_en_d,
      yt_rsc_4_16_i_q_d, yt_rsc_4_17_i_q_d, yt_rsc_4_18_i_q_d, yt_rsc_4_19_i_q_d,
      yt_rsc_4_20_i_q_d, yt_rsc_4_21_i_q_d, yt_rsc_4_22_i_q_d, yt_rsc_4_23_i_q_d,
      yt_rsc_4_24_i_q_d, yt_rsc_4_25_i_q_d, yt_rsc_4_26_i_q_d, yt_rsc_4_27_i_q_d,
      yt_rsc_4_28_i_q_d, yt_rsc_4_29_i_q_d, yt_rsc_4_30_i_q_d, yt_rsc_4_31_i_q_d,
      yt_rsc_5_0_i_clkr_en_d, yt_rsc_5_0_i_q_d, yt_rsc_5_1_i_q_d, yt_rsc_5_2_i_q_d,
      yt_rsc_5_3_i_q_d, yt_rsc_5_4_i_q_d, yt_rsc_5_5_i_q_d, yt_rsc_5_6_i_q_d, yt_rsc_5_7_i_q_d,
      yt_rsc_5_8_i_q_d, yt_rsc_5_9_i_q_d, yt_rsc_5_10_i_q_d, yt_rsc_5_11_i_q_d, yt_rsc_5_12_i_q_d,
      yt_rsc_5_13_i_q_d, yt_rsc_5_14_i_q_d, yt_rsc_5_15_i_q_d, yt_rsc_5_16_i_clkr_en_d,
      yt_rsc_5_16_i_q_d, yt_rsc_5_17_i_q_d, yt_rsc_5_18_i_q_d, yt_rsc_5_19_i_q_d,
      yt_rsc_5_20_i_q_d, yt_rsc_5_21_i_q_d, yt_rsc_5_22_i_q_d, yt_rsc_5_23_i_q_d,
      yt_rsc_5_24_i_q_d, yt_rsc_5_25_i_q_d, yt_rsc_5_26_i_q_d, yt_rsc_5_27_i_q_d,
      yt_rsc_5_28_i_q_d, yt_rsc_5_29_i_q_d, yt_rsc_5_30_i_q_d, yt_rsc_5_31_i_q_d,
      yt_rsc_6_0_i_clkr_en_d, yt_rsc_6_0_i_q_d, yt_rsc_6_1_i_q_d, yt_rsc_6_2_i_q_d,
      yt_rsc_6_3_i_q_d, yt_rsc_6_4_i_q_d, yt_rsc_6_5_i_q_d, yt_rsc_6_6_i_q_d, yt_rsc_6_7_i_q_d,
      yt_rsc_6_8_i_q_d, yt_rsc_6_9_i_q_d, yt_rsc_6_10_i_q_d, yt_rsc_6_11_i_q_d, yt_rsc_6_12_i_q_d,
      yt_rsc_6_13_i_q_d, yt_rsc_6_14_i_q_d, yt_rsc_6_15_i_q_d, yt_rsc_6_16_i_clkr_en_d,
      yt_rsc_6_16_i_q_d, yt_rsc_6_17_i_q_d, yt_rsc_6_18_i_q_d, yt_rsc_6_19_i_q_d,
      yt_rsc_6_20_i_q_d, yt_rsc_6_21_i_q_d, yt_rsc_6_22_i_q_d, yt_rsc_6_23_i_q_d,
      yt_rsc_6_24_i_q_d, yt_rsc_6_25_i_q_d, yt_rsc_6_26_i_q_d, yt_rsc_6_27_i_q_d,
      yt_rsc_6_28_i_q_d, yt_rsc_6_29_i_q_d, yt_rsc_6_30_i_q_d, yt_rsc_6_31_i_q_d,
      yt_rsc_7_0_i_clkr_en_d, yt_rsc_7_0_i_q_d, yt_rsc_7_1_i_q_d, yt_rsc_7_2_i_q_d,
      yt_rsc_7_3_i_q_d, yt_rsc_7_4_i_q_d, yt_rsc_7_5_i_q_d, yt_rsc_7_6_i_q_d, yt_rsc_7_7_i_q_d,
      yt_rsc_7_8_i_q_d, yt_rsc_7_9_i_q_d, yt_rsc_7_10_i_q_d, yt_rsc_7_11_i_q_d, yt_rsc_7_12_i_q_d,
      yt_rsc_7_13_i_q_d, yt_rsc_7_14_i_q_d, yt_rsc_7_15_i_q_d, yt_rsc_7_16_i_clkr_en_d,
      yt_rsc_7_16_i_q_d, yt_rsc_7_17_i_q_d, yt_rsc_7_18_i_q_d, yt_rsc_7_19_i_q_d,
      yt_rsc_7_20_i_q_d, yt_rsc_7_21_i_q_d, yt_rsc_7_22_i_q_d, yt_rsc_7_23_i_q_d,
      yt_rsc_7_24_i_q_d, yt_rsc_7_25_i_q_d, yt_rsc_7_26_i_q_d, yt_rsc_7_27_i_q_d,
      yt_rsc_7_28_i_q_d, yt_rsc_7_29_i_q_d, yt_rsc_7_30_i_q_d, yt_rsc_7_31_i_q_d,
      xt_rsc_0_0_i_qa_d, xt_rsc_0_1_i_qa_d, xt_rsc_0_2_i_qa_d, xt_rsc_0_3_i_qa_d,
      xt_rsc_0_4_i_qa_d, xt_rsc_0_5_i_qa_d, xt_rsc_0_6_i_qa_d, xt_rsc_0_7_i_qa_d,
      xt_rsc_0_8_i_qa_d, xt_rsc_0_9_i_qa_d, xt_rsc_0_10_i_qa_d, xt_rsc_0_11_i_qa_d,
      xt_rsc_0_12_i_qa_d, xt_rsc_0_13_i_qa_d, xt_rsc_0_14_i_qa_d, xt_rsc_0_15_i_qa_d,
      xt_rsc_0_16_i_qa_d, xt_rsc_0_17_i_qa_d, xt_rsc_0_18_i_qa_d, xt_rsc_0_19_i_qa_d,
      xt_rsc_0_20_i_qa_d, xt_rsc_0_21_i_qa_d, xt_rsc_0_22_i_qa_d, xt_rsc_0_23_i_qa_d,
      xt_rsc_0_24_i_qa_d, xt_rsc_0_25_i_qa_d, xt_rsc_0_26_i_qa_d, xt_rsc_0_27_i_qa_d,
      xt_rsc_0_28_i_qa_d, xt_rsc_0_29_i_qa_d, xt_rsc_0_30_i_qa_d, xt_rsc_0_31_i_qa_d,
      xt_rsc_1_0_i_qa_d, xt_rsc_1_1_i_qa_d, xt_rsc_1_2_i_qa_d, xt_rsc_1_3_i_qa_d,
      xt_rsc_1_4_i_qa_d, xt_rsc_1_5_i_qa_d, xt_rsc_1_6_i_qa_d, xt_rsc_1_7_i_qa_d,
      xt_rsc_1_8_i_qa_d, xt_rsc_1_9_i_qa_d, xt_rsc_1_10_i_qa_d, xt_rsc_1_11_i_qa_d,
      xt_rsc_1_12_i_qa_d, xt_rsc_1_13_i_qa_d, xt_rsc_1_14_i_qa_d, xt_rsc_1_15_i_qa_d,
      xt_rsc_1_16_i_qa_d, xt_rsc_1_17_i_qa_d, xt_rsc_1_18_i_qa_d, xt_rsc_1_19_i_qa_d,
      xt_rsc_1_20_i_qa_d, xt_rsc_1_21_i_qa_d, xt_rsc_1_22_i_qa_d, xt_rsc_1_23_i_qa_d,
      xt_rsc_1_24_i_qa_d, xt_rsc_1_25_i_qa_d, xt_rsc_1_26_i_qa_d, xt_rsc_1_27_i_qa_d,
      xt_rsc_1_28_i_qa_d, xt_rsc_1_29_i_qa_d, xt_rsc_1_30_i_qa_d, xt_rsc_1_31_i_qa_d,
      xt_rsc_2_0_i_qa_d, xt_rsc_2_1_i_qa_d, xt_rsc_2_2_i_qa_d, xt_rsc_2_3_i_qa_d,
      xt_rsc_2_4_i_qa_d, xt_rsc_2_5_i_qa_d, xt_rsc_2_6_i_qa_d, xt_rsc_2_7_i_qa_d,
      xt_rsc_2_8_i_qa_d, xt_rsc_2_9_i_qa_d, xt_rsc_2_10_i_qa_d, xt_rsc_2_11_i_qa_d,
      xt_rsc_2_12_i_qa_d, xt_rsc_2_13_i_qa_d, xt_rsc_2_14_i_qa_d, xt_rsc_2_15_i_qa_d,
      xt_rsc_2_16_i_qa_d, xt_rsc_2_17_i_qa_d, xt_rsc_2_18_i_qa_d, xt_rsc_2_19_i_qa_d,
      xt_rsc_2_20_i_qa_d, xt_rsc_2_21_i_qa_d, xt_rsc_2_22_i_qa_d, xt_rsc_2_23_i_qa_d,
      xt_rsc_2_24_i_qa_d, xt_rsc_2_25_i_qa_d, xt_rsc_2_26_i_qa_d, xt_rsc_2_27_i_qa_d,
      xt_rsc_2_28_i_qa_d, xt_rsc_2_29_i_qa_d, xt_rsc_2_30_i_qa_d, xt_rsc_2_31_i_qa_d,
      xt_rsc_3_0_i_qa_d, xt_rsc_3_1_i_qa_d, xt_rsc_3_2_i_qa_d, xt_rsc_3_3_i_qa_d,
      xt_rsc_3_4_i_qa_d, xt_rsc_3_5_i_qa_d, xt_rsc_3_6_i_qa_d, xt_rsc_3_7_i_qa_d,
      xt_rsc_3_8_i_qa_d, xt_rsc_3_9_i_qa_d, xt_rsc_3_10_i_qa_d, xt_rsc_3_11_i_qa_d,
      xt_rsc_3_12_i_qa_d, xt_rsc_3_13_i_qa_d, xt_rsc_3_14_i_qa_d, xt_rsc_3_15_i_qa_d,
      xt_rsc_3_16_i_qa_d, xt_rsc_3_17_i_qa_d, xt_rsc_3_18_i_qa_d, xt_rsc_3_19_i_qa_d,
      xt_rsc_3_20_i_qa_d, xt_rsc_3_21_i_qa_d, xt_rsc_3_22_i_qa_d, xt_rsc_3_23_i_qa_d,
      xt_rsc_3_24_i_qa_d, xt_rsc_3_25_i_qa_d, xt_rsc_3_26_i_qa_d, xt_rsc_3_27_i_qa_d,
      xt_rsc_3_28_i_qa_d, xt_rsc_3_29_i_qa_d, xt_rsc_3_30_i_qa_d, xt_rsc_3_31_i_qa_d,
      xt_rsc_4_0_i_qa_d, xt_rsc_4_1_i_qa_d, xt_rsc_4_2_i_qa_d, xt_rsc_4_3_i_qa_d,
      xt_rsc_4_4_i_qa_d, xt_rsc_4_5_i_qa_d, xt_rsc_4_6_i_qa_d, xt_rsc_4_7_i_qa_d,
      xt_rsc_4_8_i_qa_d, xt_rsc_4_9_i_qa_d, xt_rsc_4_10_i_qa_d, xt_rsc_4_11_i_qa_d,
      xt_rsc_4_12_i_qa_d, xt_rsc_4_13_i_qa_d, xt_rsc_4_14_i_qa_d, xt_rsc_4_15_i_qa_d,
      xt_rsc_4_16_i_qa_d, xt_rsc_4_17_i_qa_d, xt_rsc_4_18_i_qa_d, xt_rsc_4_19_i_qa_d,
      xt_rsc_4_20_i_qa_d, xt_rsc_4_21_i_qa_d, xt_rsc_4_22_i_qa_d, xt_rsc_4_23_i_qa_d,
      xt_rsc_4_24_i_qa_d, xt_rsc_4_25_i_qa_d, xt_rsc_4_26_i_qa_d, xt_rsc_4_27_i_qa_d,
      xt_rsc_4_28_i_qa_d, xt_rsc_4_29_i_qa_d, xt_rsc_4_30_i_qa_d, xt_rsc_4_31_i_qa_d,
      xt_rsc_5_0_i_qa_d, xt_rsc_5_1_i_qa_d, xt_rsc_5_2_i_qa_d, xt_rsc_5_3_i_qa_d,
      xt_rsc_5_4_i_qa_d, xt_rsc_5_5_i_qa_d, xt_rsc_5_6_i_qa_d, xt_rsc_5_7_i_qa_d,
      xt_rsc_5_8_i_qa_d, xt_rsc_5_9_i_qa_d, xt_rsc_5_10_i_qa_d, xt_rsc_5_11_i_qa_d,
      xt_rsc_5_12_i_qa_d, xt_rsc_5_13_i_qa_d, xt_rsc_5_14_i_qa_d, xt_rsc_5_15_i_qa_d,
      xt_rsc_5_16_i_qa_d, xt_rsc_5_17_i_qa_d, xt_rsc_5_18_i_qa_d, xt_rsc_5_19_i_qa_d,
      xt_rsc_5_20_i_qa_d, xt_rsc_5_21_i_qa_d, xt_rsc_5_22_i_qa_d, xt_rsc_5_23_i_qa_d,
      xt_rsc_5_24_i_qa_d, xt_rsc_5_25_i_qa_d, xt_rsc_5_26_i_qa_d, xt_rsc_5_27_i_qa_d,
      xt_rsc_5_28_i_qa_d, xt_rsc_5_29_i_qa_d, xt_rsc_5_30_i_qa_d, xt_rsc_5_31_i_qa_d,
      xt_rsc_6_0_i_qa_d, xt_rsc_6_1_i_qa_d, xt_rsc_6_2_i_qa_d, xt_rsc_6_3_i_qa_d,
      xt_rsc_6_4_i_qa_d, xt_rsc_6_5_i_qa_d, xt_rsc_6_6_i_qa_d, xt_rsc_6_7_i_qa_d,
      xt_rsc_6_8_i_qa_d, xt_rsc_6_9_i_qa_d, xt_rsc_6_10_i_qa_d, xt_rsc_6_11_i_qa_d,
      xt_rsc_6_12_i_qa_d, xt_rsc_6_13_i_qa_d, xt_rsc_6_14_i_qa_d, xt_rsc_6_15_i_qa_d,
      xt_rsc_6_16_i_qa_d, xt_rsc_6_17_i_qa_d, xt_rsc_6_18_i_qa_d, xt_rsc_6_19_i_qa_d,
      xt_rsc_6_20_i_qa_d, xt_rsc_6_21_i_qa_d, xt_rsc_6_22_i_qa_d, xt_rsc_6_23_i_qa_d,
      xt_rsc_6_24_i_qa_d, xt_rsc_6_25_i_qa_d, xt_rsc_6_26_i_qa_d, xt_rsc_6_27_i_qa_d,
      xt_rsc_6_28_i_qa_d, xt_rsc_6_29_i_qa_d, xt_rsc_6_30_i_qa_d, xt_rsc_6_31_i_qa_d,
      xt_rsc_7_0_i_qa_d, xt_rsc_7_1_i_qa_d, xt_rsc_7_2_i_qa_d, xt_rsc_7_3_i_qa_d,
      xt_rsc_7_4_i_qa_d, xt_rsc_7_5_i_qa_d, xt_rsc_7_6_i_qa_d, xt_rsc_7_7_i_qa_d,
      xt_rsc_7_8_i_qa_d, xt_rsc_7_9_i_qa_d, xt_rsc_7_10_i_qa_d, xt_rsc_7_11_i_qa_d,
      xt_rsc_7_12_i_qa_d, xt_rsc_7_13_i_qa_d, xt_rsc_7_14_i_qa_d, xt_rsc_7_15_i_qa_d,
      xt_rsc_7_16_i_qa_d, xt_rsc_7_17_i_qa_d, xt_rsc_7_18_i_qa_d, xt_rsc_7_19_i_qa_d,
      xt_rsc_7_20_i_qa_d, xt_rsc_7_21_i_qa_d, xt_rsc_7_22_i_qa_d, xt_rsc_7_23_i_qa_d,
      xt_rsc_7_24_i_qa_d, xt_rsc_7_25_i_qa_d, xt_rsc_7_26_i_qa_d, xt_rsc_7_27_i_qa_d,
      xt_rsc_7_28_i_qa_d, xt_rsc_7_29_i_qa_d, xt_rsc_7_30_i_qa_d, xt_rsc_7_31_i_qa_d,
      twiddle_rsc_0_0_i_adra_d, twiddle_rsc_0_0_i_qa_d, twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_adra_d, twiddle_rsc_0_1_i_qa_d, twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_adra_d, twiddle_rsc_0_2_i_qa_d, twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_adra_d, twiddle_rsc_0_3_i_qa_d, twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_adra_d, twiddle_rsc_0_4_i_qa_d, twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_adra_d, twiddle_rsc_0_5_i_qa_d, twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_adra_d, twiddle_rsc_0_6_i_qa_d, twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_adra_d, twiddle_rsc_0_7_i_qa_d, twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_adra_d, twiddle_rsc_0_8_i_qa_d, twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_adra_d, twiddle_rsc_0_9_i_qa_d, twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_adra_d, twiddle_rsc_0_10_i_qa_d, twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_adra_d, twiddle_rsc_0_11_i_qa_d, twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_adra_d, twiddle_rsc_0_12_i_qa_d, twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_adra_d, twiddle_rsc_0_13_i_qa_d, twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_adra_d, twiddle_rsc_0_14_i_qa_d, twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_adra_d, twiddle_rsc_0_15_i_qa_d, twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_0_i_adra_d, twiddle_h_rsc_0_0_i_qa_d, twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_1_i_adra_d, twiddle_h_rsc_0_1_i_qa_d, twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_2_i_adra_d, twiddle_h_rsc_0_2_i_qa_d, twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_3_i_adra_d, twiddle_h_rsc_0_3_i_qa_d, twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_4_i_adra_d, twiddle_h_rsc_0_4_i_qa_d, twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_5_i_adra_d, twiddle_h_rsc_0_5_i_qa_d, twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_6_i_adra_d, twiddle_h_rsc_0_6_i_qa_d, twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_7_i_adra_d, twiddle_h_rsc_0_7_i_qa_d, twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_8_i_adra_d, twiddle_h_rsc_0_8_i_qa_d, twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_9_i_adra_d, twiddle_h_rsc_0_9_i_qa_d, twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_10_i_adra_d, twiddle_h_rsc_0_10_i_qa_d, twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_11_i_adra_d, twiddle_h_rsc_0_11_i_qa_d, twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_12_i_adra_d, twiddle_h_rsc_0_12_i_qa_d, twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_13_i_adra_d, twiddle_h_rsc_0_13_i_qa_d, twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_14_i_adra_d, twiddle_h_rsc_0_14_i_qa_d, twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_15_i_adra_d, twiddle_h_rsc_0_15_i_qa_d, twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_0_i_d_d_pff, yt_rsc_0_0_i_radr_d_pff, yt_rsc_0_0_i_wadr_d_pff, yt_rsc_0_0_i_we_d_pff,
      yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff, yt_rsc_0_1_i_d_d_pff, yt_rsc_0_1_i_wadr_d_pff,
      yt_rsc_0_2_i_d_d_pff, yt_rsc_0_2_i_wadr_d_pff, yt_rsc_0_3_i_d_d_pff, yt_rsc_0_3_i_wadr_d_pff,
      yt_rsc_0_4_i_d_d_pff, yt_rsc_0_4_i_wadr_d_pff, yt_rsc_0_5_i_d_d_pff, yt_rsc_0_5_i_wadr_d_pff,
      yt_rsc_0_6_i_d_d_pff, yt_rsc_0_6_i_wadr_d_pff, yt_rsc_0_7_i_d_d_pff, yt_rsc_0_8_i_d_d_pff,
      yt_rsc_0_9_i_d_d_pff, yt_rsc_0_10_i_d_d_pff, yt_rsc_0_10_i_wadr_d_pff, yt_rsc_0_11_i_d_d_pff,
      yt_rsc_0_11_i_wadr_d_pff, yt_rsc_0_12_i_d_d_pff, yt_rsc_0_13_i_d_d_pff, yt_rsc_0_14_i_d_d_pff,
      yt_rsc_0_15_i_d_d_pff, yt_rsc_0_16_i_we_d_pff, yt_rsc_1_0_i_we_d_pff, yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff,
      yt_rsc_1_16_i_we_d_pff, yt_rsc_2_0_i_we_d_pff, yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff,
      yt_rsc_2_16_i_we_d_pff, yt_rsc_3_0_i_we_d_pff, yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff,
      yt_rsc_3_16_i_we_d_pff, yt_rsc_4_0_i_d_d_pff, yt_rsc_4_0_i_wadr_d_pff, yt_rsc_4_0_i_we_d_pff,
      yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff, yt_rsc_4_1_i_d_d_pff, yt_rsc_4_1_i_wadr_d_pff,
      yt_rsc_4_2_i_d_d_pff, yt_rsc_4_2_i_wadr_d_pff, yt_rsc_4_3_i_d_d_pff, yt_rsc_4_3_i_wadr_d_pff,
      yt_rsc_4_4_i_d_d_pff, yt_rsc_4_4_i_wadr_d_pff, yt_rsc_4_5_i_d_d_pff, yt_rsc_4_5_i_wadr_d_pff,
      yt_rsc_4_6_i_d_d_pff, yt_rsc_4_6_i_wadr_d_pff, yt_rsc_4_7_i_d_d_pff, yt_rsc_4_8_i_d_d_pff,
      yt_rsc_4_9_i_d_d_pff, yt_rsc_4_9_i_wadr_d_pff, yt_rsc_4_10_i_d_d_pff, yt_rsc_4_10_i_wadr_d_pff,
      yt_rsc_4_11_i_d_d_pff, yt_rsc_4_11_i_wadr_d_pff, yt_rsc_4_12_i_d_d_pff, yt_rsc_4_13_i_d_d_pff,
      yt_rsc_4_14_i_d_d_pff, yt_rsc_4_15_i_d_d_pff, yt_rsc_4_16_i_we_d_pff, yt_rsc_5_0_i_we_d_pff,
      yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff, yt_rsc_5_16_i_we_d_pff,
      yt_rsc_6_0_i_we_d_pff, yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff,
      yt_rsc_6_16_i_we_d_pff, yt_rsc_7_0_i_we_d_pff, yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff,
      yt_rsc_7_16_i_we_d_pff, xt_rsc_0_0_i_adra_d_pff, xt_rsc_0_0_i_da_d_pff, xt_rsc_0_0_i_wea_d_pff,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff, xt_rsc_0_1_i_adra_d_pff,
      xt_rsc_0_1_i_da_d_pff, xt_rsc_0_2_i_adra_d_pff, xt_rsc_0_2_i_da_d_pff, xt_rsc_0_3_i_adra_d_pff,
      xt_rsc_0_3_i_da_d_pff, xt_rsc_0_4_i_adra_d_pff, xt_rsc_0_4_i_da_d_pff, xt_rsc_0_5_i_adra_d_pff,
      xt_rsc_0_5_i_da_d_pff, xt_rsc_0_6_i_adra_d_pff, xt_rsc_0_6_i_da_d_pff, xt_rsc_0_7_i_adra_d_pff,
      xt_rsc_0_7_i_da_d_pff, xt_rsc_0_8_i_adra_d_pff, xt_rsc_0_8_i_da_d_pff, xt_rsc_0_9_i_adra_d_pff,
      xt_rsc_0_9_i_da_d_pff, xt_rsc_0_10_i_adra_d_pff, xt_rsc_0_10_i_da_d_pff, xt_rsc_0_11_i_adra_d_pff,
      xt_rsc_0_11_i_da_d_pff, xt_rsc_0_12_i_adra_d_pff, xt_rsc_0_12_i_da_d_pff, xt_rsc_0_13_i_adra_d_pff,
      xt_rsc_0_13_i_da_d_pff, xt_rsc_0_14_i_adra_d_pff, xt_rsc_0_14_i_da_d_pff, xt_rsc_0_15_i_adra_d_pff,
      xt_rsc_0_15_i_da_d_pff, xt_rsc_0_16_i_wea_d_pff, xt_rsc_1_0_i_wea_d_pff, xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff,
      xt_rsc_1_16_i_wea_d_pff, xt_rsc_2_0_i_wea_d_pff, xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff,
      xt_rsc_2_16_i_wea_d_pff, xt_rsc_3_0_i_wea_d_pff, xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff,
      xt_rsc_3_16_i_wea_d_pff, xt_rsc_4_0_i_da_d_pff, xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff,
      xt_rsc_4_1_i_adra_d_pff, xt_rsc_4_1_i_da_d_pff, xt_rsc_4_2_i_adra_d_pff, xt_rsc_4_2_i_da_d_pff,
      xt_rsc_4_3_i_da_d_pff, xt_rsc_4_4_i_da_d_pff, xt_rsc_4_5_i_da_d_pff, xt_rsc_4_6_i_da_d_pff,
      xt_rsc_4_7_i_da_d_pff, xt_rsc_4_8_i_da_d_pff, xt_rsc_4_9_i_adra_d_pff, xt_rsc_4_9_i_da_d_pff,
      xt_rsc_4_10_i_adra_d_pff, xt_rsc_4_10_i_da_d_pff, xt_rsc_4_11_i_da_d_pff, xt_rsc_4_12_i_da_d_pff,
      xt_rsc_4_13_i_da_d_pff, xt_rsc_4_14_i_da_d_pff, xt_rsc_4_15_i_da_d_pff, xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff,
      xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff, xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff
);
  input clk;
  input rst;
  output xt_rsc_triosy_0_0_lz;
  output xt_rsc_triosy_0_1_lz;
  output xt_rsc_triosy_0_2_lz;
  output xt_rsc_triosy_0_3_lz;
  output xt_rsc_triosy_0_4_lz;
  output xt_rsc_triosy_0_5_lz;
  output xt_rsc_triosy_0_6_lz;
  output xt_rsc_triosy_0_7_lz;
  output xt_rsc_triosy_0_8_lz;
  output xt_rsc_triosy_0_9_lz;
  output xt_rsc_triosy_0_10_lz;
  output xt_rsc_triosy_0_11_lz;
  output xt_rsc_triosy_0_12_lz;
  output xt_rsc_triosy_0_13_lz;
  output xt_rsc_triosy_0_14_lz;
  output xt_rsc_triosy_0_15_lz;
  output xt_rsc_triosy_0_16_lz;
  output xt_rsc_triosy_0_17_lz;
  output xt_rsc_triosy_0_18_lz;
  output xt_rsc_triosy_0_19_lz;
  output xt_rsc_triosy_0_20_lz;
  output xt_rsc_triosy_0_21_lz;
  output xt_rsc_triosy_0_22_lz;
  output xt_rsc_triosy_0_23_lz;
  output xt_rsc_triosy_0_24_lz;
  output xt_rsc_triosy_0_25_lz;
  output xt_rsc_triosy_0_26_lz;
  output xt_rsc_triosy_0_27_lz;
  output xt_rsc_triosy_0_28_lz;
  output xt_rsc_triosy_0_29_lz;
  output xt_rsc_triosy_0_30_lz;
  output xt_rsc_triosy_0_31_lz;
  output xt_rsc_triosy_1_0_lz;
  output xt_rsc_triosy_1_1_lz;
  output xt_rsc_triosy_1_2_lz;
  output xt_rsc_triosy_1_3_lz;
  output xt_rsc_triosy_1_4_lz;
  output xt_rsc_triosy_1_5_lz;
  output xt_rsc_triosy_1_6_lz;
  output xt_rsc_triosy_1_7_lz;
  output xt_rsc_triosy_1_8_lz;
  output xt_rsc_triosy_1_9_lz;
  output xt_rsc_triosy_1_10_lz;
  output xt_rsc_triosy_1_11_lz;
  output xt_rsc_triosy_1_12_lz;
  output xt_rsc_triosy_1_13_lz;
  output xt_rsc_triosy_1_14_lz;
  output xt_rsc_triosy_1_15_lz;
  output xt_rsc_triosy_1_16_lz;
  output xt_rsc_triosy_1_17_lz;
  output xt_rsc_triosy_1_18_lz;
  output xt_rsc_triosy_1_19_lz;
  output xt_rsc_triosy_1_20_lz;
  output xt_rsc_triosy_1_21_lz;
  output xt_rsc_triosy_1_22_lz;
  output xt_rsc_triosy_1_23_lz;
  output xt_rsc_triosy_1_24_lz;
  output xt_rsc_triosy_1_25_lz;
  output xt_rsc_triosy_1_26_lz;
  output xt_rsc_triosy_1_27_lz;
  output xt_rsc_triosy_1_28_lz;
  output xt_rsc_triosy_1_29_lz;
  output xt_rsc_triosy_1_30_lz;
  output xt_rsc_triosy_1_31_lz;
  output xt_rsc_triosy_2_0_lz;
  output xt_rsc_triosy_2_1_lz;
  output xt_rsc_triosy_2_2_lz;
  output xt_rsc_triosy_2_3_lz;
  output xt_rsc_triosy_2_4_lz;
  output xt_rsc_triosy_2_5_lz;
  output xt_rsc_triosy_2_6_lz;
  output xt_rsc_triosy_2_7_lz;
  output xt_rsc_triosy_2_8_lz;
  output xt_rsc_triosy_2_9_lz;
  output xt_rsc_triosy_2_10_lz;
  output xt_rsc_triosy_2_11_lz;
  output xt_rsc_triosy_2_12_lz;
  output xt_rsc_triosy_2_13_lz;
  output xt_rsc_triosy_2_14_lz;
  output xt_rsc_triosy_2_15_lz;
  output xt_rsc_triosy_2_16_lz;
  output xt_rsc_triosy_2_17_lz;
  output xt_rsc_triosy_2_18_lz;
  output xt_rsc_triosy_2_19_lz;
  output xt_rsc_triosy_2_20_lz;
  output xt_rsc_triosy_2_21_lz;
  output xt_rsc_triosy_2_22_lz;
  output xt_rsc_triosy_2_23_lz;
  output xt_rsc_triosy_2_24_lz;
  output xt_rsc_triosy_2_25_lz;
  output xt_rsc_triosy_2_26_lz;
  output xt_rsc_triosy_2_27_lz;
  output xt_rsc_triosy_2_28_lz;
  output xt_rsc_triosy_2_29_lz;
  output xt_rsc_triosy_2_30_lz;
  output xt_rsc_triosy_2_31_lz;
  output xt_rsc_triosy_3_0_lz;
  output xt_rsc_triosy_3_1_lz;
  output xt_rsc_triosy_3_2_lz;
  output xt_rsc_triosy_3_3_lz;
  output xt_rsc_triosy_3_4_lz;
  output xt_rsc_triosy_3_5_lz;
  output xt_rsc_triosy_3_6_lz;
  output xt_rsc_triosy_3_7_lz;
  output xt_rsc_triosy_3_8_lz;
  output xt_rsc_triosy_3_9_lz;
  output xt_rsc_triosy_3_10_lz;
  output xt_rsc_triosy_3_11_lz;
  output xt_rsc_triosy_3_12_lz;
  output xt_rsc_triosy_3_13_lz;
  output xt_rsc_triosy_3_14_lz;
  output xt_rsc_triosy_3_15_lz;
  output xt_rsc_triosy_3_16_lz;
  output xt_rsc_triosy_3_17_lz;
  output xt_rsc_triosy_3_18_lz;
  output xt_rsc_triosy_3_19_lz;
  output xt_rsc_triosy_3_20_lz;
  output xt_rsc_triosy_3_21_lz;
  output xt_rsc_triosy_3_22_lz;
  output xt_rsc_triosy_3_23_lz;
  output xt_rsc_triosy_3_24_lz;
  output xt_rsc_triosy_3_25_lz;
  output xt_rsc_triosy_3_26_lz;
  output xt_rsc_triosy_3_27_lz;
  output xt_rsc_triosy_3_28_lz;
  output xt_rsc_triosy_3_29_lz;
  output xt_rsc_triosy_3_30_lz;
  output xt_rsc_triosy_3_31_lz;
  output xt_rsc_triosy_4_0_lz;
  output xt_rsc_triosy_4_1_lz;
  output xt_rsc_triosy_4_2_lz;
  output xt_rsc_triosy_4_3_lz;
  output xt_rsc_triosy_4_4_lz;
  output xt_rsc_triosy_4_5_lz;
  output xt_rsc_triosy_4_6_lz;
  output xt_rsc_triosy_4_7_lz;
  output xt_rsc_triosy_4_8_lz;
  output xt_rsc_triosy_4_9_lz;
  output xt_rsc_triosy_4_10_lz;
  output xt_rsc_triosy_4_11_lz;
  output xt_rsc_triosy_4_12_lz;
  output xt_rsc_triosy_4_13_lz;
  output xt_rsc_triosy_4_14_lz;
  output xt_rsc_triosy_4_15_lz;
  output xt_rsc_triosy_4_16_lz;
  output xt_rsc_triosy_4_17_lz;
  output xt_rsc_triosy_4_18_lz;
  output xt_rsc_triosy_4_19_lz;
  output xt_rsc_triosy_4_20_lz;
  output xt_rsc_triosy_4_21_lz;
  output xt_rsc_triosy_4_22_lz;
  output xt_rsc_triosy_4_23_lz;
  output xt_rsc_triosy_4_24_lz;
  output xt_rsc_triosy_4_25_lz;
  output xt_rsc_triosy_4_26_lz;
  output xt_rsc_triosy_4_27_lz;
  output xt_rsc_triosy_4_28_lz;
  output xt_rsc_triosy_4_29_lz;
  output xt_rsc_triosy_4_30_lz;
  output xt_rsc_triosy_4_31_lz;
  output xt_rsc_triosy_5_0_lz;
  output xt_rsc_triosy_5_1_lz;
  output xt_rsc_triosy_5_2_lz;
  output xt_rsc_triosy_5_3_lz;
  output xt_rsc_triosy_5_4_lz;
  output xt_rsc_triosy_5_5_lz;
  output xt_rsc_triosy_5_6_lz;
  output xt_rsc_triosy_5_7_lz;
  output xt_rsc_triosy_5_8_lz;
  output xt_rsc_triosy_5_9_lz;
  output xt_rsc_triosy_5_10_lz;
  output xt_rsc_triosy_5_11_lz;
  output xt_rsc_triosy_5_12_lz;
  output xt_rsc_triosy_5_13_lz;
  output xt_rsc_triosy_5_14_lz;
  output xt_rsc_triosy_5_15_lz;
  output xt_rsc_triosy_5_16_lz;
  output xt_rsc_triosy_5_17_lz;
  output xt_rsc_triosy_5_18_lz;
  output xt_rsc_triosy_5_19_lz;
  output xt_rsc_triosy_5_20_lz;
  output xt_rsc_triosy_5_21_lz;
  output xt_rsc_triosy_5_22_lz;
  output xt_rsc_triosy_5_23_lz;
  output xt_rsc_triosy_5_24_lz;
  output xt_rsc_triosy_5_25_lz;
  output xt_rsc_triosy_5_26_lz;
  output xt_rsc_triosy_5_27_lz;
  output xt_rsc_triosy_5_28_lz;
  output xt_rsc_triosy_5_29_lz;
  output xt_rsc_triosy_5_30_lz;
  output xt_rsc_triosy_5_31_lz;
  output xt_rsc_triosy_6_0_lz;
  output xt_rsc_triosy_6_1_lz;
  output xt_rsc_triosy_6_2_lz;
  output xt_rsc_triosy_6_3_lz;
  output xt_rsc_triosy_6_4_lz;
  output xt_rsc_triosy_6_5_lz;
  output xt_rsc_triosy_6_6_lz;
  output xt_rsc_triosy_6_7_lz;
  output xt_rsc_triosy_6_8_lz;
  output xt_rsc_triosy_6_9_lz;
  output xt_rsc_triosy_6_10_lz;
  output xt_rsc_triosy_6_11_lz;
  output xt_rsc_triosy_6_12_lz;
  output xt_rsc_triosy_6_13_lz;
  output xt_rsc_triosy_6_14_lz;
  output xt_rsc_triosy_6_15_lz;
  output xt_rsc_triosy_6_16_lz;
  output xt_rsc_triosy_6_17_lz;
  output xt_rsc_triosy_6_18_lz;
  output xt_rsc_triosy_6_19_lz;
  output xt_rsc_triosy_6_20_lz;
  output xt_rsc_triosy_6_21_lz;
  output xt_rsc_triosy_6_22_lz;
  output xt_rsc_triosy_6_23_lz;
  output xt_rsc_triosy_6_24_lz;
  output xt_rsc_triosy_6_25_lz;
  output xt_rsc_triosy_6_26_lz;
  output xt_rsc_triosy_6_27_lz;
  output xt_rsc_triosy_6_28_lz;
  output xt_rsc_triosy_6_29_lz;
  output xt_rsc_triosy_6_30_lz;
  output xt_rsc_triosy_6_31_lz;
  output xt_rsc_triosy_7_0_lz;
  output xt_rsc_triosy_7_1_lz;
  output xt_rsc_triosy_7_2_lz;
  output xt_rsc_triosy_7_3_lz;
  output xt_rsc_triosy_7_4_lz;
  output xt_rsc_triosy_7_5_lz;
  output xt_rsc_triosy_7_6_lz;
  output xt_rsc_triosy_7_7_lz;
  output xt_rsc_triosy_7_8_lz;
  output xt_rsc_triosy_7_9_lz;
  output xt_rsc_triosy_7_10_lz;
  output xt_rsc_triosy_7_11_lz;
  output xt_rsc_triosy_7_12_lz;
  output xt_rsc_triosy_7_13_lz;
  output xt_rsc_triosy_7_14_lz;
  output xt_rsc_triosy_7_15_lz;
  output xt_rsc_triosy_7_16_lz;
  output xt_rsc_triosy_7_17_lz;
  output xt_rsc_triosy_7_18_lz;
  output xt_rsc_triosy_7_19_lz;
  output xt_rsc_triosy_7_20_lz;
  output xt_rsc_triosy_7_21_lz;
  output xt_rsc_triosy_7_22_lz;
  output xt_rsc_triosy_7_23_lz;
  output xt_rsc_triosy_7_24_lz;
  output xt_rsc_triosy_7_25_lz;
  output xt_rsc_triosy_7_26_lz;
  output xt_rsc_triosy_7_27_lz;
  output xt_rsc_triosy_7_28_lz;
  output xt_rsc_triosy_7_29_lz;
  output xt_rsc_triosy_7_30_lz;
  output xt_rsc_triosy_7_31_lz;
  input [31:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_0_0_lz;
  output twiddle_rsc_triosy_0_1_lz;
  output twiddle_rsc_triosy_0_2_lz;
  output twiddle_rsc_triosy_0_3_lz;
  output twiddle_rsc_triosy_0_4_lz;
  output twiddle_rsc_triosy_0_5_lz;
  output twiddle_rsc_triosy_0_6_lz;
  output twiddle_rsc_triosy_0_7_lz;
  output twiddle_rsc_triosy_0_8_lz;
  output twiddle_rsc_triosy_0_9_lz;
  output twiddle_rsc_triosy_0_10_lz;
  output twiddle_rsc_triosy_0_11_lz;
  output twiddle_rsc_triosy_0_12_lz;
  output twiddle_rsc_triosy_0_13_lz;
  output twiddle_rsc_triosy_0_14_lz;
  output twiddle_rsc_triosy_0_15_lz;
  output twiddle_h_rsc_triosy_0_0_lz;
  output twiddle_h_rsc_triosy_0_1_lz;
  output twiddle_h_rsc_triosy_0_2_lz;
  output twiddle_h_rsc_triosy_0_3_lz;
  output twiddle_h_rsc_triosy_0_4_lz;
  output twiddle_h_rsc_triosy_0_5_lz;
  output twiddle_h_rsc_triosy_0_6_lz;
  output twiddle_h_rsc_triosy_0_7_lz;
  output twiddle_h_rsc_triosy_0_8_lz;
  output twiddle_h_rsc_triosy_0_9_lz;
  output twiddle_h_rsc_triosy_0_10_lz;
  output twiddle_h_rsc_triosy_0_11_lz;
  output twiddle_h_rsc_triosy_0_12_lz;
  output twiddle_h_rsc_triosy_0_13_lz;
  output twiddle_h_rsc_triosy_0_14_lz;
  output twiddle_h_rsc_triosy_0_15_lz;
  output yt_rsc_0_0_i_clkr_en_d;
  input [31:0] yt_rsc_0_0_i_q_d;
  input [31:0] yt_rsc_0_1_i_q_d;
  input [31:0] yt_rsc_0_2_i_q_d;
  input [31:0] yt_rsc_0_3_i_q_d;
  input [31:0] yt_rsc_0_4_i_q_d;
  input [31:0] yt_rsc_0_5_i_q_d;
  input [31:0] yt_rsc_0_6_i_q_d;
  input [31:0] yt_rsc_0_7_i_q_d;
  input [31:0] yt_rsc_0_8_i_q_d;
  input [31:0] yt_rsc_0_9_i_q_d;
  input [31:0] yt_rsc_0_10_i_q_d;
  input [31:0] yt_rsc_0_11_i_q_d;
  input [31:0] yt_rsc_0_12_i_q_d;
  input [31:0] yt_rsc_0_13_i_q_d;
  input [31:0] yt_rsc_0_14_i_q_d;
  input [31:0] yt_rsc_0_15_i_q_d;
  output yt_rsc_0_16_i_clkr_en_d;
  input [31:0] yt_rsc_0_16_i_q_d;
  input [31:0] yt_rsc_0_17_i_q_d;
  input [31:0] yt_rsc_0_18_i_q_d;
  input [31:0] yt_rsc_0_19_i_q_d;
  input [31:0] yt_rsc_0_20_i_q_d;
  input [31:0] yt_rsc_0_21_i_q_d;
  input [31:0] yt_rsc_0_22_i_q_d;
  input [31:0] yt_rsc_0_23_i_q_d;
  input [31:0] yt_rsc_0_24_i_q_d;
  input [31:0] yt_rsc_0_25_i_q_d;
  input [31:0] yt_rsc_0_26_i_q_d;
  input [31:0] yt_rsc_0_27_i_q_d;
  input [31:0] yt_rsc_0_28_i_q_d;
  input [31:0] yt_rsc_0_29_i_q_d;
  input [31:0] yt_rsc_0_30_i_q_d;
  input [31:0] yt_rsc_0_31_i_q_d;
  output yt_rsc_1_0_i_clkr_en_d;
  input [31:0] yt_rsc_1_0_i_q_d;
  input [31:0] yt_rsc_1_1_i_q_d;
  input [31:0] yt_rsc_1_2_i_q_d;
  input [31:0] yt_rsc_1_3_i_q_d;
  input [31:0] yt_rsc_1_4_i_q_d;
  input [31:0] yt_rsc_1_5_i_q_d;
  input [31:0] yt_rsc_1_6_i_q_d;
  input [31:0] yt_rsc_1_7_i_q_d;
  input [31:0] yt_rsc_1_8_i_q_d;
  input [31:0] yt_rsc_1_9_i_q_d;
  input [31:0] yt_rsc_1_10_i_q_d;
  input [31:0] yt_rsc_1_11_i_q_d;
  input [31:0] yt_rsc_1_12_i_q_d;
  input [31:0] yt_rsc_1_13_i_q_d;
  input [31:0] yt_rsc_1_14_i_q_d;
  input [31:0] yt_rsc_1_15_i_q_d;
  output yt_rsc_1_16_i_clkr_en_d;
  input [31:0] yt_rsc_1_16_i_q_d;
  input [31:0] yt_rsc_1_17_i_q_d;
  input [31:0] yt_rsc_1_18_i_q_d;
  input [31:0] yt_rsc_1_19_i_q_d;
  input [31:0] yt_rsc_1_20_i_q_d;
  input [31:0] yt_rsc_1_21_i_q_d;
  input [31:0] yt_rsc_1_22_i_q_d;
  input [31:0] yt_rsc_1_23_i_q_d;
  input [31:0] yt_rsc_1_24_i_q_d;
  input [31:0] yt_rsc_1_25_i_q_d;
  input [31:0] yt_rsc_1_26_i_q_d;
  input [31:0] yt_rsc_1_27_i_q_d;
  input [31:0] yt_rsc_1_28_i_q_d;
  input [31:0] yt_rsc_1_29_i_q_d;
  input [31:0] yt_rsc_1_30_i_q_d;
  input [31:0] yt_rsc_1_31_i_q_d;
  output yt_rsc_2_0_i_clkr_en_d;
  input [31:0] yt_rsc_2_0_i_q_d;
  input [31:0] yt_rsc_2_1_i_q_d;
  input [31:0] yt_rsc_2_2_i_q_d;
  input [31:0] yt_rsc_2_3_i_q_d;
  input [31:0] yt_rsc_2_4_i_q_d;
  input [31:0] yt_rsc_2_5_i_q_d;
  input [31:0] yt_rsc_2_6_i_q_d;
  input [31:0] yt_rsc_2_7_i_q_d;
  input [31:0] yt_rsc_2_8_i_q_d;
  input [31:0] yt_rsc_2_9_i_q_d;
  input [31:0] yt_rsc_2_10_i_q_d;
  input [31:0] yt_rsc_2_11_i_q_d;
  input [31:0] yt_rsc_2_12_i_q_d;
  input [31:0] yt_rsc_2_13_i_q_d;
  input [31:0] yt_rsc_2_14_i_q_d;
  input [31:0] yt_rsc_2_15_i_q_d;
  output yt_rsc_2_16_i_clkr_en_d;
  input [31:0] yt_rsc_2_16_i_q_d;
  input [31:0] yt_rsc_2_17_i_q_d;
  input [31:0] yt_rsc_2_18_i_q_d;
  input [31:0] yt_rsc_2_19_i_q_d;
  input [31:0] yt_rsc_2_20_i_q_d;
  input [31:0] yt_rsc_2_21_i_q_d;
  input [31:0] yt_rsc_2_22_i_q_d;
  input [31:0] yt_rsc_2_23_i_q_d;
  input [31:0] yt_rsc_2_24_i_q_d;
  input [31:0] yt_rsc_2_25_i_q_d;
  input [31:0] yt_rsc_2_26_i_q_d;
  input [31:0] yt_rsc_2_27_i_q_d;
  input [31:0] yt_rsc_2_28_i_q_d;
  input [31:0] yt_rsc_2_29_i_q_d;
  input [31:0] yt_rsc_2_30_i_q_d;
  input [31:0] yt_rsc_2_31_i_q_d;
  output yt_rsc_3_0_i_clkr_en_d;
  input [31:0] yt_rsc_3_0_i_q_d;
  input [31:0] yt_rsc_3_1_i_q_d;
  input [31:0] yt_rsc_3_2_i_q_d;
  input [31:0] yt_rsc_3_3_i_q_d;
  input [31:0] yt_rsc_3_4_i_q_d;
  input [31:0] yt_rsc_3_5_i_q_d;
  input [31:0] yt_rsc_3_6_i_q_d;
  input [31:0] yt_rsc_3_7_i_q_d;
  input [31:0] yt_rsc_3_8_i_q_d;
  input [31:0] yt_rsc_3_9_i_q_d;
  input [31:0] yt_rsc_3_10_i_q_d;
  input [31:0] yt_rsc_3_11_i_q_d;
  input [31:0] yt_rsc_3_12_i_q_d;
  input [31:0] yt_rsc_3_13_i_q_d;
  input [31:0] yt_rsc_3_14_i_q_d;
  input [31:0] yt_rsc_3_15_i_q_d;
  output yt_rsc_3_16_i_clkr_en_d;
  input [31:0] yt_rsc_3_16_i_q_d;
  input [31:0] yt_rsc_3_17_i_q_d;
  input [31:0] yt_rsc_3_18_i_q_d;
  input [31:0] yt_rsc_3_19_i_q_d;
  input [31:0] yt_rsc_3_20_i_q_d;
  input [31:0] yt_rsc_3_21_i_q_d;
  input [31:0] yt_rsc_3_22_i_q_d;
  input [31:0] yt_rsc_3_23_i_q_d;
  input [31:0] yt_rsc_3_24_i_q_d;
  input [31:0] yt_rsc_3_25_i_q_d;
  input [31:0] yt_rsc_3_26_i_q_d;
  input [31:0] yt_rsc_3_27_i_q_d;
  input [31:0] yt_rsc_3_28_i_q_d;
  input [31:0] yt_rsc_3_29_i_q_d;
  input [31:0] yt_rsc_3_30_i_q_d;
  input [31:0] yt_rsc_3_31_i_q_d;
  output yt_rsc_4_0_i_clkr_en_d;
  input [31:0] yt_rsc_4_0_i_q_d;
  input [31:0] yt_rsc_4_1_i_q_d;
  input [31:0] yt_rsc_4_2_i_q_d;
  input [31:0] yt_rsc_4_3_i_q_d;
  input [31:0] yt_rsc_4_4_i_q_d;
  input [31:0] yt_rsc_4_5_i_q_d;
  input [31:0] yt_rsc_4_6_i_q_d;
  input [31:0] yt_rsc_4_7_i_q_d;
  input [31:0] yt_rsc_4_8_i_q_d;
  input [31:0] yt_rsc_4_9_i_q_d;
  input [31:0] yt_rsc_4_10_i_q_d;
  input [31:0] yt_rsc_4_11_i_q_d;
  input [31:0] yt_rsc_4_12_i_q_d;
  input [31:0] yt_rsc_4_13_i_q_d;
  input [31:0] yt_rsc_4_14_i_q_d;
  input [31:0] yt_rsc_4_15_i_q_d;
  output yt_rsc_4_16_i_clkr_en_d;
  input [31:0] yt_rsc_4_16_i_q_d;
  input [31:0] yt_rsc_4_17_i_q_d;
  input [31:0] yt_rsc_4_18_i_q_d;
  input [31:0] yt_rsc_4_19_i_q_d;
  input [31:0] yt_rsc_4_20_i_q_d;
  input [31:0] yt_rsc_4_21_i_q_d;
  input [31:0] yt_rsc_4_22_i_q_d;
  input [31:0] yt_rsc_4_23_i_q_d;
  input [31:0] yt_rsc_4_24_i_q_d;
  input [31:0] yt_rsc_4_25_i_q_d;
  input [31:0] yt_rsc_4_26_i_q_d;
  input [31:0] yt_rsc_4_27_i_q_d;
  input [31:0] yt_rsc_4_28_i_q_d;
  input [31:0] yt_rsc_4_29_i_q_d;
  input [31:0] yt_rsc_4_30_i_q_d;
  input [31:0] yt_rsc_4_31_i_q_d;
  output yt_rsc_5_0_i_clkr_en_d;
  input [31:0] yt_rsc_5_0_i_q_d;
  input [31:0] yt_rsc_5_1_i_q_d;
  input [31:0] yt_rsc_5_2_i_q_d;
  input [31:0] yt_rsc_5_3_i_q_d;
  input [31:0] yt_rsc_5_4_i_q_d;
  input [31:0] yt_rsc_5_5_i_q_d;
  input [31:0] yt_rsc_5_6_i_q_d;
  input [31:0] yt_rsc_5_7_i_q_d;
  input [31:0] yt_rsc_5_8_i_q_d;
  input [31:0] yt_rsc_5_9_i_q_d;
  input [31:0] yt_rsc_5_10_i_q_d;
  input [31:0] yt_rsc_5_11_i_q_d;
  input [31:0] yt_rsc_5_12_i_q_d;
  input [31:0] yt_rsc_5_13_i_q_d;
  input [31:0] yt_rsc_5_14_i_q_d;
  input [31:0] yt_rsc_5_15_i_q_d;
  output yt_rsc_5_16_i_clkr_en_d;
  input [31:0] yt_rsc_5_16_i_q_d;
  input [31:0] yt_rsc_5_17_i_q_d;
  input [31:0] yt_rsc_5_18_i_q_d;
  input [31:0] yt_rsc_5_19_i_q_d;
  input [31:0] yt_rsc_5_20_i_q_d;
  input [31:0] yt_rsc_5_21_i_q_d;
  input [31:0] yt_rsc_5_22_i_q_d;
  input [31:0] yt_rsc_5_23_i_q_d;
  input [31:0] yt_rsc_5_24_i_q_d;
  input [31:0] yt_rsc_5_25_i_q_d;
  input [31:0] yt_rsc_5_26_i_q_d;
  input [31:0] yt_rsc_5_27_i_q_d;
  input [31:0] yt_rsc_5_28_i_q_d;
  input [31:0] yt_rsc_5_29_i_q_d;
  input [31:0] yt_rsc_5_30_i_q_d;
  input [31:0] yt_rsc_5_31_i_q_d;
  output yt_rsc_6_0_i_clkr_en_d;
  input [31:0] yt_rsc_6_0_i_q_d;
  input [31:0] yt_rsc_6_1_i_q_d;
  input [31:0] yt_rsc_6_2_i_q_d;
  input [31:0] yt_rsc_6_3_i_q_d;
  input [31:0] yt_rsc_6_4_i_q_d;
  input [31:0] yt_rsc_6_5_i_q_d;
  input [31:0] yt_rsc_6_6_i_q_d;
  input [31:0] yt_rsc_6_7_i_q_d;
  input [31:0] yt_rsc_6_8_i_q_d;
  input [31:0] yt_rsc_6_9_i_q_d;
  input [31:0] yt_rsc_6_10_i_q_d;
  input [31:0] yt_rsc_6_11_i_q_d;
  input [31:0] yt_rsc_6_12_i_q_d;
  input [31:0] yt_rsc_6_13_i_q_d;
  input [31:0] yt_rsc_6_14_i_q_d;
  input [31:0] yt_rsc_6_15_i_q_d;
  output yt_rsc_6_16_i_clkr_en_d;
  input [31:0] yt_rsc_6_16_i_q_d;
  input [31:0] yt_rsc_6_17_i_q_d;
  input [31:0] yt_rsc_6_18_i_q_d;
  input [31:0] yt_rsc_6_19_i_q_d;
  input [31:0] yt_rsc_6_20_i_q_d;
  input [31:0] yt_rsc_6_21_i_q_d;
  input [31:0] yt_rsc_6_22_i_q_d;
  input [31:0] yt_rsc_6_23_i_q_d;
  input [31:0] yt_rsc_6_24_i_q_d;
  input [31:0] yt_rsc_6_25_i_q_d;
  input [31:0] yt_rsc_6_26_i_q_d;
  input [31:0] yt_rsc_6_27_i_q_d;
  input [31:0] yt_rsc_6_28_i_q_d;
  input [31:0] yt_rsc_6_29_i_q_d;
  input [31:0] yt_rsc_6_30_i_q_d;
  input [31:0] yt_rsc_6_31_i_q_d;
  output yt_rsc_7_0_i_clkr_en_d;
  input [31:0] yt_rsc_7_0_i_q_d;
  input [31:0] yt_rsc_7_1_i_q_d;
  input [31:0] yt_rsc_7_2_i_q_d;
  input [31:0] yt_rsc_7_3_i_q_d;
  input [31:0] yt_rsc_7_4_i_q_d;
  input [31:0] yt_rsc_7_5_i_q_d;
  input [31:0] yt_rsc_7_6_i_q_d;
  input [31:0] yt_rsc_7_7_i_q_d;
  input [31:0] yt_rsc_7_8_i_q_d;
  input [31:0] yt_rsc_7_9_i_q_d;
  input [31:0] yt_rsc_7_10_i_q_d;
  input [31:0] yt_rsc_7_11_i_q_d;
  input [31:0] yt_rsc_7_12_i_q_d;
  input [31:0] yt_rsc_7_13_i_q_d;
  input [31:0] yt_rsc_7_14_i_q_d;
  input [31:0] yt_rsc_7_15_i_q_d;
  output yt_rsc_7_16_i_clkr_en_d;
  input [31:0] yt_rsc_7_16_i_q_d;
  input [31:0] yt_rsc_7_17_i_q_d;
  input [31:0] yt_rsc_7_18_i_q_d;
  input [31:0] yt_rsc_7_19_i_q_d;
  input [31:0] yt_rsc_7_20_i_q_d;
  input [31:0] yt_rsc_7_21_i_q_d;
  input [31:0] yt_rsc_7_22_i_q_d;
  input [31:0] yt_rsc_7_23_i_q_d;
  input [31:0] yt_rsc_7_24_i_q_d;
  input [31:0] yt_rsc_7_25_i_q_d;
  input [31:0] yt_rsc_7_26_i_q_d;
  input [31:0] yt_rsc_7_27_i_q_d;
  input [31:0] yt_rsc_7_28_i_q_d;
  input [31:0] yt_rsc_7_29_i_q_d;
  input [31:0] yt_rsc_7_30_i_q_d;
  input [31:0] yt_rsc_7_31_i_q_d;
  input [31:0] xt_rsc_0_0_i_qa_d;
  input [31:0] xt_rsc_0_1_i_qa_d;
  input [31:0] xt_rsc_0_2_i_qa_d;
  input [31:0] xt_rsc_0_3_i_qa_d;
  input [31:0] xt_rsc_0_4_i_qa_d;
  input [31:0] xt_rsc_0_5_i_qa_d;
  input [31:0] xt_rsc_0_6_i_qa_d;
  input [31:0] xt_rsc_0_7_i_qa_d;
  input [31:0] xt_rsc_0_8_i_qa_d;
  input [31:0] xt_rsc_0_9_i_qa_d;
  input [31:0] xt_rsc_0_10_i_qa_d;
  input [31:0] xt_rsc_0_11_i_qa_d;
  input [31:0] xt_rsc_0_12_i_qa_d;
  input [31:0] xt_rsc_0_13_i_qa_d;
  input [31:0] xt_rsc_0_14_i_qa_d;
  input [31:0] xt_rsc_0_15_i_qa_d;
  input [31:0] xt_rsc_0_16_i_qa_d;
  input [31:0] xt_rsc_0_17_i_qa_d;
  input [31:0] xt_rsc_0_18_i_qa_d;
  input [31:0] xt_rsc_0_19_i_qa_d;
  input [31:0] xt_rsc_0_20_i_qa_d;
  input [31:0] xt_rsc_0_21_i_qa_d;
  input [31:0] xt_rsc_0_22_i_qa_d;
  input [31:0] xt_rsc_0_23_i_qa_d;
  input [31:0] xt_rsc_0_24_i_qa_d;
  input [31:0] xt_rsc_0_25_i_qa_d;
  input [31:0] xt_rsc_0_26_i_qa_d;
  input [31:0] xt_rsc_0_27_i_qa_d;
  input [31:0] xt_rsc_0_28_i_qa_d;
  input [31:0] xt_rsc_0_29_i_qa_d;
  input [31:0] xt_rsc_0_30_i_qa_d;
  input [31:0] xt_rsc_0_31_i_qa_d;
  input [31:0] xt_rsc_1_0_i_qa_d;
  input [31:0] xt_rsc_1_1_i_qa_d;
  input [31:0] xt_rsc_1_2_i_qa_d;
  input [31:0] xt_rsc_1_3_i_qa_d;
  input [31:0] xt_rsc_1_4_i_qa_d;
  input [31:0] xt_rsc_1_5_i_qa_d;
  input [31:0] xt_rsc_1_6_i_qa_d;
  input [31:0] xt_rsc_1_7_i_qa_d;
  input [31:0] xt_rsc_1_8_i_qa_d;
  input [31:0] xt_rsc_1_9_i_qa_d;
  input [31:0] xt_rsc_1_10_i_qa_d;
  input [31:0] xt_rsc_1_11_i_qa_d;
  input [31:0] xt_rsc_1_12_i_qa_d;
  input [31:0] xt_rsc_1_13_i_qa_d;
  input [31:0] xt_rsc_1_14_i_qa_d;
  input [31:0] xt_rsc_1_15_i_qa_d;
  input [31:0] xt_rsc_1_16_i_qa_d;
  input [31:0] xt_rsc_1_17_i_qa_d;
  input [31:0] xt_rsc_1_18_i_qa_d;
  input [31:0] xt_rsc_1_19_i_qa_d;
  input [31:0] xt_rsc_1_20_i_qa_d;
  input [31:0] xt_rsc_1_21_i_qa_d;
  input [31:0] xt_rsc_1_22_i_qa_d;
  input [31:0] xt_rsc_1_23_i_qa_d;
  input [31:0] xt_rsc_1_24_i_qa_d;
  input [31:0] xt_rsc_1_25_i_qa_d;
  input [31:0] xt_rsc_1_26_i_qa_d;
  input [31:0] xt_rsc_1_27_i_qa_d;
  input [31:0] xt_rsc_1_28_i_qa_d;
  input [31:0] xt_rsc_1_29_i_qa_d;
  input [31:0] xt_rsc_1_30_i_qa_d;
  input [31:0] xt_rsc_1_31_i_qa_d;
  input [31:0] xt_rsc_2_0_i_qa_d;
  input [31:0] xt_rsc_2_1_i_qa_d;
  input [31:0] xt_rsc_2_2_i_qa_d;
  input [31:0] xt_rsc_2_3_i_qa_d;
  input [31:0] xt_rsc_2_4_i_qa_d;
  input [31:0] xt_rsc_2_5_i_qa_d;
  input [31:0] xt_rsc_2_6_i_qa_d;
  input [31:0] xt_rsc_2_7_i_qa_d;
  input [31:0] xt_rsc_2_8_i_qa_d;
  input [31:0] xt_rsc_2_9_i_qa_d;
  input [31:0] xt_rsc_2_10_i_qa_d;
  input [31:0] xt_rsc_2_11_i_qa_d;
  input [31:0] xt_rsc_2_12_i_qa_d;
  input [31:0] xt_rsc_2_13_i_qa_d;
  input [31:0] xt_rsc_2_14_i_qa_d;
  input [31:0] xt_rsc_2_15_i_qa_d;
  input [31:0] xt_rsc_2_16_i_qa_d;
  input [31:0] xt_rsc_2_17_i_qa_d;
  input [31:0] xt_rsc_2_18_i_qa_d;
  input [31:0] xt_rsc_2_19_i_qa_d;
  input [31:0] xt_rsc_2_20_i_qa_d;
  input [31:0] xt_rsc_2_21_i_qa_d;
  input [31:0] xt_rsc_2_22_i_qa_d;
  input [31:0] xt_rsc_2_23_i_qa_d;
  input [31:0] xt_rsc_2_24_i_qa_d;
  input [31:0] xt_rsc_2_25_i_qa_d;
  input [31:0] xt_rsc_2_26_i_qa_d;
  input [31:0] xt_rsc_2_27_i_qa_d;
  input [31:0] xt_rsc_2_28_i_qa_d;
  input [31:0] xt_rsc_2_29_i_qa_d;
  input [31:0] xt_rsc_2_30_i_qa_d;
  input [31:0] xt_rsc_2_31_i_qa_d;
  input [31:0] xt_rsc_3_0_i_qa_d;
  input [31:0] xt_rsc_3_1_i_qa_d;
  input [31:0] xt_rsc_3_2_i_qa_d;
  input [31:0] xt_rsc_3_3_i_qa_d;
  input [31:0] xt_rsc_3_4_i_qa_d;
  input [31:0] xt_rsc_3_5_i_qa_d;
  input [31:0] xt_rsc_3_6_i_qa_d;
  input [31:0] xt_rsc_3_7_i_qa_d;
  input [31:0] xt_rsc_3_8_i_qa_d;
  input [31:0] xt_rsc_3_9_i_qa_d;
  input [31:0] xt_rsc_3_10_i_qa_d;
  input [31:0] xt_rsc_3_11_i_qa_d;
  input [31:0] xt_rsc_3_12_i_qa_d;
  input [31:0] xt_rsc_3_13_i_qa_d;
  input [31:0] xt_rsc_3_14_i_qa_d;
  input [31:0] xt_rsc_3_15_i_qa_d;
  input [31:0] xt_rsc_3_16_i_qa_d;
  input [31:0] xt_rsc_3_17_i_qa_d;
  input [31:0] xt_rsc_3_18_i_qa_d;
  input [31:0] xt_rsc_3_19_i_qa_d;
  input [31:0] xt_rsc_3_20_i_qa_d;
  input [31:0] xt_rsc_3_21_i_qa_d;
  input [31:0] xt_rsc_3_22_i_qa_d;
  input [31:0] xt_rsc_3_23_i_qa_d;
  input [31:0] xt_rsc_3_24_i_qa_d;
  input [31:0] xt_rsc_3_25_i_qa_d;
  input [31:0] xt_rsc_3_26_i_qa_d;
  input [31:0] xt_rsc_3_27_i_qa_d;
  input [31:0] xt_rsc_3_28_i_qa_d;
  input [31:0] xt_rsc_3_29_i_qa_d;
  input [31:0] xt_rsc_3_30_i_qa_d;
  input [31:0] xt_rsc_3_31_i_qa_d;
  input [31:0] xt_rsc_4_0_i_qa_d;
  input [31:0] xt_rsc_4_1_i_qa_d;
  input [31:0] xt_rsc_4_2_i_qa_d;
  input [31:0] xt_rsc_4_3_i_qa_d;
  input [31:0] xt_rsc_4_4_i_qa_d;
  input [31:0] xt_rsc_4_5_i_qa_d;
  input [31:0] xt_rsc_4_6_i_qa_d;
  input [31:0] xt_rsc_4_7_i_qa_d;
  input [31:0] xt_rsc_4_8_i_qa_d;
  input [31:0] xt_rsc_4_9_i_qa_d;
  input [31:0] xt_rsc_4_10_i_qa_d;
  input [31:0] xt_rsc_4_11_i_qa_d;
  input [31:0] xt_rsc_4_12_i_qa_d;
  input [31:0] xt_rsc_4_13_i_qa_d;
  input [31:0] xt_rsc_4_14_i_qa_d;
  input [31:0] xt_rsc_4_15_i_qa_d;
  input [31:0] xt_rsc_4_16_i_qa_d;
  input [31:0] xt_rsc_4_17_i_qa_d;
  input [31:0] xt_rsc_4_18_i_qa_d;
  input [31:0] xt_rsc_4_19_i_qa_d;
  input [31:0] xt_rsc_4_20_i_qa_d;
  input [31:0] xt_rsc_4_21_i_qa_d;
  input [31:0] xt_rsc_4_22_i_qa_d;
  input [31:0] xt_rsc_4_23_i_qa_d;
  input [31:0] xt_rsc_4_24_i_qa_d;
  input [31:0] xt_rsc_4_25_i_qa_d;
  input [31:0] xt_rsc_4_26_i_qa_d;
  input [31:0] xt_rsc_4_27_i_qa_d;
  input [31:0] xt_rsc_4_28_i_qa_d;
  input [31:0] xt_rsc_4_29_i_qa_d;
  input [31:0] xt_rsc_4_30_i_qa_d;
  input [31:0] xt_rsc_4_31_i_qa_d;
  input [31:0] xt_rsc_5_0_i_qa_d;
  input [31:0] xt_rsc_5_1_i_qa_d;
  input [31:0] xt_rsc_5_2_i_qa_d;
  input [31:0] xt_rsc_5_3_i_qa_d;
  input [31:0] xt_rsc_5_4_i_qa_d;
  input [31:0] xt_rsc_5_5_i_qa_d;
  input [31:0] xt_rsc_5_6_i_qa_d;
  input [31:0] xt_rsc_5_7_i_qa_d;
  input [31:0] xt_rsc_5_8_i_qa_d;
  input [31:0] xt_rsc_5_9_i_qa_d;
  input [31:0] xt_rsc_5_10_i_qa_d;
  input [31:0] xt_rsc_5_11_i_qa_d;
  input [31:0] xt_rsc_5_12_i_qa_d;
  input [31:0] xt_rsc_5_13_i_qa_d;
  input [31:0] xt_rsc_5_14_i_qa_d;
  input [31:0] xt_rsc_5_15_i_qa_d;
  input [31:0] xt_rsc_5_16_i_qa_d;
  input [31:0] xt_rsc_5_17_i_qa_d;
  input [31:0] xt_rsc_5_18_i_qa_d;
  input [31:0] xt_rsc_5_19_i_qa_d;
  input [31:0] xt_rsc_5_20_i_qa_d;
  input [31:0] xt_rsc_5_21_i_qa_d;
  input [31:0] xt_rsc_5_22_i_qa_d;
  input [31:0] xt_rsc_5_23_i_qa_d;
  input [31:0] xt_rsc_5_24_i_qa_d;
  input [31:0] xt_rsc_5_25_i_qa_d;
  input [31:0] xt_rsc_5_26_i_qa_d;
  input [31:0] xt_rsc_5_27_i_qa_d;
  input [31:0] xt_rsc_5_28_i_qa_d;
  input [31:0] xt_rsc_5_29_i_qa_d;
  input [31:0] xt_rsc_5_30_i_qa_d;
  input [31:0] xt_rsc_5_31_i_qa_d;
  input [31:0] xt_rsc_6_0_i_qa_d;
  input [31:0] xt_rsc_6_1_i_qa_d;
  input [31:0] xt_rsc_6_2_i_qa_d;
  input [31:0] xt_rsc_6_3_i_qa_d;
  input [31:0] xt_rsc_6_4_i_qa_d;
  input [31:0] xt_rsc_6_5_i_qa_d;
  input [31:0] xt_rsc_6_6_i_qa_d;
  input [31:0] xt_rsc_6_7_i_qa_d;
  input [31:0] xt_rsc_6_8_i_qa_d;
  input [31:0] xt_rsc_6_9_i_qa_d;
  input [31:0] xt_rsc_6_10_i_qa_d;
  input [31:0] xt_rsc_6_11_i_qa_d;
  input [31:0] xt_rsc_6_12_i_qa_d;
  input [31:0] xt_rsc_6_13_i_qa_d;
  input [31:0] xt_rsc_6_14_i_qa_d;
  input [31:0] xt_rsc_6_15_i_qa_d;
  input [31:0] xt_rsc_6_16_i_qa_d;
  input [31:0] xt_rsc_6_17_i_qa_d;
  input [31:0] xt_rsc_6_18_i_qa_d;
  input [31:0] xt_rsc_6_19_i_qa_d;
  input [31:0] xt_rsc_6_20_i_qa_d;
  input [31:0] xt_rsc_6_21_i_qa_d;
  input [31:0] xt_rsc_6_22_i_qa_d;
  input [31:0] xt_rsc_6_23_i_qa_d;
  input [31:0] xt_rsc_6_24_i_qa_d;
  input [31:0] xt_rsc_6_25_i_qa_d;
  input [31:0] xt_rsc_6_26_i_qa_d;
  input [31:0] xt_rsc_6_27_i_qa_d;
  input [31:0] xt_rsc_6_28_i_qa_d;
  input [31:0] xt_rsc_6_29_i_qa_d;
  input [31:0] xt_rsc_6_30_i_qa_d;
  input [31:0] xt_rsc_6_31_i_qa_d;
  input [31:0] xt_rsc_7_0_i_qa_d;
  input [31:0] xt_rsc_7_1_i_qa_d;
  input [31:0] xt_rsc_7_2_i_qa_d;
  input [31:0] xt_rsc_7_3_i_qa_d;
  input [31:0] xt_rsc_7_4_i_qa_d;
  input [31:0] xt_rsc_7_5_i_qa_d;
  input [31:0] xt_rsc_7_6_i_qa_d;
  input [31:0] xt_rsc_7_7_i_qa_d;
  input [31:0] xt_rsc_7_8_i_qa_d;
  input [31:0] xt_rsc_7_9_i_qa_d;
  input [31:0] xt_rsc_7_10_i_qa_d;
  input [31:0] xt_rsc_7_11_i_qa_d;
  input [31:0] xt_rsc_7_12_i_qa_d;
  input [31:0] xt_rsc_7_13_i_qa_d;
  input [31:0] xt_rsc_7_14_i_qa_d;
  input [31:0] xt_rsc_7_15_i_qa_d;
  input [31:0] xt_rsc_7_16_i_qa_d;
  input [31:0] xt_rsc_7_17_i_qa_d;
  input [31:0] xt_rsc_7_18_i_qa_d;
  input [31:0] xt_rsc_7_19_i_qa_d;
  input [31:0] xt_rsc_7_20_i_qa_d;
  input [31:0] xt_rsc_7_21_i_qa_d;
  input [31:0] xt_rsc_7_22_i_qa_d;
  input [31:0] xt_rsc_7_23_i_qa_d;
  input [31:0] xt_rsc_7_24_i_qa_d;
  input [31:0] xt_rsc_7_25_i_qa_d;
  input [31:0] xt_rsc_7_26_i_qa_d;
  input [31:0] xt_rsc_7_27_i_qa_d;
  input [31:0] xt_rsc_7_28_i_qa_d;
  input [31:0] xt_rsc_7_29_i_qa_d;
  input [31:0] xt_rsc_7_30_i_qa_d;
  input [31:0] xt_rsc_7_31_i_qa_d;
  output [7:0] twiddle_rsc_0_0_i_adra_d;
  input [63:0] twiddle_rsc_0_0_i_qa_d;
  output [1:0] twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_1_i_adra_d;
  input [63:0] twiddle_rsc_0_1_i_qa_d;
  output [1:0] twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_2_i_adra_d;
  input [63:0] twiddle_rsc_0_2_i_qa_d;
  output [1:0] twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_3_i_adra_d;
  input [63:0] twiddle_rsc_0_3_i_qa_d;
  output [1:0] twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_4_i_adra_d;
  input [63:0] twiddle_rsc_0_4_i_qa_d;
  output [1:0] twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_5_i_adra_d;
  input [63:0] twiddle_rsc_0_5_i_qa_d;
  output [1:0] twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_6_i_adra_d;
  input [63:0] twiddle_rsc_0_6_i_qa_d;
  output [1:0] twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_7_i_adra_d;
  input [63:0] twiddle_rsc_0_7_i_qa_d;
  output [1:0] twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_8_i_adra_d;
  input [63:0] twiddle_rsc_0_8_i_qa_d;
  output [1:0] twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_9_i_adra_d;
  input [63:0] twiddle_rsc_0_9_i_qa_d;
  output [1:0] twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_10_i_adra_d;
  input [63:0] twiddle_rsc_0_10_i_qa_d;
  output [1:0] twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_11_i_adra_d;
  input [63:0] twiddle_rsc_0_11_i_qa_d;
  output [1:0] twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_12_i_adra_d;
  input [63:0] twiddle_rsc_0_12_i_qa_d;
  output [1:0] twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_13_i_adra_d;
  input [63:0] twiddle_rsc_0_13_i_qa_d;
  output [1:0] twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_14_i_adra_d;
  input [63:0] twiddle_rsc_0_14_i_qa_d;
  output [1:0] twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_15_i_adra_d;
  input [63:0] twiddle_rsc_0_15_i_qa_d;
  output [1:0] twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_0_i_adra_d;
  input [63:0] twiddle_h_rsc_0_0_i_qa_d;
  output [1:0] twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_1_i_adra_d;
  input [63:0] twiddle_h_rsc_0_1_i_qa_d;
  output [1:0] twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_2_i_adra_d;
  input [63:0] twiddle_h_rsc_0_2_i_qa_d;
  output [1:0] twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_3_i_adra_d;
  input [63:0] twiddle_h_rsc_0_3_i_qa_d;
  output [1:0] twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_4_i_adra_d;
  input [63:0] twiddle_h_rsc_0_4_i_qa_d;
  output [1:0] twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_5_i_adra_d;
  input [63:0] twiddle_h_rsc_0_5_i_qa_d;
  output [1:0] twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_6_i_adra_d;
  input [63:0] twiddle_h_rsc_0_6_i_qa_d;
  output [1:0] twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_7_i_adra_d;
  input [63:0] twiddle_h_rsc_0_7_i_qa_d;
  output [1:0] twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_8_i_adra_d;
  input [63:0] twiddle_h_rsc_0_8_i_qa_d;
  output [1:0] twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_9_i_adra_d;
  input [63:0] twiddle_h_rsc_0_9_i_qa_d;
  output [1:0] twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_10_i_adra_d;
  input [63:0] twiddle_h_rsc_0_10_i_qa_d;
  output [1:0] twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_11_i_adra_d;
  input [63:0] twiddle_h_rsc_0_11_i_qa_d;
  output [1:0] twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_12_i_adra_d;
  input [63:0] twiddle_h_rsc_0_12_i_qa_d;
  output [1:0] twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_13_i_adra_d;
  input [63:0] twiddle_h_rsc_0_13_i_qa_d;
  output [1:0] twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_14_i_adra_d;
  input [63:0] twiddle_h_rsc_0_14_i_qa_d;
  output [1:0] twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_15_i_adra_d;
  input [63:0] twiddle_h_rsc_0_15_i_qa_d;
  output [1:0] twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [31:0] yt_rsc_0_0_i_d_d_pff;
  output [3:0] yt_rsc_0_0_i_radr_d_pff;
  output [3:0] yt_rsc_0_0_i_wadr_d_pff;
  output yt_rsc_0_0_i_we_d_pff;
  output yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output [31:0] yt_rsc_0_1_i_d_d_pff;
  output [3:0] yt_rsc_0_1_i_wadr_d_pff;
  output [31:0] yt_rsc_0_2_i_d_d_pff;
  output [3:0] yt_rsc_0_2_i_wadr_d_pff;
  output [31:0] yt_rsc_0_3_i_d_d_pff;
  output [3:0] yt_rsc_0_3_i_wadr_d_pff;
  output [31:0] yt_rsc_0_4_i_d_d_pff;
  output [3:0] yt_rsc_0_4_i_wadr_d_pff;
  output [31:0] yt_rsc_0_5_i_d_d_pff;
  output [3:0] yt_rsc_0_5_i_wadr_d_pff;
  output [31:0] yt_rsc_0_6_i_d_d_pff;
  output [3:0] yt_rsc_0_6_i_wadr_d_pff;
  output [31:0] yt_rsc_0_7_i_d_d_pff;
  output [31:0] yt_rsc_0_8_i_d_d_pff;
  output [31:0] yt_rsc_0_9_i_d_d_pff;
  output [31:0] yt_rsc_0_10_i_d_d_pff;
  output [3:0] yt_rsc_0_10_i_wadr_d_pff;
  output [31:0] yt_rsc_0_11_i_d_d_pff;
  output [3:0] yt_rsc_0_11_i_wadr_d_pff;
  output [31:0] yt_rsc_0_12_i_d_d_pff;
  output [31:0] yt_rsc_0_13_i_d_d_pff;
  output [31:0] yt_rsc_0_14_i_d_d_pff;
  output [31:0] yt_rsc_0_15_i_d_d_pff;
  output yt_rsc_0_16_i_we_d_pff;
  output yt_rsc_1_0_i_we_d_pff;
  output yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output yt_rsc_1_16_i_we_d_pff;
  output yt_rsc_2_0_i_we_d_pff;
  output yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output yt_rsc_2_16_i_we_d_pff;
  output yt_rsc_3_0_i_we_d_pff;
  output yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output yt_rsc_3_16_i_we_d_pff;
  output [31:0] yt_rsc_4_0_i_d_d_pff;
  output [3:0] yt_rsc_4_0_i_wadr_d_pff;
  output yt_rsc_4_0_i_we_d_pff;
  output yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output [31:0] yt_rsc_4_1_i_d_d_pff;
  output [3:0] yt_rsc_4_1_i_wadr_d_pff;
  output [31:0] yt_rsc_4_2_i_d_d_pff;
  output [3:0] yt_rsc_4_2_i_wadr_d_pff;
  output [31:0] yt_rsc_4_3_i_d_d_pff;
  output [3:0] yt_rsc_4_3_i_wadr_d_pff;
  output [31:0] yt_rsc_4_4_i_d_d_pff;
  output [3:0] yt_rsc_4_4_i_wadr_d_pff;
  output [31:0] yt_rsc_4_5_i_d_d_pff;
  output [3:0] yt_rsc_4_5_i_wadr_d_pff;
  output [31:0] yt_rsc_4_6_i_d_d_pff;
  output [3:0] yt_rsc_4_6_i_wadr_d_pff;
  output [31:0] yt_rsc_4_7_i_d_d_pff;
  output [31:0] yt_rsc_4_8_i_d_d_pff;
  output [31:0] yt_rsc_4_9_i_d_d_pff;
  output [3:0] yt_rsc_4_9_i_wadr_d_pff;
  output [31:0] yt_rsc_4_10_i_d_d_pff;
  output [3:0] yt_rsc_4_10_i_wadr_d_pff;
  output [31:0] yt_rsc_4_11_i_d_d_pff;
  output [3:0] yt_rsc_4_11_i_wadr_d_pff;
  output [31:0] yt_rsc_4_12_i_d_d_pff;
  output [31:0] yt_rsc_4_13_i_d_d_pff;
  output [31:0] yt_rsc_4_14_i_d_d_pff;
  output [31:0] yt_rsc_4_15_i_d_d_pff;
  output yt_rsc_4_16_i_we_d_pff;
  output yt_rsc_5_0_i_we_d_pff;
  output yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output yt_rsc_5_16_i_we_d_pff;
  output yt_rsc_6_0_i_we_d_pff;
  output yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output yt_rsc_6_16_i_we_d_pff;
  output yt_rsc_7_0_i_we_d_pff;
  output yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff;
  output yt_rsc_7_16_i_we_d_pff;
  output [3:0] xt_rsc_0_0_i_adra_d_pff;
  output [31:0] xt_rsc_0_0_i_da_d_pff;
  output xt_rsc_0_0_i_wea_d_pff;
  output xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output [3:0] xt_rsc_0_1_i_adra_d_pff;
  output [31:0] xt_rsc_0_1_i_da_d_pff;
  output [3:0] xt_rsc_0_2_i_adra_d_pff;
  output [31:0] xt_rsc_0_2_i_da_d_pff;
  output [3:0] xt_rsc_0_3_i_adra_d_pff;
  output [31:0] xt_rsc_0_3_i_da_d_pff;
  output [3:0] xt_rsc_0_4_i_adra_d_pff;
  output [31:0] xt_rsc_0_4_i_da_d_pff;
  output [3:0] xt_rsc_0_5_i_adra_d_pff;
  output [31:0] xt_rsc_0_5_i_da_d_pff;
  output [3:0] xt_rsc_0_6_i_adra_d_pff;
  output [31:0] xt_rsc_0_6_i_da_d_pff;
  output [3:0] xt_rsc_0_7_i_adra_d_pff;
  output [31:0] xt_rsc_0_7_i_da_d_pff;
  output [3:0] xt_rsc_0_8_i_adra_d_pff;
  output [31:0] xt_rsc_0_8_i_da_d_pff;
  output [3:0] xt_rsc_0_9_i_adra_d_pff;
  output [31:0] xt_rsc_0_9_i_da_d_pff;
  output [3:0] xt_rsc_0_10_i_adra_d_pff;
  output [31:0] xt_rsc_0_10_i_da_d_pff;
  output [3:0] xt_rsc_0_11_i_adra_d_pff;
  output [31:0] xt_rsc_0_11_i_da_d_pff;
  output [3:0] xt_rsc_0_12_i_adra_d_pff;
  output [31:0] xt_rsc_0_12_i_da_d_pff;
  output [3:0] xt_rsc_0_13_i_adra_d_pff;
  output [31:0] xt_rsc_0_13_i_da_d_pff;
  output [3:0] xt_rsc_0_14_i_adra_d_pff;
  output [31:0] xt_rsc_0_14_i_da_d_pff;
  output [3:0] xt_rsc_0_15_i_adra_d_pff;
  output [31:0] xt_rsc_0_15_i_da_d_pff;
  output xt_rsc_0_16_i_wea_d_pff;
  output xt_rsc_1_0_i_wea_d_pff;
  output xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output xt_rsc_1_16_i_wea_d_pff;
  output xt_rsc_2_0_i_wea_d_pff;
  output xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output xt_rsc_2_16_i_wea_d_pff;
  output xt_rsc_3_0_i_wea_d_pff;
  output xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output xt_rsc_3_16_i_wea_d_pff;
  output [31:0] xt_rsc_4_0_i_da_d_pff;
  output xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output [3:0] xt_rsc_4_1_i_adra_d_pff;
  output [31:0] xt_rsc_4_1_i_da_d_pff;
  output [3:0] xt_rsc_4_2_i_adra_d_pff;
  output [31:0] xt_rsc_4_2_i_da_d_pff;
  output [31:0] xt_rsc_4_3_i_da_d_pff;
  output [31:0] xt_rsc_4_4_i_da_d_pff;
  output [31:0] xt_rsc_4_5_i_da_d_pff;
  output [31:0] xt_rsc_4_6_i_da_d_pff;
  output [31:0] xt_rsc_4_7_i_da_d_pff;
  output [31:0] xt_rsc_4_8_i_da_d_pff;
  output [3:0] xt_rsc_4_9_i_adra_d_pff;
  output [31:0] xt_rsc_4_9_i_da_d_pff;
  output [3:0] xt_rsc_4_10_i_adra_d_pff;
  output [31:0] xt_rsc_4_10_i_da_d_pff;
  output [31:0] xt_rsc_4_11_i_da_d_pff;
  output [31:0] xt_rsc_4_12_i_da_d_pff;
  output [31:0] xt_rsc_4_13_i_da_d_pff;
  output [31:0] xt_rsc_4_14_i_da_d_pff;
  output [31:0] xt_rsc_4_15_i_da_d_pff;
  output xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;
  output xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff;


  // Interconnect Declarations
  wire [31:0] p_rsci_idat;
  wire mult_t_mul_cmp_en;
  wire [63:0] mult_t_mul_cmp_z;
  wire [63:0] mult_t_mul_cmp_1_z;
  wire [63:0] mult_t_mul_cmp_2_z;
  wire [63:0] mult_t_mul_cmp_3_z;
  wire [63:0] mult_t_mul_cmp_4_z;
  wire [63:0] mult_t_mul_cmp_5_z;
  wire [63:0] mult_t_mul_cmp_6_z;
  wire [63:0] mult_t_mul_cmp_7_z;
  wire [63:0] mult_t_mul_cmp_8_z;
  wire [63:0] mult_t_mul_cmp_9_z;
  wire [63:0] mult_t_mul_cmp_10_z;
  wire [63:0] mult_t_mul_cmp_11_z;
  wire [63:0] mult_t_mul_cmp_12_z;
  wire [63:0] mult_t_mul_cmp_13_z;
  wire [63:0] mult_t_mul_cmp_14_z;
  wire [63:0] mult_t_mul_cmp_15_z;
  wire [31:0] mult_z_mul_cmp_z;
  wire mult_z_mul_cmp_1_en;
  wire [31:0] mult_z_mul_cmp_1_z;
  wire [31:0] mult_z_mul_cmp_2_z;
  wire [31:0] mult_z_mul_cmp_3_z;
  wire [31:0] mult_z_mul_cmp_4_z;
  wire [31:0] mult_z_mul_cmp_5_z;
  wire [31:0] mult_z_mul_cmp_6_z;
  wire [31:0] mult_z_mul_cmp_7_z;
  wire [31:0] mult_z_mul_cmp_8_z;
  wire [31:0] mult_z_mul_cmp_9_z;
  wire [31:0] mult_z_mul_cmp_10_z;
  wire [31:0] mult_z_mul_cmp_11_z;
  wire [31:0] mult_z_mul_cmp_12_z;
  wire [31:0] mult_z_mul_cmp_13_z;
  wire [31:0] mult_z_mul_cmp_14_z;
  wire [31:0] mult_z_mul_cmp_15_z;
  wire [31:0] mult_z_mul_cmp_16_z;
  wire [31:0] mult_z_mul_cmp_17_z;
  wire [31:0] mult_z_mul_cmp_18_z;
  wire [31:0] mult_z_mul_cmp_19_z;
  wire [31:0] mult_z_mul_cmp_20_z;
  wire [31:0] mult_z_mul_cmp_21_z;
  wire [31:0] mult_z_mul_cmp_22_z;
  wire [31:0] mult_z_mul_cmp_23_z;
  wire [31:0] mult_z_mul_cmp_24_z;
  wire [31:0] mult_z_mul_cmp_25_z;
  wire [31:0] mult_z_mul_cmp_26_z;
  wire [31:0] mult_z_mul_cmp_27_z;
  wire [31:0] mult_z_mul_cmp_28_z;
  wire [31:0] mult_z_mul_cmp_29_z;
  wire [31:0] mult_z_mul_cmp_30_z;
  wire [31:0] mult_z_mul_cmp_31_z;
  wire [10:0] fsm_output;
  wire INNER_LOOP4_nor_tmp;
  wire or_dcpl;
  wire or_dcpl_2;
  wire or_dcpl_8;
  wire or_dcpl_10;
  wire or_dcpl_12;
  wire or_dcpl_19;
  wire or_dcpl_22;
  wire or_dcpl_25;
  wire or_dcpl_30;
  wire or_dcpl_33;
  wire or_dcpl_36;
  wire or_dcpl_63;
  wire or_dcpl_70;
  wire or_dcpl_72;
  wire or_dcpl_76;
  wire or_dcpl_78;
  wire or_dcpl_80;
  wire or_dcpl_82;
  wire or_dcpl_88;
  wire or_dcpl_89;
  wire or_dcpl_94;
  wire or_dcpl_105;
  wire or_dcpl_107;
  wire or_dcpl_109;
  wire or_dcpl_111;
  wire or_dcpl_116;
  wire or_dcpl_117;
  wire or_dcpl_119;
  wire or_dcpl_121;
  wire or_dcpl_125;
  wire or_dcpl_133;
  wire or_dcpl_135;
  wire or_dcpl_139;
  wire or_dcpl_141;
  wire or_dcpl_146;
  wire or_dcpl_148;
  wire or_dcpl_150;
  wire or_dcpl_152;
  wire or_dcpl_161;
  wire or_dcpl_163;
  wire or_dcpl_165;
  wire or_dcpl_167;
  wire or_dcpl_171;
  wire or_dcpl_173;
  wire or_dcpl_180;
  wire or_dcpl_181;
  wire or_dcpl_185;
  wire or_dcpl_187;
  wire or_dcpl_189;
  wire or_dcpl_197;
  wire or_dcpl_199;
  wire or_dcpl_201;
  wire or_dcpl_203;
  wire or_dcpl_205;
  wire or_dcpl_207;
  wire or_dcpl_210;
  wire or_dcpl_215;
  wire or_dcpl_218;
  wire or_dcpl_220;
  wire or_dcpl_224;
  wire or_dcpl_234;
  wire or_dcpl_238;
  wire or_dcpl_242;
  wire or_dcpl_246;
  wire or_dcpl_274;
  wire and_dcpl_62;
  wire or_tmp_26;
  wire or_tmp_29;
  wire mux_tmp;
  wire or_tmp_35;
  wire not_tmp_25;
  wire or_tmp_38;
  wire or_tmp_40;
  wire not_tmp_29;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire and_dcpl_73;
  wire and_dcpl_76;
  wire nor_tmp_1;
  wire or_tmp_48;
  wire or_tmp_50;
  wire mux_tmp_7;
  wire or_tmp_53;
  wire or_tmp_55;
  wire not_tmp_50;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire or_tmp_64;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire or_tmp_72;
  wire and_dcpl_89;
  wire or_tmp_75;
  wire or_tmp_77;
  wire mux_tmp_22;
  wire nor_tmp_6;
  wire or_tmp_82;
  wire nor_tmp_10;
  wire or_tmp_84;
  wire or_tmp_86;
  wire not_tmp_67;
  wire not_tmp_69;
  wire or_tmp_90;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire nor_tmp_14;
  wire nor_tmp_15;
  wire or_tmp_93;
  wire or_tmp_94;
  wire nor_tmp_19;
  wire and_dcpl_96;
  wire or_tmp_99;
  wire or_tmp_102;
  wire or_tmp_104;
  wire and_dcpl_99;
  wire nor_tmp_22;
  wire or_tmp_112;
  wire not_tmp_87;
  wire mux_tmp_45;
  wire or_tmp_120;
  wire or_tmp_122;
  wire not_tmp_91;
  wire mux_tmp_50;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_107;
  wire nor_tmp_25;
  wire mux_tmp_53;
  wire mux_tmp_56;
  wire or_tmp_133;
  wire and_dcpl_112;
  wire and_dcpl_114;
  wire and_dcpl_116;
  wire and_dcpl_123;
  wire mux_tmp_70;
  wire nor_tmp_32;
  wire or_tmp_153;
  wire not_tmp_115;
  wire or_tmp_156;
  wire and_dcpl_125;
  wire nor_tmp_36;
  wire mux_tmp_78;
  wire or_tmp_160;
  wire nor_tmp_43;
  wire nor_tmp_45;
  wire nor_tmp_46;
  wire and_dcpl_135;
  wire and_dcpl_138;
  wire and_dcpl_141;
  wire and_dcpl_145;
  wire and_dcpl_147;
  wire and_dcpl_150;
  wire and_dcpl_152;
  wire and_dcpl_154;
  wire and_dcpl_161;
  wire and_dcpl_163;
  wire and_dcpl_167;
  wire and_dcpl_169;
  wire or_dcpl_298;
  wire or_dcpl_300;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire or_dcpl_315;
  wire and_dcpl_239;
  wire or_dcpl_353;
  wire or_dcpl_361;
  wire or_tmp_3231;
  wire or_tmp_3239;
  wire or_tmp_3242;
  wire or_tmp_3250;
  wire or_tmp_3252;
  wire or_tmp_3269;
  wire or_tmp_3279;
  wire or_tmp_3345;
  wire or_tmp_3354;
  wire or_tmp_3597;
  wire or_tmp_3600;
  wire or_tmp_3650;
  wire or_tmp_3666;
  wire or_tmp_3717;
  wire or_tmp_3723;
  wire or_tmp_3732;
  wire or_tmp_3755;
  wire or_tmp_3842;
  wire and_344_cse;
  wire and_346_cse;
  wire and_715_cse;
  wire and_717_cse;
  wire and_1022_cse;
  wire and_1024_cse;
  wire and_1329_cse;
  wire and_1331_cse;
  wire and_1636_cse;
  wire and_1638_cse;
  wire and_2007_cse;
  wire and_2009_cse;
  wire and_2314_cse;
  wire and_2316_cse;
  wire and_2621_cse;
  wire and_2623_cse;
  wire and_6834_cse;
  wire and_6843_cse;
  wire and_6852_cse;
  wire and_7090_cse;
  wire and_7109_cse;
  wire and_7115_cse;
  wire and_7153_cse;
  wire and_7173_cse;
  reg [6:0] INNER_LOOP4_r_11_4_sva_6_0;
  reg [6:0] INNER_LOOP3_r_11_4_sva_6_0;
  reg [6:0] INNER_LOOP2_r_11_4_sva_6_0;
  reg [6:0] INNER_LOOP1_r_11_4_sva_6_0;
  reg [1:0] butterFly1_15_conc_2_itm_2_1;
  reg c_1_sva;
  reg INNER_LOOP1_stage_0;
  reg butterFly1_15_conc_2_itm_3_0;
  reg butterFly1_15_conc_2_itm_8_0;
  reg butterFly1_15_conc_2_itm_5_0;
  reg butterFly1_15_conc_2_itm_4_0;
  reg butterFly1_15_conc_2_itm_2_0;
  reg [1:0] butterFly2_15_conc_itm_10_2_1;
  reg [1:0] butterFly2_15_conc_2_itm_9_2_1;
  reg butterFly1_15_f1_equal_tmp_1_1;
  reg butterFly1_15_conc_2_itm_0;
  reg butterFly1_15_f1_equal_tmp_2_1;
  reg butterFly1_15_conc_2_itm_1_0;
  reg [2:0] butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1;
  reg [1:0] butterFly2_15_conc_2_itm_6_2_1;
  reg [1:0] butterFly1_15_conc_2_itm_9_2_1;
  reg butterFly1_15_conc_2_itm_9_0;
  reg INNER_LOOP1_stage_0_10;
  reg butterFly2_15_conc_2_itm_7_0;
  reg INNER_LOOP1_stage_0_11;
  reg INNER_LOOP2_stage_0_10;
  reg [1:0] butterFly2_15_conc_2_itm_8_2_1;
  reg butterFly2_15_conc_2_itm_8_0;
  reg [1:0] butterFly1_15_conc_2_itm_8_2_1;
  reg butterFly2_15_conc_2_itm_5_0;
  reg [2:0] operator_20_false_acc_cse_sva;
  reg [1:0] operator_33_true_3_lshift_psp_1_0_sva;
  reg INNER_LOOP1_stage_0_3;
  reg INNER_LOOP1_stage_0_2;
  reg butterFly2_15_conc_2_itm_0;
  reg butterFly2_15_conc_2_itm_1_0;
  reg butterFly2_15_conc_2_itm_2_0;
  reg butterFly2_15_conc_2_itm_3_0;
  reg [1:0] butterFly1_15_conc_2_itm_4_2_1;
  reg [31:0] p_sva;
  wire butterFly1_15_and_ssc;
  wire butterFly1_15_and_ssc_2;
  wire butterFly1_14_and_ssc;
  wire butterFly1_14_and_ssc_2;
  wire butterFly1_14_and_ssc_3;
  wire butterFly1_13_and_ssc;
  wire butterFly1_13_and_ssc_2;
  wire butterFly1_13_and_ssc_3;
  wire butterFly1_12_and_ssc;
  wire butterFly1_12_and_ssc_2;
  wire butterFly1_12_and_ssc_3;
  wire butterFly1_11_and_ssc;
  wire butterFly1_11_and_ssc_2;
  wire butterFly1_11_and_ssc_3;
  wire butterFly1_10_and_ssc;
  wire butterFly1_10_and_ssc_2;
  wire butterFly1_10_and_ssc_3;
  wire butterFly1_9_and_ssc;
  wire butterFly1_9_and_ssc_2;
  wire butterFly1_9_and_ssc_3;
  wire butterFly1_8_and_ssc;
  wire butterFly1_8_and_ssc_2;
  wire butterFly1_8_and_ssc_3;
  wire butterFly1_7_and_ssc;
  wire butterFly1_7_and_ssc_2;
  wire butterFly1_7_and_ssc_3;
  wire butterFly1_6_and_ssc;
  wire butterFly1_6_and_ssc_2;
  wire butterFly1_6_and_ssc_3;
  wire butterFly1_5_and_ssc;
  wire butterFly1_5_and_ssc_2;
  wire butterFly1_5_and_ssc_3;
  wire butterFly1_4_and_ssc;
  wire butterFly1_4_and_ssc_2;
  wire butterFly1_4_and_ssc_3;
  wire butterFly1_3_and_ssc;
  wire butterFly1_3_and_ssc_2;
  wire butterFly1_3_and_ssc_3;
  wire butterFly1_2_and_ssc;
  wire butterFly1_2_and_ssc_2;
  wire butterFly1_2_and_ssc_3;
  wire butterFly1_1_and_ssc;
  wire butterFly1_1_and_ssc_2;
  wire butterFly1_1_and_ssc_3;
  wire butterFly1_and_ssc;
  wire butterFly1_and_ssc_2;
  reg reg_yt_rsc_0_0_cgo_cse;
  reg reg_yt_rsc_0_16_cgo_cse;
  reg reg_yt_rsc_1_0_cgo_cse;
  reg reg_yt_rsc_1_16_cgo_cse;
  reg reg_yt_rsc_2_0_cgo_cse;
  reg reg_yt_rsc_2_16_cgo_cse;
  reg reg_yt_rsc_3_0_cgo_cse;
  reg reg_yt_rsc_3_16_cgo_cse;
  reg reg_yt_rsc_4_0_cgo_cse;
  reg reg_yt_rsc_4_16_cgo_cse;
  reg reg_yt_rsc_5_0_cgo_cse;
  reg reg_yt_rsc_5_16_cgo_cse;
  reg reg_yt_rsc_6_0_cgo_cse;
  reg reg_yt_rsc_6_16_cgo_cse;
  reg reg_yt_rsc_7_0_cgo_cse;
  reg reg_yt_rsc_7_16_cgo_cse;
  reg reg_xt_rsc_triosy_7_31_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire mult_15_t_and_49_cse;
  wire mult_15_t_and_51_cse;
  wire mult_15_t_and_53_cse;
  wire mult_15_t_and_55_cse;
  wire mult_15_t_and_44_cse;
  wire mult_15_t_and_45_cse;
  wire mult_15_t_and_46_cse;
  wire mult_15_t_and_47_cse;
  wire mult_15_t_and_48_cse;
  wire mult_15_t_and_50_cse;
  wire mult_15_t_and_52_cse;
  wire mult_15_t_and_54_cse;
  reg reg_ensig_cgo_17_cse;
  wire or_383_cse;
  wire or_398_cse;
  wire nor_27_cse;
  wire and_8912_cse;
  wire butterFly2_16_f1_nor_1_cse;
  wire nand_7_cse;
  wire and_8932_cse;
  wire and_8913_cse;
  wire and_8919_cse;
  wire butterFly2_f1_nor_cse;
  wire butterFly1_f1_nor_cse;
  wire or_329_cse;
  wire or_412_cse;
  wire nand_24_cse;
  wire butterFly2_16_f1_butterFly2_16_f1_and_6_cse;
  wire and_8941_cse;
  wire [31:0] mult_15_res_sva_1;
  wire [32:0] nl_mult_15_res_sva_1;
  wire [31:0] mult_14_res_sva_1;
  wire [32:0] nl_mult_14_res_sva_1;
  wire [31:0] mult_13_res_sva_1;
  wire [32:0] nl_mult_13_res_sva_1;
  wire [31:0] mult_12_res_sva_1;
  wire [32:0] nl_mult_12_res_sva_1;
  wire [31:0] mult_11_res_sva_1;
  wire [32:0] nl_mult_11_res_sva_1;
  wire [31:0] mult_10_res_sva_1;
  wire [32:0] nl_mult_10_res_sva_1;
  wire [31:0] mult_9_res_sva_1;
  wire [32:0] nl_mult_9_res_sva_1;
  wire [31:0] mult_8_res_sva_1;
  wire [32:0] nl_mult_8_res_sva_1;
  wire [31:0] mult_7_res_sva_1;
  wire [32:0] nl_mult_7_res_sva_1;
  wire [31:0] mult_6_res_sva_1;
  wire [32:0] nl_mult_6_res_sva_1;
  wire [31:0] mult_5_res_sva_1;
  wire [32:0] nl_mult_5_res_sva_1;
  wire [31:0] mult_4_res_sva_1;
  wire [32:0] nl_mult_4_res_sva_1;
  wire [31:0] mult_3_res_sva_1;
  wire [32:0] nl_mult_3_res_sva_1;
  wire [31:0] mult_2_res_sva_1;
  wire [32:0] nl_mult_2_res_sva_1;
  wire [31:0] mult_1_res_sva_1;
  wire [32:0] nl_mult_1_res_sva_1;
  wire [31:0] mult_res_sva_1;
  wire [32:0] nl_mult_res_sva_1;
  wire butterFly2_7_tw_nor_cse;
  wire butterFly2_7_tw_nor_1_cse;
  wire butterFly2_7_tw_nor_2_cse;
  wire mult_15_t_or_9_cse;
  wire mult_15_t_or_10_cse;
  wire mult_15_t_or_11_cse;
  wire mult_15_t_or_12_cse;
  wire mult_15_t_and_41_cse;
  wire mult_15_t_and_42_cse;
  wire mult_15_t_and_43_cse;
  wire mult_15_t_and_37_cse;
  wire mult_15_t_and_38_cse;
  wire mult_15_t_and_39_cse;
  wire mult_15_t_and_30_cse;
  wire mult_15_t_and_31_cse;
  wire mult_15_t_and_32_cse;
  wire mult_15_t_or_3_cse;
  wire mult_15_t_and_40_cse;
  wire mult_15_t_and_36_cse;
  wire mult_15_t_and_29_cse;
  wire mult_15_t_or_1_cse;
  wire mult_15_t_or_cse;
  wire or_553_rmff;
  wire or_652_rmff;
  wire or_718_rmff;
  wire or_785_rmff;
  wire or_851_rmff;
  wire or_918_rmff;
  wire or_984_rmff;
  wire or_1051_rmff;
  wire or_1117_rmff;
  wire or_1216_rmff;
  wire or_1282_rmff;
  wire or_1349_rmff;
  wire or_1415_rmff;
  wire or_1482_rmff;
  wire or_1548_rmff;
  wire or_1615_rmff;
  wire [6:0] INNER_LOOP1_tw_h_mux1h_4_rmff;
  wire and_6824_rmff;
  wire [6:0] butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  wire or_3498_rmff;
  wire or_3502_rmff;
  wire or_3506_rmff;
  wire or_3510_rmff;
  wire or_3514_rmff;
  wire or_3518_rmff;
  wire or_3522_rmff;
  wire and_6895_rmff;
  wire or_3599_rmff;
  wire or_3759_rmff;
  wire [31:0] mult_4_t_mux1h_1_rmff;
  wire [31:0] mult_t_mul_cmp_5_a_mx0w1;
  wire [31:0] mult_t_mul_cmp_5_a_mx0w4;
  wire [31:0] mult_t_mul_cmp_11_a_mx0w3;
  wire [31:0] tmp_71_lpi_3_dfm_1;
  reg [31:0] modulo_add_31_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_10_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8;
  reg [31:0] modulo_add_1_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_11_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8;
  reg [31:0] modulo_add_23_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_12_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8;
  reg [31:0] modulo_add_24_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_13_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8;
  reg [31:0] modulo_add_25_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_14_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8;
  reg [31:0] modulo_add_26_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_15_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8;
  reg [31:0] modulo_add_27_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8;
  reg [31:0] modulo_add_28_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_29_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_30_qr_lpi_3_dfm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7;
  wire [31:0] z_out;
  wire [31:0] z_out_1;
  wire [31:0] z_out_2;
  wire [31:0] z_out_3;
  wire [31:0] z_out_4;
  wire [31:0] z_out_5;
  wire [31:0] z_out_6;
  wire [31:0] z_out_7;
  wire [31:0] z_out_8;
  wire [31:0] z_out_9;
  wire [31:0] z_out_10;
  wire [31:0] z_out_11;
  wire [31:0] z_out_12;
  wire [31:0] z_out_13;
  wire [31:0] z_out_14;
  wire [31:0] z_out_15;
  wire [31:0] z_out_16;
  wire [31:0] z_out_17;
  wire [31:0] z_out_18;
  wire [31:0] z_out_19;
  wire [31:0] z_out_20;
  wire [31:0] z_out_21;
  wire [31:0] z_out_22;
  wire [31:0] z_out_23;
  wire [31:0] z_out_24;
  wire [31:0] z_out_25;
  wire [31:0] z_out_26;
  wire [31:0] z_out_27;
  wire [31:0] z_out_28;
  wire [31:0] z_out_29;
  wire [31:0] z_out_30;
  wire [31:0] z_out_31;
  wire [31:0] z_out_32;
  wire [31:0] z_out_33;
  wire [31:0] z_out_34;
  wire [31:0] z_out_35;
  wire [31:0] z_out_36;
  wire [31:0] z_out_37;
  wire [31:0] z_out_38;
  wire [31:0] z_out_39;
  wire [31:0] z_out_40;
  wire [31:0] z_out_41;
  wire [31:0] z_out_42;
  wire [31:0] z_out_43;
  wire [31:0] z_out_44;
  wire [31:0] z_out_45;
  wire [31:0] z_out_46;
  wire [31:0] z_out_47;
  wire [31:0] z_out_48;
  wire [31:0] z_out_49;
  wire [31:0] z_out_50;
  wire [31:0] z_out_51;
  wire [31:0] z_out_52;
  wire [31:0] z_out_53;
  wire [31:0] z_out_54;
  wire [31:0] z_out_55;
  wire [31:0] z_out_56;
  wire [31:0] z_out_57;
  wire [31:0] z_out_58;
  wire [31:0] z_out_59;
  wire [10:0] z_out_60;
  wire [2:0] z_out_61;
  wire [3:0] nl_z_out_61;
  wire [7:0] z_out_62;
  wire [8:0] nl_z_out_62;
  wire [31:0] z_out_68;
  wire [32:0] nl_z_out_68;
  wire [31:0] z_out_69;
  wire [32:0] nl_z_out_69;
  wire [31:0] z_out_70;
  wire [32:0] nl_z_out_70;
  wire [31:0] z_out_72;
  wire [32:0] nl_z_out_72;
  wire [31:0] z_out_73;
  wire [32:0] nl_z_out_73;
  wire [31:0] z_out_74;
  wire [32:0] nl_z_out_74;
  wire [31:0] z_out_76;
  wire [32:0] nl_z_out_76;
  wire [31:0] z_out_77;
  wire [32:0] nl_z_out_77;
  wire [31:0] z_out_78;
  wire [32:0] nl_z_out_78;
  wire [31:0] z_out_80;
  wire [32:0] nl_z_out_80;
  wire [31:0] z_out_81;
  wire [32:0] nl_z_out_81;
  wire [31:0] z_out_82;
  wire [32:0] nl_z_out_82;
  wire [31:0] z_out_84;
  wire [32:0] nl_z_out_84;
  wire [31:0] z_out_85;
  wire [32:0] nl_z_out_85;
  wire [31:0] z_out_86;
  wire [32:0] nl_z_out_86;
  wire [31:0] z_out_88;
  wire [32:0] nl_z_out_88;
  wire [31:0] z_out_89;
  wire [32:0] nl_z_out_89;
  wire [31:0] z_out_90;
  wire [32:0] nl_z_out_90;
  wire [31:0] z_out_92;
  wire [32:0] nl_z_out_92;
  wire [31:0] z_out_93;
  wire [32:0] nl_z_out_93;
  wire [31:0] z_out_94;
  wire [32:0] nl_z_out_94;
  wire [31:0] z_out_96;
  wire [32:0] nl_z_out_96;
  wire [31:0] z_out_97;
  wire [32:0] nl_z_out_97;
  wire [31:0] z_out_98;
  wire [32:0] nl_z_out_98;
  wire [31:0] z_out_100;
  wire [32:0] nl_z_out_100;
  wire [31:0] z_out_101;
  wire [32:0] nl_z_out_101;
  wire [31:0] z_out_102;
  wire [32:0] nl_z_out_102;
  wire [31:0] z_out_104;
  wire [32:0] nl_z_out_104;
  wire [31:0] z_out_105;
  wire [32:0] nl_z_out_105;
  wire [31:0] z_out_106;
  wire [32:0] nl_z_out_106;
  wire [31:0] z_out_108;
  wire [32:0] nl_z_out_108;
  wire [31:0] z_out_109;
  wire [32:0] nl_z_out_109;
  wire [31:0] z_out_111;
  wire [31:0] z_out_112;
  wire [31:0] z_out_113;
  wire [31:0] z_out_114;
  wire [31:0] z_out_115;
  wire [31:0] z_out_116;
  wire [31:0] z_out_117;
  wire [31:0] z_out_118;
  wire [31:0] z_out_119;
  wire [31:0] z_out_120;
  wire [31:0] z_out_121;
  wire [31:0] z_out_122;
  wire [31:0] z_out_123;
  wire [31:0] z_out_124;
  wire [31:0] z_out_125;
  wire [31:0] z_out_126;
  wire [31:0] z_out_127;
  wire [32:0] nl_z_out_127;
  wire [31:0] z_out_128;
  wire [32:0] nl_z_out_128;
  wire [31:0] z_out_129;
  wire [32:0] nl_z_out_129;
  wire [31:0] z_out_130;
  wire [32:0] nl_z_out_130;
  wire [31:0] z_out_131;
  wire [32:0] nl_z_out_131;
  wire [31:0] z_out_132;
  wire [32:0] nl_z_out_132;
  wire [31:0] z_out_133;
  wire [32:0] nl_z_out_133;
  wire [31:0] z_out_134;
  wire [32:0] nl_z_out_134;
  wire [31:0] z_out_135;
  wire [32:0] nl_z_out_135;
  wire [31:0] z_out_136;
  wire [32:0] nl_z_out_136;
  wire [31:0] z_out_137;
  wire [32:0] nl_z_out_137;
  wire [31:0] z_out_138;
  wire [32:0] nl_z_out_138;
  wire [31:0] z_out_139;
  wire [32:0] nl_z_out_139;
  wire [31:0] z_out_140;
  wire [32:0] nl_z_out_140;
  wire [31:0] z_out_141;
  wire [32:0] nl_z_out_141;
  wire [31:0] z_out_142;
  wire [32:0] nl_z_out_142;
  reg [5:0] operator_33_true_1_lshift_psp_9_4_sva;
  reg [2:0] butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm;
  reg [31:0] tmp_64_lpi_3_dfm_1;
  reg [31:0] tmp_66_lpi_3_dfm_1;
  reg [31:0] tmp_68_lpi_3_dfm_1;
  reg [31:0] tmp_70_lpi_3_dfm_1;
  reg [31:0] tmp_72_lpi_3_dfm_1;
  reg [31:0] tmp_74_lpi_3_dfm_1;
  reg [31:0] tmp_76_lpi_3_dfm_1;
  reg [31:0] tmp_78_lpi_3_dfm_1;
  reg [31:0] tmp_80_lpi_3_dfm_1;
  reg [31:0] tmp_82_lpi_3_dfm_1;
  reg [31:0] tmp_84_lpi_3_dfm_1;
  reg [31:0] tmp_86_lpi_3_dfm_1;
  reg [31:0] tmp_88_lpi_3_dfm_1;
  reg [31:0] tmp_90_lpi_3_dfm_1;
  reg [31:0] tmp_92_lpi_3_dfm_1;
  reg butterFly1_15_f1_equal_tmp_1;
  reg butterFly1_15_f1_equal_tmp_3_1;
  reg butterFly1_15_f1_equal_tmp_4_1;
  reg butterFly1_15_f1_equal_tmp_5_1;
  reg butterFly1_15_f1_equal_tmp_6_1;
  reg butterFly1_15_f1_equal_tmp_7_1;
  reg [31:0] tmp_94_lpi_3_dfm_1;
  reg [31:0] mult_1_z_asn_itm_1;
  reg [31:0] mult_1_z_asn_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_7;
  reg [31:0] mult_10_z_asn_itm_1;
  reg [31:0] mult_10_z_asn_itm_2;
  reg [31:0] mult_10_z_asn_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_6;
  reg [31:0] mult_11_z_asn_itm_1;
  reg [31:0] mult_11_z_asn_itm_2;
  reg [31:0] mult_11_z_asn_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_7;
  reg [31:0] mult_12_z_asn_itm_1;
  reg [31:0] mult_12_z_asn_itm_2;
  reg [31:0] mult_12_z_asn_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_7;
  reg [31:0] mult_13_z_asn_itm_1;
  reg [31:0] mult_13_z_asn_itm_2;
  reg [31:0] mult_13_z_asn_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_7;
  reg [31:0] mult_14_z_asn_itm_1;
  reg [31:0] mult_14_z_asn_itm_2;
  reg [31:0] mult_14_z_asn_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_7;
  reg [31:0] mult_15_z_asn_itm_1;
  reg [31:0] mult_15_z_asn_itm_2;
  reg [31:0] mult_15_z_asn_itm_3;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_7;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_1;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_2;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_4;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_5;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_6;
  reg [3:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_7;
  reg [31:0] tmp_lpi_3_dfm_1;
  reg [31:0] tmp_2_lpi_3_dfm_1;
  reg [31:0] tmp_4_lpi_3_dfm_1;
  reg [31:0] tmp_6_lpi_3_dfm_1;
  reg [31:0] tmp_8_lpi_3_dfm_1;
  reg [31:0] tmp_10_lpi_3_dfm_1;
  reg [31:0] tmp_10_lpi_3_dfm_2;
  reg [31:0] tmp_10_lpi_3_dfm_3;
  reg [31:0] tmp_10_lpi_3_dfm_4;
  reg [31:0] tmp_10_lpi_3_dfm_5;
  reg [31:0] tmp_10_lpi_3_dfm_6;
  reg [31:0] tmp_10_lpi_3_dfm_7;
  reg [31:0] tmp_12_lpi_3_dfm_1;
  reg [31:0] tmp_14_lpi_3_dfm_1;
  reg [31:0] tmp_16_lpi_3_dfm_1;
  reg [31:0] tmp_18_lpi_3_dfm_1;
  reg [31:0] tmp_20_lpi_3_dfm_1;
  reg [31:0] tmp_22_lpi_3_dfm_1;
  reg [31:0] tmp_24_lpi_3_dfm_1;
  reg [31:0] tmp_26_lpi_3_dfm_1;
  reg [31:0] tmp_28_lpi_3_dfm_1;
  reg [31:0] tmp_30_lpi_3_dfm_1;
  reg [31:0] mult_16_z_asn_itm_3;
  reg [31:0] mult_17_z_asn_itm_3;
  reg [31:0] mult_18_z_asn_itm_3;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_3;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_4;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_5;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_6;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_7;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_8;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_1;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_2;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_3;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_4;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_5;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_6;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_7;
  reg [3:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_8;
  reg [31:0] mult_19_z_asn_itm_3;
  reg [31:0] mult_20_z_asn_itm_3;
  reg [31:0] mult_21_z_asn_itm_3;
  reg [31:0] mult_22_z_asn_itm_3;
  reg [31:0] mult_23_z_asn_itm_1;
  reg [31:0] mult_23_z_asn_itm_2;
  reg [31:0] mult_23_z_asn_itm_3;
  reg [31:0] mult_24_z_asn_itm_1;
  reg [31:0] mult_24_z_asn_itm_2;
  reg [31:0] mult_24_z_asn_itm_3;
  reg [31:0] mult_25_z_asn_itm_1;
  reg [31:0] mult_25_z_asn_itm_2;
  reg [31:0] mult_25_z_asn_itm_3;
  reg [31:0] mult_26_z_asn_itm_1;
  reg [31:0] mult_26_z_asn_itm_2;
  reg [31:0] mult_27_z_asn_itm_1;
  reg [31:0] mult_27_z_asn_itm_2;
  reg [31:0] mult_28_z_asn_itm_1;
  reg [31:0] mult_28_z_asn_itm_2;
  reg [31:0] mult_29_z_asn_itm_1;
  reg [31:0] mult_29_z_asn_itm_2;
  reg [31:0] mult_30_z_asn_itm_1;
  reg [31:0] mult_30_z_asn_itm_2;
  reg [31:0] mult_31_z_asn_itm_1;
  reg [31:0] mult_31_z_asn_itm_2;
  reg [31:0] tmp_96_lpi_3_dfm_1;
  reg [31:0] tmp_98_lpi_3_dfm_1;
  reg [31:0] tmp_100_lpi_3_dfm_1;
  reg [31:0] tmp_102_lpi_3_dfm_1;
  reg [31:0] tmp_102_lpi_3_dfm_2;
  reg [31:0] tmp_102_lpi_3_dfm_3;
  reg [31:0] tmp_102_lpi_3_dfm_4;
  reg [31:0] tmp_102_lpi_3_dfm_5;
  reg [31:0] tmp_102_lpi_3_dfm_6;
  reg [31:0] tmp_102_lpi_3_dfm_7;
  reg [31:0] tmp_104_lpi_3_dfm_1;
  reg [31:0] tmp_104_lpi_3_dfm_2;
  reg [31:0] tmp_104_lpi_3_dfm_3;
  reg [31:0] tmp_104_lpi_3_dfm_4;
  reg [31:0] tmp_104_lpi_3_dfm_5;
  reg [31:0] tmp_104_lpi_3_dfm_6;
  reg [31:0] tmp_104_lpi_3_dfm_7;
  reg [31:0] tmp_106_lpi_3_dfm_1;
  reg [31:0] tmp_106_lpi_3_dfm_2;
  reg [31:0] tmp_106_lpi_3_dfm_3;
  reg [31:0] tmp_106_lpi_3_dfm_4;
  reg [31:0] tmp_106_lpi_3_dfm_5;
  reg [31:0] tmp_106_lpi_3_dfm_6;
  reg [31:0] tmp_106_lpi_3_dfm_7;
  reg [31:0] tmp_108_lpi_3_dfm_1;
  reg [31:0] tmp_108_lpi_3_dfm_2;
  reg [31:0] tmp_108_lpi_3_dfm_3;
  reg [31:0] tmp_108_lpi_3_dfm_4;
  reg [31:0] tmp_108_lpi_3_dfm_5;
  reg [31:0] tmp_108_lpi_3_dfm_6;
  reg [31:0] tmp_108_lpi_3_dfm_7;
  reg [31:0] tmp_110_lpi_3_dfm_1;
  reg [31:0] tmp_110_lpi_3_dfm_2;
  reg [31:0] tmp_110_lpi_3_dfm_3;
  reg [31:0] tmp_110_lpi_3_dfm_4;
  reg [31:0] tmp_110_lpi_3_dfm_5;
  reg [31:0] tmp_110_lpi_3_dfm_6;
  reg [31:0] tmp_110_lpi_3_dfm_7;
  reg [31:0] tmp_112_lpi_3_dfm_1;
  reg [31:0] tmp_112_lpi_3_dfm_2;
  reg [31:0] tmp_112_lpi_3_dfm_3;
  reg [31:0] tmp_112_lpi_3_dfm_4;
  reg [31:0] tmp_112_lpi_3_dfm_5;
  reg [31:0] tmp_112_lpi_3_dfm_6;
  reg [31:0] tmp_112_lpi_3_dfm_7;
  reg [31:0] tmp_114_lpi_3_dfm_1;
  reg [31:0] tmp_114_lpi_3_dfm_2;
  reg [31:0] tmp_114_lpi_3_dfm_3;
  reg [31:0] tmp_114_lpi_3_dfm_4;
  reg [31:0] tmp_114_lpi_3_dfm_5;
  reg [31:0] tmp_114_lpi_3_dfm_6;
  reg [31:0] tmp_114_lpi_3_dfm_7;
  reg [31:0] tmp_116_lpi_3_dfm_1;
  reg [31:0] tmp_116_lpi_3_dfm_2;
  reg [31:0] tmp_116_lpi_3_dfm_3;
  reg [31:0] tmp_116_lpi_3_dfm_4;
  reg [31:0] tmp_116_lpi_3_dfm_5;
  reg [31:0] tmp_116_lpi_3_dfm_6;
  reg [31:0] tmp_116_lpi_3_dfm_7;
  reg [31:0] tmp_118_lpi_3_dfm_1;
  reg [31:0] tmp_118_lpi_3_dfm_2;
  reg [31:0] tmp_118_lpi_3_dfm_3;
  reg [31:0] tmp_118_lpi_3_dfm_4;
  reg [31:0] tmp_118_lpi_3_dfm_5;
  reg [31:0] tmp_118_lpi_3_dfm_6;
  reg [31:0] tmp_118_lpi_3_dfm_7;
  reg [31:0] tmp_120_lpi_3_dfm_1;
  reg [31:0] tmp_120_lpi_3_dfm_2;
  reg [31:0] tmp_120_lpi_3_dfm_3;
  reg [31:0] tmp_120_lpi_3_dfm_4;
  reg [31:0] tmp_120_lpi_3_dfm_5;
  reg [31:0] tmp_120_lpi_3_dfm_6;
  reg [31:0] tmp_120_lpi_3_dfm_7;
  reg [31:0] tmp_122_lpi_3_dfm_1;
  reg [31:0] tmp_122_lpi_3_dfm_2;
  reg [31:0] tmp_122_lpi_3_dfm_3;
  reg [31:0] tmp_122_lpi_3_dfm_4;
  reg [31:0] tmp_122_lpi_3_dfm_5;
  reg [31:0] tmp_122_lpi_3_dfm_6;
  reg [31:0] tmp_122_lpi_3_dfm_7;
  reg [31:0] tmp_124_lpi_3_dfm_1;
  reg [31:0] tmp_124_lpi_3_dfm_2;
  reg [31:0] tmp_124_lpi_3_dfm_3;
  reg [31:0] tmp_124_lpi_3_dfm_4;
  reg [31:0] tmp_124_lpi_3_dfm_5;
  reg [31:0] tmp_124_lpi_3_dfm_6;
  reg [31:0] tmp_124_lpi_3_dfm_7;
  reg butterFly2_15_f1_equal_tmp_1;
  reg butterFly2_15_f1_equal_tmp_7_1;
  reg [31:0] tmp_126_lpi_3_dfm_1;
  reg [31:0] tmp_126_lpi_3_dfm_2;
  reg [31:0] tmp_126_lpi_3_dfm_3;
  reg [31:0] tmp_126_lpi_3_dfm_4;
  reg [31:0] tmp_126_lpi_3_dfm_5;
  reg [31:0] tmp_126_lpi_3_dfm_6;
  reg [31:0] tmp_126_lpi_3_dfm_7;
  reg butterFly2_15_tw_equal_tmp_1;
  reg butterFly2_15_tw_equal_tmp_3_1;
  reg butterFly2_15_tw_equal_tmp_5_1;
  reg butterFly2_15_tw_equal_tmp_6_1;
  reg butterFly2_15_tw_equal_tmp_7_1;
  reg [31:0] tmp_32_lpi_3_dfm_1;
  reg [31:0] tmp_34_lpi_3_dfm_1;
  reg [31:0] tmp_36_lpi_3_dfm_1;
  reg [31:0] tmp_38_lpi_3_dfm_1;
  reg [31:0] tmp_40_lpi_3_dfm_1;
  reg [31:0] tmp_42_lpi_3_dfm_1;
  reg [31:0] tmp_44_lpi_3_dfm_1;
  reg [31:0] tmp_46_lpi_3_dfm_1;
  reg [31:0] tmp_48_lpi_3_dfm_1;
  reg [31:0] tmp_50_lpi_3_dfm_1;
  reg [31:0] tmp_52_lpi_3_dfm_1;
  reg [31:0] tmp_54_lpi_3_dfm_1;
  reg [31:0] tmp_56_lpi_3_dfm_1;
  reg [31:0] tmp_58_lpi_3_dfm_1;
  reg [31:0] tmp_60_lpi_3_dfm_1;
  reg [31:0] tmp_60_lpi_3_dfm_2;
  reg [31:0] tmp_60_lpi_3_dfm_3;
  reg [31:0] tmp_60_lpi_3_dfm_4;
  reg [31:0] tmp_60_lpi_3_dfm_5;
  reg [31:0] tmp_60_lpi_3_dfm_6;
  reg [31:0] tmp_60_lpi_3_dfm_7;
  reg [31:0] tmp_62_lpi_3_dfm_1;
  reg [31:0] tmp_62_lpi_3_dfm_2;
  reg [31:0] tmp_62_lpi_3_dfm_3;
  reg [31:0] tmp_62_lpi_3_dfm_4;
  reg [31:0] tmp_62_lpi_3_dfm_5;
  reg [31:0] tmp_62_lpi_3_dfm_6;
  reg [31:0] tmp_62_lpi_3_dfm_7;
  reg [1:0] butterFly1_15_conc_2_itm_1_2_1;
  reg [1:0] butterFly1_15_conc_2_itm_2_2_1;
  reg [1:0] butterFly1_15_conc_2_itm_3_2_1;
  reg [1:0] butterFly1_15_conc_2_itm_5_2_1;
  reg [1:0] butterFly1_15_conc_2_itm_6_2_1;
  reg butterFly1_15_conc_2_itm_6_0;
  reg [1:0] butterFly1_15_conc_2_itm_7_2_1;
  reg butterFly1_15_conc_2_itm_7_0;
  reg butterFly2_15_conc_2_itm_4_0;
  reg [1:0] butterFly2_15_conc_2_itm_7_2_1;
  wire [1:0] operator_33_true_3_lshift_psp_1_0_sva_mx0w5;
  wire [31:0] mult_15_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_14_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_13_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_12_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_11_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_10_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_9_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_8_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_7_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_6_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_5_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_4_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_3_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_2_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_1_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_res_lpi_3_dfm_1_mx0;
  wire [6:0] INNER_LOOP2_r_11_4_sva_6_0_mx1;
  wire [2:0] operator_33_true_2_lshift_psp_2_0_sva_mx0;
  wire modulo_sub_31_qelse_and_ssc;
  wire modulo_sub_31_qelse_and_ssc_1;
  reg reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_30_qelse_and_ssc;
  wire modulo_sub_30_qelse_and_ssc_1;
  reg reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_29_qelse_and_ssc;
  wire modulo_sub_29_qelse_and_ssc_1;
  reg reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_28_qelse_and_ssc;
  wire modulo_sub_28_qelse_and_ssc_1;
  reg reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_27_qelse_and_ssc;
  wire modulo_sub_27_qelse_and_ssc_1;
  reg reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_26_qelse_and_ssc;
  wire modulo_sub_26_qelse_and_ssc_1;
  reg reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_25_qelse_and_ssc;
  wire modulo_sub_25_qelse_and_ssc_1;
  reg reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_24_qelse_and_ssc;
  wire modulo_sub_24_qelse_and_ssc_1;
  reg reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_23_qelse_and_ssc;
  wire modulo_sub_23_qelse_and_ssc_1;
  reg reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_22_qelse_and_ssc;
  wire modulo_sub_22_qelse_and_ssc_1;
  reg reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_21_qelse_and_ssc;
  wire modulo_sub_21_qelse_and_ssc_1;
  reg reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_20_qelse_and_ssc;
  wire modulo_sub_20_qelse_and_ssc_1;
  reg reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_19_qelse_and_ssc;
  wire modulo_sub_19_qelse_and_ssc_1;
  reg reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_18_qelse_and_ssc;
  wire modulo_sub_18_qelse_and_ssc_1;
  reg reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_17_qelse_and_ssc;
  wire modulo_sub_17_qelse_and_ssc_1;
  reg reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_16_qelse_and_ssc;
  wire modulo_sub_16_qelse_and_ssc_1;
  reg reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_add_1_qelse_or_m1c;
  reg [31:0] reg_mult_15_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_14_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_13_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_12_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_11_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_10_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_9_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_8_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_7_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_6_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_5_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_4_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_3_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_2_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_1_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_32_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_33_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_34_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_35_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_36_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_37_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_38_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_39_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_40_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_41_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_42_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_43_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_44_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_45_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_46_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_47_res_lpi_3_dfm_1_cse;
  wire [6:0] INNER_LOOP1_r_INNER_LOOP1_r_and_cse;
  wire [6:0] INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse;
  wire [6:0] INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse;
  wire butterFly1_15_f1_mux_cse;
  wire butterFly1_15_f1_mux_1_cse;
  wire butterFly1_15_f1_mux_2_cse;
  wire butterFly1_15_f1_mux_3_cse;
  wire butterFly1_15_f1_mux_4_cse;
  wire butterFly1_15_f1_mux_5_cse;
  wire butterFly1_15_f1_mux_6_cse;
  wire butterFly1_15_f1_mux_7_cse;
  wire butterFly1_31_f1_mux_cse;
  wire butterFly1_31_f1_mux_1_cse;
  wire butterFly1_31_f1_mux_2_cse;
  wire butterFly1_31_f1_mux_3_cse;
  wire butterFly1_31_f1_mux_4_cse;
  wire butterFly1_31_f1_mux_5_cse;
  wire butterFly1_31_f1_mux_6_cse;
  wire butterFly1_31_f1_mux_7_cse;
  wire butterFly2_f1_mux_cse;
  wire butterFly2_f1_mux_1_cse;
  wire butterFly2_f1_mux_2_cse;
  wire butterFly2_f1_mux_3_cse;
  wire butterFly2_f1_mux_4_cse;
  wire butterFly2_f1_mux_5_cse;
  wire butterFly2_f1_mux_6_cse;
  wire butterFly2_f1_mux_7_cse;
  wire butterFly2_21_f1_mux_cse;
  wire butterFly2_21_f1_mux_1_cse;
  wire butterFly2_21_f1_mux_2_cse;
  wire butterFly2_21_f1_mux_3_cse;
  wire butterFly2_21_f1_mux_4_cse;
  wire butterFly2_21_f1_mux_5_cse;
  wire butterFly2_21_f1_mux_6_cse;
  wire butterFly2_21_f1_mux_7_cse;
  wire or_4976_cse;
  wire z_out_143_32;
  wire z_out_144_32;
  wire z_out_145_32;
  wire z_out_146_32;
  wire z_out_147_32;
  wire z_out_148_32;
  wire z_out_149_32;
  wire z_out_150_32;
  wire z_out_151_32;
  wire z_out_152_32;
  wire z_out_153_32;
  wire z_out_154_32;
  wire z_out_155_32;
  wire z_out_156_32;
  wire z_out_157_32;
  wire z_out_158_32;

  wire[0:0] c_mux_nl;
  wire[0:0] butterFly2_21_tw_butterFly2_21_tw_or_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] mux_1_nl;
  wire[0:0] or_322_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] or_337_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_344_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] or_352_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] or_356_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] or_360_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] or_367_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] or_368_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] or_372_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] nor_49_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] nor_50_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] nand_1_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] mux_41_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] or_404_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] or_406_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] or_426_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] or_433_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] mux_66_nl;
  wire[0:0] or_442_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] mux_68_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] mux_72_nl;
  wire[0:0] mux_71_nl;
  wire[0:0] or_444_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] mux_80_nl;
  wire[0:0] mux_79_nl;
  wire[0:0] nor_48_nl;
  wire[0:0] mux_82_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] mux_84_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_83_nl;
  wire[0:0] mux_88_nl;
  wire[0:0] mux_87_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] mux_89_nl;
  wire[0:0] mux_92_nl;
  wire[0:0] mux_91_nl;
  wire[0:0] mult_4_t_and_nl;
  wire[0:0] mult_4_t_and_1_nl;
  wire[0:0] mult_4_t_and_2_nl;
  wire[0:0] mult_4_t_and_3_nl;
  wire[0:0] mult_4_t_and_4_nl;
  wire[0:0] mult_4_t_and_5_nl;
  wire[0:0] mult_4_t_and_6_nl;
  wire[0:0] mult_4_t_and_7_nl;
  wire[0:0] mult_4_t_and_8_nl;
  wire[0:0] mult_4_t_and_9_nl;
  wire[0:0] mult_4_t_and_10_nl;
  wire[0:0] mult_4_t_and_11_nl;
  wire[0:0] mult_4_t_and_12_nl;
  wire[0:0] mult_4_t_and_13_nl;
  wire[0:0] mult_4_t_and_14_nl;
  wire[0:0] mult_4_t_and_15_nl;
  wire[0:0] mult_4_t_and_16_nl;
  wire[0:0] mult_4_t_and_17_nl;
  wire[0:0] mult_4_t_and_18_nl;
  wire[0:0] mult_4_t_and_19_nl;
  wire[0:0] mult_4_t_and_20_nl;
  wire[0:0] mult_4_t_and_21_nl;
  wire[0:0] mult_4_t_and_22_nl;
  wire[0:0] mult_4_t_and_23_nl;
  wire[0:0] mult_4_t_and_24_nl;
  wire[0:0] mult_4_t_and_25_nl;
  wire[0:0] mult_4_t_and_26_nl;
  wire[0:0] mult_4_t_and_27_nl;
  wire[0:0] mult_4_t_and_28_nl;
  wire[0:0] mult_4_t_and_29_nl;
  wire[0:0] mult_4_t_and_30_nl;
  wire[0:0] mult_4_t_and_31_nl;
  wire[1:0] STAGE_LOOP_mux1h_nl;
  wire[32:0] acc_2_nl;
  wire[33:0] nl_acc_2_nl;
  wire[31:0] modulo_add_1_qif_mux1h_2_nl;
  wire[0:0] modulo_add_1_qelse_and_nl;
  wire[0:0] modulo_add_1_qelse_or_1_nl;
  wire[0:0] modulo_add_1_qelse_and_4_nl;
  wire[0:0] modulo_add_1_qelse_and_5_nl;
  wire[32:0] acc_3_nl;
  wire[33:0] nl_acc_3_nl;
  wire[31:0] modulo_add_10_qif_mux1h_2_nl;
  wire[0:0] modulo_add_10_qelse_and_nl;
  wire[0:0] modulo_add_10_qelse_or_nl;
  wire[0:0] modulo_add_10_qelse_and_5_nl;
  wire[0:0] modulo_add_10_qelse_and_6_nl;
  wire[0:0] modulo_add_10_qelse_and_7_nl;
  wire[32:0] acc_4_nl;
  wire[33:0] nl_acc_4_nl;
  wire[31:0] modulo_add_11_qif_mux1h_2_nl;
  wire[0:0] modulo_add_11_qelse_and_nl;
  wire[0:0] modulo_add_11_qelse_or_nl;
  wire[0:0] modulo_add_11_qelse_and_5_nl;
  wire[0:0] modulo_add_11_qelse_and_6_nl;
  wire[0:0] modulo_add_11_qelse_and_7_nl;
  wire[32:0] acc_5_nl;
  wire[33:0] nl_acc_5_nl;
  wire[31:0] modulo_add_12_qif_mux1h_2_nl;
  wire[0:0] modulo_add_12_qelse_and_nl;
  wire[0:0] modulo_add_12_qelse_or_1_nl;
  wire[0:0] modulo_add_12_qelse_and_4_nl;
  wire[0:0] modulo_add_12_qelse_and_5_nl;
  wire[32:0] acc_6_nl;
  wire[33:0] nl_acc_6_nl;
  wire[31:0] modulo_add_13_qif_mux1h_2_nl;
  wire[0:0] modulo_add_13_qelse_and_nl;
  wire[0:0] modulo_add_13_qelse_or_1_nl;
  wire[0:0] modulo_add_13_qelse_and_4_nl;
  wire[0:0] modulo_add_13_qelse_and_5_nl;
  wire[32:0] acc_10_nl;
  wire[33:0] nl_acc_10_nl;
  wire[31:0] modulo_add_14_qif_mux1h_2_nl;
  wire[0:0] modulo_add_14_qelse_and_nl;
  wire[0:0] modulo_add_14_qelse_or_1_nl;
  wire[0:0] modulo_add_14_qelse_and_4_nl;
  wire[0:0] modulo_add_14_qelse_and_5_nl;
  wire[32:0] acc_14_nl;
  wire[33:0] nl_acc_14_nl;
  wire[31:0] modulo_add_15_qif_mux1h_2_nl;
  wire[0:0] modulo_add_15_qelse_and_nl;
  wire[0:0] modulo_add_15_qelse_or_nl;
  wire[0:0] modulo_add_15_qelse_and_5_nl;
  wire[0:0] modulo_add_15_qelse_and_6_nl;
  wire[0:0] modulo_add_15_qelse_and_7_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_nor_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_nor_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_5_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_and_5_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_1_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_1_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_2_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_2_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_and_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_3_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_3_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_1_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_and_1_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_4_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_4_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_2_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_and_2_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_5_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_5_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_3_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_and_3_nl;
  wire[0:0] butterFly1_f1_butterFly1_f1_and_6_nl;
  wire[0:0] butterFly1_16_f1_butterFly1_16_f1_and_6_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_4_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_and_4_nl;
  wire[0:0] INNER_LOOP1_mux_nl;
  wire[0:0] INNER_LOOP1_mux_4_nl;
  wire[0:0] INNER_LOOP1_mux_5_nl;
  wire[0:0] INNER_LOOP1_mux_6_nl;
  wire[0:0] butterFly1_15_mux_9_nl;
  wire[0:0] butterFly1_15_mux1h_47_nl;
  wire[0:0] butterFly2_15_mux1h_3_nl;
  wire[0:0] butterFly1_15_mux_10_nl;
  wire[6:0] STAGE_LOOP_base_STAGE_LOOP_base_mux_nl;
  wire[0:0] INNER_LOOP2_r_or_nl;
  wire[32:0] acc_18_nl;
  wire[33:0] nl_acc_18_nl;
  wire[31:0] modulo_add_2_qif_mux1h_2_nl;
  wire[0:0] modulo_add_23_qelse_and_nl;
  wire[0:0] modulo_add_23_qelse_or_1_nl;
  wire[0:0] modulo_add_23_qelse_and_4_nl;
  wire[0:0] modulo_add_23_qelse_and_5_nl;
  wire[32:0] acc_22_nl;
  wire[33:0] nl_acc_22_nl;
  wire[31:0] modulo_add_3_qif_mux1h_2_nl;
  wire[0:0] modulo_add_24_qelse_and_nl;
  wire[0:0] modulo_add_24_qelse_or_1_nl;
  wire[0:0] modulo_add_24_qelse_and_4_nl;
  wire[0:0] modulo_add_24_qelse_and_5_nl;
  wire[32:0] acc_26_nl;
  wire[33:0] nl_acc_26_nl;
  wire[31:0] modulo_add_4_qif_mux1h_2_nl;
  wire[0:0] modulo_add_25_qelse_and_nl;
  wire[0:0] modulo_add_25_qelse_or_1_nl;
  wire[0:0] modulo_add_25_qelse_and_4_nl;
  wire[0:0] modulo_add_25_qelse_and_5_nl;
  wire[32:0] acc_30_nl;
  wire[33:0] nl_acc_30_nl;
  wire[31:0] modulo_add_5_qif_mux1h_2_nl;
  wire[0:0] modulo_add_26_qelse_and_nl;
  wire[0:0] modulo_add_26_qelse_or_nl;
  wire[0:0] modulo_add_26_qelse_and_5_nl;
  wire[0:0] modulo_add_26_qelse_and_6_nl;
  wire[0:0] modulo_add_26_qelse_and_7_nl;
  wire[32:0] acc_34_nl;
  wire[33:0] nl_acc_34_nl;
  wire[31:0] modulo_add_6_qif_mux1h_2_nl;
  wire[0:0] modulo_add_27_qelse_and_nl;
  wire[0:0] modulo_add_27_qelse_or_nl;
  wire[0:0] modulo_add_27_qelse_and_5_nl;
  wire[0:0] modulo_add_27_qelse_and_6_nl;
  wire[0:0] modulo_add_27_qelse_and_7_nl;
  wire[32:0] acc_38_nl;
  wire[33:0] nl_acc_38_nl;
  wire[31:0] modulo_add_7_qif_mux1h_2_nl;
  wire[0:0] modulo_add_28_qelse_and_nl;
  wire[0:0] modulo_add_28_qelse_or_nl;
  wire[0:0] modulo_add_28_qelse_and_5_nl;
  wire[0:0] modulo_add_28_qelse_and_6_nl;
  wire[0:0] modulo_add_28_qelse_and_7_nl;
  wire[32:0] acc_42_nl;
  wire[33:0] nl_acc_42_nl;
  wire[31:0] modulo_add_8_qif_mux1h_2_nl;
  wire[0:0] modulo_add_29_qelse_and_nl;
  wire[0:0] modulo_add_29_qelse_or_nl;
  wire[0:0] modulo_add_29_qelse_and_5_nl;
  wire[0:0] modulo_add_29_qelse_and_6_nl;
  wire[0:0] modulo_add_29_qelse_and_7_nl;
  wire[32:0] acc_46_nl;
  wire[33:0] nl_acc_46_nl;
  wire[31:0] modulo_add_9_qif_mux1h_2_nl;
  wire[0:0] modulo_add_30_qelse_and_nl;
  wire[0:0] modulo_add_30_qelse_or_nl;
  wire[0:0] modulo_add_30_qelse_and_5_nl;
  wire[0:0] modulo_add_30_qelse_and_6_nl;
  wire[0:0] modulo_add_30_qelse_and_7_nl;
  wire[32:0] acc_49_nl;
  wire[33:0] nl_acc_49_nl;
  wire[31:0] modulo_add_qif_mux1h_2_nl;
  wire[0:0] modulo_add_31_qelse_and_nl;
  wire[0:0] modulo_add_31_qelse_or_nl;
  wire[0:0] modulo_add_31_qelse_and_5_nl;
  wire[0:0] modulo_add_31_qelse_and_6_nl;
  wire[0:0] modulo_add_31_qelse_and_7_nl;
  wire[0:0] modulo_sub_16_qelse_or_nl;
  wire[0:0] modulo_sub_17_qelse_or_nl;
  wire[0:0] modulo_sub_18_qelse_or_nl;
  wire[0:0] modulo_sub_19_qelse_or_nl;
  wire[0:0] modulo_sub_20_qelse_or_nl;
  wire[0:0] modulo_sub_21_qelse_or_nl;
  wire[0:0] modulo_sub_22_qelse_or_nl;
  wire[0:0] modulo_sub_23_qelse_or_nl;
  wire[0:0] modulo_sub_24_qelse_or_nl;
  wire[0:0] modulo_sub_25_qelse_or_nl;
  wire[0:0] modulo_sub_26_qelse_or_nl;
  wire[0:0] modulo_sub_27_qelse_or_nl;
  wire[0:0] modulo_sub_28_qelse_or_nl;
  wire[0:0] modulo_sub_29_qelse_or_nl;
  wire[0:0] modulo_sub_30_qelse_or_nl;
  wire[0:0] modulo_sub_31_qelse_or_nl;
  wire[0:0] INNER_LOOP1_mux_7_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_nor_nl;
  wire[0:0] butterFly2_16_f1_butterFly2_16_f1_nor_nl;
  wire[0:0] butterFly2_f1_butterFly2_f1_and_6_nl;
  wire[31:0] mult_15_if_acc_nl;
  wire[32:0] nl_mult_15_if_acc_nl;
  wire[32:0] mult_31_acc_1_nl;
  wire[33:0] nl_mult_31_acc_1_nl;
  wire[31:0] mult_14_if_acc_nl;
  wire[32:0] nl_mult_14_if_acc_nl;
  wire[32:0] mult_30_acc_1_nl;
  wire[33:0] nl_mult_30_acc_1_nl;
  wire[31:0] mult_13_if_acc_nl;
  wire[32:0] nl_mult_13_if_acc_nl;
  wire[32:0] mult_29_acc_1_nl;
  wire[33:0] nl_mult_29_acc_1_nl;
  wire[31:0] mult_12_if_acc_nl;
  wire[32:0] nl_mult_12_if_acc_nl;
  wire[32:0] mult_28_acc_1_nl;
  wire[33:0] nl_mult_28_acc_1_nl;
  wire[31:0] mult_11_if_acc_nl;
  wire[32:0] nl_mult_11_if_acc_nl;
  wire[32:0] mult_27_acc_1_nl;
  wire[33:0] nl_mult_27_acc_1_nl;
  wire[31:0] mult_10_if_acc_nl;
  wire[32:0] nl_mult_10_if_acc_nl;
  wire[32:0] mult_26_acc_1_nl;
  wire[33:0] nl_mult_26_acc_1_nl;
  wire[31:0] mult_9_if_acc_nl;
  wire[32:0] nl_mult_9_if_acc_nl;
  wire[32:0] mult_25_acc_1_nl;
  wire[33:0] nl_mult_25_acc_1_nl;
  wire[31:0] mult_8_if_acc_nl;
  wire[32:0] nl_mult_8_if_acc_nl;
  wire[32:0] mult_24_acc_1_nl;
  wire[33:0] nl_mult_24_acc_1_nl;
  wire[31:0] mult_7_if_acc_nl;
  wire[32:0] nl_mult_7_if_acc_nl;
  wire[32:0] mult_23_acc_1_nl;
  wire[33:0] nl_mult_23_acc_1_nl;
  wire[31:0] mult_6_if_acc_nl;
  wire[32:0] nl_mult_6_if_acc_nl;
  wire[32:0] mult_22_acc_1_nl;
  wire[33:0] nl_mult_22_acc_1_nl;
  wire[31:0] mult_5_if_acc_nl;
  wire[32:0] nl_mult_5_if_acc_nl;
  wire[32:0] mult_21_acc_1_nl;
  wire[33:0] nl_mult_21_acc_1_nl;
  wire[31:0] mult_4_if_acc_nl;
  wire[32:0] nl_mult_4_if_acc_nl;
  wire[32:0] mult_20_acc_1_nl;
  wire[33:0] nl_mult_20_acc_1_nl;
  wire[31:0] mult_3_if_acc_nl;
  wire[32:0] nl_mult_3_if_acc_nl;
  wire[32:0] mult_19_acc_1_nl;
  wire[33:0] nl_mult_19_acc_1_nl;
  wire[31:0] mult_2_if_acc_nl;
  wire[32:0] nl_mult_2_if_acc_nl;
  wire[32:0] mult_18_acc_1_nl;
  wire[33:0] nl_mult_18_acc_1_nl;
  wire[31:0] mult_1_if_acc_nl;
  wire[32:0] nl_mult_1_if_acc_nl;
  wire[32:0] mult_17_acc_1_nl;
  wire[33:0] nl_mult_17_acc_1_nl;
  wire[31:0] mult_if_acc_nl;
  wire[32:0] nl_mult_if_acc_nl;
  wire[32:0] mult_16_acc_1_nl;
  wire[33:0] nl_mult_16_acc_1_nl;
  wire[0:0] nor_62_nl;
  wire[0:0] or_325_nl;
  wire[0:0] nor_56_nl;
  wire[0:0] or_347_nl;
  wire[0:0] and_8934_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] or_409_nl;
  wire[0:0] or_408_nl;
  wire[0:0] or_419_nl;
  wire[0:0] nor_52_nl;
  wire[0:0] or_427_nl;
  wire[0:0] or_429_nl;
  wire[0:0] or_447_nl;
  wire[0:0] mux_69_nl;
  wire[0:0] or_445_nl;
  wire[0:0] or_457_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] or_332_nl;
  wire[0:0] or_331_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] or_359_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] or_357_nl;
  wire[0:0] nor_3_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] nor_7_nl;
  wire[0:0] nor_64_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] and_8944_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] and_8943_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] or_415_nl;
  wire[0:0] or_414_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] or_434_nl;
  wire[0:0] mux_74_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] nor_63_nl;
  wire[0:0] mux_77_nl;
  wire[0:0] and_8942_nl;
  wire[0:0] mux_86_nl;
  wire[0:0] mux_85_nl;
  wire[6:0] INNER_LOOP1_tw_and_nl;
  wire[5:0] INNER_LOOP2_tw_and_nl;
  wire[0:0] butterFly1_and_4_nl;
  wire[30:0] butterFly1_mux1h_nl;
  wire[0:0] butterFly1_or_nl;
  wire[0:0] butterFly1_1_and_4_nl;
  wire[0:0] butterFly1_1_mux_nl;
  wire[30:0] butterFly1_1_mux1h_nl;
  wire[0:0] butterFly1_1_and_1_nl;
  wire[0:0] butterFly1_2_and_4_nl;
  wire[0:0] butterFly1_2_mux_nl;
  wire[30:0] butterFly1_2_mux1h_nl;
  wire[0:0] butterFly1_2_and_1_nl;
  wire[0:0] butterFly1_3_and_4_nl;
  wire[0:0] butterFly1_3_mux_nl;
  wire[30:0] butterFly1_3_mux1h_nl;
  wire[0:0] butterFly1_3_and_1_nl;
  wire[0:0] butterFly1_4_and_4_nl;
  wire[0:0] butterFly1_4_mux_nl;
  wire[30:0] butterFly1_4_mux1h_nl;
  wire[0:0] butterFly1_4_and_1_nl;
  wire[0:0] butterFly1_5_and_4_nl;
  wire[0:0] butterFly1_5_mux_nl;
  wire[30:0] butterFly1_5_mux1h_nl;
  wire[0:0] butterFly1_5_and_1_nl;
  wire[0:0] butterFly1_6_and_4_nl;
  wire[0:0] butterFly1_6_mux_nl;
  wire[30:0] butterFly1_6_mux1h_nl;
  wire[0:0] butterFly1_6_and_1_nl;
  wire[0:0] butterFly1_7_and_4_nl;
  wire[0:0] butterFly1_7_mux_nl;
  wire[30:0] butterFly1_7_mux1h_nl;
  wire[0:0] butterFly1_7_and_1_nl;
  wire[0:0] butterFly1_8_and_4_nl;
  wire[0:0] butterFly1_8_mux_nl;
  wire[30:0] butterFly1_8_mux1h_nl;
  wire[0:0] butterFly1_8_and_1_nl;
  wire[0:0] butterFly1_9_and_4_nl;
  wire[0:0] butterFly1_9_mux_nl;
  wire[30:0] butterFly1_9_mux1h_272_nl;
  wire[0:0] butterFly1_9_and_1_nl;
  wire[0:0] butterFly1_10_and_4_nl;
  wire[0:0] butterFly1_10_mux_nl;
  wire[30:0] butterFly1_10_mux1h_nl;
  wire[0:0] butterFly1_10_and_1_nl;
  wire[0:0] butterFly1_11_and_4_nl;
  wire[0:0] butterFly1_11_mux_nl;
  wire[30:0] butterFly1_11_mux1h_nl;
  wire[0:0] butterFly1_11_and_1_nl;
  wire[0:0] butterFly1_12_and_4_nl;
  wire[0:0] butterFly1_12_mux_nl;
  wire[30:0] butterFly1_12_mux1h_nl;
  wire[0:0] butterFly1_12_and_1_nl;
  wire[0:0] butterFly1_13_and_4_nl;
  wire[0:0] butterFly1_13_mux_nl;
  wire[30:0] butterFly1_13_mux1h_nl;
  wire[0:0] butterFly1_13_and_1_nl;
  wire[0:0] butterFly1_14_and_4_nl;
  wire[0:0] butterFly1_14_mux_nl;
  wire[30:0] butterFly1_14_mux1h_nl;
  wire[0:0] butterFly1_14_and_1_nl;
  wire[0:0] butterFly1_15_and_5_nl;
  wire[30:0] butterFly1_15_mux1h_nl;
  wire[0:0] butterFly1_15_or_nl;
  wire[2:0] operator_20_false_mux_2_nl;
  wire[6:0] operator_20_false_mux1h_2_nl;
  wire[30:0] modulo_sub_15_qif_mux_2_nl;
  wire[30:0] modulo_sub_31_qif_mux_2_nl;
  wire[30:0] modulo_sub_7_qif_mux_2_nl;
  wire[30:0] modulo_sub_30_qif_mux_2_nl;
  wire[30:0] modulo_sub_39_qif_mux_2_nl;
  wire[30:0] modulo_sub_29_qif_mux_2_nl;
  wire[30:0] modulo_sub_6_qif_mux_2_nl;
  wire[30:0] modulo_sub_28_qif_mux_2_nl;
  wire[30:0] modulo_sub_38_qif_mux_2_nl;
  wire[30:0] modulo_sub_27_qif_mux_2_nl;
  wire[30:0] modulo_sub_5_qif_mux_2_nl;
  wire[30:0] modulo_sub_26_qif_mux_2_nl;
  wire[30:0] modulo_sub_37_qif_mux_2_nl;
  wire[30:0] modulo_sub_25_qif_mux_2_nl;
  wire[30:0] modulo_sub_4_qif_mux_2_nl;
  wire[30:0] modulo_sub_24_qif_mux_2_nl;
  wire[30:0] modulo_sub_36_qif_mux_2_nl;
  wire[30:0] modulo_sub_23_qif_mux_2_nl;
  wire[30:0] modulo_sub_3_qif_mux_2_nl;
  wire[30:0] modulo_sub_22_qif_mux_2_nl;
  wire[30:0] modulo_sub_35_qif_mux_2_nl;
  wire[30:0] modulo_sub_21_qif_mux_2_nl;
  wire[30:0] modulo_sub_2_qif_mux_2_nl;
  wire[30:0] modulo_sub_20_qif_mux_2_nl;
  wire[30:0] modulo_sub_34_qif_mux_2_nl;
  wire[30:0] modulo_sub_19_qif_mux_2_nl;
  wire[30:0] modulo_sub_1_qif_mux_2_nl;
  wire[30:0] modulo_sub_18_qif_mux_2_nl;
  wire[30:0] modulo_sub_33_qif_mux_2_nl;
  wire[30:0] modulo_sub_17_qif_mux_2_nl;
  wire[30:0] modulo_sub_qif_mux_2_nl;
  wire[30:0] modulo_sub_16_qif_mux_2_nl;
  wire[32:0] acc_50_nl;
  wire[33:0] nl_acc_50_nl;
  wire[31:0] butterFly1_mux1h_18_nl;
  wire[32:0] acc_51_nl;
  wire[33:0] nl_acc_51_nl;
  wire[31:0] butterFly1_1_mux1h_18_nl;
  wire[32:0] acc_52_nl;
  wire[33:0] nl_acc_52_nl;
  wire[31:0] butterFly1_2_mux1h_18_nl;
  wire[32:0] acc_53_nl;
  wire[33:0] nl_acc_53_nl;
  wire[31:0] butterFly1_3_mux1h_18_nl;
  wire[32:0] acc_54_nl;
  wire[33:0] nl_acc_54_nl;
  wire[31:0] butterFly1_4_mux1h_18_nl;
  wire[32:0] acc_55_nl;
  wire[33:0] nl_acc_55_nl;
  wire[31:0] butterFly1_5_mux1h_18_nl;
  wire[32:0] acc_56_nl;
  wire[33:0] nl_acc_56_nl;
  wire[31:0] butterFly1_6_mux1h_18_nl;
  wire[32:0] acc_57_nl;
  wire[33:0] nl_acc_57_nl;
  wire[31:0] butterFly1_7_mux1h_18_nl;
  wire[32:0] acc_58_nl;
  wire[33:0] nl_acc_58_nl;
  wire[31:0] butterFly1_8_mux1h_18_nl;
  wire[32:0] acc_59_nl;
  wire[33:0] nl_acc_59_nl;
  wire[31:0] butterFly1_9_mux1h_274_nl;
  wire[32:0] acc_60_nl;
  wire[33:0] nl_acc_60_nl;
  wire[31:0] butterFly1_10_mux1h_18_nl;
  wire[32:0] acc_61_nl;
  wire[33:0] nl_acc_61_nl;
  wire[31:0] butterFly1_11_mux1h_18_nl;
  wire[32:0] acc_62_nl;
  wire[33:0] nl_acc_62_nl;
  wire[31:0] butterFly1_12_mux1h_18_nl;
  wire[32:0] acc_63_nl;
  wire[33:0] nl_acc_63_nl;
  wire[31:0] butterFly1_13_mux1h_18_nl;
  wire[32:0] acc_64_nl;
  wire[33:0] nl_acc_64_nl;
  wire[31:0] butterFly1_14_mux1h_18_nl;
  wire[32:0] acc_65_nl;
  wire[33:0] nl_acc_65_nl;
  wire[31:0] butterFly1_15_mux1h_79_nl;
  wire[31:0] butterFly1_15_mux1h_80_nl;
  wire[31:0] butterFly1_14_mux1h_19_nl;
  wire[31:0] butterFly1_13_mux1h_19_nl;
  wire[31:0] butterFly1_12_mux1h_19_nl;
  wire[31:0] butterFly1_11_mux1h_19_nl;
  wire[31:0] butterFly1_10_mux1h_19_nl;
  wire[31:0] butterFly1_9_mux1h_275_nl;
  wire[31:0] butterFly1_8_mux1h_19_nl;
  wire[31:0] butterFly1_7_mux1h_19_nl;
  wire[31:0] butterFly1_6_mux1h_19_nl;
  wire[31:0] butterFly1_5_mux1h_19_nl;
  wire[31:0] butterFly1_4_mux1h_19_nl;
  wire[31:0] butterFly1_3_mux1h_19_nl;
  wire[31:0] butterFly1_2_mux1h_19_nl;
  wire[31:0] butterFly1_1_mux1h_19_nl;
  wire[31:0] butterFly1_mux1h_19_nl;
  wire[33:0] acc_82_nl;
  wire[34:0] nl_acc_82_nl;
  wire[31:0] modulo_add_1_mux1h_3_nl;
  wire[33:0] acc_83_nl;
  wire[34:0] nl_acc_83_nl;
  wire[31:0] modulo_add_10_mux1h_3_nl;
  wire[33:0] acc_84_nl;
  wire[34:0] nl_acc_84_nl;
  wire[31:0] modulo_add_54_mux1h_3_nl;
  wire[33:0] acc_85_nl;
  wire[34:0] nl_acc_85_nl;
  wire[31:0] modulo_add_48_mux1h_3_nl;
  wire[33:0] acc_86_nl;
  wire[34:0] nl_acc_86_nl;
  wire[31:0] modulo_add_33_mux1h_3_nl;
  wire[33:0] acc_87_nl;
  wire[34:0] nl_acc_87_nl;
  wire[31:0] modulo_add_34_mux1h_3_nl;
  wire[33:0] acc_88_nl;
  wire[34:0] nl_acc_88_nl;
  wire[31:0] modulo_add_6_mux1h_3_nl;
  wire[33:0] acc_89_nl;
  wire[34:0] nl_acc_89_nl;
  wire[31:0] modulo_add_50_mux1h_3_nl;
  wire[33:0] acc_90_nl;
  wire[34:0] nl_acc_90_nl;
  wire[31:0] modulo_add_51_mux1h_3_nl;
  wire[33:0] acc_91_nl;
  wire[34:0] nl_acc_91_nl;
  wire[31:0] modulo_add_14_mux1h_3_nl;
  wire[33:0] acc_92_nl;
  wire[34:0] nl_acc_92_nl;
  wire[31:0] modulo_add_36_mux1h_3_nl;
  wire[33:0] acc_93_nl;
  wire[34:0] nl_acc_93_nl;
  wire[31:0] modulo_add_52_mux1h_3_nl;
  wire[33:0] acc_94_nl;
  wire[34:0] nl_acc_94_nl;
  wire[31:0] modulo_add_41_mux1h_3_nl;
  wire[33:0] acc_95_nl;
  wire[34:0] nl_acc_95_nl;
  wire[31:0] modulo_add_2_mux1h_3_nl;
  wire[33:0] acc_96_nl;
  wire[34:0] nl_acc_96_nl;
  wire[31:0] modulo_add_53_mux1h_3_nl;
  wire[33:0] acc_97_nl;
  wire[34:0] nl_acc_97_nl;
  wire[31:0] modulo_add_55_mux1h_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_mult_t_mul_cmp_a;
  assign nl_mult_t_mul_cmp_a = MUX1HOT_v_32_4_2(z_out_43, z_out_59, z_out_49, z_out_35,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_b;
  assign nl_mult_t_mul_cmp_b = MUX1HOT_v_32_9_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]),
      (twiddle_h_rsc_0_11_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]), (twiddle_h_rsc_0_13_i_qa_d[31:0]),
      (twiddle_h_rsc_0_14_i_qa_d[31:0]), (twiddle_h_rsc_0_15_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_44_cse , mult_15_t_and_45_cse , mult_15_t_and_46_cse , mult_15_t_and_47_cse
      , mult_15_t_or_9_cse , mult_15_t_or_10_cse , mult_15_t_or_11_cse , mult_15_t_or_12_cse});
  wire [31:0] nl_mult_t_mul_cmp_1_a;
  assign nl_mult_t_mul_cmp_1_a = MUX1HOT_v_32_4_2(z_out_49, z_out_35, z_out_42, z_out_59,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_1_b;
  assign nl_mult_t_mul_cmp_1_b = MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]),
      (twiddle_h_rsc_0_14_i_qa_d[31:0]), {or_tmp_3231 , mult_15_t_and_40_cse , mult_15_t_and_41_cse
      , mult_15_t_and_42_cse , mult_15_t_and_43_cse});
  wire [31:0] nl_mult_t_mul_cmp_2_a;
  assign nl_mult_t_mul_cmp_2_a = MUX1HOT_v_32_4_2(z_out_42, z_out_50, z_out_41, z_out_32,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_2_b;
  assign nl_mult_t_mul_cmp_2_b = MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]),
      (twiddle_h_rsc_0_13_i_qa_d[31:0]), (twiddle_h_rsc_0_1_i_qa_d[31:0]), {or_tmp_3239
      , mult_15_t_and_36_cse , mult_15_t_and_37_cse , mult_15_t_and_38_cse , mult_15_t_and_39_cse
      , or_tmp_3242});
  wire [31:0] nl_mult_t_mul_cmp_3_a;
  assign nl_mult_t_mul_cmp_3_a = MUX1HOT_v_32_4_2(z_out_41, z_out_51, z_out_40, z_out_33,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_3631_nl;
  wire [31:0] nl_mult_t_mul_cmp_3_b;
  assign or_3631_nl = and_7109_cse | modulo_add_1_qelse_or_m1c;
  assign nl_mult_t_mul_cmp_3_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_12_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]),
      {or_3631_nl , or_tmp_3250 , and_7115_cse , or_tmp_3252});
  wire [31:0] nl_mult_t_mul_cmp_4_a;
  assign nl_mult_t_mul_cmp_4_a = MUX1HOT_v_32_4_2(z_out_40, z_out_52, z_out_39, z_out_34,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_t_or_8_nl;
  wire [31:0] nl_mult_t_mul_cmp_4_b;
  assign mult_15_t_or_8_nl = modulo_add_1_qelse_or_m1c | mult_15_t_and_49_cse;
  assign nl_mult_t_mul_cmp_4_b = MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]),
      (twiddle_h_rsc_0_11_i_qa_d[31:0]), (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]),
      (twiddle_h_rsc_0_3_i_qa_d[31:0]), {mult_15_t_or_8_nl , mult_15_t_and_29_cse
      , mult_15_t_and_30_cse , mult_15_t_and_31_cse , mult_15_t_and_32_cse , mult_15_t_and_51_cse
      , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_t_mul_cmp_5_a;
  assign nl_mult_t_mul_cmp_5_a = MUX1HOT_v_32_4_2(z_out_39, mult_t_mul_cmp_5_a_mx0w1,
      z_out_38, mult_t_mul_cmp_5_a_mx0w4, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_5_b;
  assign nl_mult_t_mul_cmp_5_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_10_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]),
      {modulo_add_1_qelse_or_m1c , or_tmp_3269 , and_7153_cse , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_6_a;
  assign nl_mult_t_mul_cmp_6_a = MUX1HOT_v_32_4_2(z_out_38, z_out_53, z_out_37, z_out_54,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_6_b;
  assign nl_mult_t_mul_cmp_6_b = MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_5_i_qa_d[31:0]),
      (twiddle_h_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c , or_tmp_3279
      , and_7173_cse , or_tmp_3242 , and_7090_cse});
  wire [31:0] nl_mult_t_mul_cmp_7_a;
  assign nl_mult_t_mul_cmp_7_a = MUX1HOT_v_32_4_2(z_out_37, z_out_55, z_out_48, z_out_56,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_7_b;
  assign nl_mult_t_mul_cmp_7_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_6_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]),
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , or_tmp_3252 , and_7109_cse});
  wire [31:0] nl_mult_t_mul_cmp_8_a;
  assign nl_mult_t_mul_cmp_8_a = MUX1HOT_v_32_4_2(z_out_48, z_out_57, z_out_47, z_out_58,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_8_b;
  assign nl_mult_t_mul_cmp_8_b = MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_3_i_qa_d[31:0]),
      (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_5_i_qa_d[31:0]), (twiddle_h_rsc_0_6_i_qa_d[31:0]),
      (twiddle_h_rsc_0_7_i_qa_d[31:0]), {mult_15_t_or_3_cse , mult_15_t_and_45_cse
      , mult_15_t_and_46_cse , mult_15_t_and_47_cse , mult_15_t_or_9_cse , mult_15_t_or_10_cse
      , mult_15_t_or_11_cse , mult_15_t_or_12_cse});
  wire [31:0] nl_mult_t_mul_cmp_9_a;
  assign nl_mult_t_mul_cmp_9_a = MUX1HOT_v_32_4_2(z_out_47, z_out_58, z_out_46, z_out_57,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_t_or_2_nl;
  wire [31:0] nl_mult_t_mul_cmp_9_b;
  assign mult_15_t_or_2_nl = modulo_add_1_qelse_or_m1c | mult_15_t_and_40_cse;
  assign nl_mult_t_mul_cmp_9_b = MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_6_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), {mult_15_t_or_2_nl , mult_15_t_and_41_cse
      , mult_15_t_and_42_cse , mult_15_t_and_43_cse , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_10_a;
  assign nl_mult_t_mul_cmp_10_a = MUX1HOT_v_32_4_2(z_out_46, z_out_56, z_out_36,
      z_out_55, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_10_b;
  assign nl_mult_t_mul_cmp_10_b = MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_5_i_qa_d[31:0]),
      (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), {mult_15_t_or_1_cse
      , mult_15_t_and_37_cse , mult_15_t_and_38_cse , mult_15_t_and_39_cse , or_tmp_3242
      , and_7090_cse});
  wire [31:0] nl_mult_t_mul_cmp_11_a;
  assign nl_mult_t_mul_cmp_11_a = MUX1HOT_v_32_4_2(z_out_36, z_out_54, mult_t_mul_cmp_11_a_mx0w3,
      z_out_53, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_3709_nl;
  wire [31:0] nl_mult_t_mul_cmp_11_b;
  assign or_3709_nl = and_7115_cse | modulo_add_1_qelse_or_m1c;
  assign nl_mult_t_mul_cmp_11_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]),
      {or_3709_nl , or_tmp_3250 , or_tmp_3252 , and_7109_cse});
  wire [31:0] nl_mult_t_mul_cmp_12_b;
  assign nl_mult_t_mul_cmp_12_b = MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_3_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]),
      (twiddle_h_rsc_0_11_i_qa_d[31:0]), {mult_15_t_or_cse , mult_15_t_and_30_cse
      , mult_15_t_and_31_cse , mult_15_t_and_32_cse , mult_15_t_and_49_cse , mult_15_t_and_51_cse
      , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_t_mul_cmp_13_a;
  assign nl_mult_t_mul_cmp_13_a = MUX1HOT_v_32_4_2(tmp_71_lpi_3_dfm_1, z_out_34,
      z_out_45, z_out_52, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_13_b;
  assign nl_mult_t_mul_cmp_13_b = MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]), {or_tmp_3345
      , or_tmp_3269 , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_14_a;
  assign nl_mult_t_mul_cmp_14_a = MUX1HOT_v_32_4_2(z_out_45, z_out_33, z_out_44,
      z_out_51, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_14_b;
  assign nl_mult_t_mul_cmp_14_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_13_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]),
      {or_tmp_3354 , or_tmp_3279 , or_tmp_3242 , and_7090_cse});
  wire [31:0] nl_mult_t_mul_cmp_15_a;
  assign nl_mult_t_mul_cmp_15_a = MUX1HOT_v_32_4_2(z_out_44, z_out_32, z_out_43,
      z_out_50, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_3747_nl;
  wire [31:0] nl_mult_t_mul_cmp_15_b;
  assign or_3747_nl = modulo_add_1_qelse_or_m1c | (fsm_output[7]);
  assign nl_mult_t_mul_cmp_15_b = MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_14_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]), {or_3747_nl
      , or_tmp_3252 , and_7109_cse});
  wire[0:0] mult_t_or_nl;
  wire [31:0] nl_mult_z_mul_cmp_a;
  assign mult_t_or_nl = (fsm_output[4]) | (fsm_output[9]);
  assign nl_mult_z_mul_cmp_a = MUX1HOT_v_32_3_2(z_out_43, z_out_59, z_out_49, {(fsm_output[2])
      , mult_t_or_nl , (fsm_output[7])});
  wire [31:0] nl_mult_z_mul_cmp_b;
  assign nl_mult_z_mul_cmp_b = MUX1HOT_v_32_9_2((twiddle_rsc_0_0_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]),
      (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]), (twiddle_rsc_0_11_i_qa_d[31:0]),
      (twiddle_rsc_0_12_i_qa_d[31:0]), (twiddle_rsc_0_13_i_qa_d[31:0]), (twiddle_rsc_0_14_i_qa_d[31:0]),
      (twiddle_rsc_0_15_i_qa_d[31:0]), {or_tmp_3231 , mult_15_t_and_44_cse , mult_15_t_and_45_cse
      , mult_15_t_and_46_cse , mult_15_t_and_47_cse , mult_15_t_and_48_cse , mult_15_t_and_50_cse
      , mult_15_t_and_52_cse , mult_15_t_and_54_cse});
  wire [31:0] nl_mult_z_mul_cmp_1_a;
  assign nl_mult_z_mul_cmp_1_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_1_z[63:32]), (mult_t_mul_cmp_11_z[63:32]),
      (mult_t_mul_cmp_12_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_1_b;
  assign nl_mult_z_mul_cmp_1_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_2_a;
  assign nl_mult_z_mul_cmp_2_a = MUX1HOT_v_32_4_2(z_out_49, z_out_35, z_out_43, z_out_57,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_2_b;
  assign nl_mult_z_mul_cmp_2_b = MUX_v_32_2_2((twiddle_rsc_0_0_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]),
      fsm_output[9]);
  wire [31:0] nl_mult_z_mul_cmp_3_a;
  assign nl_mult_z_mul_cmp_3_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_2_z[63:32]), (mult_t_mul_cmp_5_z[63:32]),
      (mult_t_mul_cmp_6_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_3_b;
  assign nl_mult_z_mul_cmp_3_b = p_sva;
  wire[0:0] mult_14_t_or_nl;
  wire [31:0] nl_mult_z_mul_cmp_4_a;
  assign mult_14_t_or_nl = (fsm_output[2]) | (fsm_output[7]);
  assign nl_mult_z_mul_cmp_4_a = MUX1HOT_v_32_3_2(z_out_42, z_out_50, mult_t_mul_cmp_5_a_mx0w4,
      {mult_14_t_or_nl , (fsm_output[4]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_4_b;
  assign nl_mult_z_mul_cmp_4_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]),
      (twiddle_rsc_0_14_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_40_cse , mult_15_t_and_41_cse , mult_15_t_and_42_cse , mult_15_t_and_43_cse
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_5_a;
  assign nl_mult_z_mul_cmp_5_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_3_z[63:32]), (mult_t_mul_cmp_12_z[63:32]),
      (mult_t_mul_cmp_13_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_5_b;
  assign nl_mult_z_mul_cmp_5_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_6_a;
  assign nl_mult_z_mul_cmp_6_a = MUX1HOT_v_32_4_2(z_out_41, z_out_51, z_out_47, z_out_35,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_6_b;
  assign nl_mult_z_mul_cmp_6_b = MUX1HOT_v_32_12_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_3_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]), (twiddle_rsc_0_6_i_qa_d[31:0]),
      (twiddle_rsc_0_7_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]), (twiddle_rsc_0_13_i_qa_d[31:0]),
      (twiddle_rsc_0_14_i_qa_d[31:0]), (twiddle_rsc_0_15_i_qa_d[31:0]), {mult_15_t_or_3_cse
      , mult_15_t_and_45_cse , mult_15_t_and_46_cse , mult_15_t_and_47_cse , mult_15_t_and_48_cse
      , mult_15_t_and_50_cse , mult_15_t_and_52_cse , mult_15_t_and_54_cse , mult_15_t_and_49_cse
      , mult_15_t_and_51_cse , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_7_a;
  assign nl_mult_z_mul_cmp_7_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_4_z[63:32]), (mult_t_mul_cmp_2_z[63:32]),
      (mult_t_mul_cmp_3_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_7_b;
  assign nl_mult_z_mul_cmp_7_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_8_a;
  assign nl_mult_z_mul_cmp_8_a = MUX1HOT_v_32_4_2(z_out_40, z_out_52, z_out_44, z_out_55,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_8_b;
  assign nl_mult_z_mul_cmp_8_b = MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]),
      {or_tmp_3354 , or_tmp_3279 , or_tmp_3242 , and_7090_cse});
  wire [31:0] nl_mult_z_mul_cmp_9_a;
  assign nl_mult_z_mul_cmp_9_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_5_z[63:32]), (mult_t_mul_cmp_10_z[63:32]),
      (mult_t_mul_cmp_11_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_9_b;
  assign nl_mult_z_mul_cmp_9_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_10_a;
  assign nl_mult_z_mul_cmp_10_a = MUX1HOT_v_32_4_2(z_out_39, mult_t_mul_cmp_5_a_mx0w1,
      z_out_48, z_out_58, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_10_b;
  assign nl_mult_z_mul_cmp_10_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]),
      (twiddle_rsc_0_6_i_qa_d[31:0]), (twiddle_rsc_0_7_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , mult_15_t_and_49_cse , mult_15_t_and_51_cse , mult_15_t_and_53_cse
      , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_11_a;
  assign nl_mult_z_mul_cmp_11_a = MUX_v_32_2_2((mult_t_mul_cmp_6_z[63:32]), (mult_t_mul_cmp_7_z[63:32]),
      fsm_output[9]);
  wire [31:0] nl_mult_z_mul_cmp_11_b;
  assign nl_mult_z_mul_cmp_11_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_12_a;
  assign nl_mult_z_mul_cmp_12_a = MUX1HOT_v_32_4_2(z_out_38, z_out_53, z_out_45,
      z_out_34, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_z_or_3_nl;
  wire[0:0] mult_15_z_or_6_nl;
  wire [31:0] nl_mult_z_mul_cmp_12_b;
  assign mult_15_z_or_3_nl = or_tmp_3345 | mult_15_t_and_49_cse;
  assign mult_15_z_or_6_nl = or_tmp_3269 | mult_15_t_and_53_cse;
  assign nl_mult_z_mul_cmp_12_b = MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_3_i_qa_d[31:0]),
      {mult_15_z_or_3_nl , mult_15_z_or_6_nl , mult_15_t_and_51_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_13_a;
  assign nl_mult_z_mul_cmp_13_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_7_z[63:32]), (mult_t_mul_cmp_1_z[63:32]),
      (mult_t_mul_cmp_2_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_13_b;
  assign nl_mult_z_mul_cmp_13_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_14_a;
  assign nl_mult_z_mul_cmp_14_a = MUX1HOT_v_32_4_2(z_out_37, z_out_55, z_out_41,
      z_out_50, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_z_or_5_nl;
  wire [31:0] nl_mult_z_mul_cmp_14_b;
  assign mult_15_z_or_5_nl = mult_15_t_and_38_cse | and_7109_cse;
  assign nl_mult_z_mul_cmp_14_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]),
      (twiddle_rsc_0_13_i_qa_d[31:0]), (twiddle_rsc_0_14_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_36_cse , mult_15_t_and_37_cse , mult_15_z_or_5_nl , mult_15_t_and_39_cse
      , or_tmp_3252});
  wire [31:0] nl_mult_z_mul_cmp_15_a;
  assign nl_mult_z_mul_cmp_15_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_8_z[63:32]), (mult_t_mul_cmp_13_z[63:32]),
      (mult_t_mul_cmp_14_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_15_b;
  assign nl_mult_z_mul_cmp_15_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_16_a;
  assign nl_mult_z_mul_cmp_16_a = MUX1HOT_v_32_4_2(z_out_48, z_out_57, z_out_46,
      z_out_32, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_z_or_2_nl;
  wire [31:0] nl_mult_z_mul_cmp_16_b;
  assign mult_15_z_or_2_nl = or_tmp_3239 | mult_15_t_and_40_cse;
  assign nl_mult_z_mul_cmp_16_b = MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_6_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), {mult_15_z_or_2_nl , mult_15_t_and_41_cse ,
      mult_15_t_and_42_cse , mult_15_t_and_43_cse , or_tmp_3242});
  wire [31:0] nl_mult_z_mul_cmp_17_a;
  assign nl_mult_z_mul_cmp_17_a = MUX_v_32_2_2((mult_t_mul_cmp_9_z[63:32]), (mult_t_mul_cmp_10_z[63:32]),
      fsm_output[9]);
  wire [31:0] nl_mult_z_mul_cmp_17_b;
  assign nl_mult_z_mul_cmp_17_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_18_a;
  assign nl_mult_z_mul_cmp_18_a = MUX1HOT_v_32_4_2(z_out_47, z_out_58, z_out_37,
      z_out_53, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_3884_nl;
  wire [31:0] nl_mult_z_mul_cmp_18_b;
  assign or_3884_nl = and_7173_cse | and_7109_cse;
  assign nl_mult_z_mul_cmp_18_b = MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]),
      {modulo_add_1_qelse_or_m1c , or_tmp_3279 , or_3884_nl , or_tmp_3252});
  wire [31:0] nl_mult_z_mul_cmp_19_a;
  assign nl_mult_z_mul_cmp_19_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_10_z[63:32]),
      (mult_t_mul_cmp_4_z[63:32]), (mult_t_mul_cmp_5_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_19_b;
  assign nl_mult_z_mul_cmp_19_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_20_a;
  assign nl_mult_z_mul_cmp_20_a = MUX1HOT_v_32_4_2(z_out_46, z_out_56, z_out_40,
      z_out_54, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_20_b;
  assign nl_mult_z_mul_cmp_20_b = MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_12_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c , or_tmp_3250 ,
      and_7115_cse , or_tmp_3242 , and_7090_cse});
  wire [31:0] nl_mult_z_mul_cmp_21_a;
  assign nl_mult_z_mul_cmp_21_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_11_z[63:32]),
      (mult_t_mul_cmp_14_z[63:32]), (mult_t_mul_cmp_15_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_21_b;
  assign nl_mult_z_mul_cmp_21_b = p_sva;
  wire[0:0] mult_5_t_or_nl;
  wire [31:0] nl_mult_z_mul_cmp_22_a;
  assign mult_5_t_or_nl = (fsm_output[2]) | (fsm_output[7]);
  assign nl_mult_z_mul_cmp_22_a = MUX1HOT_v_32_3_2(z_out_36, z_out_54, z_out_51,
      {mult_5_t_or_nl , (fsm_output[4]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_22_b;
  assign nl_mult_z_mul_cmp_22_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]),
      (twiddle_rsc_0_13_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]), {mult_15_t_or_1_cse
      , mult_15_t_and_37_cse , mult_15_t_and_38_cse , mult_15_t_and_39_cse , or_tmp_3242
      , and_7090_cse});
  wire [31:0] nl_mult_z_mul_cmp_23_a;
  assign nl_mult_z_mul_cmp_23_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_12_z[63:32]),
      (mult_t_mul_cmp_3_z[63:32]), (mult_t_mul_cmp_4_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_23_b;
  assign nl_mult_z_mul_cmp_23_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_24_b;
  assign nl_mult_z_mul_cmp_24_b = MUX1HOT_v_32_8_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_3_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]),
      (twiddle_rsc_0_11_i_qa_d[31:0]), {mult_15_t_or_cse , mult_15_t_and_30_cse ,
      mult_15_t_and_31_cse , mult_15_t_and_32_cse , mult_15_t_and_49_cse , mult_15_t_and_51_cse
      , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_25_a;
  assign nl_mult_z_mul_cmp_25_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_13_z[63:32]),
      (mult_t_mul_cmp_8_z[63:32]), (mult_t_mul_cmp_9_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_25_b;
  assign nl_mult_z_mul_cmp_25_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_26_a;
  assign nl_mult_z_mul_cmp_26_a = MUX1HOT_v_32_4_2(tmp_71_lpi_3_dfm_1, z_out_34,
      z_out_38, z_out_56, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_26_b;
  assign nl_mult_z_mul_cmp_26_b = MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_10_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_6_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c , or_tmp_3269 ,
      and_7153_cse , or_tmp_3252 , and_7109_cse});
  wire [31:0] nl_mult_z_mul_cmp_27_a;
  assign nl_mult_z_mul_cmp_27_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_14_z[63:32]),
      (mult_t_mul_cmp_7_z[63:32]), (mult_t_mul_cmp_8_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_27_b;
  assign nl_mult_z_mul_cmp_27_b = p_sva;
  wire[0:0] mult_2_t_or_nl;
  wire [31:0] nl_mult_z_mul_cmp_28_a;
  assign mult_2_t_or_nl = (fsm_output[4]) | (fsm_output[9]);
  assign nl_mult_z_mul_cmp_28_a = MUX1HOT_v_32_3_2(z_out_45, z_out_33, mult_t_mul_cmp_11_a_mx0w3,
      {(fsm_output[2]) , mult_2_t_or_nl , (fsm_output[7])});
  wire[0:0] or_3957_nl;
  wire [31:0] nl_mult_z_mul_cmp_28_b;
  assign or_3957_nl = and_7115_cse | and_7109_cse | modulo_add_1_qelse_or_m1c;
  assign nl_mult_z_mul_cmp_28_b = MUX1HOT_v_32_3_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_2_i_qa_d[31:0]), {or_3957_nl
      , or_tmp_3250 , or_tmp_3252});
  wire [31:0] nl_mult_z_mul_cmp_29_a;
  assign nl_mult_z_mul_cmp_29_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_15_z[63:32]),
      (mult_t_mul_cmp_z[63:32]), (mult_t_mul_cmp_1_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_29_b;
  assign nl_mult_z_mul_cmp_29_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_30_a;
  assign nl_mult_z_mul_cmp_30_a = MUX1HOT_v_32_4_2(z_out_44, z_out_32, z_out_39,
      z_out_52, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_30_b;
  assign nl_mult_z_mul_cmp_30_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]),
      (twiddle_rsc_0_11_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_29_cse , mult_15_t_and_30_cse , mult_15_t_and_31_cse , mult_15_t_and_32_cse
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_31_a;
  assign nl_mult_z_mul_cmp_31_a = MUX_v_32_2_2((mult_t_mul_cmp_z[63:32]), (mult_t_mul_cmp_15_z[63:32]),
      fsm_output[7]);
  wire [31:0] nl_mult_z_mul_cmp_31_b;
  assign nl_mult_z_mul_cmp_31_b = p_sva;
  wire [2:0] nl_operator_33_true_3_lshift_rg_s;
  assign nl_operator_33_true_3_lshift_rg_s = {1'b0 , (~ c_1_sva) , 1'b0};
  wire[2:0] operator_33_true_mux1h_nl;
  wire[0:0] operator_33_true_operator_33_true_or_nl;
  wire [3:0] nl_operator_33_true_1_lshift_rg_s;
  assign operator_33_true_mux1h_nl = MUX1HOT_v_3_3_2(z_out_61, operator_20_false_acc_cse_sva,
      ({2'b00 , (~ c_1_sva)}), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])});
  assign operator_33_true_operator_33_true_or_nl = (~ (fsm_output[3])) | (fsm_output[1])
      | (fsm_output[6]);
  assign nl_operator_33_true_1_lshift_rg_s = {operator_33_true_mux1h_nl , operator_33_true_operator_33_true_or_nl};
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0;
  assign nl_peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0 = ~(INNER_LOOP1_stage_0
      | INNER_LOOP1_stage_0_2 | INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_0
      | butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_3_0
      | butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_5_0 | INNER_LOOP1_stage_0_10);
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0;
  assign nl_peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0 = ~(INNER_LOOP1_stage_0
      | butterFly2_15_conc_2_itm_7_0 | butterFly2_15_conc_2_itm_8_0 | butterFly2_15_conc_2_itm_0
      | butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_3_0
      | butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_5_0 | INNER_LOOP2_stage_0_10);
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0;
  assign nl_peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0 = z_out_61[2];
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1;
  assign nl_peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 = ~ INNER_LOOP4_nor_tmp;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd32)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_7_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_7_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_6_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_6_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_5_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_5_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_4_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_4_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_3_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_3_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_2_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_2_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_1_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_1_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_31_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_30_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_29_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_28_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_27_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_26_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_25_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_24_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_23_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_22_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_21_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_20_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_19_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_18_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_17_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_16_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_15_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_14_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_13_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_12_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_11_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_10_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_9_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_8_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_7_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_6_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_5_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_4_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_3_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_2_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_1_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_0_obj (
      .ld(reg_xt_rsc_triosy_7_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_0_lz)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp (
      .a(nl_mult_t_mul_cmp_a[31:0]),
      .b(nl_mult_t_mul_cmp_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_1 (
      .a(nl_mult_t_mul_cmp_1_a[31:0]),
      .b(nl_mult_t_mul_cmp_1_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_1_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_2 (
      .a(nl_mult_t_mul_cmp_2_a[31:0]),
      .b(nl_mult_t_mul_cmp_2_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_2_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_3 (
      .a(nl_mult_t_mul_cmp_3_a[31:0]),
      .b(nl_mult_t_mul_cmp_3_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_3_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_4 (
      .a(nl_mult_t_mul_cmp_4_a[31:0]),
      .b(nl_mult_t_mul_cmp_4_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_4_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_5 (
      .a(nl_mult_t_mul_cmp_5_a[31:0]),
      .b(nl_mult_t_mul_cmp_5_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_5_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_6 (
      .a(nl_mult_t_mul_cmp_6_a[31:0]),
      .b(nl_mult_t_mul_cmp_6_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_6_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_7 (
      .a(nl_mult_t_mul_cmp_7_a[31:0]),
      .b(nl_mult_t_mul_cmp_7_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_7_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_8 (
      .a(nl_mult_t_mul_cmp_8_a[31:0]),
      .b(nl_mult_t_mul_cmp_8_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_8_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_9 (
      .a(nl_mult_t_mul_cmp_9_a[31:0]),
      .b(nl_mult_t_mul_cmp_9_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_9_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_10 (
      .a(nl_mult_t_mul_cmp_10_a[31:0]),
      .b(nl_mult_t_mul_cmp_10_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_10_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_11 (
      .a(nl_mult_t_mul_cmp_11_a[31:0]),
      .b(nl_mult_t_mul_cmp_11_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_11_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_12 (
      .a(mult_4_t_mux1h_1_rmff),
      .b(nl_mult_t_mul_cmp_12_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_12_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_13 (
      .a(nl_mult_t_mul_cmp_13_a[31:0]),
      .b(nl_mult_t_mul_cmp_13_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_13_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_14 (
      .a(nl_mult_t_mul_cmp_14_a[31:0]),
      .b(nl_mult_t_mul_cmp_14_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_14_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_15 (
      .a(nl_mult_t_mul_cmp_15_a[31:0]),
      .b(nl_mult_t_mul_cmp_15_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_15_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp (
      .a(nl_mult_z_mul_cmp_a[31:0]),
      .b(nl_mult_z_mul_cmp_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_1 (
      .a(nl_mult_z_mul_cmp_1_a[31:0]),
      .b(nl_mult_z_mul_cmp_1_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_1_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_2 (
      .a(nl_mult_z_mul_cmp_2_a[31:0]),
      .b(nl_mult_z_mul_cmp_2_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_2_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_3 (
      .a(nl_mult_z_mul_cmp_3_a[31:0]),
      .b(nl_mult_z_mul_cmp_3_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_3_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_4 (
      .a(nl_mult_z_mul_cmp_4_a[31:0]),
      .b(nl_mult_z_mul_cmp_4_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_4_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_5 (
      .a(nl_mult_z_mul_cmp_5_a[31:0]),
      .b(nl_mult_z_mul_cmp_5_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_5_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_6 (
      .a(nl_mult_z_mul_cmp_6_a[31:0]),
      .b(nl_mult_z_mul_cmp_6_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_6_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_7 (
      .a(nl_mult_z_mul_cmp_7_a[31:0]),
      .b(nl_mult_z_mul_cmp_7_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_7_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_8 (
      .a(nl_mult_z_mul_cmp_8_a[31:0]),
      .b(nl_mult_z_mul_cmp_8_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_8_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_9 (
      .a(nl_mult_z_mul_cmp_9_a[31:0]),
      .b(nl_mult_z_mul_cmp_9_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_9_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_10 (
      .a(nl_mult_z_mul_cmp_10_a[31:0]),
      .b(nl_mult_z_mul_cmp_10_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_10_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_11 (
      .a(nl_mult_z_mul_cmp_11_a[31:0]),
      .b(nl_mult_z_mul_cmp_11_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_11_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_12 (
      .a(nl_mult_z_mul_cmp_12_a[31:0]),
      .b(nl_mult_z_mul_cmp_12_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_12_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_13 (
      .a(nl_mult_z_mul_cmp_13_a[31:0]),
      .b(nl_mult_z_mul_cmp_13_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_13_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_14 (
      .a(nl_mult_z_mul_cmp_14_a[31:0]),
      .b(nl_mult_z_mul_cmp_14_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_14_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_15 (
      .a(nl_mult_z_mul_cmp_15_a[31:0]),
      .b(nl_mult_z_mul_cmp_15_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_15_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_16 (
      .a(nl_mult_z_mul_cmp_16_a[31:0]),
      .b(nl_mult_z_mul_cmp_16_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_16_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_17 (
      .a(nl_mult_z_mul_cmp_17_a[31:0]),
      .b(nl_mult_z_mul_cmp_17_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_17_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_18 (
      .a(nl_mult_z_mul_cmp_18_a[31:0]),
      .b(nl_mult_z_mul_cmp_18_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_18_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_19 (
      .a(nl_mult_z_mul_cmp_19_a[31:0]),
      .b(nl_mult_z_mul_cmp_19_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_19_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_20 (
      .a(nl_mult_z_mul_cmp_20_a[31:0]),
      .b(nl_mult_z_mul_cmp_20_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_20_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_21 (
      .a(nl_mult_z_mul_cmp_21_a[31:0]),
      .b(nl_mult_z_mul_cmp_21_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_21_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_22 (
      .a(nl_mult_z_mul_cmp_22_a[31:0]),
      .b(nl_mult_z_mul_cmp_22_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_22_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_23 (
      .a(nl_mult_z_mul_cmp_23_a[31:0]),
      .b(nl_mult_z_mul_cmp_23_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_23_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_24 (
      .a(mult_4_t_mux1h_1_rmff),
      .b(nl_mult_z_mul_cmp_24_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_24_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_25 (
      .a(nl_mult_z_mul_cmp_25_a[31:0]),
      .b(nl_mult_z_mul_cmp_25_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_25_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_26 (
      .a(nl_mult_z_mul_cmp_26_a[31:0]),
      .b(nl_mult_z_mul_cmp_26_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_26_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_27 (
      .a(nl_mult_z_mul_cmp_27_a[31:0]),
      .b(nl_mult_z_mul_cmp_27_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_27_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_28 (
      .a(nl_mult_z_mul_cmp_28_a[31:0]),
      .b(nl_mult_z_mul_cmp_28_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_28_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_29 (
      .a(nl_mult_z_mul_cmp_29_a[31:0]),
      .b(nl_mult_z_mul_cmp_29_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_29_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_30 (
      .a(nl_mult_z_mul_cmp_30_a[31:0]),
      .b(nl_mult_z_mul_cmp_30_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_30_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_31 (
      .a(nl_mult_z_mul_cmp_31_a[31:0]),
      .b(nl_mult_z_mul_cmp_31_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_31_z)
    );
  mgc_shift_bl_v5 #(.width_a(32'sd1),
  .signd_a(32'sd1),
  .width_s(32'sd3),
  .width_z(32'sd2)) operator_33_true_3_lshift_rg (
      .a(1'b1),
      .s(nl_operator_33_true_3_lshift_rg_s[2:0]),
      .z(operator_33_true_3_lshift_psp_1_0_sva_mx0w5)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd11)) operator_33_true_1_lshift_rg (
      .a(1'b1),
      .s(nl_operator_33_true_1_lshift_rg_s[3:0]),
      .z(z_out_60)
    );
  peaseNTT_core_wait_dp peaseNTT_core_wait_dp_inst (
      .yt_rsc_0_0_cgo_iro(or_553_rmff),
      .yt_rsc_0_0_i_clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .yt_rsc_0_16_cgo_iro(or_652_rmff),
      .yt_rsc_0_16_i_clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .yt_rsc_1_0_cgo_iro(or_718_rmff),
      .yt_rsc_1_0_i_clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .yt_rsc_1_16_cgo_iro(or_785_rmff),
      .yt_rsc_1_16_i_clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .yt_rsc_2_0_cgo_iro(or_851_rmff),
      .yt_rsc_2_0_i_clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .yt_rsc_2_16_cgo_iro(or_918_rmff),
      .yt_rsc_2_16_i_clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .yt_rsc_3_0_cgo_iro(or_984_rmff),
      .yt_rsc_3_0_i_clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .yt_rsc_3_16_cgo_iro(or_1051_rmff),
      .yt_rsc_3_16_i_clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .yt_rsc_4_0_cgo_iro(or_1117_rmff),
      .yt_rsc_4_0_i_clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .yt_rsc_4_16_cgo_iro(or_1216_rmff),
      .yt_rsc_4_16_i_clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .yt_rsc_5_0_cgo_iro(or_1282_rmff),
      .yt_rsc_5_0_i_clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .yt_rsc_5_16_cgo_iro(or_1349_rmff),
      .yt_rsc_5_16_i_clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .yt_rsc_6_0_cgo_iro(or_1415_rmff),
      .yt_rsc_6_0_i_clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .yt_rsc_6_16_cgo_iro(or_1482_rmff),
      .yt_rsc_6_16_i_clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .yt_rsc_7_0_cgo_iro(or_1548_rmff),
      .yt_rsc_7_0_i_clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .yt_rsc_7_16_cgo_iro(or_1615_rmff),
      .yt_rsc_7_16_i_clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .ensig_cgo_iro(or_3599_rmff),
      .ensig_cgo_iro_17(or_3759_rmff),
      .yt_rsc_0_0_cgo(reg_yt_rsc_0_0_cgo_cse),
      .yt_rsc_0_16_cgo(reg_yt_rsc_0_16_cgo_cse),
      .yt_rsc_1_0_cgo(reg_yt_rsc_1_0_cgo_cse),
      .yt_rsc_1_16_cgo(reg_yt_rsc_1_16_cgo_cse),
      .yt_rsc_2_0_cgo(reg_yt_rsc_2_0_cgo_cse),
      .yt_rsc_2_16_cgo(reg_yt_rsc_2_16_cgo_cse),
      .yt_rsc_3_0_cgo(reg_yt_rsc_3_0_cgo_cse),
      .yt_rsc_3_16_cgo(reg_yt_rsc_3_16_cgo_cse),
      .yt_rsc_4_0_cgo(reg_yt_rsc_4_0_cgo_cse),
      .yt_rsc_4_16_cgo(reg_yt_rsc_4_16_cgo_cse),
      .yt_rsc_5_0_cgo(reg_yt_rsc_5_0_cgo_cse),
      .yt_rsc_5_16_cgo(reg_yt_rsc_5_16_cgo_cse),
      .yt_rsc_6_0_cgo(reg_yt_rsc_6_0_cgo_cse),
      .yt_rsc_6_16_cgo(reg_yt_rsc_6_16_cgo_cse),
      .yt_rsc_7_0_cgo(reg_yt_rsc_7_0_cgo_cse),
      .yt_rsc_7_16_cgo(reg_yt_rsc_7_16_cgo_cse),
      .ensig_cgo(reg_ensig_cgo_cse),
      .mult_t_mul_cmp_en(mult_t_mul_cmp_en),
      .ensig_cgo_17(reg_ensig_cgo_17_cse),
      .mult_z_mul_cmp_1_en(mult_z_mul_cmp_1_en)
    );
  peaseNTT_core_core_fsm peaseNTT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .INNER_LOOP1_C_0_tr0(nl_peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0[0:0]),
      .INNER_LOOP2_C_0_tr0(nl_peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0[0:0]),
      .STAGE_LOOP_C_2_tr0(nl_peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0[0:0]),
      .INNER_LOOP3_C_0_tr0(INNER_LOOP4_nor_tmp),
      .INNER_LOOP4_C_0_tr0(and_dcpl_62),
      .INNER_LOOP4_C_0_tr1(nl_peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1[0:0])
    );
  assign or_4976_cse = (fsm_output[10]) | (fsm_output[0]);
  assign mux_1_nl = MUX_s_1_2_2(mux_tmp, or_tmp_26, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign or_322_nl = (butterFly2_15_conc_2_itm_9_2_1!=2'b00) | butterFly1_15_f1_equal_tmp_1_1
      | (~ butterFly1_15_conc_2_itm_0);
  assign mux_2_nl = MUX_s_1_2_2(mux_1_nl, or_322_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign or_337_nl = (butterFly1_15_conc_2_itm_9_2_1[0]) | butterFly1_15_conc_2_itm_9_0
      | (butterFly1_15_conc_2_itm_9_2_1[1]);
  assign mux_5_nl = MUX_s_1_2_2(not_tmp_29, or_tmp_40, or_337_nl);
  assign mux_6_nl = MUX_s_1_2_2(mux_5_nl, or_tmp_38, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_553_rmff = ((~ mux_2_nl) & (fsm_output[7])) | and_344_cse | ((~ mux_6_nl)
      & (fsm_output[2])) | and_346_cse;
  assign mux_8_nl = MUX_s_1_2_2(mux_tmp_7, or_tmp_48, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign or_344_nl = (butterFly2_15_conc_2_itm_9_2_1!=2'b00) | (~ nor_tmp_1);
  assign mux_9_nl = MUX_s_1_2_2(mux_8_nl, or_344_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign or_352_nl = (butterFly1_15_conc_2_itm_9_2_1[0]) | (~ butterFly1_15_conc_2_itm_9_0)
      | (butterFly1_15_conc_2_itm_9_2_1[1]);
  assign mux_10_nl = MUX_s_1_2_2(not_tmp_50, or_tmp_55, or_352_nl);
  assign mux_11_nl = MUX_s_1_2_2(mux_10_nl, or_tmp_53, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_652_rmff = ((~ mux_9_nl) & (fsm_output[7])) | and_344_cse | ((~ mux_11_nl)
      & (fsm_output[2])) | and_346_cse;
  assign or_356_nl = (butterFly2_15_conc_2_itm_9_2_1!=2'b01) | butterFly1_15_f1_equal_tmp_1_1
      | (~ butterFly1_15_conc_2_itm_0);
  assign mux_12_nl = MUX_s_1_2_2(or_tmp_26, mux_tmp, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_13_nl = MUX_s_1_2_2(or_356_nl, mux_12_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign or_360_nl = (~ (butterFly1_15_conc_2_itm_9_2_1[0])) | butterFly1_15_conc_2_itm_9_0
      | (butterFly1_15_conc_2_itm_9_2_1[1]);
  assign mux_16_nl = MUX_s_1_2_2(not_tmp_29, or_tmp_40, or_360_nl);
  assign mux_17_nl = MUX_s_1_2_2(or_tmp_64, mux_16_nl, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_718_rmff = ((~ mux_13_nl) & (fsm_output[7])) | and_715_cse | ((~ mux_17_nl)
      & (fsm_output[2])) | and_717_cse;
  assign or_367_nl = (butterFly2_15_conc_2_itm_9_2_1!=2'b01) | (~ nor_tmp_1);
  assign mux_18_nl = MUX_s_1_2_2(or_tmp_48, mux_tmp_7, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_19_nl = MUX_s_1_2_2(or_367_nl, mux_18_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign or_368_nl = (~ (butterFly1_15_conc_2_itm_9_2_1[0])) | (~ butterFly1_15_conc_2_itm_9_0)
      | (butterFly1_15_conc_2_itm_9_2_1[1]);
  assign mux_20_nl = MUX_s_1_2_2(not_tmp_50, or_tmp_55, or_368_nl);
  assign mux_21_nl = MUX_s_1_2_2(or_tmp_72, mux_20_nl, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_785_rmff = ((~ mux_19_nl) & (fsm_output[7])) | and_715_cse | ((~ mux_21_nl)
      & (fsm_output[2])) | and_717_cse;
  assign mux_23_nl = MUX_s_1_2_2(mux_tmp_22, or_tmp_75, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign or_372_nl = (butterFly2_15_conc_2_itm_9_2_1!=2'b10) | butterFly1_15_f1_equal_tmp_1_1
      | (~ butterFly1_15_conc_2_itm_0);
  assign mux_24_nl = MUX_s_1_2_2(mux_23_nl, or_372_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign mux_27_nl = MUX_s_1_2_2(not_tmp_67, or_tmp_86, or_383_cse);
  assign mux_28_nl = MUX_s_1_2_2(mux_27_nl, or_tmp_84, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_851_rmff = ((~ mux_24_nl) & (fsm_output[7])) | and_1022_cse | ((~ mux_28_nl)
      & (fsm_output[2])) | and_1024_cse;
  assign mux_30_nl = MUX_s_1_2_2(or_tmp_93, nor_tmp_15, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign nor_49_nl = ~((butterFly2_15_conc_2_itm_9_2_1[0]) | (~ nor_tmp_14));
  assign mux_31_nl = MUX_s_1_2_2(mux_30_nl, nor_49_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign nor_50_nl = ~(((~ (butterFly1_15_conc_2_itm_9_2_1[0])) & butterFly1_15_conc_2_itm_9_0
      & (butterFly1_15_conc_2_itm_9_2_1[1]) & INNER_LOOP1_stage_0_10) | nor_tmp_19);
  assign mux_32_nl = MUX_s_1_2_2(nor_50_nl, or_tmp_94, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_918_rmff = (mux_31_nl & (fsm_output[7])) | and_1022_cse | ((~ mux_32_nl)
      & (fsm_output[2])) | and_1024_cse;
  assign nand_1_nl = ~((butterFly2_15_conc_2_itm_9_2_1==2'b11) & (~ butterFly1_15_f1_equal_tmp_1_1)
      & butterFly1_15_conc_2_itm_0);
  assign mux_33_nl = MUX_s_1_2_2(or_tmp_75, mux_tmp_22, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_34_nl = MUX_s_1_2_2(nand_1_nl, mux_33_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign mux_38_nl = MUX_s_1_2_2(not_tmp_67, or_tmp_86, or_398_cse);
  assign mux_39_nl = MUX_s_1_2_2(or_tmp_102, mux_38_nl, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_984_rmff = ((~ mux_34_nl) & (fsm_output[7])) | and_1329_cse | ((~ mux_39_nl)
      & (fsm_output[2])) | and_1331_cse;
  assign mux_41_nl = MUX_s_1_2_2(nor_tmp_15, or_tmp_93, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_42_nl = MUX_s_1_2_2(nor_tmp_22, mux_41_nl, butterFly2_15_conc_itm_10_2_1[0]);
  assign or_404_nl = and_8913_cse | nor_tmp_19;
  assign mux_43_nl = MUX_s_1_2_2(and_8913_cse, or_404_nl, butterFly2_15_conc_2_itm_6_2_1[0]);
  assign or_1051_rmff = (mux_42_nl & (fsm_output[7])) | and_1329_cse | (mux_43_nl
      & (fsm_output[2])) | and_1331_cse;
  assign mux_46_nl = MUX_s_1_2_2(mux_tmp_45, or_tmp_29, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign or_406_nl = (butterFly2_15_conc_2_itm_8_2_1!=2'b00) | butterFly2_15_conc_2_itm_8_0
      | (~ butterFly1_15_conc_2_itm_9_0);
  assign mux_47_nl = MUX_s_1_2_2(mux_46_nl, or_406_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_51_nl = MUX_s_1_2_2(mux_tmp_50, or_tmp_120, or_383_cse);
  assign mux_52_nl = MUX_s_1_2_2(mux_51_nl, or_tmp_38, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1117_rmff = ((~ mux_47_nl) & (fsm_output[7])) | and_1636_cse | ((~ mux_52_nl)
      & (fsm_output[2])) | and_1638_cse;
  assign mux_54_nl = MUX_s_1_2_2(mux_tmp_53, or_tmp_50, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign or_426_nl = (butterFly2_15_conc_2_itm_8_2_1!=2'b00) | (~ nor_tmp_25);
  assign mux_55_nl = MUX_s_1_2_2(mux_54_nl, or_426_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_57_nl = MUX_s_1_2_2(or_tmp_133, mux_tmp_56, nor_27_cse);
  assign mux_58_nl = MUX_s_1_2_2(mux_57_nl, or_tmp_53, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1216_rmff = ((~ mux_55_nl) & (fsm_output[7])) | and_1636_cse | ((~ mux_58_nl)
      & (fsm_output[2])) | and_1638_cse;
  assign or_433_nl = (butterFly2_15_conc_2_itm_8_2_1!=2'b01) | butterFly2_15_conc_2_itm_8_0
      | (~ butterFly1_15_conc_2_itm_9_0);
  assign mux_59_nl = MUX_s_1_2_2(or_tmp_29, mux_tmp_45, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign mux_60_nl = MUX_s_1_2_2(or_433_nl, mux_59_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_63_nl = MUX_s_1_2_2(mux_tmp_50, or_tmp_120, or_398_cse);
  assign mux_64_nl = MUX_s_1_2_2(or_tmp_64, mux_63_nl, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1282_rmff = ((~ mux_60_nl) & (fsm_output[7])) | and_2007_cse | ((~ mux_64_nl)
      & (fsm_output[2])) | and_2009_cse;
  assign or_442_nl = (butterFly2_15_conc_2_itm_8_2_1!=2'b01) | (~ nor_tmp_25);
  assign mux_65_nl = MUX_s_1_2_2(or_tmp_50, mux_tmp_53, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign mux_66_nl = MUX_s_1_2_2(or_442_nl, mux_65_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_67_nl = MUX_s_1_2_2(or_tmp_133, mux_tmp_56, and_8912_cse);
  assign mux_68_nl = MUX_s_1_2_2(or_tmp_72, mux_67_nl, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1349_rmff = ((~ mux_66_nl) & (fsm_output[7])) | and_2007_cse | ((~ mux_68_nl)
      & (fsm_output[2])) | and_2009_cse;
  assign mux_71_nl = MUX_s_1_2_2(mux_tmp_70, or_tmp_77, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign or_444_nl = (butterFly2_15_conc_2_itm_8_2_1!=2'b10) | butterFly2_15_conc_2_itm_8_0
      | (~ butterFly1_15_conc_2_itm_9_0);
  assign mux_72_nl = MUX_s_1_2_2(mux_71_nl, or_444_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_75_nl = MUX_s_1_2_2(not_tmp_115, or_tmp_153, or_383_cse);
  assign mux_76_nl = MUX_s_1_2_2(mux_75_nl, or_tmp_84, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1415_rmff = ((~ mux_72_nl) & (fsm_output[7])) | and_2314_cse | ((~ mux_76_nl)
      & (fsm_output[2])) | and_2316_cse;
  assign mux_79_nl = MUX_s_1_2_2(mux_tmp_78, nor_tmp_14, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign nor_48_nl = ~((butterFly2_15_conc_2_itm_8_2_1[0]) | (~ nor_tmp_36));
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, nor_48_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_81_nl = MUX_s_1_2_2(and_8919_cse, or_tmp_160, nor_27_cse);
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, (~ or_tmp_94), butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1482_rmff = (mux_80_nl & (fsm_output[7])) | and_2314_cse | (mux_82_nl
      & (fsm_output[2])) | and_2316_cse;
  assign nand_nl = ~((butterFly2_15_conc_2_itm_8_2_1==2'b11) & (~ butterFly2_15_conc_2_itm_8_0)
      & butterFly1_15_conc_2_itm_9_0);
  assign mux_83_nl = MUX_s_1_2_2(or_tmp_77, mux_tmp_70, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign mux_84_nl = MUX_s_1_2_2(nand_nl, mux_83_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_87_nl = MUX_s_1_2_2(not_tmp_115, or_tmp_153, or_398_cse);
  assign mux_88_nl = MUX_s_1_2_2(or_tmp_102, mux_87_nl, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1548_rmff = ((~ mux_84_nl) & (fsm_output[7])) | and_2621_cse | ((~ mux_88_nl)
      & (fsm_output[2])) | and_2623_cse;
  assign mux_89_nl = MUX_s_1_2_2(nor_tmp_14, mux_tmp_78, butterFly2_15_conc_2_itm_8_2_1[0]);
  assign mux_90_nl = MUX_s_1_2_2(nor_tmp_46, mux_89_nl, butterFly2_15_conc_2_itm_9_2_1[0]);
  assign mux_91_nl = MUX_s_1_2_2(and_8919_cse, or_tmp_160, and_8912_cse);
  assign mux_92_nl = MUX_s_1_2_2(and_8913_cse, mux_91_nl, butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_1615_rmff = (mux_90_nl & (fsm_output[7])) | and_2621_cse | (mux_92_nl
      & (fsm_output[2])) | and_2623_cse;
  assign and_6824_rmff = INNER_LOOP1_stage_0 & or_dcpl_300;
  assign butterFly2_1_tw_butterFly2_1_tw_mux_rmff = MUX_v_7_2_2(INNER_LOOP3_r_11_4_sva_6_0,
      INNER_LOOP4_r_11_4_sva_6_0, fsm_output[9]);
  assign or_3498_rmff = (and_dcpl_173 & (fsm_output[7])) | and_6834_cse;
  assign or_3502_rmff = (and_dcpl_175 & (fsm_output[7])) | and_6843_cse;
  assign or_3506_rmff = (and_dcpl_175 & (operator_20_false_acc_cse_sva[0]) & (fsm_output[7]))
      | and_6852_cse;
  assign or_3510_rmff = (INNER_LOOP1_stage_0 & (operator_20_false_acc_cse_sva[2])
      & (fsm_output[7])) | (INNER_LOOP1_stage_0 & (fsm_output[9]));
  assign or_3514_rmff = (and_dcpl_173 & (operator_20_false_acc_cse_sva[2]) & (fsm_output[7]))
      | and_6834_cse;
  assign or_3518_rmff = (and_dcpl_175 & (operator_20_false_acc_cse_sva[2]) & (fsm_output[7]))
      | and_6843_cse;
  assign or_3522_rmff = (and_dcpl_175 & (operator_20_false_acc_cse_sva[0]) & (operator_20_false_acc_cse_sva[2])
      & (fsm_output[7])) | and_6852_cse;
  assign and_6895_rmff = INNER_LOOP1_stage_0 & or_dcpl_298;
  assign or_3599_rmff = ((butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_4_0
      | butterFly1_15_conc_2_itm_3_0) & or_dcpl_298) | ((INNER_LOOP1_stage_0_3 |
      INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_0) & (fsm_output[2])) | ((butterFly2_15_conc_2_itm_0
      | butterFly2_15_conc_2_itm_8_0 | butterFly2_15_conc_2_itm_7_0) & (fsm_output[4]));
  assign mult_15_t_and_49_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b00) &
      (fsm_output[9]);
  assign mult_15_t_and_51_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b01) &
      (fsm_output[9]);
  assign mult_15_t_and_53_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b10) &
      (fsm_output[9]);
  assign mult_15_t_and_55_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b11) &
      (fsm_output[9]);
  assign mult_15_t_and_44_cse = butterFly2_15_tw_equal_tmp_1 & (fsm_output[7]);
  assign butterFly2_7_tw_nor_cse = ~((operator_20_false_acc_cse_sva[2:1]!=2'b00));
  assign mult_15_t_and_45_cse = (operator_20_false_acc_cse_sva[0]) & butterFly2_7_tw_nor_cse
      & (fsm_output[7]);
  assign butterFly2_7_tw_nor_1_cse = ~((operator_20_false_acc_cse_sva[2]) | (operator_20_false_acc_cse_sva[0]));
  assign mult_15_t_and_46_cse = (operator_20_false_acc_cse_sva[1]) & butterFly2_7_tw_nor_1_cse
      & (fsm_output[7]);
  assign mult_15_t_and_47_cse = butterFly2_15_tw_equal_tmp_3_1 & (fsm_output[7]);
  assign butterFly2_7_tw_nor_2_cse = ~((operator_20_false_acc_cse_sva[1:0]!=2'b00));
  assign mult_15_t_and_48_cse = (operator_20_false_acc_cse_sva[2]) & butterFly2_7_tw_nor_2_cse
      & (fsm_output[7]);
  assign mult_15_t_and_50_cse = butterFly2_15_tw_equal_tmp_5_1 & (fsm_output[7]);
  assign mult_15_t_and_52_cse = butterFly2_15_tw_equal_tmp_6_1 & (fsm_output[7]);
  assign mult_15_t_and_54_cse = butterFly2_15_tw_equal_tmp_7_1 & (fsm_output[7]);
  assign mult_15_t_or_9_cse = mult_15_t_and_48_cse | mult_15_t_and_49_cse;
  assign mult_15_t_or_10_cse = mult_15_t_and_50_cse | mult_15_t_and_51_cse;
  assign mult_15_t_or_11_cse = mult_15_t_and_52_cse | mult_15_t_and_53_cse;
  assign mult_15_t_or_12_cse = mult_15_t_and_54_cse | mult_15_t_and_55_cse;
  assign mult_15_t_and_41_cse = (operator_20_false_acc_cse_sva[2:1]==2'b01) & (fsm_output[7]);
  assign mult_15_t_and_42_cse = (operator_20_false_acc_cse_sva[2:1]==2'b10) & (fsm_output[7]);
  assign mult_15_t_and_43_cse = (operator_20_false_acc_cse_sva[2:1]==2'b11) & (fsm_output[7]);
  assign mult_15_t_and_40_cse = butterFly2_7_tw_nor_cse & (fsm_output[7]);
  assign mult_15_t_and_37_cse = (operator_20_false_acc_cse_sva[0]) & (~ (operator_20_false_acc_cse_sva[2]))
      & (fsm_output[7]);
  assign mult_15_t_and_38_cse = (operator_20_false_acc_cse_sva[2]) & (~ (operator_20_false_acc_cse_sva[0]))
      & (fsm_output[7]);
  assign mult_15_t_and_39_cse = (operator_20_false_acc_cse_sva[2]) & (operator_20_false_acc_cse_sva[0])
      & (fsm_output[7]);
  assign mult_15_t_and_36_cse = butterFly2_7_tw_nor_1_cse & (fsm_output[7]);
  assign mult_15_t_and_30_cse = (operator_20_false_acc_cse_sva[1:0]==2'b01) & (fsm_output[7]);
  assign mult_15_t_and_31_cse = (operator_20_false_acc_cse_sva[1:0]==2'b10) & (fsm_output[7]);
  assign mult_15_t_and_32_cse = (operator_20_false_acc_cse_sva[1:0]==2'b11) & (fsm_output[7]);
  assign mult_15_t_and_29_cse = butterFly2_7_tw_nor_2_cse & (fsm_output[7]);
  assign mult_15_t_or_3_cse = modulo_add_1_qelse_or_m1c | mult_15_t_and_44_cse;
  assign mult_15_t_or_1_cse = modulo_add_1_qelse_or_m1c | mult_15_t_and_36_cse;
  assign mult_4_t_and_nl = butterFly1_15_f1_equal_tmp_1 & (fsm_output[2]);
  assign mult_4_t_and_1_nl = butterFly1_15_f1_equal_tmp_1_1 & (fsm_output[2]);
  assign mult_4_t_and_2_nl = butterFly1_15_f1_equal_tmp_2_1 & (fsm_output[2]);
  assign mult_4_t_and_3_nl = butterFly1_15_f1_equal_tmp_3_1 & (fsm_output[2]);
  assign mult_4_t_and_4_nl = butterFly1_15_f1_equal_tmp_4_1 & (fsm_output[2]);
  assign mult_4_t_and_5_nl = butterFly1_15_f1_equal_tmp_5_1 & (fsm_output[2]);
  assign mult_4_t_and_6_nl = butterFly1_15_f1_equal_tmp_6_1 & (fsm_output[2]);
  assign mult_4_t_and_7_nl = butterFly1_15_f1_equal_tmp_7_1 & (fsm_output[2]);
  assign mult_4_t_and_8_nl = butterFly1_15_f1_equal_tmp_1 & (fsm_output[4]);
  assign mult_4_t_and_9_nl = butterFly1_15_f1_equal_tmp_1_1 & (fsm_output[4]);
  assign mult_4_t_and_10_nl = butterFly1_15_f1_equal_tmp_2_1 & (fsm_output[4]);
  assign mult_4_t_and_11_nl = butterFly1_15_f1_equal_tmp_3_1 & (fsm_output[4]);
  assign mult_4_t_and_12_nl = butterFly1_15_f1_equal_tmp_4_1 & (fsm_output[4]);
  assign mult_4_t_and_13_nl = butterFly1_15_f1_equal_tmp_5_1 & (fsm_output[4]);
  assign mult_4_t_and_14_nl = butterFly1_15_f1_equal_tmp_6_1 & (fsm_output[4]);
  assign mult_4_t_and_15_nl = butterFly1_15_f1_equal_tmp_7_1 & (fsm_output[4]);
  assign mult_4_t_and_16_nl = butterFly2_15_f1_equal_tmp_1 & (fsm_output[7]);
  assign mult_4_t_and_17_nl = butterFly1_15_f1_equal_tmp_3_1 & (fsm_output[7]);
  assign mult_4_t_and_18_nl = butterFly1_15_f1_equal_tmp_4_1 & (fsm_output[7]);
  assign mult_4_t_and_19_nl = butterFly1_15_f1_equal_tmp_5_1 & (fsm_output[7]);
  assign mult_4_t_and_20_nl = butterFly1_15_f1_equal_tmp_6_1 & (fsm_output[7]);
  assign mult_4_t_and_21_nl = butterFly1_15_f1_equal_tmp_7_1 & (fsm_output[7]);
  assign mult_4_t_and_22_nl = butterFly1_15_f1_equal_tmp_1 & (fsm_output[7]);
  assign mult_4_t_and_23_nl = butterFly2_15_f1_equal_tmp_7_1 & (fsm_output[7]);
  assign mult_4_t_and_24_nl = butterFly2_15_f1_equal_tmp_1 & (fsm_output[9]);
  assign mult_4_t_and_25_nl = butterFly1_15_f1_equal_tmp_3_1 & (fsm_output[9]);
  assign mult_4_t_and_26_nl = butterFly1_15_f1_equal_tmp_4_1 & (fsm_output[9]);
  assign mult_4_t_and_27_nl = butterFly1_15_f1_equal_tmp_5_1 & (fsm_output[9]);
  assign mult_4_t_and_28_nl = butterFly1_15_f1_equal_tmp_6_1 & (fsm_output[9]);
  assign mult_4_t_and_29_nl = butterFly1_15_f1_equal_tmp_7_1 & (fsm_output[9]);
  assign mult_4_t_and_30_nl = butterFly1_15_f1_equal_tmp_1 & (fsm_output[9]);
  assign mult_4_t_and_31_nl = butterFly2_15_f1_equal_tmp_7_1 & (fsm_output[9]);
  assign mult_4_t_mux1h_1_rmff = MUX1HOT_v_32_32_2(xt_rsc_0_9_i_qa_d, xt_rsc_1_9_i_qa_d,
      xt_rsc_2_9_i_qa_d, xt_rsc_3_9_i_qa_d, xt_rsc_4_9_i_qa_d, xt_rsc_5_9_i_qa_d,
      xt_rsc_6_9_i_qa_d, xt_rsc_7_9_i_qa_d, yt_rsc_0_9_i_q_d, yt_rsc_1_9_i_q_d, yt_rsc_2_9_i_q_d,
      yt_rsc_3_9_i_q_d, yt_rsc_4_9_i_q_d, yt_rsc_5_9_i_q_d, yt_rsc_6_9_i_q_d, yt_rsc_7_9_i_q_d,
      xt_rsc_0_7_i_qa_d, xt_rsc_1_7_i_qa_d, xt_rsc_2_7_i_qa_d, xt_rsc_3_7_i_qa_d,
      xt_rsc_4_7_i_qa_d, xt_rsc_5_7_i_qa_d, xt_rsc_6_7_i_qa_d, xt_rsc_7_7_i_qa_d,
      yt_rsc_0_23_i_q_d, yt_rsc_1_23_i_q_d, yt_rsc_2_23_i_q_d, yt_rsc_3_23_i_q_d,
      yt_rsc_4_23_i_q_d, yt_rsc_5_23_i_q_d, yt_rsc_6_23_i_q_d, yt_rsc_7_23_i_q_d,
      {mult_4_t_and_nl , mult_4_t_and_1_nl , mult_4_t_and_2_nl , mult_4_t_and_3_nl
      , mult_4_t_and_4_nl , mult_4_t_and_5_nl , mult_4_t_and_6_nl , mult_4_t_and_7_nl
      , mult_4_t_and_8_nl , mult_4_t_and_9_nl , mult_4_t_and_10_nl , mult_4_t_and_11_nl
      , mult_4_t_and_12_nl , mult_4_t_and_13_nl , mult_4_t_and_14_nl , mult_4_t_and_15_nl
      , mult_4_t_and_16_nl , mult_4_t_and_17_nl , mult_4_t_and_18_nl , mult_4_t_and_19_nl
      , mult_4_t_and_20_nl , mult_4_t_and_21_nl , mult_4_t_and_22_nl , mult_4_t_and_23_nl
      , mult_4_t_and_24_nl , mult_4_t_and_25_nl , mult_4_t_and_26_nl , mult_4_t_and_27_nl
      , mult_4_t_and_28_nl , mult_4_t_and_29_nl , mult_4_t_and_30_nl , mult_4_t_and_31_nl});
  assign mult_15_t_or_cse = modulo_add_1_qelse_or_m1c | mult_15_t_and_29_cse;
  assign or_3759_rmff = ((butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_6_0
      | butterFly1_15_conc_2_itm_5_0) & or_dcpl_298) | ((butterFly2_15_conc_2_itm_1_0
      | butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_3_0) & modulo_add_1_qelse_or_m1c);
  assign modulo_add_1_qelse_or_m1c = (fsm_output[2]) | (fsm_output[4]);
  assign butterFly1_f1_nor_cse = ~((INNER_LOOP1_r_11_4_sva_6_0[6:5]!=2'b00));
  assign butterFly2_f1_nor_cse = ~((INNER_LOOP3_r_11_4_sva_6_0[6:5]!=2'b00));
  assign butterFly2_16_f1_nor_1_cse = ~((INNER_LOOP4_r_11_4_sva_6_0[6]) | (INNER_LOOP4_r_11_4_sva_6_0[4]));
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_cse = MUX_v_7_2_2(7'b0000000, (z_out_62[6:0]),
      (fsm_output[2]));
  assign modulo_sub_16_qelse_and_ssc = ~((z_out_126[31]) | (fsm_output[9]));
  assign modulo_sub_16_qelse_and_ssc_1 = (~ (z_out_111[31])) & (fsm_output[9]);
  assign modulo_sub_17_qelse_and_ssc = ~((z_out_116[31]) | (fsm_output[9]));
  assign modulo_sub_17_qelse_and_ssc_1 = (~ (z_out_112[31])) & (fsm_output[9]);
  assign modulo_sub_18_qelse_and_ssc = ~((z_out_123[31]) | (fsm_output[9]));
  assign modulo_sub_18_qelse_and_ssc_1 = (~ (z_out_113[31])) & (fsm_output[9]);
  assign modulo_sub_19_qelse_and_ssc = ~((z_out_124[31]) | (fsm_output[9]));
  assign modulo_sub_19_qelse_and_ssc_1 = (~ (z_out_114[31])) & (fsm_output[9]);
  assign modulo_sub_20_qelse_and_ssc = ~((z_out_125[31]) | (fsm_output[9]));
  assign modulo_sub_20_qelse_and_ssc_1 = (~ (z_out_115[31])) & (fsm_output[9]);
  assign modulo_sub_21_qelse_and_ssc = ~((z_out_111[31]) | (fsm_output[9]));
  assign modulo_sub_21_qelse_and_ssc_1 = (~ (z_out_116[31])) & (fsm_output[9]);
  assign modulo_sub_22_qelse_and_ssc = ~((z_out_112[31]) | (fsm_output[9]));
  assign modulo_sub_22_qelse_and_ssc_1 = (~ (z_out_117[31])) & (fsm_output[9]);
  assign modulo_sub_23_qelse_and_ssc = ~((z_out_113[31]) | (fsm_output[9]));
  assign modulo_sub_23_qelse_and_ssc_1 = (~ (z_out_118[31])) & (fsm_output[9]);
  assign modulo_sub_24_qelse_and_ssc = ~((z_out_114[31]) | (fsm_output[9]));
  assign modulo_sub_24_qelse_and_ssc_1 = (~ (z_out_119[31])) & (fsm_output[9]);
  assign modulo_sub_25_qelse_and_ssc = ~((z_out_115[31]) | (fsm_output[9]));
  assign modulo_sub_25_qelse_and_ssc_1 = (~ (z_out_120[31])) & (fsm_output[9]);
  assign modulo_sub_26_qelse_and_ssc = ~((z_out_117[31]) | (fsm_output[9]));
  assign modulo_sub_26_qelse_and_ssc_1 = (~ (z_out_121[31])) & (fsm_output[9]);
  assign modulo_sub_27_qelse_and_ssc = ~((z_out_118[31]) | (fsm_output[9]));
  assign modulo_sub_27_qelse_and_ssc_1 = (~ (z_out_122[31])) & (fsm_output[9]);
  assign modulo_sub_28_qelse_and_ssc = ~((z_out_119[31]) | (fsm_output[9]));
  assign modulo_sub_28_qelse_and_ssc_1 = (~ (z_out_123[31])) & (fsm_output[9]);
  assign modulo_sub_29_qelse_and_ssc = ~((z_out_120[31]) | (fsm_output[9]));
  assign modulo_sub_29_qelse_and_ssc_1 = (~ (z_out_124[31])) & (fsm_output[9]);
  assign modulo_sub_30_qelse_and_ssc = ~((z_out_121[31]) | (fsm_output[9]));
  assign modulo_sub_30_qelse_and_ssc_1 = (~ (z_out_125[31])) & (fsm_output[9]);
  assign modulo_sub_31_qelse_and_ssc = ~((z_out_122[31]) | (fsm_output[9]));
  assign modulo_sub_31_qelse_and_ssc_1 = (~ (z_out_126[31])) & (fsm_output[9]);
  assign butterFly2_16_f1_butterFly2_16_f1_and_6_cse = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b111);
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse = MUX_v_7_2_2(7'b0000000, (z_out_62[6:0]),
      (fsm_output[7]));
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse = MUX_v_7_2_2(7'b0000000, (z_out_62[6:0]),
      (fsm_output[9]));
  assign or_383_cse = (butterFly1_15_conc_2_itm_9_2_1[0]) | butterFly1_15_conc_2_itm_9_0;
  assign or_398_cse = (~ (butterFly1_15_conc_2_itm_9_2_1[0])) | butterFly1_15_conc_2_itm_9_0;
  assign and_8913_cse = (butterFly1_15_conc_2_itm_9_2_1[0]) & butterFly1_15_conc_2_itm_9_0
      & (butterFly1_15_conc_2_itm_9_2_1[1]) & INNER_LOOP1_stage_0_10;
  assign nor_27_cse = ~((butterFly1_15_conc_2_itm_9_2_1[0]) | (~ butterFly1_15_conc_2_itm_9_0));
  assign and_8912_cse = (butterFly1_15_conc_2_itm_9_2_1[0]) & butterFly1_15_conc_2_itm_9_0;
  assign mult_t_mul_cmp_5_a_mx0w1 = MUX1HOT_v_32_8_2(yt_rsc_0_23_i_q_d, yt_rsc_1_23_i_q_d,
      yt_rsc_2_23_i_q_d, yt_rsc_3_23_i_q_d, yt_rsc_4_23_i_q_d, yt_rsc_5_23_i_q_d,
      yt_rsc_6_23_i_q_d, yt_rsc_7_23_i_q_d, {butterFly1_15_f1_equal_tmp_1 , butterFly1_15_f1_equal_tmp_1_1
      , butterFly1_15_f1_equal_tmp_2_1 , butterFly1_15_f1_equal_tmp_3_1 , butterFly1_15_f1_equal_tmp_4_1
      , butterFly1_15_f1_equal_tmp_5_1 , butterFly1_15_f1_equal_tmp_6_1 , butterFly1_15_f1_equal_tmp_7_1});
  assign mult_t_mul_cmp_5_a_mx0w4 = MUX1HOT_v_32_8_2(yt_rsc_0_9_i_q_d, yt_rsc_1_9_i_q_d,
      yt_rsc_2_9_i_q_d, yt_rsc_3_9_i_q_d, yt_rsc_4_9_i_q_d, yt_rsc_5_9_i_q_d, yt_rsc_6_9_i_q_d,
      yt_rsc_7_9_i_q_d, {butterFly2_15_f1_equal_tmp_1 , butterFly1_15_f1_equal_tmp_3_1
      , butterFly1_15_f1_equal_tmp_4_1 , butterFly1_15_f1_equal_tmp_5_1 , butterFly1_15_f1_equal_tmp_6_1
      , butterFly1_15_f1_equal_tmp_7_1 , butterFly1_15_f1_equal_tmp_1 , butterFly2_15_f1_equal_tmp_7_1});
  assign mult_t_mul_cmp_11_a_mx0w3 = MUX1HOT_v_32_8_2(xt_rsc_0_9_i_qa_d, xt_rsc_1_9_i_qa_d,
      xt_rsc_2_9_i_qa_d, xt_rsc_3_9_i_qa_d, xt_rsc_4_9_i_qa_d, xt_rsc_5_9_i_qa_d,
      xt_rsc_6_9_i_qa_d, xt_rsc_7_9_i_qa_d, {butterFly2_15_f1_equal_tmp_1 , butterFly1_15_f1_equal_tmp_3_1
      , butterFly1_15_f1_equal_tmp_4_1 , butterFly1_15_f1_equal_tmp_5_1 , butterFly1_15_f1_equal_tmp_6_1
      , butterFly1_15_f1_equal_tmp_7_1 , butterFly1_15_f1_equal_tmp_1 , butterFly2_15_f1_equal_tmp_7_1});
  assign nl_mult_15_if_acc_nl = mult_15_res_sva_1 - p_sva;
  assign mult_15_if_acc_nl = nl_mult_15_if_acc_nl[31:0];
  assign nl_mult_31_acc_1_nl = ({1'b1 , mult_15_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_31_acc_1_nl = nl_mult_31_acc_1_nl[32:0];
  assign mult_15_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_15_if_acc_nl, mult_15_res_sva_1,
      readslicef_33_1_32(mult_31_acc_1_nl));
  assign nl_mult_14_if_acc_nl = mult_14_res_sva_1 - p_sva;
  assign mult_14_if_acc_nl = nl_mult_14_if_acc_nl[31:0];
  assign nl_mult_30_acc_1_nl = ({1'b1 , mult_14_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_30_acc_1_nl = nl_mult_30_acc_1_nl[32:0];
  assign mult_14_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_14_if_acc_nl, mult_14_res_sva_1,
      readslicef_33_1_32(mult_30_acc_1_nl));
  assign nl_mult_13_if_acc_nl = mult_13_res_sva_1 - p_sva;
  assign mult_13_if_acc_nl = nl_mult_13_if_acc_nl[31:0];
  assign nl_mult_29_acc_1_nl = ({1'b1 , mult_13_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_29_acc_1_nl = nl_mult_29_acc_1_nl[32:0];
  assign mult_13_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_13_if_acc_nl, mult_13_res_sva_1,
      readslicef_33_1_32(mult_29_acc_1_nl));
  assign nl_mult_12_if_acc_nl = mult_12_res_sva_1 - p_sva;
  assign mult_12_if_acc_nl = nl_mult_12_if_acc_nl[31:0];
  assign nl_mult_28_acc_1_nl = ({1'b1 , mult_12_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_28_acc_1_nl = nl_mult_28_acc_1_nl[32:0];
  assign mult_12_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_12_if_acc_nl, mult_12_res_sva_1,
      readslicef_33_1_32(mult_28_acc_1_nl));
  assign nl_mult_11_if_acc_nl = mult_11_res_sva_1 - p_sva;
  assign mult_11_if_acc_nl = nl_mult_11_if_acc_nl[31:0];
  assign nl_mult_27_acc_1_nl = ({1'b1 , mult_11_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_27_acc_1_nl = nl_mult_27_acc_1_nl[32:0];
  assign mult_11_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_11_if_acc_nl, mult_11_res_sva_1,
      readslicef_33_1_32(mult_27_acc_1_nl));
  assign nl_mult_10_if_acc_nl = mult_10_res_sva_1 - p_sva;
  assign mult_10_if_acc_nl = nl_mult_10_if_acc_nl[31:0];
  assign nl_mult_26_acc_1_nl = ({1'b1 , mult_10_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_26_acc_1_nl = nl_mult_26_acc_1_nl[32:0];
  assign mult_10_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_10_if_acc_nl, mult_10_res_sva_1,
      readslicef_33_1_32(mult_26_acc_1_nl));
  assign nl_mult_9_if_acc_nl = mult_9_res_sva_1 - p_sva;
  assign mult_9_if_acc_nl = nl_mult_9_if_acc_nl[31:0];
  assign nl_mult_25_acc_1_nl = ({1'b1 , mult_9_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_25_acc_1_nl = nl_mult_25_acc_1_nl[32:0];
  assign mult_9_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_9_if_acc_nl, mult_9_res_sva_1,
      readslicef_33_1_32(mult_25_acc_1_nl));
  assign nl_mult_8_if_acc_nl = mult_8_res_sva_1 - p_sva;
  assign mult_8_if_acc_nl = nl_mult_8_if_acc_nl[31:0];
  assign nl_mult_24_acc_1_nl = ({1'b1 , mult_8_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_24_acc_1_nl = nl_mult_24_acc_1_nl[32:0];
  assign mult_8_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_8_if_acc_nl, mult_8_res_sva_1,
      readslicef_33_1_32(mult_24_acc_1_nl));
  assign nl_mult_7_if_acc_nl = mult_7_res_sva_1 - p_sva;
  assign mult_7_if_acc_nl = nl_mult_7_if_acc_nl[31:0];
  assign nl_mult_23_acc_1_nl = ({1'b1 , mult_7_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_23_acc_1_nl = nl_mult_23_acc_1_nl[32:0];
  assign mult_7_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_7_if_acc_nl, mult_7_res_sva_1,
      readslicef_33_1_32(mult_23_acc_1_nl));
  assign nl_mult_6_if_acc_nl = mult_6_res_sva_1 - p_sva;
  assign mult_6_if_acc_nl = nl_mult_6_if_acc_nl[31:0];
  assign nl_mult_22_acc_1_nl = ({1'b1 , mult_6_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_22_acc_1_nl = nl_mult_22_acc_1_nl[32:0];
  assign mult_6_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_6_if_acc_nl, mult_6_res_sva_1,
      readslicef_33_1_32(mult_22_acc_1_nl));
  assign nl_mult_5_if_acc_nl = mult_5_res_sva_1 - p_sva;
  assign mult_5_if_acc_nl = nl_mult_5_if_acc_nl[31:0];
  assign nl_mult_21_acc_1_nl = ({1'b1 , mult_5_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_21_acc_1_nl = nl_mult_21_acc_1_nl[32:0];
  assign mult_5_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_5_if_acc_nl, mult_5_res_sva_1,
      readslicef_33_1_32(mult_21_acc_1_nl));
  assign nl_mult_4_if_acc_nl = mult_4_res_sva_1 - p_sva;
  assign mult_4_if_acc_nl = nl_mult_4_if_acc_nl[31:0];
  assign nl_mult_20_acc_1_nl = ({1'b1 , mult_4_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_20_acc_1_nl = nl_mult_20_acc_1_nl[32:0];
  assign mult_4_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_4_if_acc_nl, mult_4_res_sva_1,
      readslicef_33_1_32(mult_20_acc_1_nl));
  assign nl_mult_3_if_acc_nl = mult_3_res_sva_1 - p_sva;
  assign mult_3_if_acc_nl = nl_mult_3_if_acc_nl[31:0];
  assign nl_mult_19_acc_1_nl = ({1'b1 , mult_3_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_19_acc_1_nl = nl_mult_19_acc_1_nl[32:0];
  assign mult_3_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_3_if_acc_nl, mult_3_res_sva_1,
      readslicef_33_1_32(mult_19_acc_1_nl));
  assign nl_mult_2_if_acc_nl = mult_2_res_sva_1 - p_sva;
  assign mult_2_if_acc_nl = nl_mult_2_if_acc_nl[31:0];
  assign nl_mult_18_acc_1_nl = ({1'b1 , mult_2_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_18_acc_1_nl = nl_mult_18_acc_1_nl[32:0];
  assign mult_2_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_2_if_acc_nl, mult_2_res_sva_1,
      readslicef_33_1_32(mult_18_acc_1_nl));
  assign nl_mult_1_if_acc_nl = mult_1_res_sva_1 - p_sva;
  assign mult_1_if_acc_nl = nl_mult_1_if_acc_nl[31:0];
  assign nl_mult_17_acc_1_nl = ({1'b1 , mult_1_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_17_acc_1_nl = nl_mult_17_acc_1_nl[32:0];
  assign mult_1_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_1_if_acc_nl, mult_1_res_sva_1,
      readslicef_33_1_32(mult_17_acc_1_nl));
  assign nl_mult_if_acc_nl = mult_res_sva_1 - p_sva;
  assign mult_if_acc_nl = nl_mult_if_acc_nl[31:0];
  assign nl_mult_16_acc_1_nl = ({1'b1 , mult_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_16_acc_1_nl = nl_mult_16_acc_1_nl[32:0];
  assign mult_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_if_acc_nl, mult_res_sva_1,
      readslicef_33_1_32(mult_16_acc_1_nl));
  assign INNER_LOOP2_r_11_4_sva_6_0_mx1 = MUX_v_7_2_2(7'b0000000, (z_out_62[6:0]),
      (fsm_output[4]));
  assign nl_mult_15_res_sva_1 = mult_15_z_asn_itm_3 - mult_z_mul_cmp_1_z;
  assign mult_15_res_sva_1 = nl_mult_15_res_sva_1[31:0];
  assign nl_mult_14_res_sva_1 = mult_14_z_asn_itm_3 - mult_z_mul_cmp_3_z;
  assign mult_14_res_sva_1 = nl_mult_14_res_sva_1[31:0];
  assign nl_mult_13_res_sva_1 = mult_13_z_asn_itm_3 - mult_z_mul_cmp_5_z;
  assign mult_13_res_sva_1 = nl_mult_13_res_sva_1[31:0];
  assign nl_mult_12_res_sva_1 = mult_12_z_asn_itm_3 - mult_z_mul_cmp_7_z;
  assign mult_12_res_sva_1 = nl_mult_12_res_sva_1[31:0];
  assign nl_mult_11_res_sva_1 = mult_11_z_asn_itm_3 - mult_z_mul_cmp_9_z;
  assign mult_11_res_sva_1 = nl_mult_11_res_sva_1[31:0];
  assign nl_mult_10_res_sva_1 = mult_10_z_asn_itm_3 - mult_z_mul_cmp_11_z;
  assign mult_10_res_sva_1 = nl_mult_10_res_sva_1[31:0];
  assign nl_mult_9_res_sva_1 = mult_25_z_asn_itm_3 - mult_z_mul_cmp_13_z;
  assign mult_9_res_sva_1 = nl_mult_9_res_sva_1[31:0];
  assign nl_mult_8_res_sva_1 = mult_24_z_asn_itm_3 - mult_z_mul_cmp_15_z;
  assign mult_8_res_sva_1 = nl_mult_8_res_sva_1[31:0];
  assign nl_mult_7_res_sva_1 = mult_23_z_asn_itm_3 - mult_z_mul_cmp_17_z;
  assign mult_7_res_sva_1 = nl_mult_7_res_sva_1[31:0];
  assign nl_mult_6_res_sva_1 = mult_22_z_asn_itm_3 - mult_z_mul_cmp_19_z;
  assign mult_6_res_sva_1 = nl_mult_6_res_sva_1[31:0];
  assign nl_mult_5_res_sva_1 = mult_21_z_asn_itm_3 - mult_z_mul_cmp_21_z;
  assign mult_5_res_sva_1 = nl_mult_5_res_sva_1[31:0];
  assign nl_mult_4_res_sva_1 = mult_20_z_asn_itm_3 - mult_z_mul_cmp_23_z;
  assign mult_4_res_sva_1 = nl_mult_4_res_sva_1[31:0];
  assign nl_mult_3_res_sva_1 = mult_19_z_asn_itm_3 - mult_z_mul_cmp_25_z;
  assign mult_3_res_sva_1 = nl_mult_3_res_sva_1[31:0];
  assign nl_mult_2_res_sva_1 = mult_18_z_asn_itm_3 - mult_z_mul_cmp_27_z;
  assign mult_2_res_sva_1 = nl_mult_2_res_sva_1[31:0];
  assign nl_mult_1_res_sva_1 = mult_17_z_asn_itm_3 - mult_z_mul_cmp_29_z;
  assign mult_1_res_sva_1 = nl_mult_1_res_sva_1[31:0];
  assign nl_mult_res_sva_1 = mult_16_z_asn_itm_3 - mult_z_mul_cmp_31_z;
  assign mult_res_sva_1 = nl_mult_res_sva_1[31:0];
  assign tmp_71_lpi_3_dfm_1 = MUX1HOT_v_32_8_2(xt_rsc_0_7_i_qa_d, xt_rsc_1_7_i_qa_d,
      xt_rsc_2_7_i_qa_d, xt_rsc_3_7_i_qa_d, xt_rsc_4_7_i_qa_d, xt_rsc_5_7_i_qa_d,
      xt_rsc_6_7_i_qa_d, xt_rsc_7_7_i_qa_d, {butterFly1_15_f1_equal_tmp_1 , butterFly1_15_f1_equal_tmp_1_1
      , butterFly1_15_f1_equal_tmp_2_1 , butterFly1_15_f1_equal_tmp_3_1 , butterFly1_15_f1_equal_tmp_4_1
      , butterFly1_15_f1_equal_tmp_5_1 , butterFly1_15_f1_equal_tmp_6_1 , butterFly1_15_f1_equal_tmp_7_1});
  assign operator_33_true_2_lshift_psp_2_0_sva_mx0 = MUX_v_3_2_2((z_out_60[2:0]),
      operator_20_false_acc_cse_sva, fsm_output[7]);
  assign INNER_LOOP4_nor_tmp = ~(INNER_LOOP1_stage_0 | butterFly1_15_conc_2_itm_2_0
      | butterFly1_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_4_0 | butterFly1_15_conc_2_itm_5_0
      | butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_8_0
      | butterFly1_15_conc_2_itm_9_0 | butterFly1_15_conc_2_itm_0);
  assign or_dcpl = butterFly1_15_conc_2_itm_5_0 | butterFly2_15_conc_2_itm_1_0;
  assign or_dcpl_2 = butterFly1_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_0;
  assign or_dcpl_8 = butterFly1_15_conc_2_itm_8_0 | butterFly2_15_conc_2_itm_4_0;
  assign or_dcpl_10 = butterFly1_15_conc_2_itm_7_0 | butterFly2_15_conc_2_itm_3_0;
  assign or_dcpl_12 = butterFly1_15_conc_2_itm_6_0 | butterFly2_15_conc_2_itm_2_0;
  assign or_dcpl_19 = butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_0;
  assign or_dcpl_22 = butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_8_0;
  assign or_dcpl_25 = butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_7_0;
  assign or_dcpl_30 = butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_3_0;
  assign or_dcpl_33 = butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_2_0;
  assign or_dcpl_36 = butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_1_0;
  assign or_dcpl_63 = butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_8_0;
  assign or_dcpl_70 = butterFly1_15_conc_2_itm_8_0 | butterFly1_15_conc_2_itm_9_0;
  assign or_dcpl_72 = butterFly2_15_conc_2_itm_3_0 | butterFly2_15_conc_2_itm_5_0;
  assign or_dcpl_76 = butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_8_0;
  assign or_dcpl_78 = butterFly2_15_conc_2_itm_3_0 | butterFly2_15_conc_2_itm_7_0;
  assign or_dcpl_80 = butterFly1_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_8_0;
  assign or_dcpl_82 = butterFly2_15_conc_2_itm_3_0 | butterFly2_15_conc_2_itm_8_0;
  assign or_dcpl_88 = butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_8_0;
  assign or_dcpl_89 = butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_3_0;
  assign or_dcpl_94 = butterFly1_15_conc_2_itm_7_0 | butterFly2_15_conc_2_itm_2_0;
  assign or_dcpl_105 = butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_9_0;
  assign or_dcpl_107 = butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_5_0;
  assign or_dcpl_109 = butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_7_0;
  assign or_dcpl_111 = butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_7_0;
  assign or_dcpl_116 = butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_7_0;
  assign or_dcpl_117 = butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_6_0;
  assign or_dcpl_119 = butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_3_0;
  assign or_dcpl_121 = butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_8_0;
  assign or_dcpl_125 = butterFly1_15_conc_2_itm_6_0 | butterFly2_15_conc_2_itm_1_0;
  assign or_dcpl_133 = butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_6_0;
  assign or_dcpl_135 = butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_3_0;
  assign or_dcpl_139 = butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_9_0;
  assign or_dcpl_141 = butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_5_0;
  assign or_dcpl_146 = butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_5_0;
  assign or_dcpl_148 = butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_7_0;
  assign or_dcpl_150 = butterFly1_15_conc_2_itm_5_0 | butterFly1_15_conc_2_itm_3_0;
  assign or_dcpl_152 = butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_8_0;
  assign or_dcpl_161 = butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_5_0;
  assign or_dcpl_163 = butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_2_0;
  assign or_dcpl_165 = butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_5_0;
  assign or_dcpl_167 = butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_3_0;
  assign or_dcpl_171 = butterFly1_15_conc_2_itm_5_0 | butterFly1_15_conc_2_itm_9_0;
  assign or_dcpl_173 = butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_5_0;
  assign or_dcpl_180 = INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_5_0;
  assign or_dcpl_181 = butterFly1_15_conc_2_itm_4_0 | butterFly1_15_conc_2_itm_9_0;
  assign or_dcpl_185 = butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_4_0;
  assign or_dcpl_187 = INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_7_0;
  assign or_dcpl_189 = butterFly1_15_conc_2_itm_4_0 | butterFly1_15_conc_2_itm_3_0;
  assign or_dcpl_197 = butterFly1_15_conc_2_itm_5_0 | butterFly1_15_conc_2_itm_4_0;
  assign or_dcpl_199 = INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_1_0;
  assign or_dcpl_201 = butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_4_0;
  assign or_dcpl_203 = INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_2_0;
  assign or_dcpl_205 = butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_4_0;
  assign or_dcpl_207 = INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_3_0;
  assign or_dcpl_210 = INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_4_0;
  assign or_dcpl_215 = INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_4_0;
  assign or_dcpl_218 = butterFly1_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_9_0;
  assign or_dcpl_220 = INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_5_0;
  assign or_dcpl_224 = butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_3_0;
  assign or_dcpl_234 = INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_0;
  assign or_dcpl_238 = INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_1_0;
  assign or_dcpl_242 = INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_2_0;
  assign or_dcpl_246 = INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_3_0;
  assign or_dcpl_274 = butterFly1_15_conc_2_itm_9_0 | butterFly2_15_conc_2_itm_5_0;
  assign and_dcpl_62 = INNER_LOOP4_nor_tmp & c_1_sva;
  assign or_tmp_26 = butterFly1_15_f1_equal_tmp_2_1 | (butterFly2_15_conc_itm_10_2_1[1])
      | (~ butterFly1_15_conc_2_itm_1_0);
  assign or_tmp_29 = (butterFly2_15_conc_2_itm_9_2_1[1]) | butterFly1_15_f1_equal_tmp_1_1
      | (~ butterFly1_15_conc_2_itm_0);
  assign nor_62_nl = ~(butterFly1_15_conc_2_itm_1_0 | (~ or_tmp_29));
  assign or_325_nl = butterFly1_15_f1_equal_tmp_2_1 | (butterFly2_15_conc_itm_10_2_1[1]);
  assign mux_tmp = MUX_s_1_2_2(nor_62_nl, or_tmp_29, or_325_nl);
  assign or_tmp_35 = (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1]) | (~
      butterFly1_15_conc_2_itm_2_0);
  assign not_tmp_25 = ~((~((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])
      | (~ butterFly1_15_conc_2_itm_2_0))) | INNER_LOOP1_stage_0);
  assign or_tmp_38 = (butterFly1_15_conc_2_itm_9_2_1[0]) | butterFly1_15_conc_2_itm_9_0
      | (butterFly1_15_conc_2_itm_9_2_1[1]) | (~ INNER_LOOP1_stage_0_10);
  assign or_tmp_40 = (butterFly2_15_conc_2_itm_6_2_1[1]) | (~ INNER_LOOP1_stage_0_11)
      | INNER_LOOP2_stage_0_10;
  assign not_tmp_29 = ~(INNER_LOOP1_stage_0_10 | (~ or_tmp_40));
  assign and_dcpl_66 = ~((butterFly2_15_conc_2_itm_9_2_1!=2'b00));
  assign and_dcpl_67 = butterFly1_15_conc_2_itm_0 & (~ butterFly1_15_f1_equal_tmp_1_1);
  assign and_dcpl_68 = and_dcpl_67 & and_dcpl_66;
  assign and_dcpl_69 = ~(butterFly1_15_conc_2_itm_9_0 | (butterFly1_15_conc_2_itm_9_2_1[0]));
  assign and_dcpl_70 = INNER_LOOP1_stage_0_10 & (~ (butterFly1_15_conc_2_itm_9_2_1[1]));
  assign and_dcpl_73 = INNER_LOOP1_stage_0 & (~ (INNER_LOOP4_r_11_4_sva_6_0[5]));
  assign and_dcpl_76 = INNER_LOOP1_stage_0 & (~ (INNER_LOOP2_r_11_4_sva_6_0[5]));
  assign nor_tmp_1 = butterFly1_15_f1_equal_tmp_1_1 & butterFly1_15_conc_2_itm_0;
  assign or_tmp_48 = (~ butterFly1_15_f1_equal_tmp_2_1) | (butterFly2_15_conc_itm_10_2_1[1])
      | (~ butterFly1_15_conc_2_itm_1_0);
  assign or_tmp_50 = (butterFly2_15_conc_2_itm_9_2_1[1]) | (~ nor_tmp_1);
  assign nor_56_nl = ~(butterFly1_15_conc_2_itm_1_0 | (~ or_tmp_50));
  assign or_347_nl = (~ butterFly1_15_f1_equal_tmp_2_1) | (butterFly2_15_conc_itm_10_2_1[1]);
  assign mux_tmp_7 = MUX_s_1_2_2(nor_56_nl, or_tmp_50, or_347_nl);
  assign or_tmp_53 = (butterFly1_15_conc_2_itm_9_2_1[0]) | (~ butterFly1_15_conc_2_itm_9_0)
      | (butterFly1_15_conc_2_itm_9_2_1[1]) | (~ INNER_LOOP1_stage_0_10);
  assign or_tmp_55 = (butterFly2_15_conc_2_itm_6_2_1[1]) | (~(INNER_LOOP1_stage_0_11
      & INNER_LOOP2_stage_0_10));
  assign not_tmp_50 = ~(INNER_LOOP1_stage_0_10 | (~ or_tmp_55));
  assign and_dcpl_78 = nor_tmp_1 & and_dcpl_66;
  assign and_dcpl_79 = butterFly1_15_conc_2_itm_9_0 & (~ (butterFly1_15_conc_2_itm_9_2_1[0]));
  assign or_tmp_64 = (~ (butterFly1_15_conc_2_itm_9_2_1[0])) | butterFly1_15_conc_2_itm_9_0
      | (butterFly1_15_conc_2_itm_9_2_1[1]) | (~ INNER_LOOP1_stage_0_10);
  assign and_dcpl_81 = (butterFly2_15_conc_2_itm_9_2_1==2'b01);
  assign and_dcpl_82 = and_dcpl_67 & and_dcpl_81;
  assign and_dcpl_83 = (~ butterFly1_15_conc_2_itm_9_0) & (butterFly1_15_conc_2_itm_9_2_1[0]);
  assign or_tmp_72 = ~((butterFly1_15_conc_2_itm_9_2_1[0]) & butterFly1_15_conc_2_itm_9_0
      & (~ (butterFly1_15_conc_2_itm_9_2_1[1])) & INNER_LOOP1_stage_0_10);
  assign and_dcpl_89 = nor_tmp_1 & and_dcpl_81;
  assign nand_7_cse = ~((butterFly2_15_conc_itm_10_2_1[1]) & butterFly1_15_conc_2_itm_1_0);
  assign or_tmp_75 = butterFly1_15_f1_equal_tmp_2_1 | nand_7_cse;
  assign or_tmp_77 = (~ (butterFly2_15_conc_2_itm_9_2_1[1])) | butterFly1_15_f1_equal_tmp_1_1
      | (~ butterFly1_15_conc_2_itm_0);
  assign and_8934_nl = nand_7_cse & or_tmp_77;
  assign mux_tmp_22 = MUX_s_1_2_2(and_8934_nl, or_tmp_77, butterFly1_15_f1_equal_tmp_2_1);
  assign nor_tmp_6 = (INNER_LOOP4_r_11_4_sva_6_0[5]) & INNER_LOOP1_stage_0;
  assign and_8932_cse = (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1]) &
      butterFly1_15_conc_2_itm_2_0;
  assign or_tmp_82 = and_8932_cse | INNER_LOOP1_stage_0;
  assign nor_tmp_10 = (butterFly1_15_conc_2_itm_9_2_1[1]) & INNER_LOOP1_stage_0_10;
  assign or_tmp_84 = (butterFly1_15_conc_2_itm_9_2_1[0]) | butterFly1_15_conc_2_itm_9_0
      | (~ nor_tmp_10);
  assign or_tmp_86 = (~ (butterFly2_15_conc_2_itm_6_2_1[1])) | (~ INNER_LOOP1_stage_0_11)
      | INNER_LOOP2_stage_0_10;
  assign not_tmp_67 = (~((butterFly1_15_conc_2_itm_9_2_1[1]) & INNER_LOOP1_stage_0_10))
      & or_tmp_86;
  assign not_tmp_69 = ~((INNER_LOOP2_r_11_4_sva_6_0[5]) & INNER_LOOP1_stage_0);
  assign or_tmp_90 = (INNER_LOOP2_r_11_4_sva_6_0[4]) | (INNER_LOOP2_r_11_4_sva_6_0[6])
      | not_tmp_69;
  assign and_dcpl_92 = (butterFly2_15_conc_2_itm_9_2_1==2'b10);
  assign and_dcpl_93 = and_dcpl_67 & and_dcpl_92;
  assign nor_tmp_14 = (butterFly2_15_conc_2_itm_9_2_1[1]) & butterFly1_15_f1_equal_tmp_1_1
      & butterFly1_15_conc_2_itm_0;
  assign nor_tmp_15 = butterFly1_15_f1_equal_tmp_2_1 & (butterFly2_15_conc_itm_10_2_1[1])
      & butterFly1_15_conc_2_itm_1_0;
  assign or_tmp_93 = nor_tmp_15 | nor_tmp_14;
  assign or_tmp_94 = (butterFly1_15_conc_2_itm_9_2_1[0]) | (~(butterFly1_15_conc_2_itm_9_0
      & (butterFly1_15_conc_2_itm_9_2_1[1]) & INNER_LOOP1_stage_0_10));
  assign nor_tmp_19 = (butterFly2_15_conc_2_itm_6_2_1[1]) & INNER_LOOP1_stage_0_11
      & INNER_LOOP2_stage_0_10;
  assign and_dcpl_96 = nor_tmp_1 & and_dcpl_92;
  assign or_tmp_99 = (~ (INNER_LOOP4_r_11_4_sva_6_0[4])) | (INNER_LOOP4_r_11_4_sva_6_0[6])
      | (~ nor_tmp_6);
  assign or_tmp_102 = (~ (butterFly1_15_conc_2_itm_9_2_1[0])) | butterFly1_15_conc_2_itm_9_0
      | (~ nor_tmp_10);
  assign or_tmp_104 = (~ (INNER_LOOP2_r_11_4_sva_6_0[4])) | (INNER_LOOP2_r_11_4_sva_6_0[6])
      | not_tmp_69;
  assign and_dcpl_99 = and_dcpl_67 & (butterFly2_15_conc_2_itm_9_2_1==2'b11);
  assign nor_tmp_22 = (butterFly2_15_conc_2_itm_9_2_1==2'b11) & butterFly1_15_f1_equal_tmp_1_1
      & butterFly1_15_conc_2_itm_0;
  assign or_tmp_112 = butterFly1_15_f1_equal_tmp_1_1 | (~ butterFly1_15_conc_2_itm_0);
  assign not_tmp_87 = ~(butterFly1_15_conc_2_itm_9_0 | and_dcpl_67);
  assign or_409_nl = (butterFly2_15_conc_2_itm_8_2_1[1]) | butterFly2_15_conc_2_itm_8_0;
  assign mux_44_nl = MUX_s_1_2_2(not_tmp_87, or_tmp_112, or_409_nl);
  assign or_408_nl = (butterFly2_15_conc_2_itm_8_2_1[1]) | butterFly2_15_conc_2_itm_8_0
      | (~ butterFly1_15_conc_2_itm_9_0);
  assign mux_tmp_45 = MUX_s_1_2_2(mux_44_nl, or_408_nl, butterFly2_15_conc_2_itm_9_2_1[1]);
  assign or_tmp_120 = butterFly1_15_conc_2_itm_8_0 | (butterFly1_15_conc_2_itm_8_2_1[1])
      | (~ butterFly2_15_conc_2_itm_5_0);
  assign or_tmp_122 = (butterFly1_15_conc_2_itm_9_2_1[1]) | (~ INNER_LOOP1_stage_0_10);
  assign not_tmp_91 = ~(butterFly2_15_conc_2_itm_5_0 | and_dcpl_70);
  assign or_419_nl = butterFly1_15_conc_2_itm_8_0 | (butterFly1_15_conc_2_itm_8_2_1[1]);
  assign mux_tmp_50 = MUX_s_1_2_2(not_tmp_91, or_tmp_122, or_419_nl);
  assign and_dcpl_101 = ~((butterFly2_15_conc_2_itm_8_2_1!=2'b00));
  assign and_dcpl_102 = butterFly1_15_conc_2_itm_9_0 & (~ butterFly2_15_conc_2_itm_8_0);
  assign and_dcpl_104 = ~(butterFly1_15_conc_2_itm_8_0 | (butterFly1_15_conc_2_itm_8_2_1[0]));
  assign and_dcpl_105 = butterFly2_15_conc_2_itm_5_0 & (~ (butterFly1_15_conc_2_itm_8_2_1[1]));
  assign and_dcpl_107 = (INNER_LOOP4_r_11_4_sva_6_0[6]) & (~ (INNER_LOOP4_r_11_4_sva_6_0[4]));
  assign nor_tmp_25 = butterFly2_15_conc_2_itm_8_0 & butterFly1_15_conc_2_itm_9_0;
  assign nor_52_nl = ~((~((butterFly2_15_conc_2_itm_8_2_1[1]) | (~ butterFly2_15_conc_2_itm_8_0)
      | (~ butterFly1_15_conc_2_itm_9_0))) | nor_tmp_1);
  assign or_427_nl = (butterFly2_15_conc_2_itm_8_2_1[1]) | (~ nor_tmp_25);
  assign mux_tmp_53 = MUX_s_1_2_2(nor_52_nl, or_427_nl, butterFly2_15_conc_2_itm_9_2_1[1]);
  assign or_429_nl = (~ butterFly1_15_conc_2_itm_8_0) | (butterFly1_15_conc_2_itm_8_2_1[1]);
  assign mux_tmp_56 = MUX_s_1_2_2(not_tmp_91, or_tmp_122, or_429_nl);
  assign or_tmp_133 = (~ butterFly1_15_conc_2_itm_8_0) | (butterFly1_15_conc_2_itm_8_2_1[1])
      | (~ butterFly2_15_conc_2_itm_5_0);
  assign and_dcpl_112 = butterFly1_15_conc_2_itm_8_0 & (~ (butterFly1_15_conc_2_itm_8_2_1[0]));
  assign and_dcpl_114 = (butterFly2_15_conc_2_itm_8_2_1==2'b01);
  assign and_dcpl_116 = (~ butterFly1_15_conc_2_itm_8_0) & (butterFly1_15_conc_2_itm_8_2_1[0]);
  assign and_dcpl_123 = butterFly1_15_conc_2_itm_8_0 & (butterFly1_15_conc_2_itm_8_2_1[0]);
  assign or_447_nl = (~ (butterFly2_15_conc_2_itm_8_2_1[1])) | butterFly2_15_conc_2_itm_8_0
      | (~ butterFly1_15_conc_2_itm_9_0);
  assign or_445_nl = (~ (butterFly2_15_conc_2_itm_8_2_1[1])) | butterFly2_15_conc_2_itm_8_0;
  assign mux_69_nl = MUX_s_1_2_2(not_tmp_87, or_tmp_112, or_445_nl);
  assign mux_tmp_70 = MUX_s_1_2_2(or_447_nl, mux_69_nl, butterFly2_15_conc_2_itm_9_2_1[1]);
  assign nor_tmp_32 = (butterFly1_15_conc_2_itm_8_2_1[1]) & butterFly2_15_conc_2_itm_5_0;
  assign or_tmp_153 = butterFly1_15_conc_2_itm_8_0 | (~ nor_tmp_32);
  assign not_tmp_115 = ~((~(butterFly1_15_conc_2_itm_8_0 | (~ (butterFly1_15_conc_2_itm_8_2_1[1]))
      | (~ butterFly2_15_conc_2_itm_5_0))) | nor_tmp_10);
  assign or_tmp_156 = (INNER_LOOP2_r_11_4_sva_6_0[4]) | (~((INNER_LOOP2_r_11_4_sva_6_0[6:5]==2'b11)
      & INNER_LOOP1_stage_0));
  assign and_dcpl_125 = (butterFly2_15_conc_2_itm_8_2_1==2'b10);
  assign nor_tmp_36 = (butterFly2_15_conc_2_itm_8_2_1[1]) & butterFly2_15_conc_2_itm_8_0
      & butterFly1_15_conc_2_itm_9_0;
  assign or_457_nl = nor_tmp_36 | nor_tmp_1;
  assign mux_tmp_78 = MUX_s_1_2_2(nor_tmp_36, or_457_nl, butterFly2_15_conc_2_itm_9_2_1[1]);
  assign and_8919_cse = butterFly1_15_conc_2_itm_8_0 & (butterFly1_15_conc_2_itm_8_2_1[1])
      & butterFly2_15_conc_2_itm_5_0;
  assign or_tmp_160 = and_8919_cse | nor_tmp_10;
  assign nor_tmp_43 = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b111) & INNER_LOOP1_stage_0;
  assign nor_tmp_45 = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b111) & INNER_LOOP1_stage_0;
  assign nor_tmp_46 = (butterFly2_15_conc_2_itm_8_2_1==2'b11) & butterFly2_15_conc_2_itm_8_0
      & butterFly1_15_conc_2_itm_9_0;
  assign and_dcpl_135 = INNER_LOOP2_stage_0_10 & (~ (butterFly1_15_conc_2_itm_9_2_1[1]));
  assign and_dcpl_138 = INNER_LOOP1_stage_0 & (~ (INNER_LOOP3_r_11_4_sva_6_0[4]));
  assign and_dcpl_141 = INNER_LOOP1_stage_0 & (~ (INNER_LOOP1_r_11_4_sva_6_0[4]));
  assign and_dcpl_145 = INNER_LOOP1_stage_0 & (INNER_LOOP3_r_11_4_sva_6_0[4]);
  assign and_dcpl_147 = INNER_LOOP1_stage_0 & (INNER_LOOP1_r_11_4_sva_6_0[4]);
  assign and_dcpl_150 = INNER_LOOP2_stage_0_10 & (butterFly1_15_conc_2_itm_9_2_1[1]);
  assign and_dcpl_152 = (INNER_LOOP3_r_11_4_sva_6_0[6:5]==2'b01);
  assign and_dcpl_154 = (INNER_LOOP1_r_11_4_sva_6_0[6:5]==2'b01);
  assign and_dcpl_161 = (INNER_LOOP3_r_11_4_sva_6_0[6:5]==2'b10);
  assign and_dcpl_163 = (INNER_LOOP1_r_11_4_sva_6_0[6:5]==2'b10);
  assign and_dcpl_167 = (INNER_LOOP3_r_11_4_sva_6_0[6:5]==2'b11);
  assign and_dcpl_169 = (INNER_LOOP1_r_11_4_sva_6_0[6:5]==2'b11);
  assign or_dcpl_298 = (fsm_output[7]) | (fsm_output[9]);
  assign or_dcpl_300 = modulo_add_1_qelse_or_m1c | or_dcpl_298;
  assign and_dcpl_173 = INNER_LOOP1_stage_0 & (operator_20_false_acc_cse_sva[0]);
  assign and_dcpl_175 = INNER_LOOP1_stage_0 & (operator_20_false_acc_cse_sva[1]);
  assign and_dcpl_176 = INNER_LOOP1_stage_0 & (operator_33_true_3_lshift_psp_1_0_sva[1]);
  assign or_dcpl_315 = (fsm_output[4:3]!=2'b00);
  assign and_dcpl_239 = ~((fsm_output[4]) | (fsm_output[2]));
  assign or_dcpl_353 = (fsm_output[2]) | (fsm_output[7]);
  assign or_dcpl_361 = (fsm_output[4]) | (fsm_output[7]);
  assign or_329_cse = (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]) | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]);
  assign or_332_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b000);
  assign mux_3_nl = MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_332_nl);
  assign or_331_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b000) | (~ INNER_LOOP1_stage_0);
  assign mux_4_nl = MUX_s_1_2_2(mux_3_nl, or_331_nl, or_329_cse);
  assign and_344_cse = (~ mux_4_nl) & (fsm_output[9]);
  assign and_346_cse = (~(((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2])
      | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]) | (~ butterFly2_15_conc_2_itm_7_0)
      | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])) & ((INNER_LOOP2_r_11_4_sva_6_0[6:4]!=3'b000)
      | (~ INNER_LOOP1_stage_0)))) & (fsm_output[4]);
  assign or_359_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b001) | (~ INNER_LOOP1_stage_0);
  assign or_357_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b001);
  assign mux_14_nl = MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_357_nl);
  assign nor_3_nl = ~((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]) | (~
      (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0])));
  assign mux_15_nl = MUX_s_1_2_2(or_359_nl, mux_14_nl, nor_3_nl);
  assign and_715_cse = (~ mux_15_nl) & (fsm_output[9]);
  assign and_717_cse = (~(((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2])
      | (~ (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0])) | (~ butterFly2_15_conc_2_itm_7_0)
      | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])) & ((INNER_LOOP2_r_11_4_sva_6_0[6:4]!=3'b001)
      | (~ INNER_LOOP1_stage_0)))) & (fsm_output[4]);
  assign nor_7_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b010));
  assign mux_25_nl = MUX_s_1_2_2(and_8932_cse, or_tmp_82, nor_7_nl);
  assign nor_64_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[4]) | (INNER_LOOP4_r_11_4_sva_6_0[6])
      | (~ nor_tmp_6));
  assign mux_26_nl = MUX_s_1_2_2(mux_25_nl, nor_64_nl, or_329_cse);
  assign and_1022_cse = mux_26_nl & (fsm_output[9]);
  assign nand_24_cse = ~(butterFly2_15_conc_2_itm_7_0 & (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1]));
  assign and_8944_nl = nand_24_cse & or_tmp_90;
  assign mux_29_nl = MUX_s_1_2_2(and_8944_nl, or_tmp_90, or_329_cse);
  assign and_1024_cse = (~ mux_29_nl) & (fsm_output[4]);
  assign nor_20_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b011));
  assign mux_35_nl = MUX_s_1_2_2(and_8932_cse, or_tmp_82, nor_20_nl);
  assign mux_36_nl = MUX_s_1_2_2((~ or_tmp_99), mux_35_nl, butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]);
  assign mux_37_nl = MUX_s_1_2_2(mux_36_nl, (~ or_tmp_99), butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]);
  assign and_1329_cse = mux_37_nl & (fsm_output[9]);
  assign and_8943_nl = (~((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0])
      & butterFly2_15_conc_2_itm_7_0 & (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])))
      & or_tmp_104;
  assign mux_40_nl = MUX_s_1_2_2(and_8943_nl, or_tmp_104, butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]);
  assign and_1331_cse = (~ mux_40_nl) & (fsm_output[4]);
  assign or_412_cse = (~ (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]))
      | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]);
  assign or_415_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b100);
  assign mux_48_nl = MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_415_nl);
  assign or_414_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b100) | (~ INNER_LOOP1_stage_0);
  assign mux_49_nl = MUX_s_1_2_2(mux_48_nl, or_414_nl, or_412_cse);
  assign and_1636_cse = (~ mux_49_nl) & (fsm_output[9]);
  assign and_1638_cse = (~(((~ (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]))
      | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]) | (~ butterFly2_15_conc_2_itm_7_0)
      | (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])) & ((INNER_LOOP2_r_11_4_sva_6_0[6:4]!=3'b100)
      | (~ INNER_LOOP1_stage_0)))) & (fsm_output[4]);
  assign and_8941_cse = (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2]) &
      (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]);
  assign nand_17_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b101) & INNER_LOOP1_stage_0);
  assign or_434_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b101);
  assign mux_61_nl = MUX_s_1_2_2(not_tmp_25, or_tmp_35, or_434_nl);
  assign mux_62_nl = MUX_s_1_2_2(nand_17_nl, mux_61_nl, and_8941_cse);
  assign and_2007_cse = (~ mux_62_nl) & (fsm_output[9]);
  assign and_2009_cse = (~((~((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2])
      & (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]) & butterFly2_15_conc_2_itm_7_0
      & (~ (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])))) & (~((INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b101)
      & INNER_LOOP1_stage_0)))) & (fsm_output[4]);
  assign nor_31_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b110));
  assign mux_73_nl = MUX_s_1_2_2(and_8932_cse, or_tmp_82, nor_31_nl);
  assign nor_63_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[4]) | (~((INNER_LOOP4_r_11_4_sva_6_0[6:5]==2'b11)
      & INNER_LOOP1_stage_0)));
  assign mux_74_nl = MUX_s_1_2_2(mux_73_nl, nor_63_nl, or_412_cse);
  assign and_2314_cse = mux_74_nl & (fsm_output[9]);
  assign and_8942_nl = nand_24_cse & or_tmp_156;
  assign mux_77_nl = MUX_s_1_2_2(and_8942_nl, or_tmp_156, or_412_cse);
  assign and_2316_cse = (~ mux_77_nl) & (fsm_output[4]);
  assign mux_85_nl = MUX_s_1_2_2(and_8932_cse, or_tmp_82, butterFly2_16_f1_butterFly2_16_f1_and_6_cse);
  assign mux_86_nl = MUX_s_1_2_2(nor_tmp_43, mux_85_nl, and_8941_cse);
  assign and_2621_cse = mux_86_nl & (fsm_output[9]);
  assign and_2623_cse = (((butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[2])
      & (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[0]) & butterFly2_15_conc_2_itm_7_0
      & (butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1[1])) | nor_tmp_45) & (fsm_output[4]);
  assign and_6834_cse = INNER_LOOP1_stage_0 & (operator_33_true_3_lshift_psp_1_0_sva[0])
      & (fsm_output[9]);
  assign and_6843_cse = and_dcpl_176 & (fsm_output[9]);
  assign and_6852_cse = and_dcpl_176 & (operator_33_true_3_lshift_psp_1_0_sva[0])
      & (fsm_output[9]);
  assign or_tmp_3231 = modulo_add_1_qelse_or_m1c | (fsm_output[9]);
  assign and_7090_cse = (~ (operator_33_true_3_lshift_psp_1_0_sva[0])) & (fsm_output[9]);
  assign or_tmp_3239 = and_7090_cse | modulo_add_1_qelse_or_m1c;
  assign or_tmp_3242 = (operator_33_true_3_lshift_psp_1_0_sva[0]) & (fsm_output[9]);
  assign and_7109_cse = (~ (operator_33_true_3_lshift_psp_1_0_sva[1])) & (fsm_output[9]);
  assign or_tmp_3250 = (operator_20_false_acc_cse_sva[2]) & (fsm_output[7]);
  assign and_7115_cse = (~ (operator_20_false_acc_cse_sva[2])) & (fsm_output[7]);
  assign or_tmp_3252 = (operator_33_true_3_lshift_psp_1_0_sva[1]) & (fsm_output[9]);
  assign or_tmp_3269 = (operator_20_false_acc_cse_sva[1]) & (fsm_output[7]);
  assign and_7153_cse = (~ (operator_20_false_acc_cse_sva[1])) & (fsm_output[7]);
  assign or_tmp_3279 = (operator_20_false_acc_cse_sva[0]) & (fsm_output[7]);
  assign and_7173_cse = (~ (operator_20_false_acc_cse_sva[0])) & (fsm_output[7]);
  assign or_tmp_3345 = and_7153_cse | modulo_add_1_qelse_or_m1c;
  assign or_tmp_3354 = and_7173_cse | modulo_add_1_qelse_or_m1c;
  assign or_tmp_3597 = (fsm_output[2:1]!=2'b00);
  assign or_tmp_3600 = (fsm_output[7:6]!=2'b00);
  assign or_tmp_3650 = and_dcpl_239 & (~ (fsm_output[7])) & (~ (fsm_output[9]));
  assign or_tmp_3666 = (fsm_output[2]) | (fsm_output[9]);
  assign or_tmp_3717 = ~((fsm_output[2]) | (fsm_output[7]));
  assign or_tmp_3723 = ~((fsm_output[6]) | (fsm_output[2]) | (fsm_output[7]));
  assign or_tmp_3732 = (fsm_output[9:8]!=2'b00);
  assign or_tmp_3755 = (fsm_output[4]) | (fsm_output[9]);
  assign or_tmp_3842 = or_dcpl_361 | (fsm_output[9]);
  assign INNER_LOOP1_tw_and_nl = INNER_LOOP2_r_11_4_sva_6_0 & INNER_LOOP1_r_11_4_sva_6_0;
  assign INNER_LOOP2_tw_and_nl = operator_33_true_1_lshift_psp_9_4_sva & (INNER_LOOP2_r_11_4_sva_6_0[5:0]);
  assign INNER_LOOP1_tw_h_mux1h_4_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_tw_and_nl, ({(INNER_LOOP2_r_11_4_sva_6_0[6])
      , INNER_LOOP2_tw_and_nl}), INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_and_ssc = ~((z_out_111[31]) | (fsm_output[7]));
  assign butterFly1_and_ssc_2 = (~ (z_out_125[31])) & (fsm_output[7]);
  assign butterFly1_1_and_ssc = ~((z_out_112[31]) | (fsm_output[7]));
  assign butterFly1_1_and_ssc_2 = (~ (z_out_126[31])) & (fsm_output[7]);
  assign butterFly1_1_and_ssc_3 = (z_out_126[31]) & (fsm_output[7]);
  assign butterFly1_2_and_ssc = ~((z_out_113[31]) | (fsm_output[7]));
  assign butterFly1_2_and_ssc_2 = (~ (z_out_111[31])) & (fsm_output[7]);
  assign butterFly1_2_and_ssc_3 = (z_out_111[31]) & (fsm_output[7]);
  assign butterFly1_3_and_ssc = ~((z_out_114[31]) | (fsm_output[7]));
  assign butterFly1_3_and_ssc_2 = (~ (z_out_112[31])) & (fsm_output[7]);
  assign butterFly1_3_and_ssc_3 = (z_out_112[31]) & (fsm_output[7]);
  assign butterFly1_4_and_ssc = ~((z_out_115[31]) | (fsm_output[7]));
  assign butterFly1_4_and_ssc_2 = (~ (z_out_113[31])) & (fsm_output[7]);
  assign butterFly1_4_and_ssc_3 = (z_out_113[31]) & (fsm_output[7]);
  assign butterFly1_5_and_ssc = ~((z_out_116[31]) | (fsm_output[7]));
  assign butterFly1_5_and_ssc_2 = (~ (z_out_114[31])) & (fsm_output[7]);
  assign butterFly1_5_and_ssc_3 = (z_out_114[31]) & (fsm_output[7]);
  assign butterFly1_6_and_ssc = ~((z_out_117[31]) | (fsm_output[7]));
  assign butterFly1_6_and_ssc_2 = (~ (z_out_115[31])) & (fsm_output[7]);
  assign butterFly1_6_and_ssc_3 = (z_out_115[31]) & (fsm_output[7]);
  assign butterFly1_7_and_ssc = ~((z_out_118[31]) | (fsm_output[7]));
  assign butterFly1_7_and_ssc_2 = (~ (z_out_116[31])) & (fsm_output[7]);
  assign butterFly1_7_and_ssc_3 = (z_out_116[31]) & (fsm_output[7]);
  assign butterFly1_8_and_ssc = ~((z_out_119[31]) | (fsm_output[7]));
  assign butterFly1_8_and_ssc_2 = (~ (z_out_117[31])) & (fsm_output[7]);
  assign butterFly1_8_and_ssc_3 = (z_out_117[31]) & (fsm_output[7]);
  assign butterFly1_9_and_ssc = ~((z_out_120[31]) | (fsm_output[7]));
  assign butterFly1_9_and_ssc_2 = (~ (z_out_118[31])) & (fsm_output[7]);
  assign butterFly1_9_and_ssc_3 = (z_out_118[31]) & (fsm_output[7]);
  assign butterFly1_10_and_ssc = ~((z_out_121[31]) | (fsm_output[7]));
  assign butterFly1_10_and_ssc_2 = (~ (z_out_119[31])) & (fsm_output[7]);
  assign butterFly1_10_and_ssc_3 = (z_out_119[31]) & (fsm_output[7]);
  assign butterFly1_11_and_ssc = ~((z_out_122[31]) | (fsm_output[7]));
  assign butterFly1_11_and_ssc_2 = (~ (z_out_120[31])) & (fsm_output[7]);
  assign butterFly1_11_and_ssc_3 = (z_out_120[31]) & (fsm_output[7]);
  assign butterFly1_12_and_ssc = ~((z_out_123[31]) | (fsm_output[7]));
  assign butterFly1_12_and_ssc_2 = (~ (z_out_121[31])) & (fsm_output[7]);
  assign butterFly1_12_and_ssc_3 = (z_out_121[31]) & (fsm_output[7]);
  assign butterFly1_13_and_ssc = ~((z_out_124[31]) | (fsm_output[7]));
  assign butterFly1_13_and_ssc_2 = (~ (z_out_122[31])) & (fsm_output[7]);
  assign butterFly1_13_and_ssc_3 = (z_out_122[31]) & (fsm_output[7]);
  assign butterFly1_14_and_ssc = ~((z_out_125[31]) | (fsm_output[7]));
  assign butterFly1_14_and_ssc_2 = (~ (z_out_123[31])) & (fsm_output[7]);
  assign butterFly1_14_and_ssc_3 = (z_out_123[31]) & (fsm_output[7]);
  assign butterFly1_15_and_ssc = ~((z_out_126[31]) | (fsm_output[7]));
  assign butterFly1_15_and_ssc_2 = (~ (z_out_124[31])) & (fsm_output[7]);
  assign yt_rsc_0_0_i_d_d_pff = MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1, modulo_add_10_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_0_i_radr_d_pff = MUX_v_4_2_2((INNER_LOOP2_r_11_4_sva_6_0[3:0]),
      (INNER_LOOP4_r_11_4_sva_6_0[3:0]), fsm_output[9]);
  assign yt_rsc_0_0_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8, fsm_output[7]);
  assign yt_rsc_0_0_i_we_d_pff = (and_dcpl_68 & (fsm_output[7])) | (and_dcpl_70 &
      and_dcpl_69 & (fsm_output[2]));
  assign yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_73 & butterFly2_16_f1_nor_1_cse
      & (fsm_output[9])) | (and_dcpl_76 & (~ (INNER_LOOP2_r_11_4_sva_6_0[6])) & (~
      (INNER_LOOP2_r_11_4_sva_6_0[4])) & (fsm_output[4]));
  assign yt_rsc_0_1_i_d_d_pff = MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1, modulo_add_11_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_1_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8, fsm_output[7]);
  assign yt_rsc_0_2_i_d_d_pff = MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1, modulo_add_12_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_2_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8, fsm_output[7]);
  assign yt_rsc_0_3_i_d_d_pff = MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1, modulo_add_13_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_3_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8, fsm_output[7]);
  assign yt_rsc_0_4_i_d_d_pff = MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1, modulo_add_14_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_4_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8, fsm_output[7]);
  assign yt_rsc_0_5_i_d_d_pff = MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1, modulo_add_15_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_5_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8, fsm_output[7]);
  assign yt_rsc_0_6_i_d_d_pff = MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1, modulo_add_1_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_6_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8, fsm_output[7]);
  assign yt_rsc_0_7_i_d_d_pff = MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1, modulo_add_23_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_8_i_d_d_pff = MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1, modulo_add_24_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_9_i_d_d_pff = MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1, modulo_add_25_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_10_i_d_d_pff = MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1, modulo_add_26_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_10_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8, fsm_output[7]);
  assign yt_rsc_0_11_i_d_d_pff = MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1, modulo_add_27_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_11_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8, fsm_output[7]);
  assign yt_rsc_0_12_i_d_d_pff = MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1, modulo_add_28_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_13_i_d_d_pff = MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1, modulo_add_29_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_14_i_d_d_pff = MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1, modulo_add_30_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_15_i_d_d_pff = MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1, modulo_add_31_qr_lpi_3_dfm_1,
      fsm_output[7]);
  assign yt_rsc_0_16_i_we_d_pff = (and_dcpl_78 & (fsm_output[7])) | (and_dcpl_70
      & and_dcpl_79 & (fsm_output[2]));
  assign yt_rsc_1_0_i_we_d_pff = (and_dcpl_82 & (fsm_output[7])) | (and_dcpl_70 &
      and_dcpl_83 & (fsm_output[2]));
  assign yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_73 & (~ (INNER_LOOP4_r_11_4_sva_6_0[6]))
      & (INNER_LOOP4_r_11_4_sva_6_0[4]) & (fsm_output[9])) | (and_dcpl_76 & (~ (INNER_LOOP2_r_11_4_sva_6_0[6]))
      & (INNER_LOOP2_r_11_4_sva_6_0[4]) & (fsm_output[4]));
  assign yt_rsc_1_16_i_we_d_pff = (and_dcpl_89 & (fsm_output[7])) | (and_dcpl_70
      & and_8912_cse & (fsm_output[2]));
  assign yt_rsc_2_0_i_we_d_pff = (and_dcpl_93 & (fsm_output[7])) | (nor_tmp_10 &
      and_dcpl_69 & (fsm_output[2]));
  assign yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (nor_tmp_6 & butterFly2_16_f1_nor_1_cse
      & (fsm_output[9])) | ((~ or_tmp_90) & (fsm_output[4]));
  assign yt_rsc_2_16_i_we_d_pff = (and_dcpl_96 & (fsm_output[7])) | (nor_tmp_10 &
      and_dcpl_79 & (fsm_output[2]));
  assign yt_rsc_3_0_i_we_d_pff = (and_dcpl_99 & (fsm_output[7])) | (nor_tmp_10 &
      and_dcpl_83 & (fsm_output[2]));
  assign yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = ((~ or_tmp_99) & (fsm_output[9]))
      | ((~ or_tmp_104) & (fsm_output[4]));
  assign yt_rsc_3_16_i_we_d_pff = (nor_tmp_22 & (fsm_output[7])) | (and_8913_cse
      & (fsm_output[2]));
  assign butterFly1_and_4_nl = (z_out_108[31]) & (~(butterFly1_and_ssc | butterFly1_and_ssc_2));
  assign butterFly1_or_nl = ((z_out_111[31]) & (~ (fsm_output[7]))) | ((z_out_125[31])
      & (fsm_output[7]));
  assign butterFly1_mux1h_nl = MUX1HOT_v_31_3_2((z_out_111[30:0]), (z_out_108[30:0]),
      (z_out_125[30:0]), {butterFly1_and_ssc , butterFly1_or_nl , butterFly1_and_ssc_2});
  assign yt_rsc_4_0_i_d_d_pff = {butterFly1_and_4_nl , butterFly1_mux1h_nl};
  assign yt_rsc_4_0_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8, fsm_output[7]);
  assign yt_rsc_4_0_i_we_d_pff = (and_dcpl_102 & and_dcpl_101 & (fsm_output[7]))
      | (and_dcpl_105 & and_dcpl_104 & (fsm_output[2]));
  assign yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_73 & and_dcpl_107
      & (fsm_output[9])) | (and_dcpl_76 & (INNER_LOOP2_r_11_4_sva_6_0[6]) & (~ (INNER_LOOP2_r_11_4_sva_6_0[4]))
      & (fsm_output[4]));
  assign butterFly1_1_mux_nl = MUX_s_1_2_2((z_out_102[31]), (z_out_105[31]), butterFly1_1_and_ssc_3);
  assign butterFly1_1_and_4_nl = butterFly1_1_mux_nl & (~(butterFly1_1_and_ssc |
      butterFly1_1_and_ssc_2));
  assign butterFly1_1_and_1_nl = (z_out_112[31]) & (~ (fsm_output[7]));
  assign butterFly1_1_mux1h_nl = MUX1HOT_v_31_4_2((z_out_112[30:0]), (z_out_102[30:0]),
      (z_out_126[30:0]), (z_out_105[30:0]), {butterFly1_1_and_ssc , butterFly1_1_and_1_nl
      , butterFly1_1_and_ssc_2 , butterFly1_1_and_ssc_3});
  assign yt_rsc_4_1_i_d_d_pff = {butterFly1_1_and_4_nl , butterFly1_1_mux1h_nl};
  assign yt_rsc_4_1_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8, fsm_output[7]);
  assign butterFly1_2_mux_nl = MUX_s_1_2_2((z_out_97[31]), (z_out_100[31]), butterFly1_2_and_ssc_3);
  assign butterFly1_2_and_4_nl = butterFly1_2_mux_nl & (~(butterFly1_2_and_ssc |
      butterFly1_2_and_ssc_2));
  assign butterFly1_2_and_1_nl = (z_out_113[31]) & (~ (fsm_output[7]));
  assign butterFly1_2_mux1h_nl = MUX1HOT_v_31_4_2((z_out_113[30:0]), (z_out_97[30:0]),
      (z_out_111[30:0]), (z_out_100[30:0]), {butterFly1_2_and_ssc , butterFly1_2_and_1_nl
      , butterFly1_2_and_ssc_2 , butterFly1_2_and_ssc_3});
  assign yt_rsc_4_2_i_d_d_pff = {butterFly1_2_and_4_nl , butterFly1_2_mux1h_nl};
  assign yt_rsc_4_2_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8, fsm_output[7]);
  assign butterFly1_3_mux_nl = MUX_s_1_2_2((z_out_92[31]), (z_out_94[31]), butterFly1_3_and_ssc_3);
  assign butterFly1_3_and_4_nl = butterFly1_3_mux_nl & (~(butterFly1_3_and_ssc |
      butterFly1_3_and_ssc_2));
  assign butterFly1_3_and_1_nl = (z_out_114[31]) & (~ (fsm_output[7]));
  assign butterFly1_3_mux1h_nl = MUX1HOT_v_31_4_2((z_out_114[30:0]), (z_out_92[30:0]),
      (z_out_112[30:0]), (z_out_94[30:0]), {butterFly1_3_and_ssc , butterFly1_3_and_1_nl
      , butterFly1_3_and_ssc_2 , butterFly1_3_and_ssc_3});
  assign yt_rsc_4_3_i_d_d_pff = {butterFly1_3_and_4_nl , butterFly1_3_mux1h_nl};
  assign yt_rsc_4_3_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8, fsm_output[7]);
  assign butterFly1_4_mux_nl = MUX_s_1_2_2((z_out_86[31]), (z_out_89[31]), butterFly1_4_and_ssc_3);
  assign butterFly1_4_and_4_nl = butterFly1_4_mux_nl & (~(butterFly1_4_and_ssc |
      butterFly1_4_and_ssc_2));
  assign butterFly1_4_and_1_nl = (z_out_115[31]) & (~ (fsm_output[7]));
  assign butterFly1_4_mux1h_nl = MUX1HOT_v_31_4_2((z_out_115[30:0]), (z_out_86[30:0]),
      (z_out_113[30:0]), (z_out_89[30:0]), {butterFly1_4_and_ssc , butterFly1_4_and_1_nl
      , butterFly1_4_and_ssc_2 , butterFly1_4_and_ssc_3});
  assign yt_rsc_4_4_i_d_d_pff = {butterFly1_4_and_4_nl , butterFly1_4_mux1h_nl};
  assign yt_rsc_4_4_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8, fsm_output[7]);
  assign butterFly1_5_mux_nl = MUX_s_1_2_2((z_out_81[31]), (z_out_84[31]), butterFly1_5_and_ssc_3);
  assign butterFly1_5_and_4_nl = butterFly1_5_mux_nl & (~(butterFly1_5_and_ssc |
      butterFly1_5_and_ssc_2));
  assign butterFly1_5_and_1_nl = (z_out_116[31]) & (~ (fsm_output[7]));
  assign butterFly1_5_mux1h_nl = MUX1HOT_v_31_4_2((z_out_116[30:0]), (z_out_81[30:0]),
      (z_out_114[30:0]), (z_out_84[30:0]), {butterFly1_5_and_ssc , butterFly1_5_and_1_nl
      , butterFly1_5_and_ssc_2 , butterFly1_5_and_ssc_3});
  assign yt_rsc_4_5_i_d_d_pff = {butterFly1_5_and_4_nl , butterFly1_5_mux1h_nl};
  assign yt_rsc_4_5_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8, fsm_output[7]);
  assign butterFly1_6_mux_nl = MUX_s_1_2_2((z_out_76[31]), (z_out_78[31]), butterFly1_6_and_ssc_3);
  assign butterFly1_6_and_4_nl = butterFly1_6_mux_nl & (~(butterFly1_6_and_ssc |
      butterFly1_6_and_ssc_2));
  assign butterFly1_6_and_1_nl = (z_out_117[31]) & (~ (fsm_output[7]));
  assign butterFly1_6_mux1h_nl = MUX1HOT_v_31_4_2((z_out_117[30:0]), (z_out_76[30:0]),
      (z_out_115[30:0]), (z_out_78[30:0]), {butterFly1_6_and_ssc , butterFly1_6_and_1_nl
      , butterFly1_6_and_ssc_2 , butterFly1_6_and_ssc_3});
  assign yt_rsc_4_6_i_d_d_pff = {butterFly1_6_and_4_nl , butterFly1_6_mux1h_nl};
  assign yt_rsc_4_6_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8, fsm_output[7]);
  assign butterFly1_7_mux_nl = MUX_s_1_2_2((z_out_70[31]), (z_out_73[31]), butterFly1_7_and_ssc_3);
  assign butterFly1_7_and_4_nl = butterFly1_7_mux_nl & (~(butterFly1_7_and_ssc |
      butterFly1_7_and_ssc_2));
  assign butterFly1_7_and_1_nl = (z_out_118[31]) & (~ (fsm_output[7]));
  assign butterFly1_7_mux1h_nl = MUX1HOT_v_31_4_2((z_out_118[30:0]), (z_out_70[30:0]),
      (z_out_116[30:0]), (z_out_73[30:0]), {butterFly1_7_and_ssc , butterFly1_7_and_1_nl
      , butterFly1_7_and_ssc_2 , butterFly1_7_and_ssc_3});
  assign yt_rsc_4_7_i_d_d_pff = {butterFly1_7_and_4_nl , butterFly1_7_mux1h_nl};
  assign butterFly1_8_mux_nl = MUX_s_1_2_2((z_out_105[31]), (z_out_102[31]), butterFly1_8_and_ssc_3);
  assign butterFly1_8_and_4_nl = butterFly1_8_mux_nl & (~(butterFly1_8_and_ssc |
      butterFly1_8_and_ssc_2));
  assign butterFly1_8_and_1_nl = (z_out_119[31]) & (~ (fsm_output[7]));
  assign butterFly1_8_mux1h_nl = MUX1HOT_v_31_4_2((z_out_119[30:0]), (z_out_105[30:0]),
      (z_out_117[30:0]), (z_out_102[30:0]), {butterFly1_8_and_ssc , butterFly1_8_and_1_nl
      , butterFly1_8_and_ssc_2 , butterFly1_8_and_ssc_3});
  assign yt_rsc_4_8_i_d_d_pff = {butterFly1_8_and_4_nl , butterFly1_8_mux1h_nl};
  assign butterFly1_9_mux_nl = MUX_s_1_2_2((z_out_100[31]), (z_out_97[31]), butterFly1_9_and_ssc_3);
  assign butterFly1_9_and_4_nl = butterFly1_9_mux_nl & (~(butterFly1_9_and_ssc |
      butterFly1_9_and_ssc_2));
  assign butterFly1_9_and_1_nl = (z_out_120[31]) & (~ (fsm_output[7]));
  assign butterFly1_9_mux1h_272_nl = MUX1HOT_v_31_4_2((z_out_120[30:0]), (z_out_100[30:0]),
      (z_out_118[30:0]), (z_out_97[30:0]), {butterFly1_9_and_ssc , butterFly1_9_and_1_nl
      , butterFly1_9_and_ssc_2 , butterFly1_9_and_ssc_3});
  assign yt_rsc_4_9_i_d_d_pff = {butterFly1_9_and_4_nl , butterFly1_9_mux1h_272_nl};
  assign yt_rsc_4_9_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8, fsm_output[7]);
  assign butterFly1_10_mux_nl = MUX_s_1_2_2((z_out_94[31]), (z_out_92[31]), butterFly1_10_and_ssc_3);
  assign butterFly1_10_and_4_nl = butterFly1_10_mux_nl & (~(butterFly1_10_and_ssc
      | butterFly1_10_and_ssc_2));
  assign butterFly1_10_and_1_nl = (z_out_121[31]) & (~ (fsm_output[7]));
  assign butterFly1_10_mux1h_nl = MUX1HOT_v_31_4_2((z_out_121[30:0]), (z_out_94[30:0]),
      (z_out_119[30:0]), (z_out_92[30:0]), {butterFly1_10_and_ssc , butterFly1_10_and_1_nl
      , butterFly1_10_and_ssc_2 , butterFly1_10_and_ssc_3});
  assign yt_rsc_4_10_i_d_d_pff = {butterFly1_10_and_4_nl , butterFly1_10_mux1h_nl};
  assign yt_rsc_4_10_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8, fsm_output[7]);
  assign butterFly1_11_mux_nl = MUX_s_1_2_2((z_out_89[31]), (z_out_86[31]), butterFly1_11_and_ssc_3);
  assign butterFly1_11_and_4_nl = butterFly1_11_mux_nl & (~(butterFly1_11_and_ssc
      | butterFly1_11_and_ssc_2));
  assign butterFly1_11_and_1_nl = (z_out_122[31]) & (~ (fsm_output[7]));
  assign butterFly1_11_mux1h_nl = MUX1HOT_v_31_4_2((z_out_122[30:0]), (z_out_89[30:0]),
      (z_out_120[30:0]), (z_out_86[30:0]), {butterFly1_11_and_ssc , butterFly1_11_and_1_nl
      , butterFly1_11_and_ssc_2 , butterFly1_11_and_ssc_3});
  assign yt_rsc_4_11_i_d_d_pff = {butterFly1_11_and_4_nl , butterFly1_11_mux1h_nl};
  assign yt_rsc_4_11_i_wadr_d_pff = MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8, fsm_output[7]);
  assign butterFly1_12_mux_nl = MUX_s_1_2_2((z_out_84[31]), (z_out_81[31]), butterFly1_12_and_ssc_3);
  assign butterFly1_12_and_4_nl = butterFly1_12_mux_nl & (~(butterFly1_12_and_ssc
      | butterFly1_12_and_ssc_2));
  assign butterFly1_12_and_1_nl = (z_out_123[31]) & (~ (fsm_output[7]));
  assign butterFly1_12_mux1h_nl = MUX1HOT_v_31_4_2((z_out_123[30:0]), (z_out_84[30:0]),
      (z_out_121[30:0]), (z_out_81[30:0]), {butterFly1_12_and_ssc , butterFly1_12_and_1_nl
      , butterFly1_12_and_ssc_2 , butterFly1_12_and_ssc_3});
  assign yt_rsc_4_12_i_d_d_pff = {butterFly1_12_and_4_nl , butterFly1_12_mux1h_nl};
  assign butterFly1_13_mux_nl = MUX_s_1_2_2((z_out_78[31]), (z_out_76[31]), butterFly1_13_and_ssc_3);
  assign butterFly1_13_and_4_nl = butterFly1_13_mux_nl & (~(butterFly1_13_and_ssc
      | butterFly1_13_and_ssc_2));
  assign butterFly1_13_and_1_nl = (z_out_124[31]) & (~ (fsm_output[7]));
  assign butterFly1_13_mux1h_nl = MUX1HOT_v_31_4_2((z_out_124[30:0]), (z_out_78[30:0]),
      (z_out_122[30:0]), (z_out_76[30:0]), {butterFly1_13_and_ssc , butterFly1_13_and_1_nl
      , butterFly1_13_and_ssc_2 , butterFly1_13_and_ssc_3});
  assign yt_rsc_4_13_i_d_d_pff = {butterFly1_13_and_4_nl , butterFly1_13_mux1h_nl};
  assign butterFly1_14_mux_nl = MUX_s_1_2_2((z_out_73[31]), (z_out_70[31]), butterFly1_14_and_ssc_3);
  assign butterFly1_14_and_4_nl = butterFly1_14_mux_nl & (~(butterFly1_14_and_ssc
      | butterFly1_14_and_ssc_2));
  assign butterFly1_14_and_1_nl = (z_out_125[31]) & (~ (fsm_output[7]));
  assign butterFly1_14_mux1h_nl = MUX1HOT_v_31_4_2((z_out_125[30:0]), (z_out_73[30:0]),
      (z_out_123[30:0]), (z_out_70[30:0]), {butterFly1_14_and_ssc , butterFly1_14_and_1_nl
      , butterFly1_14_and_ssc_2 , butterFly1_14_and_ssc_3});
  assign yt_rsc_4_14_i_d_d_pff = {butterFly1_14_and_4_nl , butterFly1_14_mux1h_nl};
  assign butterFly1_15_and_5_nl = (z_out_68[31]) & (~(butterFly1_15_and_ssc | butterFly1_15_and_ssc_2));
  assign butterFly1_15_or_nl = ((z_out_126[31]) & (~ (fsm_output[7]))) | ((z_out_124[31])
      & (fsm_output[7]));
  assign butterFly1_15_mux1h_nl = MUX1HOT_v_31_3_2((z_out_126[30:0]), (z_out_68[30:0]),
      (z_out_124[30:0]), {butterFly1_15_and_ssc , butterFly1_15_or_nl , butterFly1_15_and_ssc_2});
  assign yt_rsc_4_15_i_d_d_pff = {butterFly1_15_and_5_nl , butterFly1_15_mux1h_nl};
  assign yt_rsc_4_16_i_we_d_pff = (nor_tmp_25 & and_dcpl_101 & (fsm_output[7])) |
      (and_dcpl_105 & and_dcpl_112 & (fsm_output[2]));
  assign yt_rsc_5_0_i_we_d_pff = (and_dcpl_102 & and_dcpl_114 & (fsm_output[7]))
      | (and_dcpl_105 & and_dcpl_116 & (fsm_output[2]));
  assign yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_73 & (INNER_LOOP4_r_11_4_sva_6_0[6])
      & (INNER_LOOP4_r_11_4_sva_6_0[4]) & (fsm_output[9])) | (and_dcpl_76 & (INNER_LOOP2_r_11_4_sva_6_0[6])
      & (INNER_LOOP2_r_11_4_sva_6_0[4]) & (fsm_output[4]));
  assign yt_rsc_5_16_i_we_d_pff = (nor_tmp_25 & and_dcpl_114 & (fsm_output[7])) |
      (and_dcpl_105 & and_dcpl_123 & (fsm_output[2]));
  assign yt_rsc_6_0_i_we_d_pff = (and_dcpl_102 & and_dcpl_125 & (fsm_output[7]))
      | (nor_tmp_32 & and_dcpl_104 & (fsm_output[2]));
  assign yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (nor_tmp_6 & and_dcpl_107
      & (fsm_output[9])) | ((~ or_tmp_156) & (fsm_output[4]));
  assign yt_rsc_6_16_i_we_d_pff = (nor_tmp_25 & and_dcpl_125 & (fsm_output[7])) |
      (nor_tmp_32 & and_dcpl_112 & (fsm_output[2]));
  assign yt_rsc_7_0_i_we_d_pff = (and_dcpl_102 & (butterFly2_15_conc_2_itm_8_2_1==2'b11)
      & (fsm_output[7])) | (nor_tmp_32 & and_dcpl_116 & (fsm_output[2]));
  assign yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff = (nor_tmp_43 & (fsm_output[9]))
      | (nor_tmp_45 & (fsm_output[4]));
  assign yt_rsc_7_16_i_we_d_pff = (nor_tmp_46 & (fsm_output[7])) | (nor_tmp_32 &
      and_dcpl_123 & (fsm_output[2]));
  assign xt_rsc_0_0_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_0_i_da_d_pff = modulo_add_10_qr_lpi_3_dfm_1;
  assign xt_rsc_0_0_i_wea_d_pff = (and_dcpl_68 & (fsm_output[9])) | (and_dcpl_135
      & and_dcpl_69 & (fsm_output[4]));
  assign xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_138 & butterFly2_f1_nor_cse
      & (fsm_output[7])) | (and_dcpl_141 & butterFly1_f1_nor_cse & (fsm_output[2]));
  assign xt_rsc_0_1_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_1_i_da_d_pff = modulo_add_11_qr_lpi_3_dfm_1;
  assign xt_rsc_0_2_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_2_i_da_d_pff = modulo_add_12_qr_lpi_3_dfm_1;
  assign xt_rsc_0_3_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_3_i_da_d_pff = modulo_add_13_qr_lpi_3_dfm_1;
  assign xt_rsc_0_4_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_4_i_da_d_pff = modulo_add_14_qr_lpi_3_dfm_1;
  assign xt_rsc_0_5_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_5_i_da_d_pff = modulo_add_15_qr_lpi_3_dfm_1;
  assign xt_rsc_0_6_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_6_i_da_d_pff = modulo_add_1_qr_lpi_3_dfm_1;
  assign xt_rsc_0_7_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_7_i_da_d_pff = modulo_add_23_qr_lpi_3_dfm_1;
  assign xt_rsc_0_8_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_8_i_da_d_pff = modulo_add_24_qr_lpi_3_dfm_1;
  assign xt_rsc_0_9_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_9_i_da_d_pff = modulo_add_25_qr_lpi_3_dfm_1;
  assign xt_rsc_0_10_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_10_i_da_d_pff = modulo_add_26_qr_lpi_3_dfm_1;
  assign xt_rsc_0_11_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_11_i_da_d_pff = modulo_add_27_qr_lpi_3_dfm_1;
  assign xt_rsc_0_12_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_12_i_da_d_pff = modulo_add_28_qr_lpi_3_dfm_1;
  assign xt_rsc_0_13_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_13_i_da_d_pff = modulo_add_29_qr_lpi_3_dfm_1;
  assign xt_rsc_0_14_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_14_i_da_d_pff = modulo_add_30_qr_lpi_3_dfm_1;
  assign xt_rsc_0_15_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_0_15_i_da_d_pff = modulo_add_31_qr_lpi_3_dfm_1;
  assign xt_rsc_0_16_i_wea_d_pff = (and_dcpl_78 & (fsm_output[9])) | (and_dcpl_135
      & and_dcpl_79 & (fsm_output[4]));
  assign xt_rsc_1_0_i_wea_d_pff = (and_dcpl_82 & (fsm_output[9])) | (and_dcpl_135
      & and_dcpl_83 & (fsm_output[4]));
  assign xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_145 & butterFly2_f1_nor_cse
      & (fsm_output[7])) | (and_dcpl_147 & butterFly1_f1_nor_cse & (fsm_output[2]));
  assign xt_rsc_1_16_i_wea_d_pff = (and_dcpl_89 & (fsm_output[9])) | (and_dcpl_135
      & and_8912_cse & (fsm_output[4]));
  assign xt_rsc_2_0_i_wea_d_pff = (and_dcpl_93 & (fsm_output[9])) | (and_dcpl_150
      & and_dcpl_69 & (fsm_output[4]));
  assign xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_138 & and_dcpl_152
      & (fsm_output[7])) | (and_dcpl_141 & and_dcpl_154 & (fsm_output[2]));
  assign xt_rsc_2_16_i_wea_d_pff = (and_dcpl_96 & (fsm_output[9])) | (and_dcpl_150
      & and_dcpl_79 & (fsm_output[4]));
  assign xt_rsc_3_0_i_wea_d_pff = (and_dcpl_99 & (fsm_output[9])) | (and_dcpl_150
      & and_dcpl_83 & (fsm_output[4]));
  assign xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_145 & and_dcpl_152
      & (fsm_output[7])) | (and_dcpl_147 & and_dcpl_154 & (fsm_output[2]));
  assign xt_rsc_3_16_i_wea_d_pff = (nor_tmp_22 & (fsm_output[9])) | (and_dcpl_150
      & and_8912_cse & (fsm_output[4]));
  assign xt_rsc_4_0_i_da_d_pff = {reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_138 & and_dcpl_161
      & (fsm_output[7])) | (and_dcpl_141 & and_dcpl_163 & (fsm_output[2]));
  assign xt_rsc_4_1_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_4_1_i_da_d_pff = {reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_2_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_4_2_i_da_d_pff = {reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_3_i_da_d_pff = {reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_4_i_da_d_pff = {reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_5_i_da_d_pff = {reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_6_i_da_d_pff = {reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_7_i_da_d_pff = {reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_8_i_da_d_pff = {reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_9_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_4_9_i_da_d_pff = {reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_10_i_adra_d_pff = MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[3:0]),
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8, {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign xt_rsc_4_10_i_da_d_pff = {reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_11_i_da_d_pff = {reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_12_i_da_d_pff = {reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_13_i_da_d_pff = {reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_14_i_da_d_pff = {reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_4_15_i_da_d_pff = {reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1};
  assign xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_145 & and_dcpl_161
      & (fsm_output[7])) | (and_dcpl_147 & and_dcpl_163 & (fsm_output[2]));
  assign xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_138 & and_dcpl_167
      & (fsm_output[7])) | (and_dcpl_141 & and_dcpl_169 & (fsm_output[2]));
  assign xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff = (and_dcpl_145 & and_dcpl_167
      & (fsm_output[7])) | (and_dcpl_147 & and_dcpl_169 & (fsm_output[2]));
  assign twiddle_rsc_0_0_i_adra_d = {1'b0 , INNER_LOOP1_tw_h_mux1h_4_rmff};
  assign twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_6824_rmff};
  assign twiddle_rsc_0_1_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3498_rmff};
  assign twiddle_rsc_0_2_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3502_rmff};
  assign twiddle_rsc_0_3_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3506_rmff};
  assign twiddle_rsc_0_4_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3510_rmff};
  assign twiddle_rsc_0_5_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3514_rmff};
  assign twiddle_rsc_0_6_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3518_rmff};
  assign twiddle_rsc_0_7_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3522_rmff};
  assign twiddle_rsc_0_8_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_6895_rmff};
  assign twiddle_rsc_0_9_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3498_rmff};
  assign twiddle_rsc_0_10_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3502_rmff};
  assign twiddle_rsc_0_11_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3506_rmff};
  assign twiddle_rsc_0_12_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3510_rmff};
  assign twiddle_rsc_0_13_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3514_rmff};
  assign twiddle_rsc_0_14_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3518_rmff};
  assign twiddle_rsc_0_15_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3522_rmff};
  assign twiddle_h_rsc_0_0_i_adra_d = {1'b0 , INNER_LOOP1_tw_h_mux1h_4_rmff};
  assign twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_6824_rmff};
  assign twiddle_h_rsc_0_1_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3498_rmff};
  assign twiddle_h_rsc_0_2_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3502_rmff};
  assign twiddle_h_rsc_0_3_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3506_rmff};
  assign twiddle_h_rsc_0_4_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3510_rmff};
  assign twiddle_h_rsc_0_5_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3514_rmff};
  assign twiddle_h_rsc_0_6_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3518_rmff};
  assign twiddle_h_rsc_0_7_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3522_rmff};
  assign twiddle_h_rsc_0_8_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_6895_rmff};
  assign twiddle_h_rsc_0_9_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3498_rmff};
  assign twiddle_h_rsc_0_10_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3502_rmff};
  assign twiddle_h_rsc_0_11_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3506_rmff};
  assign twiddle_h_rsc_0_12_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3510_rmff};
  assign twiddle_h_rsc_0_13_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3514_rmff};
  assign twiddle_h_rsc_0_14_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3518_rmff};
  assign twiddle_h_rsc_0_15_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_3522_rmff};
  assign butterFly1_15_f1_mux_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly2_15_f1_equal_tmp_1,
      fsm_output[7]);
  assign butterFly1_15_f1_mux_1_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1_1,
      butterFly1_15_f1_equal_tmp_3_1, fsm_output[7]);
  assign butterFly1_15_f1_mux_2_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_2_1,
      butterFly1_15_f1_equal_tmp_4_1, fsm_output[7]);
  assign butterFly1_15_f1_mux_3_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1,
      butterFly1_15_f1_equal_tmp_5_1, fsm_output[7]);
  assign butterFly1_15_f1_mux_4_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1,
      butterFly1_15_f1_equal_tmp_6_1, fsm_output[7]);
  assign butterFly1_15_f1_mux_5_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1,
      butterFly1_15_f1_equal_tmp_7_1, fsm_output[7]);
  assign butterFly1_15_f1_mux_6_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1,
      butterFly1_15_f1_equal_tmp_1, fsm_output[7]);
  assign butterFly1_15_f1_mux_7_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1,
      butterFly2_15_f1_equal_tmp_7_1, fsm_output[7]);
  assign butterFly1_31_f1_mux_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly2_15_f1_equal_tmp_1,
      fsm_output[9]);
  assign butterFly1_31_f1_mux_1_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1_1,
      butterFly1_15_f1_equal_tmp_3_1, fsm_output[9]);
  assign butterFly1_31_f1_mux_2_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_2_1,
      butterFly1_15_f1_equal_tmp_4_1, fsm_output[9]);
  assign butterFly1_31_f1_mux_3_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1,
      butterFly1_15_f1_equal_tmp_5_1, fsm_output[9]);
  assign butterFly1_31_f1_mux_4_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1,
      butterFly1_15_f1_equal_tmp_6_1, fsm_output[9]);
  assign butterFly1_31_f1_mux_5_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1,
      butterFly1_15_f1_equal_tmp_7_1, fsm_output[9]);
  assign butterFly1_31_f1_mux_6_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1,
      butterFly1_15_f1_equal_tmp_1, fsm_output[9]);
  assign butterFly1_31_f1_mux_7_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1,
      butterFly2_15_f1_equal_tmp_7_1, fsm_output[9]);
  assign butterFly2_f1_mux_cse = MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_1_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1, butterFly1_15_f1_equal_tmp_1_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_2_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1, butterFly1_15_f1_equal_tmp_2_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_3_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1, butterFly1_15_f1_equal_tmp_3_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_4_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1, butterFly1_15_f1_equal_tmp_4_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_5_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1, butterFly1_15_f1_equal_tmp_5_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_6_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_6_1,
      fsm_output[2]);
  assign butterFly2_f1_mux_7_cse = MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_7_1, butterFly1_15_f1_equal_tmp_7_1,
      fsm_output[2]);
  assign butterFly2_21_f1_mux_cse = MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_1,
      fsm_output[4]);
  assign butterFly2_21_f1_mux_1_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_3_1,
      butterFly1_15_f1_equal_tmp_1_1, fsm_output[4]);
  assign butterFly2_21_f1_mux_2_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_4_1,
      butterFly1_15_f1_equal_tmp_2_1, fsm_output[4]);
  assign butterFly2_21_f1_mux_3_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_5_1,
      butterFly1_15_f1_equal_tmp_3_1, fsm_output[4]);
  assign butterFly2_21_f1_mux_4_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_6_1,
      butterFly1_15_f1_equal_tmp_4_1, fsm_output[4]);
  assign butterFly2_21_f1_mux_5_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_7_1,
      butterFly1_15_f1_equal_tmp_5_1, fsm_output[4]);
  assign butterFly2_21_f1_mux_6_cse = MUX_s_1_2_2(butterFly1_15_f1_equal_tmp_1, butterFly1_15_f1_equal_tmp_6_1,
      fsm_output[4]);
  assign butterFly2_21_f1_mux_7_cse = MUX_s_1_2_2(butterFly2_15_f1_equal_tmp_7_1,
      butterFly1_15_f1_equal_tmp_7_1, fsm_output[4]);
  always @(posedge clk) begin
    if ( or_4976_cse ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      c_1_sva <= 1'b0;
    end
    else if ( (fsm_output[0]) | (fsm_output[5]) | (fsm_output[9]) ) begin
      c_1_sva <= c_mux_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_yt_rsc_0_0_cgo_cse <= 1'b0;
      reg_yt_rsc_0_16_cgo_cse <= 1'b0;
      reg_yt_rsc_1_0_cgo_cse <= 1'b0;
      reg_yt_rsc_1_16_cgo_cse <= 1'b0;
      reg_yt_rsc_2_0_cgo_cse <= 1'b0;
      reg_yt_rsc_2_16_cgo_cse <= 1'b0;
      reg_yt_rsc_3_0_cgo_cse <= 1'b0;
      reg_yt_rsc_3_16_cgo_cse <= 1'b0;
      reg_yt_rsc_4_0_cgo_cse <= 1'b0;
      reg_yt_rsc_4_16_cgo_cse <= 1'b0;
      reg_yt_rsc_5_0_cgo_cse <= 1'b0;
      reg_yt_rsc_5_16_cgo_cse <= 1'b0;
      reg_yt_rsc_6_0_cgo_cse <= 1'b0;
      reg_yt_rsc_6_16_cgo_cse <= 1'b0;
      reg_yt_rsc_7_0_cgo_cse <= 1'b0;
      reg_yt_rsc_7_16_cgo_cse <= 1'b0;
      reg_xt_rsc_triosy_7_31_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      reg_ensig_cgo_17_cse <= 1'b0;
      butterFly1_15_conc_2_itm_2_1 <= 2'b00;
      butterFly1_15_conc_2_itm_9_0 <= 1'b0;
      butterFly1_15_conc_2_itm_8_0 <= 1'b0;
      butterFly1_15_f1_equal_tmp_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_1_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_2_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_3_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_4_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_5_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_6_1 <= 1'b0;
      butterFly1_15_f1_equal_tmp_7_1 <= 1'b0;
      INNER_LOOP1_stage_0 <= 1'b0;
      INNER_LOOP1_r_11_4_sva_6_0 <= 7'b0000000;
      INNER_LOOP1_stage_0_2 <= 1'b0;
      INNER_LOOP1_stage_0_3 <= 1'b0;
      INNER_LOOP1_stage_0_10 <= 1'b0;
      INNER_LOOP1_stage_0_11 <= 1'b0;
      butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm <= 3'b000;
      butterFly1_15_conc_2_itm_7_0 <= 1'b0;
      butterFly1_15_conc_2_itm_6_0 <= 1'b0;
      butterFly1_15_conc_2_itm_5_0 <= 1'b0;
      butterFly1_15_conc_2_itm_4_2_1 <= 2'b00;
      butterFly1_15_conc_2_itm_4_0 <= 1'b0;
      butterFly1_15_conc_2_itm_3_0 <= 1'b0;
      butterFly1_15_conc_2_itm_2_2_1 <= 2'b00;
      butterFly1_15_conc_2_itm_2_0 <= 1'b0;
      butterFly1_15_conc_2_itm_1_0 <= 1'b0;
      butterFly1_15_conc_2_itm_0 <= 1'b0;
      butterFly2_15_conc_2_itm_0 <= 1'b0;
      butterFly2_15_conc_2_itm_1_0 <= 1'b0;
      butterFly2_15_conc_2_itm_2_0 <= 1'b0;
      butterFly2_15_conc_2_itm_3_0 <= 1'b0;
      butterFly2_15_conc_2_itm_4_0 <= 1'b0;
      butterFly2_15_conc_2_itm_5_0 <= 1'b0;
      INNER_LOOP2_stage_0_10 <= 1'b0;
      butterFly2_15_conc_2_itm_7_0 <= 1'b0;
      butterFly2_15_conc_2_itm_8_0 <= 1'b0;
      butterFly2_15_conc_itm_10_2_1 <= 2'b00;
      butterFly2_15_f1_equal_tmp_1 <= 1'b0;
      butterFly2_15_f1_equal_tmp_7_1 <= 1'b0;
      INNER_LOOP3_r_11_4_sva_6_0 <= 7'b0000000;
      INNER_LOOP4_r_11_4_sva_6_0 <= 7'b0000000;
    end
    else begin
      reg_yt_rsc_0_0_cgo_cse <= or_553_rmff;
      reg_yt_rsc_0_16_cgo_cse <= or_652_rmff;
      reg_yt_rsc_1_0_cgo_cse <= or_718_rmff;
      reg_yt_rsc_1_16_cgo_cse <= or_785_rmff;
      reg_yt_rsc_2_0_cgo_cse <= or_851_rmff;
      reg_yt_rsc_2_16_cgo_cse <= or_918_rmff;
      reg_yt_rsc_3_0_cgo_cse <= or_984_rmff;
      reg_yt_rsc_3_16_cgo_cse <= or_1051_rmff;
      reg_yt_rsc_4_0_cgo_cse <= or_1117_rmff;
      reg_yt_rsc_4_16_cgo_cse <= or_1216_rmff;
      reg_yt_rsc_5_0_cgo_cse <= or_1282_rmff;
      reg_yt_rsc_5_16_cgo_cse <= or_1349_rmff;
      reg_yt_rsc_6_0_cgo_cse <= or_1415_rmff;
      reg_yt_rsc_6_16_cgo_cse <= or_1482_rmff;
      reg_yt_rsc_7_0_cgo_cse <= or_1548_rmff;
      reg_yt_rsc_7_16_cgo_cse <= or_1615_rmff;
      reg_xt_rsc_triosy_7_31_obj_ld_cse <= and_dcpl_62 & (fsm_output[9]);
      reg_ensig_cgo_cse <= or_3599_rmff;
      reg_ensig_cgo_17_cse <= or_3759_rmff;
      butterFly1_15_conc_2_itm_2_1 <= MUX_v_2_2_2(STAGE_LOOP_mux1h_nl, 2'b11, or_4976_cse);
      butterFly1_15_conc_2_itm_9_0 <= butterFly1_15_conc_2_itm_8_0 & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_8_0 <= butterFly1_15_conc_2_itm_7_0 & (~ or_tmp_3650);
      butterFly1_15_f1_equal_tmp_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_nor_nl,
          butterFly1_16_f1_butterFly1_16_f1_nor_nl, butterFly2_f1_butterFly2_f1_and_5_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_5_nl, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9])});
      butterFly1_15_f1_equal_tmp_1_1 <= MUX1HOT_s_1_3_2(butterFly1_f1_butterFly1_f1_and_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_nl, butterFly2_15_conc_2_itm_8_0,
          {(fsm_output[2]) , (fsm_output[4]) , or_dcpl_298});
      butterFly1_15_f1_equal_tmp_2_1 <= MUX1HOT_s_1_3_2(butterFly1_f1_butterFly1_f1_and_1_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_1_nl, butterFly1_15_f1_equal_tmp_1_1,
          {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])});
      butterFly1_15_f1_equal_tmp_3_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_2_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_2_nl, butterFly2_f1_butterFly2_f1_and_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_nl, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9])});
      butterFly1_15_f1_equal_tmp_4_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_3_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_3_nl, butterFly2_f1_butterFly2_f1_and_1_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_1_nl, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9])});
      butterFly1_15_f1_equal_tmp_5_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_4_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_4_nl, butterFly2_f1_butterFly2_f1_and_2_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_2_nl, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9])});
      butterFly1_15_f1_equal_tmp_6_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_5_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_5_nl, butterFly2_f1_butterFly2_f1_and_3_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_3_nl, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9])});
      butterFly1_15_f1_equal_tmp_7_1 <= MUX1HOT_s_1_4_2(butterFly1_f1_butterFly1_f1_and_6_nl,
          butterFly1_16_f1_butterFly1_16_f1_and_6_nl, butterFly2_f1_butterFly2_f1_and_4_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_4_nl, {(fsm_output[2]) , (fsm_output[4])
          , (fsm_output[7]) , (fsm_output[9])});
      INNER_LOOP1_stage_0 <= (INNER_LOOP1_stage_0 & (~ (z_out_62[7]))) | or_tmp_3650;
      INNER_LOOP1_r_11_4_sva_6_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_cse;
      INNER_LOOP1_stage_0_2 <= INNER_LOOP1_mux_nl & (~ or_tmp_3717);
      INNER_LOOP1_stage_0_3 <= INNER_LOOP1_mux_4_nl & (~ or_tmp_3717);
      INNER_LOOP1_stage_0_10 <= INNER_LOOP1_mux_5_nl & (~ or_tmp_3723);
      INNER_LOOP1_stage_0_11 <= INNER_LOOP1_mux_6_nl & (~ or_tmp_3723);
      butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm <= MUX1HOT_v_3_4_2((INNER_LOOP1_r_INNER_LOOP1_r_and_cse[6:4]),
          (INNER_LOOP2_r_11_4_sva_6_0_mx1[6:4]), (INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse[6:4]),
          (INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse[6:4]), {or_tmp_3597 , or_dcpl_315
          , or_tmp_3600 , or_tmp_3732});
      butterFly1_15_conc_2_itm_7_0 <= butterFly1_15_conc_2_itm_6_0 & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_6_0 <= butterFly1_15_conc_2_itm_5_0 & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_5_0 <= butterFly1_15_conc_2_itm_4_0 & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_4_2_1 <= MUX1HOT_v_2_3_2(butterFly1_15_conc_2_itm_3_2_1,
          (INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse[6:5]), (INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse[6:5]),
          {modulo_add_1_qelse_or_m1c , or_tmp_3600 , or_tmp_3732});
      butterFly1_15_conc_2_itm_4_0 <= butterFly1_15_conc_2_itm_3_0 & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_3_0 <= butterFly1_15_conc_2_itm_2_0 & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_2_2_1 <= MUX1HOT_v_2_4_2(butterFly1_15_conc_2_itm_1_2_1,
          (operator_33_true_2_lshift_psp_2_0_sva_mx0[2:1]), operator_33_true_3_lshift_psp_1_0_sva_mx0w5,
          operator_33_true_3_lshift_psp_1_0_sva, {modulo_add_1_qelse_or_m1c , or_tmp_3600
          , (fsm_output[8]) , (fsm_output[9])});
      butterFly1_15_conc_2_itm_2_0 <= butterFly1_15_mux_9_nl & (~ or_tmp_3650);
      butterFly1_15_conc_2_itm_1_0 <= butterFly1_15_conc_2_itm_0 & (~(and_dcpl_239
          & (~ (fsm_output[7]))));
      butterFly1_15_conc_2_itm_0 <= butterFly1_15_mux1h_47_nl & (~(or_4976_cse |
          (fsm_output[5]) | (fsm_output[6]) | (fsm_output[8])));
      butterFly2_15_conc_2_itm_0 <= butterFly2_15_mux1h_3_nl & (~((fsm_output[3])
          | (fsm_output[10]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5])));
      butterFly2_15_conc_2_itm_1_0 <= butterFly2_15_conc_2_itm_0 & or_dcpl_300;
      butterFly2_15_conc_2_itm_2_0 <= butterFly2_15_conc_2_itm_1_0 & or_dcpl_300;
      butterFly2_15_conc_2_itm_3_0 <= butterFly2_15_conc_2_itm_2_0 & or_dcpl_300;
      butterFly2_15_conc_2_itm_4_0 <= butterFly2_15_conc_2_itm_3_0 & or_dcpl_300;
      butterFly2_15_conc_2_itm_5_0 <= butterFly2_15_conc_2_itm_4_0 & or_dcpl_300;
      INNER_LOOP2_stage_0_10 <= butterFly1_15_mux_10_nl & (~ or_tmp_3650);
      butterFly2_15_conc_2_itm_7_0 <= INNER_LOOP1_mux_7_nl & ((fsm_output[4]) | (fsm_output[7])
          | (fsm_output[9]));
      butterFly2_15_conc_2_itm_8_0 <= butterFly2_15_conc_2_itm_7_0 & or_tmp_3842;
      butterFly2_15_conc_itm_10_2_1 <= MUX1HOT_v_2_3_2(butterFly2_15_conc_2_itm_9_2_1,
          operator_33_true_3_lshift_psp_1_0_sva_mx0w5, operator_33_true_3_lshift_psp_1_0_sva,
          {(fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])});
      butterFly2_15_f1_equal_tmp_1 <= MUX_s_1_2_2(butterFly2_f1_butterFly2_f1_nor_nl,
          butterFly2_16_f1_butterFly2_16_f1_nor_nl, fsm_output[9]);
      butterFly2_15_f1_equal_tmp_7_1 <= MUX_s_1_2_2(butterFly2_f1_butterFly2_f1_and_6_nl,
          butterFly2_16_f1_butterFly2_16_f1_and_6_cse, fsm_output[9]);
      INNER_LOOP3_r_11_4_sva_6_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse;
      INNER_LOOP4_r_11_4_sva_6_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse;
    end
  end
  always @(posedge clk) begin
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    modulo_add_1_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_141, (readslicef_33_32_1(acc_2_nl)),
        z_out_138, z_out_136, {modulo_add_1_qelse_and_nl , modulo_add_1_qelse_or_1_nl
        , modulo_add_1_qelse_and_4_nl , modulo_add_1_qelse_and_5_nl});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    modulo_add_10_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_132, (readslicef_33_32_1(acc_3_nl)),
        z_out_127, z_out_128, z_out_142, {modulo_add_10_qelse_and_nl , modulo_add_10_qelse_or_nl
        , modulo_add_10_qelse_and_5_nl , modulo_add_10_qelse_and_6_nl , modulo_add_10_qelse_and_7_nl});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9 <= MUX_v_4_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8,
        (INNER_LOOP3_r_11_4_sva_6_0[4:1]), fsm_output[7]);
    modulo_add_11_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_131, (readslicef_33_32_1(acc_4_nl)),
        z_out_137, z_out_127, z_out_141, {modulo_add_11_qelse_and_nl , modulo_add_11_qelse_or_nl
        , modulo_add_11_qelse_and_5_nl , modulo_add_11_qelse_and_6_nl , modulo_add_11_qelse_and_7_nl});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9 <= MUX1HOT_v_4_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP3_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    modulo_add_12_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_130, (readslicef_33_32_1(acc_5_nl)),
        z_out_142, z_out_140, {modulo_add_12_qelse_and_nl , modulo_add_12_qelse_or_1_nl
        , modulo_add_12_qelse_and_4_nl , modulo_add_12_qelse_and_5_nl});
    modulo_add_13_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_129, (readslicef_33_32_1(acc_6_nl)),
        z_out_141, z_out_139, {modulo_add_13_qelse_and_nl , modulo_add_13_qelse_or_1_nl
        , modulo_add_13_qelse_and_4_nl , modulo_add_13_qelse_and_5_nl});
    modulo_add_14_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_128, (readslicef_33_32_1(acc_10_nl)),
        z_out_140, z_out_138, {modulo_add_14_qelse_and_nl , modulo_add_14_qelse_or_1_nl
        , modulo_add_14_qelse_and_4_nl , modulo_add_14_qelse_and_5_nl});
    modulo_add_15_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_127, (readslicef_33_32_1(acc_14_nl)),
        z_out_142, z_out_139, z_out_137, {modulo_add_15_qelse_and_nl , modulo_add_15_qelse_or_nl
        , modulo_add_15_qelse_and_5_nl , modulo_add_15_qelse_and_6_nl , modulo_add_15_qelse_and_7_nl});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    mult_15_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_15_z_asn_itm_2, mult_31_z_asn_itm_2,
        mult_14_z_asn_itm_2, mult_27_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_14_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_14_z_asn_itm_2, mult_30_z_asn_itm_2,
        mult_26_z_asn_itm_2, mult_15_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_13_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_13_z_asn_itm_2, mult_29_z_asn_itm_2,
        mult_28_z_asn_itm_2, {or_dcpl_353 , (fsm_output[4]) , (fsm_output[9])});
    mult_12_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_12_z_asn_itm_2, mult_28_z_asn_itm_2,
        mult_29_z_asn_itm_2, {or_tmp_3666 , (fsm_output[4]) , (fsm_output[7])});
    mult_11_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_11_z_asn_itm_2, mult_27_z_asn_itm_2,
        mult_15_z_asn_itm_2, mult_26_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_10_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_10_z_asn_itm_2, mult_26_z_asn_itm_2,
        mult_25_z_asn_itm_2, mult_1_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_8 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_7 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    mult_15_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_2_z, mult_z_mul_cmp_22_z,
        mult_z_mul_cmp_20_z, {(fsm_output[2]) , or_dcpl_361 , (fsm_output[9])});
    mult_14_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_4_z, mult_z_mul_cmp_24_z,
        mult_z_mul_cmp_28_z, {or_tmp_3666 , (fsm_output[4]) , (fsm_output[7])});
    mult_13_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_6_z, mult_z_mul_cmp_26_z,
        mult_z_mul_cmp_24_z, mult_z_mul_cmp_12_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_12_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_8_z, mult_z_mul_cmp_28_z,
        mult_z_mul_cmp_12_z, {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    mult_11_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_10_z, mult_z_mul_cmp_30_z,
        mult_z_mul_cmp_8_z, mult_z_mul_cmp_16_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_10_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_12_z, mult_z_mul_cmp_z,
        mult_z_mul_cmp_2_z, {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_7 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_6 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    mult_1_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_30_z, mult_z_mul_cmp_20_z,
        mult_z_mul_cmp_16_z, mult_z_mul_cmp_26_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_6 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_5 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_4 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_5 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_4 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_3 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_3 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_2 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11516_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11005_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10494_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_2 <= MUX1HOT_v_4_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1,
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {or_dcpl_353
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_1 <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10015_itm_9,
        (INNER_LOOP4_r_11_4_sva_6_0[4:1]), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
        , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9472_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8961_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_1 <= MUX_v_4_2_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8450_itm_9, or_tmp_3842);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_1 <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        (INNER_LOOP2_r_11_4_sva_6_0[4:1]), (INNER_LOOP3_r_11_4_sva_6_0[4:1]), (INNER_LOOP4_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_1 <= MUX1HOT_v_4_3_2((INNER_LOOP1_r_11_4_sva_6_0[4:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8, (INNER_LOOP3_r_11_4_sva_6_0[4:1]),
        {(fsm_output[2]) , or_tmp_3755 , (fsm_output[7])});
    mult_16_z_asn_itm_3 <= MUX_v_32_2_2(mult_31_z_asn_itm_2, mult_10_z_asn_itm_2,
        or_dcpl_361);
    mult_17_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_1_z_asn_itm_2, mult_11_z_asn_itm_2,
        mult_31_z_asn_itm_2, mult_10_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_18_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_23_z_asn_itm_2, mult_12_z_asn_itm_2,
        mult_24_z_asn_itm_2, {or_tmp_3666 , (fsm_output[4]) , (fsm_output[7])});
    mult_19_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_24_z_asn_itm_2, mult_13_z_asn_itm_2,
        mult_23_z_asn_itm_2, {or_tmp_3666 , (fsm_output[4]) , (fsm_output[7])});
    mult_20_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_25_z_asn_itm_2, mult_14_z_asn_itm_2,
        mult_28_z_asn_itm_2, mult_13_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_21_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_26_z_asn_itm_2, mult_15_z_asn_itm_2,
        mult_11_z_asn_itm_2, mult_30_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_22_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_27_z_asn_itm_2, mult_1_z_asn_itm_2,
        mult_14_z_asn_itm_2, {or_dcpl_353 , (fsm_output[4]) , (fsm_output[9])});
    mult_23_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_28_z_asn_itm_2, mult_23_z_asn_itm_2,
        mult_1_z_asn_itm_2, mult_25_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_24_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_29_z_asn_itm_2, mult_24_z_asn_itm_2,
        mult_12_z_asn_itm_2, {or_tmp_3666 , (fsm_output[4]) , (fsm_output[7])});
    mult_25_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_30_z_asn_itm_2, mult_25_z_asn_itm_2,
        mult_11_z_asn_itm_2, {or_dcpl_353 , (fsm_output[4]) , (fsm_output[9])});
    modulo_add_23_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_140, (readslicef_33_32_1(acc_18_nl)),
        z_out_137, z_out_135, {modulo_add_23_qelse_and_nl , modulo_add_23_qelse_or_1_nl
        , modulo_add_23_qelse_and_4_nl , modulo_add_23_qelse_and_5_nl});
    modulo_add_24_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_139, (readslicef_33_32_1(acc_22_nl)),
        z_out_136, z_out_134, {modulo_add_24_qelse_and_nl , modulo_add_24_qelse_or_1_nl
        , modulo_add_24_qelse_and_4_nl , modulo_add_24_qelse_and_5_nl});
    modulo_add_25_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_138, (readslicef_33_32_1(acc_26_nl)),
        z_out_135, z_out_133, {modulo_add_25_qelse_and_nl , modulo_add_25_qelse_or_1_nl
        , modulo_add_25_qelse_and_4_nl , modulo_add_25_qelse_and_5_nl});
    modulo_add_26_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_137, (readslicef_33_32_1(acc_30_nl)),
        z_out_136, z_out_134, z_out_132, {modulo_add_26_qelse_and_nl , modulo_add_26_qelse_or_nl
        , modulo_add_26_qelse_and_5_nl , modulo_add_26_qelse_and_6_nl , modulo_add_26_qelse_and_7_nl});
    modulo_add_27_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_136, (readslicef_33_32_1(acc_34_nl)),
        z_out_135, z_out_133, z_out_131, {modulo_add_27_qelse_and_nl , modulo_add_27_qelse_or_nl
        , modulo_add_27_qelse_and_5_nl , modulo_add_27_qelse_and_6_nl , modulo_add_27_qelse_and_7_nl});
    modulo_add_28_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_135, (readslicef_33_32_1(acc_38_nl)),
        z_out_134, z_out_132, z_out_130, {modulo_add_28_qelse_and_nl , modulo_add_28_qelse_or_nl
        , modulo_add_28_qelse_and_5_nl , modulo_add_28_qelse_and_6_nl , modulo_add_28_qelse_and_7_nl});
    modulo_add_29_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_134, (readslicef_33_32_1(acc_42_nl)),
        z_out_133, z_out_131, z_out_129, {modulo_add_29_qelse_and_nl , modulo_add_29_qelse_or_nl
        , modulo_add_29_qelse_and_5_nl , modulo_add_29_qelse_and_6_nl , modulo_add_29_qelse_and_7_nl});
    modulo_add_30_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_133, (readslicef_33_32_1(acc_46_nl)),
        z_out_132, z_out_130, z_out_128, {modulo_add_30_qelse_and_nl , modulo_add_30_qelse_or_nl
        , modulo_add_30_qelse_and_5_nl , modulo_add_30_qelse_and_6_nl , modulo_add_30_qelse_and_7_nl});
    modulo_add_31_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_142, (readslicef_33_32_1(acc_49_nl)),
        z_out_131, z_out_129, z_out_127, {modulo_add_31_qelse_and_nl , modulo_add_31_qelse_or_nl
        , modulo_add_31_qelse_and_5_nl , modulo_add_31_qelse_and_6_nl , modulo_add_31_qelse_and_7_nl});
    mult_23_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_28_z, mult_z_mul_cmp_18_z,
        mult_z_mul_cmp_6_z, mult_z_mul_cmp_10_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_24_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_26_z, mult_z_mul_cmp_16_z,
        mult_z_mul_cmp_10_z, mult_z_mul_cmp_2_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_25_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_24_z, mult_z_mul_cmp_14_z,
        mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_26_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_22_z, mult_z_mul_cmp_12_z,
        mult_z_mul_cmp_26_z, mult_z_mul_cmp_18_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_27_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_20_z, mult_z_mul_cmp_10_z,
        mult_z_mul_cmp_30_z, mult_z_mul_cmp_24_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_28_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z,
        mult_z_mul_cmp_20_z, mult_z_mul_cmp_30_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_29_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_16_z, mult_z_mul_cmp_6_z,
        mult_z_mul_cmp_14_z, mult_z_mul_cmp_22_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_30_z_asn_itm_1 <= MUX_v_32_2_2(mult_z_mul_cmp_14_z, mult_z_mul_cmp_4_z,
        or_dcpl_361);
    mult_31_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_z, mult_z_mul_cmp_2_z,
        mult_z_mul_cmp_6_z, {or_dcpl_353 , (fsm_output[4]) , (fsm_output[9])});
    tmp_10_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_64_lpi_3_dfm_1, tmp_10_lpi_3_dfm_1,
        tmp_100_lpi_3_dfm_1, tmp_32_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_102_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_66_lpi_3_dfm_1, tmp_12_lpi_3_dfm_1,
        tmp_102_lpi_3_dfm_1, tmp_34_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_104_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_68_lpi_3_dfm_1, tmp_14_lpi_3_dfm_1,
        tmp_104_lpi_3_dfm_1, tmp_36_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_106_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_70_lpi_3_dfm_1, tmp_16_lpi_3_dfm_1,
        tmp_106_lpi_3_dfm_1, tmp_38_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_108_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_72_lpi_3_dfm_1, tmp_18_lpi_3_dfm_1,
        tmp_108_lpi_3_dfm_1, tmp_40_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_110_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_74_lpi_3_dfm_1, tmp_2_lpi_3_dfm_1,
        tmp_110_lpi_3_dfm_1, tmp_42_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_112_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_76_lpi_3_dfm_1, tmp_20_lpi_3_dfm_1,
        tmp_112_lpi_3_dfm_1, tmp_44_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_114_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_78_lpi_3_dfm_1, tmp_22_lpi_3_dfm_1,
        tmp_114_lpi_3_dfm_1, tmp_46_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_116_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_80_lpi_3_dfm_1, tmp_24_lpi_3_dfm_1,
        tmp_116_lpi_3_dfm_1, tmp_48_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_118_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_82_lpi_3_dfm_1, tmp_26_lpi_3_dfm_1,
        tmp_118_lpi_3_dfm_1, tmp_50_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_120_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_84_lpi_3_dfm_1, tmp_28_lpi_3_dfm_1,
        tmp_120_lpi_3_dfm_1, tmp_52_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_122_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_86_lpi_3_dfm_1, tmp_30_lpi_3_dfm_1,
        tmp_122_lpi_3_dfm_1, tmp_54_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_124_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_88_lpi_3_dfm_1, tmp_4_lpi_3_dfm_1,
        tmp_124_lpi_3_dfm_1, tmp_56_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_126_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_90_lpi_3_dfm_1, tmp_6_lpi_3_dfm_1,
        tmp_126_lpi_3_dfm_1, tmp_58_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_60_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_92_lpi_3_dfm_1, tmp_8_lpi_3_dfm_1,
        tmp_96_lpi_3_dfm_1, tmp_60_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    tmp_62_lpi_3_dfm_2 <= MUX1HOT_v_32_4_2(tmp_94_lpi_3_dfm_1, tmp_lpi_3_dfm_1, tmp_98_lpi_3_dfm_1,
        tmp_62_lpi_3_dfm_1, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
        , (fsm_output[9])});
    reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd <= (z_out_109[31]) & (~(modulo_sub_16_qelse_and_ssc
        | modulo_sub_16_qelse_and_ssc_1));
    reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_126[30:0]),
        (z_out_109[30:0]), (z_out_111[30:0]), {modulo_sub_16_qelse_and_ssc , modulo_sub_16_qelse_or_nl
        , modulo_sub_16_qelse_and_ssc_1});
    reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd <= (z_out_106[31]) & (~(modulo_sub_17_qelse_and_ssc
        | modulo_sub_17_qelse_and_ssc_1));
    reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_116[30:0]),
        (z_out_106[30:0]), (z_out_112[30:0]), {modulo_sub_17_qelse_and_ssc , modulo_sub_17_qelse_or_nl
        , modulo_sub_17_qelse_and_ssc_1});
    reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd <= (z_out_104[31]) & (~(modulo_sub_18_qelse_and_ssc
        | modulo_sub_18_qelse_and_ssc_1));
    reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_123[30:0]),
        (z_out_104[30:0]), (z_out_113[30:0]), {modulo_sub_18_qelse_and_ssc , modulo_sub_18_qelse_or_nl
        , modulo_sub_18_qelse_and_ssc_1});
    reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd <= (z_out_101[31]) & (~(modulo_sub_19_qelse_and_ssc
        | modulo_sub_19_qelse_and_ssc_1));
    reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_124[30:0]),
        (z_out_101[30:0]), (z_out_114[30:0]), {modulo_sub_19_qelse_and_ssc , modulo_sub_19_qelse_or_nl
        , modulo_sub_19_qelse_and_ssc_1});
    reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd <= (z_out_98[31]) & (~(modulo_sub_20_qelse_and_ssc
        | modulo_sub_20_qelse_and_ssc_1));
    reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_125[30:0]),
        (z_out_98[30:0]), (z_out_115[30:0]), {modulo_sub_20_qelse_and_ssc , modulo_sub_20_qelse_or_nl
        , modulo_sub_20_qelse_and_ssc_1});
    reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd <= (z_out_96[31]) & (~(modulo_sub_21_qelse_and_ssc
        | modulo_sub_21_qelse_and_ssc_1));
    reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_111[30:0]),
        (z_out_96[30:0]), (z_out_116[30:0]), {modulo_sub_21_qelse_and_ssc , modulo_sub_21_qelse_or_nl
        , modulo_sub_21_qelse_and_ssc_1});
    reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd <= (z_out_93[31]) & (~(modulo_sub_22_qelse_and_ssc
        | modulo_sub_22_qelse_and_ssc_1));
    reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_112[30:0]),
        (z_out_93[30:0]), (z_out_117[30:0]), {modulo_sub_22_qelse_and_ssc , modulo_sub_22_qelse_or_nl
        , modulo_sub_22_qelse_and_ssc_1});
    reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd <= (z_out_90[31]) & (~(modulo_sub_23_qelse_and_ssc
        | modulo_sub_23_qelse_and_ssc_1));
    reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_113[30:0]),
        (z_out_90[30:0]), (z_out_118[30:0]), {modulo_sub_23_qelse_and_ssc , modulo_sub_23_qelse_or_nl
        , modulo_sub_23_qelse_and_ssc_1});
    reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd <= (z_out_88[31]) & (~(modulo_sub_24_qelse_and_ssc
        | modulo_sub_24_qelse_and_ssc_1));
    reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_114[30:0]),
        (z_out_88[30:0]), (z_out_119[30:0]), {modulo_sub_24_qelse_and_ssc , modulo_sub_24_qelse_or_nl
        , modulo_sub_24_qelse_and_ssc_1});
    reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd <= (z_out_85[31]) & (~(modulo_sub_25_qelse_and_ssc
        | modulo_sub_25_qelse_and_ssc_1));
    reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_115[30:0]),
        (z_out_85[30:0]), (z_out_120[30:0]), {modulo_sub_25_qelse_and_ssc , modulo_sub_25_qelse_or_nl
        , modulo_sub_25_qelse_and_ssc_1});
    reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd <= (z_out_82[31]) & (~(modulo_sub_26_qelse_and_ssc
        | modulo_sub_26_qelse_and_ssc_1));
    reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_117[30:0]),
        (z_out_82[30:0]), (z_out_121[30:0]), {modulo_sub_26_qelse_and_ssc , modulo_sub_26_qelse_or_nl
        , modulo_sub_26_qelse_and_ssc_1});
    reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd <= (z_out_80[31]) & (~(modulo_sub_27_qelse_and_ssc
        | modulo_sub_27_qelse_and_ssc_1));
    reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_118[30:0]),
        (z_out_80[30:0]), (z_out_122[30:0]), {modulo_sub_27_qelse_and_ssc , modulo_sub_27_qelse_or_nl
        , modulo_sub_27_qelse_and_ssc_1});
    reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd <= (z_out_77[31]) & (~(modulo_sub_28_qelse_and_ssc
        | modulo_sub_28_qelse_and_ssc_1));
    reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_119[30:0]),
        (z_out_77[30:0]), (z_out_123[30:0]), {modulo_sub_28_qelse_and_ssc , modulo_sub_28_qelse_or_nl
        , modulo_sub_28_qelse_and_ssc_1});
    reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd <= (z_out_74[31]) & (~(modulo_sub_29_qelse_and_ssc
        | modulo_sub_29_qelse_and_ssc_1));
    reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_120[30:0]),
        (z_out_74[30:0]), (z_out_124[30:0]), {modulo_sub_29_qelse_and_ssc , modulo_sub_29_qelse_or_nl
        , modulo_sub_29_qelse_and_ssc_1});
    reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd <= (z_out_72[31]) & (~(modulo_sub_30_qelse_and_ssc
        | modulo_sub_30_qelse_and_ssc_1));
    reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_121[30:0]),
        (z_out_72[30:0]), (z_out_125[30:0]), {modulo_sub_30_qelse_and_ssc , modulo_sub_30_qelse_or_nl
        , modulo_sub_30_qelse_and_ssc_1});
    reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd <= (z_out_69[31]) & (~(modulo_sub_31_qelse_and_ssc
        | modulo_sub_31_qelse_and_ssc_1));
    reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_122[30:0]),
        (z_out_69[30:0]), (z_out_126[30:0]), {modulo_sub_31_qelse_and_ssc , modulo_sub_31_qelse_or_nl
        , modulo_sub_31_qelse_and_ssc_1});
    INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8;
    INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_1 <= MUX_v_4_2_2((INNER_LOOP2_r_11_4_sva_6_0[4:1]),
        (INNER_LOOP4_r_11_4_sva_6_0[4:1]), fsm_output[9]);
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_conc_2_itm_9_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_5_0 | butterFly2_15_conc_2_itm_5_0 ) begin
      butterFly1_15_conc_2_itm_9_2_1 <= butterFly1_15_conc_2_itm_8_2_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_4_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_19
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_8833_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_22
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9344_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_25
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_9855_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_8_0 | butterFly1_15_conc_2_itm_9_0 | butterFly2_15_conc_2_itm_4_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10366_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_30
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_10877_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_33
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11388_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_5_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_36
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_11899_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_9_0 | butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_5_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_conc_2_itm_8_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_4_0 ) begin
      butterFly1_15_conc_2_itm_8_2_1 <= butterFly1_15_conc_2_itm_7_2_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly2_15_conc_2_itm_4_0 ) begin
      reg_mult_15_res_lpi_3_dfm_1_cse <= mult_15_res_lpi_3_dfm_1_mx0;
      reg_mult_14_res_lpi_3_dfm_1_cse <= mult_14_res_lpi_3_dfm_1_mx0;
      reg_mult_13_res_lpi_3_dfm_1_cse <= mult_13_res_lpi_3_dfm_1_mx0;
      reg_mult_12_res_lpi_3_dfm_1_cse <= mult_12_res_lpi_3_dfm_1_mx0;
      reg_mult_11_res_lpi_3_dfm_1_cse <= mult_11_res_lpi_3_dfm_1_mx0;
      reg_mult_10_res_lpi_3_dfm_1_cse <= mult_10_res_lpi_3_dfm_1_mx0;
      reg_mult_9_res_lpi_3_dfm_1_cse <= mult_9_res_lpi_3_dfm_1_mx0;
      reg_mult_8_res_lpi_3_dfm_1_cse <= mult_8_res_lpi_3_dfm_1_mx0;
      reg_mult_7_res_lpi_3_dfm_1_cse <= mult_7_res_lpi_3_dfm_1_mx0;
      reg_mult_6_res_lpi_3_dfm_1_cse <= mult_6_res_lpi_3_dfm_1_mx0;
      reg_mult_5_res_lpi_3_dfm_1_cse <= mult_5_res_lpi_3_dfm_1_mx0;
      reg_mult_4_res_lpi_3_dfm_1_cse <= mult_4_res_lpi_3_dfm_1_mx0;
      reg_mult_3_res_lpi_3_dfm_1_cse <= mult_3_res_lpi_3_dfm_1_mx0;
      reg_mult_2_res_lpi_3_dfm_1_cse <= mult_2_res_lpi_3_dfm_1_mx0;
      reg_mult_1_res_lpi_3_dfm_1_cse <= mult_1_res_lpi_3_dfm_1_mx0;
      reg_mult_res_lpi_3_dfm_1_cse <= mult_res_lpi_3_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1 <= 3'b000;
      butterFly1_15_conc_2_itm_1_2_1 <= 2'b00;
      butterFly2_15_tw_equal_tmp_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_3_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_5_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_6_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_7_1 <= 1'b0;
    end
    else if ( INNER_LOOP1_stage_0 ) begin
      butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm_1 <= butterFly1_15_f1_slc_INNER_LOOP1_r_11_4_6_4_itm;
      butterFly1_15_conc_2_itm_1_2_1 <= butterFly1_15_conc_2_itm_2_1;
      butterFly2_15_tw_equal_tmp_1 <= ~((operator_20_false_acc_cse_sva!=3'b000));
      butterFly2_15_tw_equal_tmp_3_1 <= (operator_20_false_acc_cse_sva==3'b011);
      butterFly2_15_tw_equal_tmp_5_1 <= (operator_20_false_acc_cse_sva==3'b101);
      butterFly2_15_tw_equal_tmp_6_1 <= (operator_20_false_acc_cse_sva==3'b110);
      butterFly2_15_tw_equal_tmp_7_1 <= (operator_20_false_acc_cse_sva==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_20_false_acc_cse_sva <= 3'b000;
    end
    else if ( ~(or_dcpl_315 | or_dcpl_353) ) begin
      operator_20_false_acc_cse_sva <= MUX_v_3_2_2(z_out_61, (z_out_60[2:0]), fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_conc_2_itm_7_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_3_0 | butterFly2_15_conc_2_itm_3_0 ) begin
      butterFly1_15_conc_2_itm_7_2_1 <= butterFly1_15_conc_2_itm_6_2_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_8_0
        | butterFly2_15_conc_2_itm_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_5_0 | butterFly1_15_conc_2_itm_8_0 | or_dcpl_36
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_12 ) begin
      mult_15_z_asn_itm_2 <= mult_15_z_asn_itm_1;
      mult_14_z_asn_itm_2 <= mult_14_z_asn_itm_1;
      mult_13_z_asn_itm_2 <= mult_13_z_asn_itm_1;
      mult_12_z_asn_itm_2 <= mult_12_z_asn_itm_1;
      mult_11_z_asn_itm_2 <= mult_11_z_asn_itm_1;
      mult_10_z_asn_itm_2 <= mult_10_z_asn_itm_1;
      mult_1_z_asn_itm_2 <= mult_1_z_asn_itm_1;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_5;
      mult_23_z_asn_itm_2 <= mult_23_z_asn_itm_1;
      mult_24_z_asn_itm_2 <= mult_24_z_asn_itm_1;
      mult_25_z_asn_itm_2 <= mult_25_z_asn_itm_1;
      mult_26_z_asn_itm_2 <= mult_26_z_asn_itm_1;
      mult_27_z_asn_itm_2 <= mult_27_z_asn_itm_1;
      mult_28_z_asn_itm_2 <= mult_28_z_asn_itm_1;
      mult_29_z_asn_itm_2 <= mult_29_z_asn_itm_1;
      mult_30_z_asn_itm_2 <= mult_30_z_asn_itm_1;
      mult_31_z_asn_itm_2 <= mult_31_z_asn_itm_1;
      tmp_10_lpi_3_dfm_5 <= tmp_10_lpi_3_dfm_4;
      tmp_102_lpi_3_dfm_5 <= tmp_102_lpi_3_dfm_4;
      tmp_104_lpi_3_dfm_5 <= tmp_104_lpi_3_dfm_4;
      tmp_106_lpi_3_dfm_5 <= tmp_106_lpi_3_dfm_4;
      tmp_108_lpi_3_dfm_5 <= tmp_108_lpi_3_dfm_4;
      tmp_110_lpi_3_dfm_5 <= tmp_110_lpi_3_dfm_4;
      tmp_112_lpi_3_dfm_5 <= tmp_112_lpi_3_dfm_4;
      tmp_114_lpi_3_dfm_5 <= tmp_114_lpi_3_dfm_4;
      tmp_116_lpi_3_dfm_5 <= tmp_116_lpi_3_dfm_4;
      tmp_118_lpi_3_dfm_5 <= tmp_118_lpi_3_dfm_4;
      tmp_120_lpi_3_dfm_5 <= tmp_120_lpi_3_dfm_4;
      tmp_122_lpi_3_dfm_5 <= tmp_122_lpi_3_dfm_4;
      tmp_124_lpi_3_dfm_5 <= tmp_124_lpi_3_dfm_4;
      tmp_126_lpi_3_dfm_5 <= tmp_126_lpi_3_dfm_4;
      tmp_60_lpi_3_dfm_5 <= tmp_60_lpi_3_dfm_4;
      tmp_62_lpi_3_dfm_5 <= tmp_62_lpi_3_dfm_4;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_5;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_5_0 | butterFly2_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_8_0
        | butterFly2_15_conc_2_itm_1_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_8_0 | or_dcpl_33
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_6_0 | butterFly2_15_conc_2_itm_3_0 | butterFly1_15_conc_2_itm_8_0
        | butterFly2_15_conc_2_itm_2_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_63 | or_dcpl_30 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_63 | butterFly2_15_conc_2_itm_3_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_8 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_7;
      tmp_10_lpi_3_dfm_7 <= tmp_10_lpi_3_dfm_6;
      tmp_102_lpi_3_dfm_7 <= tmp_102_lpi_3_dfm_6;
      tmp_104_lpi_3_dfm_7 <= tmp_104_lpi_3_dfm_6;
      tmp_106_lpi_3_dfm_7 <= tmp_106_lpi_3_dfm_6;
      tmp_108_lpi_3_dfm_7 <= tmp_108_lpi_3_dfm_6;
      tmp_110_lpi_3_dfm_7 <= tmp_110_lpi_3_dfm_6;
      tmp_112_lpi_3_dfm_7 <= tmp_112_lpi_3_dfm_6;
      tmp_114_lpi_3_dfm_7 <= tmp_114_lpi_3_dfm_6;
      tmp_116_lpi_3_dfm_7 <= tmp_116_lpi_3_dfm_6;
      tmp_118_lpi_3_dfm_7 <= tmp_118_lpi_3_dfm_6;
      tmp_120_lpi_3_dfm_7 <= tmp_120_lpi_3_dfm_6;
      tmp_122_lpi_3_dfm_7 <= tmp_122_lpi_3_dfm_6;
      tmp_124_lpi_3_dfm_7 <= tmp_124_lpi_3_dfm_6;
      tmp_126_lpi_3_dfm_7 <= tmp_126_lpi_3_dfm_6;
      tmp_60_lpi_3_dfm_7 <= tmp_60_lpi_3_dfm_6;
      tmp_62_lpi_3_dfm_7 <= tmp_62_lpi_3_dfm_6;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_7;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_8_0 | butterFly2_15_conc_2_itm_3_0 | butterFly2_15_conc_2_itm_4_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_70 | butterFly2_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_5_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_70 | or_dcpl_72 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_76 | or_dcpl_25 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_76 | or_dcpl_78 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_80 | or_dcpl_22 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_80 | or_dcpl_82 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_4_0 | butterFly1_15_conc_2_itm_8_0 | or_dcpl_19
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_conc_2_itm_6_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_2_0 ) begin
      butterFly1_15_conc_2_itm_6_2_1 <= butterFly1_15_conc_2_itm_5_2_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_89 | or_dcpl_88 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_10 | or_dcpl_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_94 | or_dcpl_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_10 | or_dcpl ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_94 | or_dcpl ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_10 | or_dcpl_12 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_7_0 | butterFly1_15_conc_2_itm_6_0 | butterFly2_15_conc_2_itm_2_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_10 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_6;
      tmp_10_lpi_3_dfm_6 <= tmp_10_lpi_3_dfm_5;
      tmp_102_lpi_3_dfm_6 <= tmp_102_lpi_3_dfm_5;
      tmp_104_lpi_3_dfm_6 <= tmp_104_lpi_3_dfm_5;
      tmp_106_lpi_3_dfm_6 <= tmp_106_lpi_3_dfm_5;
      tmp_108_lpi_3_dfm_6 <= tmp_108_lpi_3_dfm_5;
      tmp_110_lpi_3_dfm_6 <= tmp_110_lpi_3_dfm_5;
      tmp_112_lpi_3_dfm_6 <= tmp_112_lpi_3_dfm_5;
      tmp_114_lpi_3_dfm_6 <= tmp_114_lpi_3_dfm_5;
      tmp_116_lpi_3_dfm_6 <= tmp_116_lpi_3_dfm_5;
      tmp_118_lpi_3_dfm_6 <= tmp_118_lpi_3_dfm_5;
      tmp_120_lpi_3_dfm_6 <= tmp_120_lpi_3_dfm_5;
      tmp_122_lpi_3_dfm_6 <= tmp_122_lpi_3_dfm_5;
      tmp_124_lpi_3_dfm_6 <= tmp_124_lpi_3_dfm_5;
      tmp_126_lpi_3_dfm_6 <= tmp_126_lpi_3_dfm_5;
      tmp_60_lpi_3_dfm_6 <= tmp_60_lpi_3_dfm_5;
      tmp_62_lpi_3_dfm_6 <= tmp_62_lpi_3_dfm_5;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_6;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_7_0 | butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_3_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_10 | or_dcpl_8 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_94 | or_dcpl_8 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_105 | or_dcpl_72 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_105 | or_dcpl_107 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_109 | or_dcpl_78 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_109 | or_dcpl_111 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_89 | or_dcpl_82 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_conc_2_itm_5_2_1 <= 2'b00;
    end
    else if ( INNER_LOOP1_stage_0 | butterFly2_15_conc_2_itm_1_0 ) begin
      butterFly1_15_conc_2_itm_5_2_1 <= butterFly1_15_conc_2_itm_4_2_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_117 | or_dcpl_116 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_119 | or_dcpl_88 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_119 | or_dcpl_121 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_12 | or_dcpl_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_125 | or_dcpl_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_12 | or_dcpl ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_6_0 | butterFly1_15_conc_2_itm_5_0 | butterFly2_15_conc_2_itm_1_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_6_0 | butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_2_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_133 | butterFly2_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_3_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_133 | or_dcpl_135 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_12 | or_dcpl_8 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_125 | or_dcpl_8 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_139 | or_dcpl_107 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_139 | or_dcpl_141 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_117 | or_dcpl_111 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_146 | or_dcpl_116 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_146 | or_dcpl_148 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_150 | or_dcpl_121 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_150 | or_dcpl_152 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl | or_dcpl_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_5_0 | butterFly1_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_4;
      tmp_10_lpi_3_dfm_4 <= tmp_10_lpi_3_dfm_3;
      tmp_102_lpi_3_dfm_4 <= tmp_102_lpi_3_dfm_3;
      tmp_104_lpi_3_dfm_4 <= tmp_104_lpi_3_dfm_3;
      tmp_106_lpi_3_dfm_4 <= tmp_106_lpi_3_dfm_3;
      tmp_108_lpi_3_dfm_4 <= tmp_108_lpi_3_dfm_3;
      tmp_110_lpi_3_dfm_4 <= tmp_110_lpi_3_dfm_3;
      tmp_112_lpi_3_dfm_4 <= tmp_112_lpi_3_dfm_3;
      tmp_114_lpi_3_dfm_4 <= tmp_114_lpi_3_dfm_3;
      tmp_116_lpi_3_dfm_4 <= tmp_116_lpi_3_dfm_3;
      tmp_118_lpi_3_dfm_4 <= tmp_118_lpi_3_dfm_3;
      tmp_120_lpi_3_dfm_4 <= tmp_120_lpi_3_dfm_3;
      tmp_122_lpi_3_dfm_4 <= tmp_122_lpi_3_dfm_3;
      tmp_124_lpi_3_dfm_4 <= tmp_124_lpi_3_dfm_3;
      tmp_126_lpi_3_dfm_4 <= tmp_126_lpi_3_dfm_3;
      tmp_60_lpi_3_dfm_4 <= tmp_60_lpi_3_dfm_3;
      tmp_62_lpi_3_dfm_4 <= tmp_62_lpi_3_dfm_3;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_4;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_5_0 | butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_1_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_161 | butterFly2_15_conc_2_itm_1_0 | butterFly2_15_conc_2_itm_2_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_161 | or_dcpl_163 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_165 | or_dcpl_135 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_165 | or_dcpl_167 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl | or_dcpl_8 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_5_0 | butterFly2_15_conc_2_itm_0 | or_dcpl_8 )
        begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_171 | or_dcpl_141 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_171 | or_dcpl_173 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly1_15_conc_2_itm_3_2_1 <= 2'b00;
    end
    else if ( INNER_LOOP1_stage_0 | INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_8_0
        ) begin
      butterFly1_15_conc_2_itm_3_2_1 <= butterFly1_15_conc_2_itm_2_2_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_181 | or_dcpl_180 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_185 | or_dcpl_148 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_185 | or_dcpl_187 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15476_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_189 | or_dcpl_152 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_189 | INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_8_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_3;
      tmp_10_lpi_3_dfm_3 <= tmp_10_lpi_3_dfm_2;
      tmp_102_lpi_3_dfm_3 <= tmp_102_lpi_3_dfm_2;
      tmp_104_lpi_3_dfm_3 <= tmp_104_lpi_3_dfm_2;
      tmp_106_lpi_3_dfm_3 <= tmp_106_lpi_3_dfm_2;
      tmp_108_lpi_3_dfm_3 <= tmp_108_lpi_3_dfm_2;
      tmp_110_lpi_3_dfm_3 <= tmp_110_lpi_3_dfm_2;
      tmp_112_lpi_3_dfm_3 <= tmp_112_lpi_3_dfm_2;
      tmp_114_lpi_3_dfm_3 <= tmp_114_lpi_3_dfm_2;
      tmp_116_lpi_3_dfm_3 <= tmp_116_lpi_3_dfm_2;
      tmp_118_lpi_3_dfm_3 <= tmp_118_lpi_3_dfm_2;
      tmp_120_lpi_3_dfm_3 <= tmp_120_lpi_3_dfm_2;
      tmp_122_lpi_3_dfm_3 <= tmp_122_lpi_3_dfm_2;
      tmp_124_lpi_3_dfm_3 <= tmp_124_lpi_3_dfm_2;
      tmp_126_lpi_3_dfm_3 <= tmp_126_lpi_3_dfm_2;
      tmp_60_lpi_3_dfm_3 <= tmp_60_lpi_3_dfm_2;
      tmp_62_lpi_3_dfm_3 <= tmp_62_lpi_3_dfm_2;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_3;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_4_0 | INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_197 | butterFly2_15_conc_2_itm_0 | butterFly2_15_conc_2_itm_1_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_197 | or_dcpl_199 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_201 | or_dcpl_163 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_201 | or_dcpl_203 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_205 | or_dcpl_167 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_205 | or_dcpl_207 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_4_0 | butterFly2_15_conc_2_itm_0 | or_dcpl_8 )
        begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_4_0 | butterFly1_15_conc_2_itm_8_0 | or_dcpl_210
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_181 | or_dcpl_173 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_80 | or_dcpl_215 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16498_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_218 | or_dcpl_180 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_218 | or_dcpl_220 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15987_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_224 | or_dcpl_187 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15093_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_224 | INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_7_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14965_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_3_0 | INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_8_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_3_0 | INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_8_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14454_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_189 | INNER_LOOP1_stage_0_3 | butterFly2_15_conc_2_itm_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_189 | or_dcpl_234 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13943_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_150 | or_dcpl_199 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_150 | or_dcpl_238 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13432_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_119 | or_dcpl_203 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_119 | or_dcpl_242 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12921_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_89 | or_dcpl_207 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_89 | or_dcpl_246 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12410_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_80 | or_dcpl_210 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_stage_0_2 ) begin
      tmp_94_lpi_3_dfm_1 <= z_out;
      tmp_92_lpi_3_dfm_1 <= z_out_1;
      tmp_90_lpi_3_dfm_1 <= z_out_2;
      tmp_88_lpi_3_dfm_1 <= z_out_3;
      tmp_86_lpi_3_dfm_1 <= z_out_4;
      tmp_84_lpi_3_dfm_1 <= z_out_5;
      tmp_82_lpi_3_dfm_1 <= z_out_6;
      tmp_80_lpi_3_dfm_1 <= z_out_7;
      tmp_78_lpi_3_dfm_1 <= z_out_8;
      tmp_76_lpi_3_dfm_1 <= z_out_9;
      tmp_74_lpi_3_dfm_1 <= z_out_10;
      tmp_72_lpi_3_dfm_1 <= z_out_11;
      tmp_70_lpi_3_dfm_1 <= z_out_12;
      tmp_68_lpi_3_dfm_1 <= z_out_13;
      tmp_66_lpi_3_dfm_1 <= z_out_14;
      tmp_64_lpi_3_dfm_1 <= z_out_15;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_8_0 | or_dcpl_215
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_16115_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_9_0 | or_dcpl_220
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_15604_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | INNER_LOOP1_stage_0_2 | butterFly2_15_conc_2_itm_7_0
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14582_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_3_0 | INNER_LOOP1_stage_0_2
        | butterFly2_15_conc_2_itm_8_0 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_14071_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_4_0 | or_dcpl_234
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13560_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_5_0 | or_dcpl_238
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_13049_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_6_0 | or_dcpl_242
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12538_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly1_15_conc_2_itm_7_0 | or_dcpl_246
        ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_12027_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      INNER_LOOP2_r_11_4_sva_6_0 <= 7'b0000000;
    end
    else if ( ~ (fsm_output[2]) ) begin
      INNER_LOOP2_r_11_4_sva_6_0 <= MUX_v_7_2_2(7'b0000000, STAGE_LOOP_base_STAGE_LOOP_base_mux_nl,
          INNER_LOOP2_r_or_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly2_15_conc_2_itm_6_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_6_0 | INNER_LOOP1_stage_0_10 ) begin
      butterFly2_15_conc_2_itm_6_2_1 <= butterFly1_15_conc_2_itm_9_2_1;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_274 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9472_itm_8;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( ~ (fsm_output[4]) ) begin
      operator_33_true_1_lshift_psp_9_4_sva <= z_out_60[9:4];
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_3_0 | butterFly2_15_conc_2_itm_8_0 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( butterFly2_15_conc_2_itm_7_0 ) begin
      tmp_30_lpi_3_dfm_1 <= z_out_16;
      tmp_28_lpi_3_dfm_1 <= z_out_17;
      tmp_26_lpi_3_dfm_1 <= z_out_18;
      tmp_24_lpi_3_dfm_1 <= z_out_19;
      tmp_22_lpi_3_dfm_1 <= z_out_20;
      tmp_20_lpi_3_dfm_1 <= z_out_21;
      tmp_18_lpi_3_dfm_1 <= z_out_22;
      tmp_16_lpi_3_dfm_1 <= z_out_23;
      tmp_14_lpi_3_dfm_1 <= z_out_24;
      tmp_12_lpi_3_dfm_1 <= z_out_25;
      tmp_10_lpi_3_dfm_1 <= z_out_26;
      tmp_8_lpi_3_dfm_1 <= z_out_27;
      tmp_6_lpi_3_dfm_1 <= z_out_28;
      tmp_4_lpi_3_dfm_1 <= z_out_29;
      tmp_2_lpi_3_dfm_1 <= z_out_30;
      tmp_lpi_3_dfm_1 <= z_out_31;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 | butterFly2_15_conc_2_itm_7_0 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_9855_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly2_15_conc_2_itm_9_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_9_0 ) begin
      butterFly2_15_conc_2_itm_9_2_1 <= butterFly2_15_conc_2_itm_8_2_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_8_0 ) begin
      reg_mult_47_res_lpi_3_dfm_1_cse <= mult_1_res_lpi_3_dfm_1_mx0;
      reg_mult_46_res_lpi_3_dfm_1_cse <= mult_9_res_lpi_3_dfm_1_mx0;
      reg_mult_45_res_lpi_3_dfm_1_cse <= mult_12_res_lpi_3_dfm_1_mx0;
      reg_mult_44_res_lpi_3_dfm_1_cse <= mult_4_res_lpi_3_dfm_1_mx0;
      reg_mult_43_res_lpi_3_dfm_1_cse <= mult_6_res_lpi_3_dfm_1_mx0;
      reg_mult_42_res_lpi_3_dfm_1_cse <= mult_14_res_lpi_3_dfm_1_mx0;
      reg_mult_41_res_lpi_3_dfm_1_cse <= mult_10_res_lpi_3_dfm_1_mx0;
      reg_mult_40_res_lpi_3_dfm_1_cse <= mult_2_res_lpi_3_dfm_1_mx0;
      reg_mult_39_res_lpi_3_dfm_1_cse <= mult_3_res_lpi_3_dfm_1_mx0;
      reg_mult_38_res_lpi_3_dfm_1_cse <= mult_7_res_lpi_3_dfm_1_mx0;
      reg_mult_37_res_lpi_3_dfm_1_cse <= mult_11_res_lpi_3_dfm_1_mx0;
      reg_mult_36_res_lpi_3_dfm_1_cse <= mult_15_res_lpi_3_dfm_1_mx0;
      reg_mult_35_res_lpi_3_dfm_1_cse <= mult_13_res_lpi_3_dfm_1_mx0;
      reg_mult_34_res_lpi_3_dfm_1_cse <= mult_8_res_lpi_3_dfm_1_mx0;
      reg_mult_33_res_lpi_3_dfm_1_cse <= mult_5_res_lpi_3_dfm_1_mx0;
      reg_mult_32_res_lpi_3_dfm_1_cse <= mult_res_lpi_3_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly2_15_conc_2_itm_8_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_8_0 ) begin
      butterFly2_15_conc_2_itm_8_2_1 <= butterFly2_15_conc_2_itm_7_2_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly2_15_conc_2_itm_7_2_1 <= 2'b00;
    end
    else if ( butterFly1_15_conc_2_itm_7_0 ) begin
      butterFly2_15_conc_2_itm_7_2_1 <= butterFly2_15_conc_2_itm_6_2_1;
    end
  end
  always @(posedge clk) begin
    if ( butterFly1_15_conc_2_itm_2_0 ) begin
      tmp_126_lpi_3_dfm_1 <= z_out;
      tmp_124_lpi_3_dfm_1 <= z_out_1;
      tmp_122_lpi_3_dfm_1 <= z_out_2;
      tmp_120_lpi_3_dfm_1 <= z_out_3;
      tmp_118_lpi_3_dfm_1 <= z_out_4;
      tmp_116_lpi_3_dfm_1 <= z_out_5;
      tmp_114_lpi_3_dfm_1 <= z_out_6;
      tmp_112_lpi_3_dfm_1 <= z_out_7;
      tmp_110_lpi_3_dfm_1 <= z_out_8;
      tmp_108_lpi_3_dfm_1 <= z_out_9;
      tmp_106_lpi_3_dfm_1 <= z_out_10;
      tmp_104_lpi_3_dfm_1 <= z_out_11;
      tmp_102_lpi_3_dfm_1 <= z_out_12;
      tmp_100_lpi_3_dfm_1 <= z_out_13;
      tmp_98_lpi_3_dfm_1 <= z_out_14;
      tmp_96_lpi_3_dfm_1 <= z_out_15;
      tmp_62_lpi_3_dfm_1 <= z_out_16;
      tmp_60_lpi_3_dfm_1 <= z_out_17;
      tmp_58_lpi_3_dfm_1 <= z_out_18;
      tmp_56_lpi_3_dfm_1 <= z_out_19;
      tmp_54_lpi_3_dfm_1 <= z_out_20;
      tmp_52_lpi_3_dfm_1 <= z_out_21;
      tmp_50_lpi_3_dfm_1 <= z_out_22;
      tmp_48_lpi_3_dfm_1 <= z_out_23;
      tmp_46_lpi_3_dfm_1 <= z_out_24;
      tmp_44_lpi_3_dfm_1 <= z_out_25;
      tmp_42_lpi_3_dfm_1 <= z_out_26;
      tmp_40_lpi_3_dfm_1 <= z_out_27;
      tmp_38_lpi_3_dfm_1 <= z_out_28;
      tmp_36_lpi_3_dfm_1 <= z_out_29;
      tmp_34_lpi_3_dfm_1 <= z_out_30;
      tmp_32_lpi_3_dfm_1 <= z_out_31;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_33_true_3_lshift_psp_1_0_sva <= 2'b00;
    end
    else if ( ~ (fsm_output[9]) ) begin
      operator_33_true_3_lshift_psp_1_0_sva <= operator_33_true_3_lshift_psp_1_0_sva_mx0w5;
    end
  end
  assign butterFly2_21_tw_butterFly2_21_tw_or_nl = c_1_sva | INNER_LOOP4_nor_tmp;
  assign c_mux_nl = MUX_s_1_2_2((operator_20_false_acc_cse_sva[0]), butterFly2_21_tw_butterFly2_21_tw_or_nl,
      fsm_output[9]);
  assign STAGE_LOOP_mux1h_nl = MUX1HOT_v_2_6_2((INNER_LOOP1_r_INNER_LOOP1_r_and_cse[6:5]),
      (INNER_LOOP2_r_11_4_sva_6_0_mx1[6:5]), (operator_20_false_acc_cse_sva[2:1]),
      (operator_33_true_2_lshift_psp_2_0_sva_mx0[1:0]), operator_33_true_3_lshift_psp_1_0_sva_mx0w5,
      operator_33_true_3_lshift_psp_1_0_sva, {or_tmp_3597 , or_dcpl_315 , (fsm_output[5])
      , or_tmp_3600 , (fsm_output[8]) , (fsm_output[9])});
  assign modulo_add_1_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_141, z_out_138, z_out_136,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_2_nl = ({modulo_add_1_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[32:0];
  assign modulo_add_1_qelse_and_nl = (~ z_out_143_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_1_qelse_or_1_nl = (z_out_143_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_143_32 & (fsm_output[7])) | (z_out_145_32 & (fsm_output[9]));
  assign modulo_add_1_qelse_and_4_nl = (~ z_out_143_32) & (fsm_output[7]);
  assign modulo_add_1_qelse_and_5_nl = (~ z_out_145_32) & (fsm_output[9]);
  assign modulo_add_10_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_132, z_out_127, z_out_128,
      z_out_142, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_3_nl = ({modulo_add_10_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[32:0];
  assign modulo_add_10_qelse_and_nl = (~ z_out_144_32) & (fsm_output[2]);
  assign modulo_add_10_qelse_or_nl = (z_out_144_32 & (fsm_output[2])) | (z_out_144_32
      & (fsm_output[4])) | (z_out_144_32 & (fsm_output[7])) | (z_out_146_32 & (fsm_output[9]));
  assign modulo_add_10_qelse_and_5_nl = (~ z_out_144_32) & (fsm_output[4]);
  assign modulo_add_10_qelse_and_6_nl = (~ z_out_144_32) & (fsm_output[7]);
  assign modulo_add_10_qelse_and_7_nl = (~ z_out_146_32) & (fsm_output[9]);
  assign modulo_add_11_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_131, z_out_137, z_out_127,
      z_out_141, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_4_nl = ({modulo_add_11_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[32:0];
  assign modulo_add_11_qelse_and_nl = (~ z_out_146_32) & (fsm_output[2]);
  assign modulo_add_11_qelse_or_nl = (z_out_146_32 & (fsm_output[2])) | (z_out_146_32
      & (fsm_output[4])) | (z_out_147_32 & (fsm_output[7])) | (z_out_147_32 & (fsm_output[9]));
  assign modulo_add_11_qelse_and_5_nl = (~ z_out_146_32) & (fsm_output[4]);
  assign modulo_add_11_qelse_and_6_nl = (~ z_out_147_32) & (fsm_output[7]);
  assign modulo_add_11_qelse_and_7_nl = (~ z_out_147_32) & (fsm_output[9]);
  assign modulo_add_12_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_130, z_out_142, z_out_140,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_5_nl = ({modulo_add_12_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[32:0];
  assign modulo_add_12_qelse_and_nl = (~ z_out_147_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_12_qelse_or_1_nl = (z_out_147_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_148_32 & (fsm_output[7])) | (z_out_150_32 & (fsm_output[9]));
  assign modulo_add_12_qelse_and_4_nl = (~ z_out_148_32) & (fsm_output[7]);
  assign modulo_add_12_qelse_and_5_nl = (~ z_out_150_32) & (fsm_output[9]);
  assign modulo_add_13_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_129, z_out_141, z_out_139,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_6_nl = ({modulo_add_13_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[32:0];
  assign modulo_add_13_qelse_and_nl = (~ z_out_150_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_13_qelse_or_1_nl = (z_out_150_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_150_32 & (fsm_output[7])) | (z_out_151_32 & (fsm_output[9]));
  assign modulo_add_13_qelse_and_4_nl = (~ z_out_150_32) & (fsm_output[7]);
  assign modulo_add_13_qelse_and_5_nl = (~ z_out_151_32) & (fsm_output[9]);
  assign modulo_add_14_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_128, z_out_140, z_out_138,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_10_nl = ({modulo_add_14_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[32:0];
  assign modulo_add_14_qelse_and_nl = (~ z_out_152_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_14_qelse_or_1_nl = (z_out_152_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_153_32 & (fsm_output[7])) | (z_out_154_32 & (fsm_output[9]));
  assign modulo_add_14_qelse_and_4_nl = (~ z_out_153_32) & (fsm_output[7]);
  assign modulo_add_14_qelse_and_5_nl = (~ z_out_154_32) & (fsm_output[9]);
  assign modulo_add_15_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_127, z_out_142, z_out_139,
      z_out_137, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_14_nl = ({modulo_add_15_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[32:0];
  assign modulo_add_15_qelse_and_nl = (~ z_out_153_32) & (fsm_output[2]);
  assign modulo_add_15_qelse_or_nl = (z_out_153_32 & (fsm_output[2])) | (z_out_153_32
      & (fsm_output[4])) | (z_out_154_32 & (fsm_output[7])) | (z_out_157_32 & (fsm_output[9]));
  assign modulo_add_15_qelse_and_5_nl = (~ z_out_153_32) & (fsm_output[4]);
  assign modulo_add_15_qelse_and_6_nl = (~ z_out_154_32) & (fsm_output[7]);
  assign modulo_add_15_qelse_and_7_nl = (~ z_out_157_32) & (fsm_output[9]);
  assign butterFly1_f1_butterFly1_f1_nor_nl = ~((INNER_LOOP1_r_11_4_sva_6_0[6:4]!=3'b000));
  assign butterFly1_16_f1_butterFly1_16_f1_nor_nl = ~((INNER_LOOP2_r_11_4_sva_6_0[6:4]!=3'b000));
  assign butterFly2_f1_butterFly2_f1_and_5_nl = (INNER_LOOP3_r_11_4_sva_6_0[6:4]==3'b110);
  assign butterFly2_16_f1_butterFly2_16_f1_and_5_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b110);
  assign butterFly1_f1_butterFly1_f1_and_nl = (INNER_LOOP1_r_11_4_sva_6_0[4]) & butterFly1_f1_nor_cse;
  assign butterFly1_16_f1_butterFly1_16_f1_and_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b001);
  assign butterFly1_f1_butterFly1_f1_and_1_nl = (INNER_LOOP1_r_11_4_sva_6_0[6:4]==3'b010);
  assign butterFly1_16_f1_butterFly1_16_f1_and_1_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b010);
  assign butterFly1_f1_butterFly1_f1_and_2_nl = (INNER_LOOP1_r_11_4_sva_6_0[6:4]==3'b011);
  assign butterFly1_16_f1_butterFly1_16_f1_and_2_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b011);
  assign butterFly2_f1_butterFly2_f1_and_nl = (INNER_LOOP3_r_11_4_sva_6_0[4]) & butterFly2_f1_nor_cse;
  assign butterFly2_16_f1_butterFly2_16_f1_and_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b001);
  assign butterFly1_f1_butterFly1_f1_and_3_nl = (INNER_LOOP1_r_11_4_sva_6_0[6:4]==3'b100);
  assign butterFly1_16_f1_butterFly1_16_f1_and_3_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b100);
  assign butterFly2_f1_butterFly2_f1_and_1_nl = (INNER_LOOP3_r_11_4_sva_6_0[6:4]==3'b010);
  assign butterFly2_16_f1_butterFly2_16_f1_and_1_nl = (INNER_LOOP4_r_11_4_sva_6_0[5])
      & butterFly2_16_f1_nor_1_cse;
  assign butterFly1_f1_butterFly1_f1_and_4_nl = (INNER_LOOP1_r_11_4_sva_6_0[6:4]==3'b101);
  assign butterFly1_16_f1_butterFly1_16_f1_and_4_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b101);
  assign butterFly2_f1_butterFly2_f1_and_2_nl = (INNER_LOOP3_r_11_4_sva_6_0[6:4]==3'b011);
  assign butterFly2_16_f1_butterFly2_16_f1_and_2_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b011);
  assign butterFly1_f1_butterFly1_f1_and_5_nl = (INNER_LOOP1_r_11_4_sva_6_0[6:4]==3'b110);
  assign butterFly1_16_f1_butterFly1_16_f1_and_5_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b110);
  assign butterFly2_f1_butterFly2_f1_and_3_nl = (INNER_LOOP3_r_11_4_sva_6_0[6:4]==3'b100);
  assign butterFly2_16_f1_butterFly2_16_f1_and_3_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b100);
  assign butterFly1_f1_butterFly1_f1_and_6_nl = (INNER_LOOP1_r_11_4_sva_6_0[6:4]==3'b111);
  assign butterFly1_16_f1_butterFly1_16_f1_and_6_nl = (INNER_LOOP2_r_11_4_sva_6_0[6:4]==3'b111);
  assign butterFly2_f1_butterFly2_f1_and_4_nl = (INNER_LOOP3_r_11_4_sva_6_0[6:4]==3'b101);
  assign butterFly2_16_f1_butterFly2_16_f1_and_4_nl = (INNER_LOOP4_r_11_4_sva_6_0[6:4]==3'b101);
  assign INNER_LOOP1_mux_nl = MUX_s_1_2_2(INNER_LOOP1_stage_0, INNER_LOOP1_stage_0_10,
      fsm_output[7]);
  assign INNER_LOOP1_mux_4_nl = MUX_s_1_2_2(INNER_LOOP1_stage_0_2, INNER_LOOP1_stage_0_11,
      fsm_output[7]);
  assign INNER_LOOP1_mux_5_nl = MUX_s_1_2_2(butterFly2_15_conc_2_itm_5_0, (operator_33_true_2_lshift_psp_2_0_sva_mx0[0]),
      or_tmp_3600);
  assign INNER_LOOP1_mux_6_nl = MUX_s_1_2_2(INNER_LOOP1_stage_0_10, (operator_33_true_2_lshift_psp_2_0_sva_mx0[2]),
      or_tmp_3600);
  assign butterFly1_15_mux_9_nl = MUX_s_1_2_2(butterFly1_15_conc_2_itm_1_0, INNER_LOOP1_stage_0,
      or_dcpl_298);
  assign butterFly1_15_mux1h_47_nl = MUX1HOT_s_1_3_2((INNER_LOOP1_r_INNER_LOOP1_r_and_cse[0]),
      (INNER_LOOP2_r_11_4_sva_6_0_mx1[0]), butterFly1_15_conc_2_itm_9_0, {or_tmp_3597
      , or_dcpl_315 , or_dcpl_298});
  assign butterFly2_15_mux1h_3_nl = MUX1HOT_s_1_4_2(INNER_LOOP1_stage_0_3, butterFly2_15_conc_2_itm_8_0,
      (INNER_LOOP1_r_INNER_LOOP1_r_and_3_cse[0]), (INNER_LOOP1_r_INNER_LOOP1_r_and_5_cse[0]),
      {(fsm_output[2]) , (fsm_output[4]) , or_tmp_3600 , or_tmp_3732});
  assign butterFly1_15_mux_10_nl = MUX_s_1_2_2(butterFly1_15_conc_2_itm_9_0, butterFly2_15_conc_2_itm_5_0,
      or_tmp_3842);
  assign modulo_add_2_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_140, z_out_137, z_out_135,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_18_nl = ({modulo_add_2_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[32:0];
  assign modulo_add_23_qelse_and_nl = (~ z_out_156_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_23_qelse_or_1_nl = (z_out_156_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_156_32 & (fsm_output[7])) | (z_out_158_32 & (fsm_output[9]));
  assign modulo_add_23_qelse_and_4_nl = (~ z_out_156_32) & (fsm_output[7]);
  assign modulo_add_23_qelse_and_5_nl = (~ z_out_158_32) & (fsm_output[9]);
  assign modulo_add_3_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_139, z_out_136, z_out_134,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_22_nl = ({modulo_add_3_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[32:0];
  assign modulo_add_24_qelse_and_nl = (~ z_out_158_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_24_qelse_or_1_nl = (z_out_158_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_157_32 & (fsm_output[7])) | (z_out_156_32 & (fsm_output[9]));
  assign modulo_add_24_qelse_and_4_nl = (~ z_out_157_32) & (fsm_output[7]);
  assign modulo_add_24_qelse_and_5_nl = (~ z_out_156_32) & (fsm_output[9]);
  assign modulo_add_4_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_138, z_out_135, z_out_133,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_26_nl = ({modulo_add_4_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_26_nl = nl_acc_26_nl[32:0];
  assign modulo_add_25_qelse_and_nl = (~ z_out_157_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_25_qelse_or_1_nl = (z_out_157_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_155_32 & (fsm_output[7])) | (z_out_152_32 & (fsm_output[9]));
  assign modulo_add_25_qelse_and_4_nl = (~ z_out_155_32) & (fsm_output[7]);
  assign modulo_add_25_qelse_and_5_nl = (~ z_out_152_32) & (fsm_output[9]);
  assign modulo_add_5_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_137, z_out_136, z_out_134,
      z_out_132, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_30_nl = ({modulo_add_5_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_30_nl = nl_acc_30_nl[32:0];
  assign modulo_add_26_qelse_and_nl = (~ z_out_151_32) & (fsm_output[2]);
  assign modulo_add_26_qelse_or_nl = (z_out_151_32 & (fsm_output[2])) | (z_out_151_32
      & (fsm_output[4])) | (z_out_151_32 & (fsm_output[7])) | (z_out_148_32 & (fsm_output[9]));
  assign modulo_add_26_qelse_and_5_nl = (~ z_out_151_32) & (fsm_output[4]);
  assign modulo_add_26_qelse_and_6_nl = (~ z_out_151_32) & (fsm_output[7]);
  assign modulo_add_26_qelse_and_7_nl = (~ z_out_148_32) & (fsm_output[9]);
  assign modulo_add_6_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_136, z_out_135, z_out_133,
      z_out_131, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_34_nl = ({modulo_add_6_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_34_nl = nl_acc_34_nl[32:0];
  assign modulo_add_27_qelse_and_nl = (~ z_out_149_32) & (fsm_output[2]);
  assign modulo_add_27_qelse_or_nl = (z_out_149_32 & (fsm_output[2])) | (z_out_149_32
      & (fsm_output[4])) | (z_out_145_32 & (fsm_output[7])) | (z_out_144_32 & (fsm_output[9]));
  assign modulo_add_27_qelse_and_5_nl = (~ z_out_149_32) & (fsm_output[4]);
  assign modulo_add_27_qelse_and_6_nl = (~ z_out_145_32) & (fsm_output[7]);
  assign modulo_add_27_qelse_and_7_nl = (~ z_out_144_32) & (fsm_output[9]);
  assign modulo_add_7_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_135, z_out_134, z_out_132,
      z_out_130, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_38_nl = ({modulo_add_7_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_38_nl = nl_acc_38_nl[32:0];
  assign modulo_add_28_qelse_and_nl = (~ z_out_145_32) & (fsm_output[2]);
  assign modulo_add_28_qelse_or_nl = (z_out_145_32 & (fsm_output[2])) | (z_out_145_32
      & (fsm_output[4])) | (z_out_149_32 & (fsm_output[7])) | (z_out_153_32 & (fsm_output[9]));
  assign modulo_add_28_qelse_and_5_nl = (~ z_out_145_32) & (fsm_output[4]);
  assign modulo_add_28_qelse_and_6_nl = (~ z_out_149_32) & (fsm_output[7]);
  assign modulo_add_28_qelse_and_7_nl = (~ z_out_153_32) & (fsm_output[9]);
  assign modulo_add_8_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_134, z_out_133, z_out_131,
      z_out_129, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_42_nl = ({modulo_add_8_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_42_nl = nl_acc_42_nl[32:0];
  assign modulo_add_29_qelse_and_nl = (~ z_out_155_32) & (fsm_output[2]);
  assign modulo_add_29_qelse_or_nl = (z_out_155_32 & (fsm_output[2])) | (z_out_155_32
      & (fsm_output[4])) | (z_out_158_32 & (fsm_output[7])) | (z_out_155_32 & (fsm_output[9]));
  assign modulo_add_29_qelse_and_5_nl = (~ z_out_155_32) & (fsm_output[4]);
  assign modulo_add_29_qelse_and_6_nl = (~ z_out_158_32) & (fsm_output[7]);
  assign modulo_add_29_qelse_and_7_nl = (~ z_out_155_32) & (fsm_output[9]);
  assign modulo_add_9_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_133, z_out_132, z_out_130,
      z_out_128, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_46_nl = ({modulo_add_9_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_46_nl = nl_acc_46_nl[32:0];
  assign modulo_add_30_qelse_and_nl = (~ z_out_154_32) & (fsm_output[2]);
  assign modulo_add_30_qelse_or_nl = (z_out_154_32 & (fsm_output[2])) | (z_out_154_32
      & (fsm_output[4])) | (z_out_152_32 & (fsm_output[7])) | (z_out_149_32 & (fsm_output[9]));
  assign modulo_add_30_qelse_and_5_nl = (~ z_out_154_32) & (fsm_output[4]);
  assign modulo_add_30_qelse_and_6_nl = (~ z_out_152_32) & (fsm_output[7]);
  assign modulo_add_30_qelse_and_7_nl = (~ z_out_149_32) & (fsm_output[9]);
  assign modulo_add_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_142, z_out_131, z_out_129,
      z_out_127, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_49_nl = ({modulo_add_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_49_nl = nl_acc_49_nl[32:0];
  assign modulo_add_31_qelse_and_nl = (~ z_out_148_32) & (fsm_output[2]);
  assign modulo_add_31_qelse_or_nl = (z_out_148_32 & (fsm_output[2])) | (z_out_148_32
      & (fsm_output[4])) | (z_out_146_32 & (fsm_output[7])) | (z_out_143_32 & (fsm_output[9]));
  assign modulo_add_31_qelse_and_5_nl = (~ z_out_148_32) & (fsm_output[4]);
  assign modulo_add_31_qelse_and_6_nl = (~ z_out_146_32) & (fsm_output[7]);
  assign modulo_add_31_qelse_and_7_nl = (~ z_out_143_32) & (fsm_output[9]);
  assign modulo_sub_16_qelse_or_nl = ((z_out_126[31]) & (~ (fsm_output[9]))) | ((z_out_111[31])
      & (fsm_output[9]));
  assign modulo_sub_17_qelse_or_nl = ((z_out_116[31]) & (~ (fsm_output[9]))) | ((z_out_112[31])
      & (fsm_output[9]));
  assign modulo_sub_18_qelse_or_nl = ((z_out_123[31]) & (~ (fsm_output[9]))) | ((z_out_113[31])
      & (fsm_output[9]));
  assign modulo_sub_19_qelse_or_nl = ((z_out_124[31]) & (~ (fsm_output[9]))) | ((z_out_114[31])
      & (fsm_output[9]));
  assign modulo_sub_20_qelse_or_nl = ((z_out_125[31]) & (~ (fsm_output[9]))) | ((z_out_115[31])
      & (fsm_output[9]));
  assign modulo_sub_21_qelse_or_nl = ((z_out_111[31]) & (~ (fsm_output[9]))) | ((z_out_116[31])
      & (fsm_output[9]));
  assign modulo_sub_22_qelse_or_nl = ((z_out_112[31]) & (~ (fsm_output[9]))) | ((z_out_117[31])
      & (fsm_output[9]));
  assign modulo_sub_23_qelse_or_nl = ((z_out_113[31]) & (~ (fsm_output[9]))) | ((z_out_118[31])
      & (fsm_output[9]));
  assign modulo_sub_24_qelse_or_nl = ((z_out_114[31]) & (~ (fsm_output[9]))) | ((z_out_119[31])
      & (fsm_output[9]));
  assign modulo_sub_25_qelse_or_nl = ((z_out_115[31]) & (~ (fsm_output[9]))) | ((z_out_120[31])
      & (fsm_output[9]));
  assign modulo_sub_26_qelse_or_nl = ((z_out_117[31]) & (~ (fsm_output[9]))) | ((z_out_121[31])
      & (fsm_output[9]));
  assign modulo_sub_27_qelse_or_nl = ((z_out_118[31]) & (~ (fsm_output[9]))) | ((z_out_122[31])
      & (fsm_output[9]));
  assign modulo_sub_28_qelse_or_nl = ((z_out_119[31]) & (~ (fsm_output[9]))) | ((z_out_123[31])
      & (fsm_output[9]));
  assign modulo_sub_29_qelse_or_nl = ((z_out_120[31]) & (~ (fsm_output[9]))) | ((z_out_124[31])
      & (fsm_output[9]));
  assign modulo_sub_30_qelse_or_nl = ((z_out_121[31]) & (~ (fsm_output[9]))) | ((z_out_125[31])
      & (fsm_output[9]));
  assign modulo_sub_31_qelse_or_nl = ((z_out_122[31]) & (~ (fsm_output[9]))) | ((z_out_126[31])
      & (fsm_output[9]));
  assign INNER_LOOP1_mux_7_nl = MUX_s_1_2_2(INNER_LOOP1_stage_0, INNER_LOOP2_stage_0_10,
      or_dcpl_298);
  assign butterFly2_f1_butterFly2_f1_nor_nl = ~((INNER_LOOP3_r_11_4_sva_6_0[6:4]!=3'b000));
  assign butterFly2_16_f1_butterFly2_16_f1_nor_nl = ~((INNER_LOOP4_r_11_4_sva_6_0[6:4]!=3'b000));
  assign butterFly2_f1_butterFly2_f1_and_6_nl = (INNER_LOOP3_r_11_4_sva_6_0[6:4]==3'b111);
  assign STAGE_LOOP_base_STAGE_LOOP_base_mux_nl = MUX_v_7_2_2((z_out_60[10:4]), (z_out_62[6:0]),
      fsm_output[4]);
  assign INNER_LOOP2_r_or_nl = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[2]);
  assign operator_20_false_mux_2_nl = MUX_v_3_2_2(({butterFly1_15_conc_2_itm_2_1
      , c_1_sva}), operator_20_false_acc_cse_sva, fsm_output[5]);
  assign nl_z_out_61 = operator_20_false_mux_2_nl + ({1'b1 , (~ (fsm_output[5]))
      , 1'b1});
  assign z_out_61 = nl_z_out_61[2:0];
  assign operator_20_false_mux1h_2_nl = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      INNER_LOOP2_r_11_4_sva_6_0, INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_62 = conv_u2u_7_8(operator_20_false_mux1h_2_nl) + 8'b00000001;
  assign z_out_62 = nl_z_out_62[7:0];
  assign modulo_sub_15_qif_mux_2_nl = MUX_v_31_2_2((z_out_126[30:0]), (z_out_124[30:0]),
      fsm_output[7]);
  assign nl_z_out_68 = ({1'b1 , modulo_sub_15_qif_mux_2_nl}) + p_sva;
  assign z_out_68 = nl_z_out_68[31:0];
  assign modulo_sub_31_qif_mux_2_nl = MUX_v_31_2_2((z_out_122[30:0]), (z_out_126[30:0]),
      fsm_output[9]);
  assign nl_z_out_69 = ({1'b1 , modulo_sub_31_qif_mux_2_nl}) + p_sva;
  assign z_out_69 = nl_z_out_69[31:0];
  assign modulo_sub_7_qif_mux_2_nl = MUX_v_31_2_2((z_out_118[30:0]), (z_out_123[30:0]),
      fsm_output[7]);
  assign nl_z_out_70 = ({1'b1 , modulo_sub_7_qif_mux_2_nl}) + p_sva;
  assign z_out_70 = nl_z_out_70[31:0];
  assign modulo_sub_30_qif_mux_2_nl = MUX_v_31_2_2((z_out_121[30:0]), (z_out_125[30:0]),
      fsm_output[9]);
  assign nl_z_out_72 = ({1'b1 , modulo_sub_30_qif_mux_2_nl}) + p_sva;
  assign z_out_72 = nl_z_out_72[31:0];
  assign modulo_sub_39_qif_mux_2_nl = MUX_v_31_2_2((z_out_116[30:0]), (z_out_125[30:0]),
      fsm_output[2]);
  assign nl_z_out_73 = ({1'b1 , modulo_sub_39_qif_mux_2_nl}) + p_sva;
  assign z_out_73 = nl_z_out_73[31:0];
  assign modulo_sub_29_qif_mux_2_nl = MUX_v_31_2_2((z_out_120[30:0]), (z_out_124[30:0]),
      fsm_output[9]);
  assign nl_z_out_74 = ({1'b1 , modulo_sub_29_qif_mux_2_nl}) + p_sva;
  assign z_out_74 = nl_z_out_74[31:0];
  assign modulo_sub_6_qif_mux_2_nl = MUX_v_31_2_2((z_out_117[30:0]), (z_out_122[30:0]),
      fsm_output[7]);
  assign nl_z_out_76 = ({1'b1 , modulo_sub_6_qif_mux_2_nl}) + p_sva;
  assign z_out_76 = nl_z_out_76[31:0];
  assign modulo_sub_28_qif_mux_2_nl = MUX_v_31_2_2((z_out_119[30:0]), (z_out_123[30:0]),
      fsm_output[9]);
  assign nl_z_out_77 = ({1'b1 , modulo_sub_28_qif_mux_2_nl}) + p_sva;
  assign z_out_77 = nl_z_out_77[31:0];
  assign modulo_sub_38_qif_mux_2_nl = MUX_v_31_2_2((z_out_115[30:0]), (z_out_124[30:0]),
      fsm_output[2]);
  assign nl_z_out_78 = ({1'b1 , modulo_sub_38_qif_mux_2_nl}) + p_sva;
  assign z_out_78 = nl_z_out_78[31:0];
  assign modulo_sub_27_qif_mux_2_nl = MUX_v_31_2_2((z_out_118[30:0]), (z_out_122[30:0]),
      fsm_output[9]);
  assign nl_z_out_80 = ({1'b1 , modulo_sub_27_qif_mux_2_nl}) + p_sva;
  assign z_out_80 = nl_z_out_80[31:0];
  assign modulo_sub_5_qif_mux_2_nl = MUX_v_31_2_2((z_out_116[30:0]), (z_out_121[30:0]),
      fsm_output[7]);
  assign nl_z_out_81 = ({1'b1 , modulo_sub_5_qif_mux_2_nl}) + p_sva;
  assign z_out_81 = nl_z_out_81[31:0];
  assign modulo_sub_26_qif_mux_2_nl = MUX_v_31_2_2((z_out_117[30:0]), (z_out_121[30:0]),
      fsm_output[9]);
  assign nl_z_out_82 = ({1'b1 , modulo_sub_26_qif_mux_2_nl}) + p_sva;
  assign z_out_82 = nl_z_out_82[31:0];
  assign modulo_sub_37_qif_mux_2_nl = MUX_v_31_2_2((z_out_114[30:0]), (z_out_123[30:0]),
      fsm_output[2]);
  assign nl_z_out_84 = ({1'b1 , modulo_sub_37_qif_mux_2_nl}) + p_sva;
  assign z_out_84 = nl_z_out_84[31:0];
  assign modulo_sub_25_qif_mux_2_nl = MUX_v_31_2_2((z_out_115[30:0]), (z_out_120[30:0]),
      fsm_output[9]);
  assign nl_z_out_85 = ({1'b1 , modulo_sub_25_qif_mux_2_nl}) + p_sva;
  assign z_out_85 = nl_z_out_85[31:0];
  assign modulo_sub_4_qif_mux_2_nl = MUX_v_31_2_2((z_out_115[30:0]), (z_out_120[30:0]),
      fsm_output[7]);
  assign nl_z_out_86 = ({1'b1 , modulo_sub_4_qif_mux_2_nl}) + p_sva;
  assign z_out_86 = nl_z_out_86[31:0];
  assign modulo_sub_24_qif_mux_2_nl = MUX_v_31_2_2((z_out_114[30:0]), (z_out_119[30:0]),
      fsm_output[9]);
  assign nl_z_out_88 = ({1'b1 , modulo_sub_24_qif_mux_2_nl}) + p_sva;
  assign z_out_88 = nl_z_out_88[31:0];
  assign modulo_sub_36_qif_mux_2_nl = MUX_v_31_2_2((z_out_113[30:0]), (z_out_122[30:0]),
      fsm_output[2]);
  assign nl_z_out_89 = ({1'b1 , modulo_sub_36_qif_mux_2_nl}) + p_sva;
  assign z_out_89 = nl_z_out_89[31:0];
  assign modulo_sub_23_qif_mux_2_nl = MUX_v_31_2_2((z_out_113[30:0]), (z_out_118[30:0]),
      fsm_output[9]);
  assign nl_z_out_90 = ({1'b1 , modulo_sub_23_qif_mux_2_nl}) + p_sva;
  assign z_out_90 = nl_z_out_90[31:0];
  assign modulo_sub_3_qif_mux_2_nl = MUX_v_31_2_2((z_out_114[30:0]), (z_out_119[30:0]),
      fsm_output[7]);
  assign nl_z_out_92 = ({1'b1 , modulo_sub_3_qif_mux_2_nl}) + p_sva;
  assign z_out_92 = nl_z_out_92[31:0];
  assign modulo_sub_22_qif_mux_2_nl = MUX_v_31_2_2((z_out_112[30:0]), (z_out_117[30:0]),
      fsm_output[9]);
  assign nl_z_out_93 = ({1'b1 , modulo_sub_22_qif_mux_2_nl}) + p_sva;
  assign z_out_93 = nl_z_out_93[31:0];
  assign modulo_sub_35_qif_mux_2_nl = MUX_v_31_2_2((z_out_112[30:0]), (z_out_121[30:0]),
      fsm_output[2]);
  assign nl_z_out_94 = ({1'b1 , modulo_sub_35_qif_mux_2_nl}) + p_sva;
  assign z_out_94 = nl_z_out_94[31:0];
  assign modulo_sub_21_qif_mux_2_nl = MUX_v_31_2_2((z_out_111[30:0]), (z_out_116[30:0]),
      fsm_output[9]);
  assign nl_z_out_96 = ({1'b1 , modulo_sub_21_qif_mux_2_nl}) + p_sva;
  assign z_out_96 = nl_z_out_96[31:0];
  assign modulo_sub_2_qif_mux_2_nl = MUX_v_31_2_2((z_out_113[30:0]), (z_out_118[30:0]),
      fsm_output[7]);
  assign nl_z_out_97 = ({1'b1 , modulo_sub_2_qif_mux_2_nl}) + p_sva;
  assign z_out_97 = nl_z_out_97[31:0];
  assign modulo_sub_20_qif_mux_2_nl = MUX_v_31_2_2((z_out_125[30:0]), (z_out_115[30:0]),
      fsm_output[9]);
  assign nl_z_out_98 = ({1'b1 , modulo_sub_20_qif_mux_2_nl}) + p_sva;
  assign z_out_98 = nl_z_out_98[31:0];
  assign modulo_sub_34_qif_mux_2_nl = MUX_v_31_2_2((z_out_111[30:0]), (z_out_120[30:0]),
      fsm_output[2]);
  assign nl_z_out_100 = ({1'b1 , modulo_sub_34_qif_mux_2_nl}) + p_sva;
  assign z_out_100 = nl_z_out_100[31:0];
  assign modulo_sub_19_qif_mux_2_nl = MUX_v_31_2_2((z_out_124[30:0]), (z_out_114[30:0]),
      fsm_output[9]);
  assign nl_z_out_101 = ({1'b1 , modulo_sub_19_qif_mux_2_nl}) + p_sva;
  assign z_out_101 = nl_z_out_101[31:0];
  assign modulo_sub_1_qif_mux_2_nl = MUX_v_31_2_2((z_out_112[30:0]), (z_out_117[30:0]),
      fsm_output[7]);
  assign nl_z_out_102 = ({1'b1 , modulo_sub_1_qif_mux_2_nl}) + p_sva;
  assign z_out_102 = nl_z_out_102[31:0];
  assign modulo_sub_18_qif_mux_2_nl = MUX_v_31_2_2((z_out_123[30:0]), (z_out_113[30:0]),
      fsm_output[9]);
  assign nl_z_out_104 = ({1'b1 , modulo_sub_18_qif_mux_2_nl}) + p_sva;
  assign z_out_104 = nl_z_out_104[31:0];
  assign modulo_sub_33_qif_mux_2_nl = MUX_v_31_2_2((z_out_126[30:0]), (z_out_119[30:0]),
      fsm_output[2]);
  assign nl_z_out_105 = ({1'b1 , modulo_sub_33_qif_mux_2_nl}) + p_sva;
  assign z_out_105 = nl_z_out_105[31:0];
  assign modulo_sub_17_qif_mux_2_nl = MUX_v_31_2_2((z_out_116[30:0]), (z_out_112[30:0]),
      fsm_output[9]);
  assign nl_z_out_106 = ({1'b1 , modulo_sub_17_qif_mux_2_nl}) + p_sva;
  assign z_out_106 = nl_z_out_106[31:0];
  assign modulo_sub_qif_mux_2_nl = MUX_v_31_2_2((z_out_111[30:0]), (z_out_125[30:0]),
      fsm_output[7]);
  assign nl_z_out_108 = ({1'b1 , modulo_sub_qif_mux_2_nl}) + p_sva;
  assign z_out_108 = nl_z_out_108[31:0];
  assign modulo_sub_16_qif_mux_2_nl = MUX_v_31_2_2((z_out_126[30:0]), (z_out_111[30:0]),
      fsm_output[9]);
  assign nl_z_out_109 = ({1'b1 , modulo_sub_16_qif_mux_2_nl}) + p_sva;
  assign z_out_109 = nl_z_out_109[31:0];
  assign butterFly1_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_res_lpi_3_dfm_1_cse),
      (~ reg_mult_5_res_lpi_3_dfm_1_cse), (~ reg_mult_34_res_lpi_3_dfm_1_cse), (~
      reg_mult_47_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_50_nl = ({tmp_10_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_mux1h_18_nl
      , 1'b1});
  assign acc_50_nl = nl_acc_50_nl[32:0];
  assign z_out_111 = readslicef_33_32_1(acc_50_nl);
  assign butterFly1_1_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_1_res_lpi_3_dfm_1_cse),
      (~ reg_mult_6_res_lpi_3_dfm_1_cse), (~ reg_mult_35_res_lpi_3_dfm_1_cse), (~
      reg_mult_46_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_51_nl = ({tmp_102_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_1_mux1h_18_nl
      , 1'b1});
  assign acc_51_nl = nl_acc_51_nl[32:0];
  assign z_out_112 = readslicef_33_32_1(acc_51_nl);
  assign butterFly1_2_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_2_res_lpi_3_dfm_1_cse),
      (~ reg_mult_7_res_lpi_3_dfm_1_cse), (~ reg_mult_36_res_lpi_3_dfm_1_cse), (~
      reg_mult_45_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_52_nl = ({tmp_104_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_2_mux1h_18_nl
      , 1'b1});
  assign acc_52_nl = nl_acc_52_nl[32:0];
  assign z_out_113 = readslicef_33_32_1(acc_52_nl);
  assign butterFly1_3_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_3_res_lpi_3_dfm_1_cse),
      (~ reg_mult_8_res_lpi_3_dfm_1_cse), (~ reg_mult_37_res_lpi_3_dfm_1_cse), (~
      reg_mult_44_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_53_nl = ({tmp_106_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_3_mux1h_18_nl
      , 1'b1});
  assign acc_53_nl = nl_acc_53_nl[32:0];
  assign z_out_114 = readslicef_33_32_1(acc_53_nl);
  assign butterFly1_4_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_4_res_lpi_3_dfm_1_cse),
      (~ reg_mult_9_res_lpi_3_dfm_1_cse), (~ reg_mult_38_res_lpi_3_dfm_1_cse), (~
      reg_mult_43_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_54_nl = ({tmp_108_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_4_mux1h_18_nl
      , 1'b1});
  assign acc_54_nl = nl_acc_54_nl[32:0];
  assign z_out_115 = readslicef_33_32_1(acc_54_nl);
  assign butterFly1_5_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_5_res_lpi_3_dfm_1_cse),
      (~ reg_mult_1_res_lpi_3_dfm_1_cse), (~ reg_mult_39_res_lpi_3_dfm_1_cse), (~
      reg_mult_42_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_55_nl = ({tmp_110_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_5_mux1h_18_nl
      , 1'b1});
  assign acc_55_nl = nl_acc_55_nl[32:0];
  assign z_out_116 = readslicef_33_32_1(acc_55_nl);
  assign butterFly1_6_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_6_res_lpi_3_dfm_1_cse),
      (~ reg_mult_10_res_lpi_3_dfm_1_cse), (~ reg_mult_40_res_lpi_3_dfm_1_cse), (~
      reg_mult_41_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_56_nl = ({tmp_112_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_6_mux1h_18_nl
      , 1'b1});
  assign acc_56_nl = nl_acc_56_nl[32:0];
  assign z_out_117 = readslicef_33_32_1(acc_56_nl);
  assign butterFly1_7_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_7_res_lpi_3_dfm_1_cse),
      (~ reg_mult_11_res_lpi_3_dfm_1_cse), (~ reg_mult_41_res_lpi_3_dfm_1_cse), (~
      reg_mult_40_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_57_nl = ({tmp_114_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_7_mux1h_18_nl
      , 1'b1});
  assign acc_57_nl = nl_acc_57_nl[32:0];
  assign z_out_118 = readslicef_33_32_1(acc_57_nl);
  assign butterFly1_8_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_8_res_lpi_3_dfm_1_cse),
      (~ reg_mult_12_res_lpi_3_dfm_1_cse), (~ reg_mult_42_res_lpi_3_dfm_1_cse), (~
      reg_mult_39_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_58_nl = ({tmp_116_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_8_mux1h_18_nl
      , 1'b1});
  assign acc_58_nl = nl_acc_58_nl[32:0];
  assign z_out_119 = readslicef_33_32_1(acc_58_nl);
  assign butterFly1_9_mux1h_274_nl = MUX1HOT_v_32_4_2((~ reg_mult_9_res_lpi_3_dfm_1_cse),
      (~ reg_mult_13_res_lpi_3_dfm_1_cse), (~ reg_mult_43_res_lpi_3_dfm_1_cse), (~
      reg_mult_38_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_59_nl = ({tmp_118_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_9_mux1h_274_nl
      , 1'b1});
  assign acc_59_nl = nl_acc_59_nl[32:0];
  assign z_out_120 = readslicef_33_32_1(acc_59_nl);
  assign butterFly1_10_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_10_res_lpi_3_dfm_1_cse),
      (~ reg_mult_14_res_lpi_3_dfm_1_cse), (~ reg_mult_44_res_lpi_3_dfm_1_cse), (~
      reg_mult_37_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_60_nl = ({tmp_120_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_10_mux1h_18_nl
      , 1'b1});
  assign acc_60_nl = nl_acc_60_nl[32:0];
  assign z_out_121 = readslicef_33_32_1(acc_60_nl);
  assign butterFly1_11_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_11_res_lpi_3_dfm_1_cse),
      (~ reg_mult_15_res_lpi_3_dfm_1_cse), (~ reg_mult_45_res_lpi_3_dfm_1_cse), (~
      reg_mult_36_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_61_nl = ({tmp_122_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_11_mux1h_18_nl
      , 1'b1});
  assign acc_61_nl = nl_acc_61_nl[32:0];
  assign z_out_122 = readslicef_33_32_1(acc_61_nl);
  assign butterFly1_12_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_12_res_lpi_3_dfm_1_cse),
      (~ reg_mult_2_res_lpi_3_dfm_1_cse), (~ reg_mult_46_res_lpi_3_dfm_1_cse), (~
      reg_mult_35_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_62_nl = ({tmp_124_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_12_mux1h_18_nl
      , 1'b1});
  assign acc_62_nl = nl_acc_62_nl[32:0];
  assign z_out_123 = readslicef_33_32_1(acc_62_nl);
  assign butterFly1_13_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_13_res_lpi_3_dfm_1_cse),
      (~ reg_mult_3_res_lpi_3_dfm_1_cse), (~ reg_mult_47_res_lpi_3_dfm_1_cse), (~
      reg_mult_34_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_63_nl = ({tmp_126_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_13_mux1h_18_nl
      , 1'b1});
  assign acc_63_nl = nl_acc_63_nl[32:0];
  assign z_out_124 = readslicef_33_32_1(acc_63_nl);
  assign butterFly1_14_mux1h_18_nl = MUX1HOT_v_32_4_2((~ reg_mult_14_res_lpi_3_dfm_1_cse),
      (~ reg_mult_4_res_lpi_3_dfm_1_cse), (~ reg_mult_32_res_lpi_3_dfm_1_cse), (~
      reg_mult_33_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_64_nl = ({tmp_60_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_14_mux1h_18_nl
      , 1'b1});
  assign acc_64_nl = nl_acc_64_nl[32:0];
  assign z_out_125 = readslicef_33_32_1(acc_64_nl);
  assign butterFly1_15_mux1h_79_nl = MUX1HOT_v_32_4_2((~ reg_mult_15_res_lpi_3_dfm_1_cse),
      (~ reg_mult_res_lpi_3_dfm_1_cse), (~ reg_mult_33_res_lpi_3_dfm_1_cse), (~ reg_mult_32_res_lpi_3_dfm_1_cse),
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_65_nl = ({tmp_62_lpi_3_dfm_7 , 1'b1}) + ({butterFly1_15_mux1h_79_nl
      , 1'b1});
  assign acc_65_nl = nl_acc_65_nl[32:0];
  assign z_out_126 = readslicef_33_32_1(acc_65_nl);
  assign butterFly1_15_mux1h_80_nl = MUX1HOT_v_32_4_2(reg_mult_15_res_lpi_3_dfm_1_cse,
      reg_mult_res_lpi_3_dfm_1_cse, reg_mult_33_res_lpi_3_dfm_1_cse, reg_mult_32_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_127 = tmp_62_lpi_3_dfm_7 + butterFly1_15_mux1h_80_nl;
  assign z_out_127 = nl_z_out_127[31:0];
  assign butterFly1_14_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_14_res_lpi_3_dfm_1_cse,
      reg_mult_4_res_lpi_3_dfm_1_cse, reg_mult_32_res_lpi_3_dfm_1_cse, reg_mult_33_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_128 = tmp_60_lpi_3_dfm_7 + butterFly1_14_mux1h_19_nl;
  assign z_out_128 = nl_z_out_128[31:0];
  assign butterFly1_13_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_13_res_lpi_3_dfm_1_cse,
      reg_mult_3_res_lpi_3_dfm_1_cse, reg_mult_47_res_lpi_3_dfm_1_cse, reg_mult_34_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_129 = tmp_126_lpi_3_dfm_7 + butterFly1_13_mux1h_19_nl;
  assign z_out_129 = nl_z_out_129[31:0];
  assign butterFly1_12_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_12_res_lpi_3_dfm_1_cse,
      reg_mult_2_res_lpi_3_dfm_1_cse, reg_mult_46_res_lpi_3_dfm_1_cse, reg_mult_35_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_130 = tmp_124_lpi_3_dfm_7 + butterFly1_12_mux1h_19_nl;
  assign z_out_130 = nl_z_out_130[31:0];
  assign butterFly1_11_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_11_res_lpi_3_dfm_1_cse,
      reg_mult_15_res_lpi_3_dfm_1_cse, reg_mult_45_res_lpi_3_dfm_1_cse, reg_mult_36_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_131 = tmp_122_lpi_3_dfm_7 + butterFly1_11_mux1h_19_nl;
  assign z_out_131 = nl_z_out_131[31:0];
  assign butterFly1_10_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_10_res_lpi_3_dfm_1_cse,
      reg_mult_14_res_lpi_3_dfm_1_cse, reg_mult_44_res_lpi_3_dfm_1_cse, reg_mult_37_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_132 = tmp_120_lpi_3_dfm_7 + butterFly1_10_mux1h_19_nl;
  assign z_out_132 = nl_z_out_132[31:0];
  assign butterFly1_9_mux1h_275_nl = MUX1HOT_v_32_4_2(reg_mult_9_res_lpi_3_dfm_1_cse,
      reg_mult_13_res_lpi_3_dfm_1_cse, reg_mult_43_res_lpi_3_dfm_1_cse, reg_mult_38_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_133 = tmp_118_lpi_3_dfm_7 + butterFly1_9_mux1h_275_nl;
  assign z_out_133 = nl_z_out_133[31:0];
  assign butterFly1_8_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_8_res_lpi_3_dfm_1_cse,
      reg_mult_12_res_lpi_3_dfm_1_cse, reg_mult_42_res_lpi_3_dfm_1_cse, reg_mult_39_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_134 = tmp_116_lpi_3_dfm_7 + butterFly1_8_mux1h_19_nl;
  assign z_out_134 = nl_z_out_134[31:0];
  assign butterFly1_7_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_7_res_lpi_3_dfm_1_cse,
      reg_mult_11_res_lpi_3_dfm_1_cse, reg_mult_41_res_lpi_3_dfm_1_cse, reg_mult_40_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_135 = tmp_114_lpi_3_dfm_7 + butterFly1_7_mux1h_19_nl;
  assign z_out_135 = nl_z_out_135[31:0];
  assign butterFly1_6_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_6_res_lpi_3_dfm_1_cse,
      reg_mult_10_res_lpi_3_dfm_1_cse, reg_mult_40_res_lpi_3_dfm_1_cse, reg_mult_41_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_136 = tmp_112_lpi_3_dfm_7 + butterFly1_6_mux1h_19_nl;
  assign z_out_136 = nl_z_out_136[31:0];
  assign butterFly1_5_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_5_res_lpi_3_dfm_1_cse,
      reg_mult_1_res_lpi_3_dfm_1_cse, reg_mult_39_res_lpi_3_dfm_1_cse, reg_mult_42_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_137 = tmp_110_lpi_3_dfm_7 + butterFly1_5_mux1h_19_nl;
  assign z_out_137 = nl_z_out_137[31:0];
  assign butterFly1_4_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_4_res_lpi_3_dfm_1_cse,
      reg_mult_9_res_lpi_3_dfm_1_cse, reg_mult_38_res_lpi_3_dfm_1_cse, reg_mult_43_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_138 = tmp_108_lpi_3_dfm_7 + butterFly1_4_mux1h_19_nl;
  assign z_out_138 = nl_z_out_138[31:0];
  assign butterFly1_3_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_3_res_lpi_3_dfm_1_cse,
      reg_mult_8_res_lpi_3_dfm_1_cse, reg_mult_37_res_lpi_3_dfm_1_cse, reg_mult_44_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_139 = tmp_106_lpi_3_dfm_7 + butterFly1_3_mux1h_19_nl;
  assign z_out_139 = nl_z_out_139[31:0];
  assign butterFly1_2_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_2_res_lpi_3_dfm_1_cse,
      reg_mult_7_res_lpi_3_dfm_1_cse, reg_mult_36_res_lpi_3_dfm_1_cse, reg_mult_45_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_140 = tmp_104_lpi_3_dfm_7 + butterFly1_2_mux1h_19_nl;
  assign z_out_140 = nl_z_out_140[31:0];
  assign butterFly1_1_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_1_res_lpi_3_dfm_1_cse,
      reg_mult_6_res_lpi_3_dfm_1_cse, reg_mult_35_res_lpi_3_dfm_1_cse, reg_mult_46_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_141 = tmp_102_lpi_3_dfm_7 + butterFly1_1_mux1h_19_nl;
  assign z_out_141 = nl_z_out_141[31:0];
  assign butterFly1_mux1h_19_nl = MUX1HOT_v_32_4_2(reg_mult_res_lpi_3_dfm_1_cse,
      reg_mult_5_res_lpi_3_dfm_1_cse, reg_mult_34_res_lpi_3_dfm_1_cse, reg_mult_47_res_lpi_3_dfm_1_cse,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_142 = tmp_10_lpi_3_dfm_7 + butterFly1_mux1h_19_nl;
  assign z_out_142 = nl_z_out_142[31:0];
  assign modulo_add_1_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_141), (~ z_out_138),
      (~ z_out_127), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_82_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_1_mux1h_3_nl
      , 1'b1});
  assign acc_82_nl = nl_acc_82_nl[33:0];
  assign z_out_143_32 = readslicef_34_1_33(acc_82_nl);
  assign modulo_add_10_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_132), (~ z_out_127),
      (~ z_out_128), (~ z_out_131), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_83_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_10_mux1h_3_nl
      , 1'b1});
  assign acc_83_nl = nl_acc_83_nl[33:0];
  assign z_out_144_32 = readslicef_34_1_33(acc_83_nl);
  assign modulo_add_54_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_136), (~ z_out_133),
      (~ z_out_135), (~ z_out_134), {(fsm_output[9]) , (fsm_output[7]) , (fsm_output[2])
      , (fsm_output[4])});
  assign nl_acc_84_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_54_mux1h_3_nl
      , 1'b1});
  assign acc_84_nl = nl_acc_84_nl[33:0];
  assign z_out_145_32 = readslicef_34_1_33(acc_84_nl);
  assign modulo_add_48_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_142), (~ z_out_131),
      (~ z_out_137), (~ z_out_129), {(fsm_output[9]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7])});
  assign nl_acc_85_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_48_mux1h_3_nl
      , 1'b1});
  assign acc_85_nl = nl_acc_85_nl[33:0];
  assign z_out_146_32 = readslicef_34_1_33(acc_85_nl);
  assign modulo_add_33_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_127), (~ z_out_141),
      (~ z_out_130), {(fsm_output[7]) , (fsm_output[9]) , modulo_add_1_qelse_or_m1c});
  assign nl_acc_86_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_33_mux1h_3_nl
      , 1'b1});
  assign acc_86_nl = nl_acc_86_nl[33:0];
  assign z_out_147_32 = readslicef_34_1_33(acc_86_nl);
  assign modulo_add_34_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_142), (~ z_out_132),
      (~ z_out_131), {or_dcpl_353 , (fsm_output[9]) , (fsm_output[4])});
  assign nl_acc_87_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_34_mux1h_3_nl
      , 1'b1});
  assign acc_87_nl = nl_acc_87_nl[33:0];
  assign z_out_148_32 = readslicef_34_1_33(acc_87_nl);
  assign modulo_add_6_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_136), (~ z_out_135),
      (~ z_out_132), (~ z_out_128), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_88_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_6_mux1h_3_nl
      , 1'b1});
  assign acc_88_nl = nl_acc_88_nl[33:0];
  assign z_out_149_32 = readslicef_34_1_33(acc_88_nl);
  assign modulo_add_50_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_140), (~ z_out_129),
      (~ z_out_141), {(fsm_output[9]) , modulo_add_1_qelse_or_m1c , (fsm_output[7])});
  assign nl_acc_89_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_50_mux1h_3_nl
      , 1'b1});
  assign acc_89_nl = nl_acc_89_nl[33:0];
  assign z_out_150_32 = readslicef_34_1_33(acc_89_nl);
  assign modulo_add_51_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_139), (~ z_out_137),
      (~ z_out_136), (~ z_out_134), {(fsm_output[9]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7])});
  assign nl_acc_90_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_51_mux1h_3_nl
      , 1'b1});
  assign acc_90_nl = nl_acc_90_nl[33:0];
  assign z_out_151_32 = readslicef_34_1_33(acc_90_nl);
  assign modulo_add_14_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_128), (~ z_out_133),
      (~ z_out_130), {modulo_add_1_qelse_or_m1c , (fsm_output[9]) , (fsm_output[7])});
  assign nl_acc_91_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_14_mux1h_3_nl
      , 1'b1});
  assign acc_91_nl = nl_acc_91_nl[33:0];
  assign z_out_152_32 = readslicef_34_1_33(acc_91_nl);
  assign modulo_add_36_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_140), (~ z_out_127),
      (~ z_out_142), (~ z_out_130), {(fsm_output[7]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[9])});
  assign nl_acc_92_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_36_mux1h_3_nl
      , 1'b1});
  assign acc_92_nl = nl_acc_92_nl[33:0];
  assign z_out_153_32 = readslicef_34_1_33(acc_92_nl);
  assign modulo_add_52_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_138), (~ z_out_139),
      (~ z_out_133), (~ z_out_132), {(fsm_output[9]) , (fsm_output[7]) , (fsm_output[2])
      , (fsm_output[4])});
  assign nl_acc_93_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_52_mux1h_3_nl
      , 1'b1});
  assign acc_93_nl = nl_acc_93_nl[33:0];
  assign z_out_154_32 = readslicef_34_1_33(acc_93_nl);
  assign modulo_add_41_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_135), (~ z_out_134),
      (~ z_out_133), (~ z_out_129), {(fsm_output[7]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[9])});
  assign nl_acc_94_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_41_mux1h_3_nl
      , 1'b1});
  assign acc_94_nl = nl_acc_94_nl[33:0];
  assign z_out_155_32 = readslicef_34_1_33(acc_94_nl);
  assign modulo_add_2_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_140), (~ z_out_137),
      (~ z_out_134), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_95_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_2_mux1h_3_nl
      , 1'b1});
  assign acc_95_nl = nl_acc_95_nl[33:0];
  assign z_out_156_32 = readslicef_34_1_33(acc_95_nl);
  assign modulo_add_53_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_137), (~ z_out_136),
      (~ z_out_138), {(fsm_output[9]) , (fsm_output[7]) , modulo_add_1_qelse_or_m1c});
  assign nl_acc_96_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_53_mux1h_3_nl
      , 1'b1});
  assign acc_96_nl = nl_acc_96_nl[33:0];
  assign z_out_157_32 = readslicef_34_1_33(acc_96_nl);
  assign modulo_add_55_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_135), (~ z_out_139),
      (~ z_out_131), {(fsm_output[9]) , modulo_add_1_qelse_or_m1c , (fsm_output[7])});
  assign nl_acc_97_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_55_mux1h_3_nl
      , 1'b1});
  assign acc_97_nl = nl_acc_97_nl[33:0];
  assign z_out_158_32 = readslicef_34_1_33(acc_97_nl);
  assign z_out = MUX1HOT_v_32_8_2(xt_rsc_0_30_i_qa_d, xt_rsc_1_30_i_qa_d, xt_rsc_2_30_i_qa_d,
      xt_rsc_3_30_i_qa_d, xt_rsc_4_30_i_qa_d, xt_rsc_5_30_i_qa_d, xt_rsc_6_30_i_qa_d,
      xt_rsc_7_30_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_1 = MUX1HOT_v_32_8_2(xt_rsc_0_28_i_qa_d, xt_rsc_1_28_i_qa_d, xt_rsc_2_28_i_qa_d,
      xt_rsc_3_28_i_qa_d, xt_rsc_4_28_i_qa_d, xt_rsc_5_28_i_qa_d, xt_rsc_6_28_i_qa_d,
      xt_rsc_7_28_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_2 = MUX1HOT_v_32_8_2(xt_rsc_0_26_i_qa_d, xt_rsc_1_26_i_qa_d, xt_rsc_2_26_i_qa_d,
      xt_rsc_3_26_i_qa_d, xt_rsc_4_26_i_qa_d, xt_rsc_5_26_i_qa_d, xt_rsc_6_26_i_qa_d,
      xt_rsc_7_26_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_3 = MUX1HOT_v_32_8_2(xt_rsc_0_24_i_qa_d, xt_rsc_1_24_i_qa_d, xt_rsc_2_24_i_qa_d,
      xt_rsc_3_24_i_qa_d, xt_rsc_4_24_i_qa_d, xt_rsc_5_24_i_qa_d, xt_rsc_6_24_i_qa_d,
      xt_rsc_7_24_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_4 = MUX1HOT_v_32_8_2(xt_rsc_0_22_i_qa_d, xt_rsc_1_22_i_qa_d, xt_rsc_2_22_i_qa_d,
      xt_rsc_3_22_i_qa_d, xt_rsc_4_22_i_qa_d, xt_rsc_5_22_i_qa_d, xt_rsc_6_22_i_qa_d,
      xt_rsc_7_22_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_5 = MUX1HOT_v_32_8_2(xt_rsc_0_20_i_qa_d, xt_rsc_1_20_i_qa_d, xt_rsc_2_20_i_qa_d,
      xt_rsc_3_20_i_qa_d, xt_rsc_4_20_i_qa_d, xt_rsc_5_20_i_qa_d, xt_rsc_6_20_i_qa_d,
      xt_rsc_7_20_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_6 = MUX1HOT_v_32_8_2(xt_rsc_0_18_i_qa_d, xt_rsc_1_18_i_qa_d, xt_rsc_2_18_i_qa_d,
      xt_rsc_3_18_i_qa_d, xt_rsc_4_18_i_qa_d, xt_rsc_5_18_i_qa_d, xt_rsc_6_18_i_qa_d,
      xt_rsc_7_18_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_7 = MUX1HOT_v_32_8_2(xt_rsc_0_16_i_qa_d, xt_rsc_1_16_i_qa_d, xt_rsc_2_16_i_qa_d,
      xt_rsc_3_16_i_qa_d, xt_rsc_4_16_i_qa_d, xt_rsc_5_16_i_qa_d, xt_rsc_6_16_i_qa_d,
      xt_rsc_7_16_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_8 = MUX1HOT_v_32_8_2(xt_rsc_0_14_i_qa_d, xt_rsc_1_14_i_qa_d, xt_rsc_2_14_i_qa_d,
      xt_rsc_3_14_i_qa_d, xt_rsc_4_14_i_qa_d, xt_rsc_5_14_i_qa_d, xt_rsc_6_14_i_qa_d,
      xt_rsc_7_14_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_9 = MUX1HOT_v_32_8_2(xt_rsc_0_12_i_qa_d, xt_rsc_1_12_i_qa_d, xt_rsc_2_12_i_qa_d,
      xt_rsc_3_12_i_qa_d, xt_rsc_4_12_i_qa_d, xt_rsc_5_12_i_qa_d, xt_rsc_6_12_i_qa_d,
      xt_rsc_7_12_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_10 = MUX1HOT_v_32_8_2(xt_rsc_0_10_i_qa_d, xt_rsc_1_10_i_qa_d, xt_rsc_2_10_i_qa_d,
      xt_rsc_3_10_i_qa_d, xt_rsc_4_10_i_qa_d, xt_rsc_5_10_i_qa_d, xt_rsc_6_10_i_qa_d,
      xt_rsc_7_10_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_11 = MUX1HOT_v_32_8_2(xt_rsc_0_8_i_qa_d, xt_rsc_1_8_i_qa_d, xt_rsc_2_8_i_qa_d,
      xt_rsc_3_8_i_qa_d, xt_rsc_4_8_i_qa_d, xt_rsc_5_8_i_qa_d, xt_rsc_6_8_i_qa_d,
      xt_rsc_7_8_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse ,
      butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_12 = MUX1HOT_v_32_8_2(xt_rsc_0_6_i_qa_d, xt_rsc_1_6_i_qa_d, xt_rsc_2_6_i_qa_d,
      xt_rsc_3_6_i_qa_d, xt_rsc_4_6_i_qa_d, xt_rsc_5_6_i_qa_d, xt_rsc_6_6_i_qa_d,
      xt_rsc_7_6_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse ,
      butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_13 = MUX1HOT_v_32_8_2(xt_rsc_0_4_i_qa_d, xt_rsc_1_4_i_qa_d, xt_rsc_2_4_i_qa_d,
      xt_rsc_3_4_i_qa_d, xt_rsc_4_4_i_qa_d, xt_rsc_5_4_i_qa_d, xt_rsc_6_4_i_qa_d,
      xt_rsc_7_4_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse ,
      butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_14 = MUX1HOT_v_32_8_2(xt_rsc_0_2_i_qa_d, xt_rsc_1_2_i_qa_d, xt_rsc_2_2_i_qa_d,
      xt_rsc_3_2_i_qa_d, xt_rsc_4_2_i_qa_d, xt_rsc_5_2_i_qa_d, xt_rsc_6_2_i_qa_d,
      xt_rsc_7_2_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse ,
      butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_15 = MUX1HOT_v_32_8_2(xt_rsc_0_0_i_qa_d, xt_rsc_1_0_i_qa_d, xt_rsc_2_0_i_qa_d,
      xt_rsc_3_0_i_qa_d, xt_rsc_4_0_i_qa_d, xt_rsc_5_0_i_qa_d, xt_rsc_6_0_i_qa_d,
      xt_rsc_7_0_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse ,
      butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_16 = MUX1HOT_v_32_8_2(yt_rsc_0_30_i_q_d, yt_rsc_1_30_i_q_d, yt_rsc_2_30_i_q_d,
      yt_rsc_3_30_i_q_d, yt_rsc_4_30_i_q_d, yt_rsc_5_30_i_q_d, yt_rsc_6_30_i_q_d,
      yt_rsc_7_30_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_17 = MUX1HOT_v_32_8_2(yt_rsc_0_28_i_q_d, yt_rsc_1_28_i_q_d, yt_rsc_2_28_i_q_d,
      yt_rsc_3_28_i_q_d, yt_rsc_4_28_i_q_d, yt_rsc_5_28_i_q_d, yt_rsc_6_28_i_q_d,
      yt_rsc_7_28_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_18 = MUX1HOT_v_32_8_2(yt_rsc_0_26_i_q_d, yt_rsc_1_26_i_q_d, yt_rsc_2_26_i_q_d,
      yt_rsc_3_26_i_q_d, yt_rsc_4_26_i_q_d, yt_rsc_5_26_i_q_d, yt_rsc_6_26_i_q_d,
      yt_rsc_7_26_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_19 = MUX1HOT_v_32_8_2(yt_rsc_0_24_i_q_d, yt_rsc_1_24_i_q_d, yt_rsc_2_24_i_q_d,
      yt_rsc_3_24_i_q_d, yt_rsc_4_24_i_q_d, yt_rsc_5_24_i_q_d, yt_rsc_6_24_i_q_d,
      yt_rsc_7_24_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_20 = MUX1HOT_v_32_8_2(yt_rsc_0_22_i_q_d, yt_rsc_1_22_i_q_d, yt_rsc_2_22_i_q_d,
      yt_rsc_3_22_i_q_d, yt_rsc_4_22_i_q_d, yt_rsc_5_22_i_q_d, yt_rsc_6_22_i_q_d,
      yt_rsc_7_22_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_21 = MUX1HOT_v_32_8_2(yt_rsc_0_20_i_q_d, yt_rsc_1_20_i_q_d, yt_rsc_2_20_i_q_d,
      yt_rsc_3_20_i_q_d, yt_rsc_4_20_i_q_d, yt_rsc_5_20_i_q_d, yt_rsc_6_20_i_q_d,
      yt_rsc_7_20_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_22 = MUX1HOT_v_32_8_2(yt_rsc_0_18_i_q_d, yt_rsc_1_18_i_q_d, yt_rsc_2_18_i_q_d,
      yt_rsc_3_18_i_q_d, yt_rsc_4_18_i_q_d, yt_rsc_5_18_i_q_d, yt_rsc_6_18_i_q_d,
      yt_rsc_7_18_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_23 = MUX1HOT_v_32_8_2(yt_rsc_0_16_i_q_d, yt_rsc_1_16_i_q_d, yt_rsc_2_16_i_q_d,
      yt_rsc_3_16_i_q_d, yt_rsc_4_16_i_q_d, yt_rsc_5_16_i_q_d, yt_rsc_6_16_i_q_d,
      yt_rsc_7_16_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_24 = MUX1HOT_v_32_8_2(yt_rsc_0_14_i_q_d, yt_rsc_1_14_i_q_d, yt_rsc_2_14_i_q_d,
      yt_rsc_3_14_i_q_d, yt_rsc_4_14_i_q_d, yt_rsc_5_14_i_q_d, yt_rsc_6_14_i_q_d,
      yt_rsc_7_14_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_25 = MUX1HOT_v_32_8_2(yt_rsc_0_12_i_q_d, yt_rsc_1_12_i_q_d, yt_rsc_2_12_i_q_d,
      yt_rsc_3_12_i_q_d, yt_rsc_4_12_i_q_d, yt_rsc_5_12_i_q_d, yt_rsc_6_12_i_q_d,
      yt_rsc_7_12_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_26 = MUX1HOT_v_32_8_2(yt_rsc_0_10_i_q_d, yt_rsc_1_10_i_q_d, yt_rsc_2_10_i_q_d,
      yt_rsc_3_10_i_q_d, yt_rsc_4_10_i_q_d, yt_rsc_5_10_i_q_d, yt_rsc_6_10_i_q_d,
      yt_rsc_7_10_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_27 = MUX1HOT_v_32_8_2(yt_rsc_0_8_i_q_d, yt_rsc_1_8_i_q_d, yt_rsc_2_8_i_q_d,
      yt_rsc_3_8_i_q_d, yt_rsc_4_8_i_q_d, yt_rsc_5_8_i_q_d, yt_rsc_6_8_i_q_d, yt_rsc_7_8_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_28 = MUX1HOT_v_32_8_2(yt_rsc_0_6_i_q_d, yt_rsc_1_6_i_q_d, yt_rsc_2_6_i_q_d,
      yt_rsc_3_6_i_q_d, yt_rsc_4_6_i_q_d, yt_rsc_5_6_i_q_d, yt_rsc_6_6_i_q_d, yt_rsc_7_6_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_29 = MUX1HOT_v_32_8_2(yt_rsc_0_4_i_q_d, yt_rsc_1_4_i_q_d, yt_rsc_2_4_i_q_d,
      yt_rsc_3_4_i_q_d, yt_rsc_4_4_i_q_d, yt_rsc_5_4_i_q_d, yt_rsc_6_4_i_q_d, yt_rsc_7_4_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_30 = MUX1HOT_v_32_8_2(yt_rsc_0_2_i_q_d, yt_rsc_1_2_i_q_d, yt_rsc_2_2_i_q_d,
      yt_rsc_3_2_i_q_d, yt_rsc_4_2_i_q_d, yt_rsc_5_2_i_q_d, yt_rsc_6_2_i_q_d, yt_rsc_7_2_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_31 = MUX1HOT_v_32_8_2(yt_rsc_0_0_i_q_d, yt_rsc_1_0_i_q_d, yt_rsc_2_0_i_q_d,
      yt_rsc_3_0_i_q_d, yt_rsc_4_0_i_q_d, yt_rsc_5_0_i_q_d, yt_rsc_6_0_i_q_d, yt_rsc_7_0_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_32 = MUX1HOT_v_32_8_2(yt_rsc_0_3_i_q_d, yt_rsc_1_3_i_q_d, yt_rsc_2_3_i_q_d,
      yt_rsc_3_3_i_q_d, yt_rsc_4_3_i_q_d, yt_rsc_5_3_i_q_d, yt_rsc_6_3_i_q_d, yt_rsc_7_3_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_33 = MUX1HOT_v_32_8_2(yt_rsc_0_5_i_q_d, yt_rsc_1_5_i_q_d, yt_rsc_2_5_i_q_d,
      yt_rsc_3_5_i_q_d, yt_rsc_4_5_i_q_d, yt_rsc_5_5_i_q_d, yt_rsc_6_5_i_q_d, yt_rsc_7_5_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_34 = MUX1HOT_v_32_8_2(yt_rsc_0_7_i_q_d, yt_rsc_1_7_i_q_d, yt_rsc_2_7_i_q_d,
      yt_rsc_3_7_i_q_d, yt_rsc_4_7_i_q_d, yt_rsc_5_7_i_q_d, yt_rsc_6_7_i_q_d, yt_rsc_7_7_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_35 = MUX1HOT_v_32_8_2(yt_rsc_0_31_i_q_d, yt_rsc_1_31_i_q_d, yt_rsc_2_31_i_q_d,
      yt_rsc_3_31_i_q_d, yt_rsc_4_31_i_q_d, yt_rsc_5_31_i_q_d, yt_rsc_6_31_i_q_d,
      yt_rsc_7_31_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_36 = MUX1HOT_v_32_8_2(xt_rsc_0_11_i_qa_d, xt_rsc_1_11_i_qa_d, xt_rsc_2_11_i_qa_d,
      xt_rsc_3_11_i_qa_d, xt_rsc_4_11_i_qa_d, xt_rsc_5_11_i_qa_d, xt_rsc_6_11_i_qa_d,
      xt_rsc_7_11_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_37 = MUX1HOT_v_32_8_2(xt_rsc_0_19_i_qa_d, xt_rsc_1_19_i_qa_d, xt_rsc_2_19_i_qa_d,
      xt_rsc_3_19_i_qa_d, xt_rsc_4_19_i_qa_d, xt_rsc_5_19_i_qa_d, xt_rsc_6_19_i_qa_d,
      xt_rsc_7_19_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_38 = MUX1HOT_v_32_8_2(xt_rsc_0_21_i_qa_d, xt_rsc_1_21_i_qa_d, xt_rsc_2_21_i_qa_d,
      xt_rsc_3_21_i_qa_d, xt_rsc_4_21_i_qa_d, xt_rsc_5_21_i_qa_d, xt_rsc_6_21_i_qa_d,
      xt_rsc_7_21_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_39 = MUX1HOT_v_32_8_2(xt_rsc_0_23_i_qa_d, xt_rsc_1_23_i_qa_d, xt_rsc_2_23_i_qa_d,
      xt_rsc_3_23_i_qa_d, xt_rsc_4_23_i_qa_d, xt_rsc_5_23_i_qa_d, xt_rsc_6_23_i_qa_d,
      xt_rsc_7_23_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_40 = MUX1HOT_v_32_8_2(xt_rsc_0_25_i_qa_d, xt_rsc_1_25_i_qa_d, xt_rsc_2_25_i_qa_d,
      xt_rsc_3_25_i_qa_d, xt_rsc_4_25_i_qa_d, xt_rsc_5_25_i_qa_d, xt_rsc_6_25_i_qa_d,
      xt_rsc_7_25_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_41 = MUX1HOT_v_32_8_2(xt_rsc_0_27_i_qa_d, xt_rsc_1_27_i_qa_d, xt_rsc_2_27_i_qa_d,
      xt_rsc_3_27_i_qa_d, xt_rsc_4_27_i_qa_d, xt_rsc_5_27_i_qa_d, xt_rsc_6_27_i_qa_d,
      xt_rsc_7_27_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_42 = MUX1HOT_v_32_8_2(xt_rsc_0_29_i_qa_d, xt_rsc_1_29_i_qa_d, xt_rsc_2_29_i_qa_d,
      xt_rsc_3_29_i_qa_d, xt_rsc_4_29_i_qa_d, xt_rsc_5_29_i_qa_d, xt_rsc_6_29_i_qa_d,
      xt_rsc_7_29_i_qa_d, {butterFly1_15_f1_mux_cse , butterFly1_15_f1_mux_1_cse
      , butterFly1_15_f1_mux_2_cse , butterFly1_15_f1_mux_3_cse , butterFly1_15_f1_mux_4_cse
      , butterFly1_15_f1_mux_5_cse , butterFly1_15_f1_mux_6_cse , butterFly1_15_f1_mux_7_cse});
  assign z_out_43 = MUX1HOT_v_32_8_2(xt_rsc_0_1_i_qa_d, xt_rsc_1_1_i_qa_d, xt_rsc_2_1_i_qa_d,
      xt_rsc_3_1_i_qa_d, xt_rsc_4_1_i_qa_d, xt_rsc_5_1_i_qa_d, xt_rsc_6_1_i_qa_d,
      xt_rsc_7_1_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_44 = MUX1HOT_v_32_8_2(xt_rsc_0_3_i_qa_d, xt_rsc_1_3_i_qa_d, xt_rsc_2_3_i_qa_d,
      xt_rsc_3_3_i_qa_d, xt_rsc_4_3_i_qa_d, xt_rsc_5_3_i_qa_d, xt_rsc_6_3_i_qa_d,
      xt_rsc_7_3_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_45 = MUX1HOT_v_32_8_2(xt_rsc_0_5_i_qa_d, xt_rsc_1_5_i_qa_d, xt_rsc_2_5_i_qa_d,
      xt_rsc_3_5_i_qa_d, xt_rsc_4_5_i_qa_d, xt_rsc_5_5_i_qa_d, xt_rsc_6_5_i_qa_d,
      xt_rsc_7_5_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_46 = MUX1HOT_v_32_8_2(xt_rsc_0_13_i_qa_d, xt_rsc_1_13_i_qa_d, xt_rsc_2_13_i_qa_d,
      xt_rsc_3_13_i_qa_d, xt_rsc_4_13_i_qa_d, xt_rsc_5_13_i_qa_d, xt_rsc_6_13_i_qa_d,
      xt_rsc_7_13_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_47 = MUX1HOT_v_32_8_2(xt_rsc_0_15_i_qa_d, xt_rsc_1_15_i_qa_d, xt_rsc_2_15_i_qa_d,
      xt_rsc_3_15_i_qa_d, xt_rsc_4_15_i_qa_d, xt_rsc_5_15_i_qa_d, xt_rsc_6_15_i_qa_d,
      xt_rsc_7_15_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_48 = MUX1HOT_v_32_8_2(xt_rsc_0_17_i_qa_d, xt_rsc_1_17_i_qa_d, xt_rsc_2_17_i_qa_d,
      xt_rsc_3_17_i_qa_d, xt_rsc_4_17_i_qa_d, xt_rsc_5_17_i_qa_d, xt_rsc_6_17_i_qa_d,
      xt_rsc_7_17_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_49 = MUX1HOT_v_32_8_2(xt_rsc_0_31_i_qa_d, xt_rsc_1_31_i_qa_d, xt_rsc_2_31_i_qa_d,
      xt_rsc_3_31_i_qa_d, xt_rsc_4_31_i_qa_d, xt_rsc_5_31_i_qa_d, xt_rsc_6_31_i_qa_d,
      xt_rsc_7_31_i_qa_d, {butterFly2_f1_mux_cse , butterFly2_f1_mux_1_cse , butterFly2_f1_mux_2_cse
      , butterFly2_f1_mux_3_cse , butterFly2_f1_mux_4_cse , butterFly2_f1_mux_5_cse
      , butterFly2_f1_mux_6_cse , butterFly2_f1_mux_7_cse});
  assign z_out_50 = MUX1HOT_v_32_8_2(yt_rsc_0_29_i_q_d, yt_rsc_1_29_i_q_d, yt_rsc_2_29_i_q_d,
      yt_rsc_3_29_i_q_d, yt_rsc_4_29_i_q_d, yt_rsc_5_29_i_q_d, yt_rsc_6_29_i_q_d,
      yt_rsc_7_29_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_51 = MUX1HOT_v_32_8_2(yt_rsc_0_27_i_q_d, yt_rsc_1_27_i_q_d, yt_rsc_2_27_i_q_d,
      yt_rsc_3_27_i_q_d, yt_rsc_4_27_i_q_d, yt_rsc_5_27_i_q_d, yt_rsc_6_27_i_q_d,
      yt_rsc_7_27_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_52 = MUX1HOT_v_32_8_2(yt_rsc_0_25_i_q_d, yt_rsc_1_25_i_q_d, yt_rsc_2_25_i_q_d,
      yt_rsc_3_25_i_q_d, yt_rsc_4_25_i_q_d, yt_rsc_5_25_i_q_d, yt_rsc_6_25_i_q_d,
      yt_rsc_7_25_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_53 = MUX1HOT_v_32_8_2(yt_rsc_0_21_i_q_d, yt_rsc_1_21_i_q_d, yt_rsc_2_21_i_q_d,
      yt_rsc_3_21_i_q_d, yt_rsc_4_21_i_q_d, yt_rsc_5_21_i_q_d, yt_rsc_6_21_i_q_d,
      yt_rsc_7_21_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_54 = MUX1HOT_v_32_8_2(yt_rsc_0_11_i_q_d, yt_rsc_1_11_i_q_d, yt_rsc_2_11_i_q_d,
      yt_rsc_3_11_i_q_d, yt_rsc_4_11_i_q_d, yt_rsc_5_11_i_q_d, yt_rsc_6_11_i_q_d,
      yt_rsc_7_11_i_q_d, {butterFly2_21_f1_mux_cse , butterFly2_21_f1_mux_1_cse ,
      butterFly2_21_f1_mux_2_cse , butterFly2_21_f1_mux_3_cse , butterFly2_21_f1_mux_4_cse
      , butterFly2_21_f1_mux_5_cse , butterFly2_21_f1_mux_6_cse , butterFly2_21_f1_mux_7_cse});
  assign z_out_55 = MUX1HOT_v_32_8_2(yt_rsc_0_19_i_q_d, yt_rsc_1_19_i_q_d, yt_rsc_2_19_i_q_d,
      yt_rsc_3_19_i_q_d, yt_rsc_4_19_i_q_d, yt_rsc_5_19_i_q_d, yt_rsc_6_19_i_q_d,
      yt_rsc_7_19_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_56 = MUX1HOT_v_32_8_2(yt_rsc_0_13_i_q_d, yt_rsc_1_13_i_q_d, yt_rsc_2_13_i_q_d,
      yt_rsc_3_13_i_q_d, yt_rsc_4_13_i_q_d, yt_rsc_5_13_i_q_d, yt_rsc_6_13_i_q_d,
      yt_rsc_7_13_i_q_d, {butterFly2_21_f1_mux_cse , butterFly2_21_f1_mux_1_cse ,
      butterFly2_21_f1_mux_2_cse , butterFly2_21_f1_mux_3_cse , butterFly2_21_f1_mux_4_cse
      , butterFly2_21_f1_mux_5_cse , butterFly2_21_f1_mux_6_cse , butterFly2_21_f1_mux_7_cse});
  assign z_out_57 = MUX1HOT_v_32_8_2(yt_rsc_0_17_i_q_d, yt_rsc_1_17_i_q_d, yt_rsc_2_17_i_q_d,
      yt_rsc_3_17_i_q_d, yt_rsc_4_17_i_q_d, yt_rsc_5_17_i_q_d, yt_rsc_6_17_i_q_d,
      yt_rsc_7_17_i_q_d, {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse ,
      butterFly1_31_f1_mux_2_cse , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse
      , butterFly1_31_f1_mux_5_cse , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});
  assign z_out_58 = MUX1HOT_v_32_8_2(yt_rsc_0_15_i_q_d, yt_rsc_1_15_i_q_d, yt_rsc_2_15_i_q_d,
      yt_rsc_3_15_i_q_d, yt_rsc_4_15_i_q_d, yt_rsc_5_15_i_q_d, yt_rsc_6_15_i_q_d,
      yt_rsc_7_15_i_q_d, {butterFly2_21_f1_mux_cse , butterFly2_21_f1_mux_1_cse ,
      butterFly2_21_f1_mux_2_cse , butterFly2_21_f1_mux_3_cse , butterFly2_21_f1_mux_4_cse
      , butterFly2_21_f1_mux_5_cse , butterFly2_21_f1_mux_6_cse , butterFly2_21_f1_mux_7_cse});
  assign z_out_59 = MUX1HOT_v_32_8_2(yt_rsc_0_1_i_q_d, yt_rsc_1_1_i_q_d, yt_rsc_2_1_i_q_d,
      yt_rsc_3_1_i_q_d, yt_rsc_4_1_i_q_d, yt_rsc_5_1_i_q_d, yt_rsc_6_1_i_q_d, yt_rsc_7_1_i_q_d,
      {butterFly1_31_f1_mux_cse , butterFly1_31_f1_mux_1_cse , butterFly1_31_f1_mux_2_cse
      , butterFly1_31_f1_mux_3_cse , butterFly1_31_f1_mux_4_cse , butterFly1_31_f1_mux_5_cse
      , butterFly1_31_f1_mux_6_cse , butterFly1_31_f1_mux_7_cse});

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    result = result | ( input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_3_2;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [2:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | ( input_1 & {31{sel[1]}});
    result = result | ( input_2 & {31{sel[2]}});
    MUX1HOT_v_31_3_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_4_2;
    input [30:0] input_3;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [3:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | ( input_1 & {31{sel[1]}});
    result = result | ( input_2 & {31{sel[2]}});
    result = result | ( input_3 & {31{sel[3]}});
    MUX1HOT_v_31_4_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_12_2;
    input [31:0] input_11;
    input [31:0] input_10;
    input [31:0] input_9;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [11:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    result = result | ( input_9 & {32{sel[9]}});
    result = result | ( input_10 & {32{sel[10]}});
    result = result | ( input_11 & {32{sel[11]}});
    MUX1HOT_v_32_12_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_32_2;
    input [31:0] input_31;
    input [31:0] input_30;
    input [31:0] input_29;
    input [31:0] input_28;
    input [31:0] input_27;
    input [31:0] input_26;
    input [31:0] input_25;
    input [31:0] input_24;
    input [31:0] input_23;
    input [31:0] input_22;
    input [31:0] input_21;
    input [31:0] input_20;
    input [31:0] input_19;
    input [31:0] input_18;
    input [31:0] input_17;
    input [31:0] input_16;
    input [31:0] input_15;
    input [31:0] input_14;
    input [31:0] input_13;
    input [31:0] input_12;
    input [31:0] input_11;
    input [31:0] input_10;
    input [31:0] input_9;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [31:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    result = result | ( input_9 & {32{sel[9]}});
    result = result | ( input_10 & {32{sel[10]}});
    result = result | ( input_11 & {32{sel[11]}});
    result = result | ( input_12 & {32{sel[12]}});
    result = result | ( input_13 & {32{sel[13]}});
    result = result | ( input_14 & {32{sel[14]}});
    result = result | ( input_15 & {32{sel[15]}});
    result = result | ( input_16 & {32{sel[16]}});
    result = result | ( input_17 & {32{sel[17]}});
    result = result | ( input_18 & {32{sel[18]}});
    result = result | ( input_19 & {32{sel[19]}});
    result = result | ( input_20 & {32{sel[20]}});
    result = result | ( input_21 & {32{sel[21]}});
    result = result | ( input_22 & {32{sel[22]}});
    result = result | ( input_23 & {32{sel[23]}});
    result = result | ( input_24 & {32{sel[24]}});
    result = result | ( input_25 & {32{sel[25]}});
    result = result | ( input_26 & {32{sel[26]}});
    result = result | ( input_27 & {32{sel[27]}});
    result = result | ( input_28 & {32{sel[28]}});
    result = result | ( input_29 & {32{sel[29]}});
    result = result | ( input_30 & {32{sel[30]}});
    result = result | ( input_31 & {32{sel[31]}});
    MUX1HOT_v_32_32_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_5_2;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [4:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    MUX1HOT_v_32_5_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_6_2;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [5:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    MUX1HOT_v_32_6_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_8_2;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [7:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    MUX1HOT_v_32_8_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_9_2;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [8:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    MUX1HOT_v_32_9_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_4_2;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [3:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    MUX1HOT_v_3_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT
// ------------------------------------------------------------------


module peaseNTT (
  clk, rst, xt_rsc_0_0_adra, xt_rsc_0_0_da, xt_rsc_0_0_wea, xt_rsc_0_0_qa, xt_rsc_triosy_0_0_lz,
      xt_rsc_0_1_adra, xt_rsc_0_1_da, xt_rsc_0_1_wea, xt_rsc_0_1_qa, xt_rsc_triosy_0_1_lz,
      xt_rsc_0_2_adra, xt_rsc_0_2_da, xt_rsc_0_2_wea, xt_rsc_0_2_qa, xt_rsc_triosy_0_2_lz,
      xt_rsc_0_3_adra, xt_rsc_0_3_da, xt_rsc_0_3_wea, xt_rsc_0_3_qa, xt_rsc_triosy_0_3_lz,
      xt_rsc_0_4_adra, xt_rsc_0_4_da, xt_rsc_0_4_wea, xt_rsc_0_4_qa, xt_rsc_triosy_0_4_lz,
      xt_rsc_0_5_adra, xt_rsc_0_5_da, xt_rsc_0_5_wea, xt_rsc_0_5_qa, xt_rsc_triosy_0_5_lz,
      xt_rsc_0_6_adra, xt_rsc_0_6_da, xt_rsc_0_6_wea, xt_rsc_0_6_qa, xt_rsc_triosy_0_6_lz,
      xt_rsc_0_7_adra, xt_rsc_0_7_da, xt_rsc_0_7_wea, xt_rsc_0_7_qa, xt_rsc_triosy_0_7_lz,
      xt_rsc_0_8_adra, xt_rsc_0_8_da, xt_rsc_0_8_wea, xt_rsc_0_8_qa, xt_rsc_triosy_0_8_lz,
      xt_rsc_0_9_adra, xt_rsc_0_9_da, xt_rsc_0_9_wea, xt_rsc_0_9_qa, xt_rsc_triosy_0_9_lz,
      xt_rsc_0_10_adra, xt_rsc_0_10_da, xt_rsc_0_10_wea, xt_rsc_0_10_qa, xt_rsc_triosy_0_10_lz,
      xt_rsc_0_11_adra, xt_rsc_0_11_da, xt_rsc_0_11_wea, xt_rsc_0_11_qa, xt_rsc_triosy_0_11_lz,
      xt_rsc_0_12_adra, xt_rsc_0_12_da, xt_rsc_0_12_wea, xt_rsc_0_12_qa, xt_rsc_triosy_0_12_lz,
      xt_rsc_0_13_adra, xt_rsc_0_13_da, xt_rsc_0_13_wea, xt_rsc_0_13_qa, xt_rsc_triosy_0_13_lz,
      xt_rsc_0_14_adra, xt_rsc_0_14_da, xt_rsc_0_14_wea, xt_rsc_0_14_qa, xt_rsc_triosy_0_14_lz,
      xt_rsc_0_15_adra, xt_rsc_0_15_da, xt_rsc_0_15_wea, xt_rsc_0_15_qa, xt_rsc_triosy_0_15_lz,
      xt_rsc_0_16_adra, xt_rsc_0_16_da, xt_rsc_0_16_wea, xt_rsc_0_16_qa, xt_rsc_triosy_0_16_lz,
      xt_rsc_0_17_adra, xt_rsc_0_17_da, xt_rsc_0_17_wea, xt_rsc_0_17_qa, xt_rsc_triosy_0_17_lz,
      xt_rsc_0_18_adra, xt_rsc_0_18_da, xt_rsc_0_18_wea, xt_rsc_0_18_qa, xt_rsc_triosy_0_18_lz,
      xt_rsc_0_19_adra, xt_rsc_0_19_da, xt_rsc_0_19_wea, xt_rsc_0_19_qa, xt_rsc_triosy_0_19_lz,
      xt_rsc_0_20_adra, xt_rsc_0_20_da, xt_rsc_0_20_wea, xt_rsc_0_20_qa, xt_rsc_triosy_0_20_lz,
      xt_rsc_0_21_adra, xt_rsc_0_21_da, xt_rsc_0_21_wea, xt_rsc_0_21_qa, xt_rsc_triosy_0_21_lz,
      xt_rsc_0_22_adra, xt_rsc_0_22_da, xt_rsc_0_22_wea, xt_rsc_0_22_qa, xt_rsc_triosy_0_22_lz,
      xt_rsc_0_23_adra, xt_rsc_0_23_da, xt_rsc_0_23_wea, xt_rsc_0_23_qa, xt_rsc_triosy_0_23_lz,
      xt_rsc_0_24_adra, xt_rsc_0_24_da, xt_rsc_0_24_wea, xt_rsc_0_24_qa, xt_rsc_triosy_0_24_lz,
      xt_rsc_0_25_adra, xt_rsc_0_25_da, xt_rsc_0_25_wea, xt_rsc_0_25_qa, xt_rsc_triosy_0_25_lz,
      xt_rsc_0_26_adra, xt_rsc_0_26_da, xt_rsc_0_26_wea, xt_rsc_0_26_qa, xt_rsc_triosy_0_26_lz,
      xt_rsc_0_27_adra, xt_rsc_0_27_da, xt_rsc_0_27_wea, xt_rsc_0_27_qa, xt_rsc_triosy_0_27_lz,
      xt_rsc_0_28_adra, xt_rsc_0_28_da, xt_rsc_0_28_wea, xt_rsc_0_28_qa, xt_rsc_triosy_0_28_lz,
      xt_rsc_0_29_adra, xt_rsc_0_29_da, xt_rsc_0_29_wea, xt_rsc_0_29_qa, xt_rsc_triosy_0_29_lz,
      xt_rsc_0_30_adra, xt_rsc_0_30_da, xt_rsc_0_30_wea, xt_rsc_0_30_qa, xt_rsc_triosy_0_30_lz,
      xt_rsc_0_31_adra, xt_rsc_0_31_da, xt_rsc_0_31_wea, xt_rsc_0_31_qa, xt_rsc_triosy_0_31_lz,
      xt_rsc_1_0_adra, xt_rsc_1_0_da, xt_rsc_1_0_wea, xt_rsc_1_0_qa, xt_rsc_triosy_1_0_lz,
      xt_rsc_1_1_adra, xt_rsc_1_1_da, xt_rsc_1_1_wea, xt_rsc_1_1_qa, xt_rsc_triosy_1_1_lz,
      xt_rsc_1_2_adra, xt_rsc_1_2_da, xt_rsc_1_2_wea, xt_rsc_1_2_qa, xt_rsc_triosy_1_2_lz,
      xt_rsc_1_3_adra, xt_rsc_1_3_da, xt_rsc_1_3_wea, xt_rsc_1_3_qa, xt_rsc_triosy_1_3_lz,
      xt_rsc_1_4_adra, xt_rsc_1_4_da, xt_rsc_1_4_wea, xt_rsc_1_4_qa, xt_rsc_triosy_1_4_lz,
      xt_rsc_1_5_adra, xt_rsc_1_5_da, xt_rsc_1_5_wea, xt_rsc_1_5_qa, xt_rsc_triosy_1_5_lz,
      xt_rsc_1_6_adra, xt_rsc_1_6_da, xt_rsc_1_6_wea, xt_rsc_1_6_qa, xt_rsc_triosy_1_6_lz,
      xt_rsc_1_7_adra, xt_rsc_1_7_da, xt_rsc_1_7_wea, xt_rsc_1_7_qa, xt_rsc_triosy_1_7_lz,
      xt_rsc_1_8_adra, xt_rsc_1_8_da, xt_rsc_1_8_wea, xt_rsc_1_8_qa, xt_rsc_triosy_1_8_lz,
      xt_rsc_1_9_adra, xt_rsc_1_9_da, xt_rsc_1_9_wea, xt_rsc_1_9_qa, xt_rsc_triosy_1_9_lz,
      xt_rsc_1_10_adra, xt_rsc_1_10_da, xt_rsc_1_10_wea, xt_rsc_1_10_qa, xt_rsc_triosy_1_10_lz,
      xt_rsc_1_11_adra, xt_rsc_1_11_da, xt_rsc_1_11_wea, xt_rsc_1_11_qa, xt_rsc_triosy_1_11_lz,
      xt_rsc_1_12_adra, xt_rsc_1_12_da, xt_rsc_1_12_wea, xt_rsc_1_12_qa, xt_rsc_triosy_1_12_lz,
      xt_rsc_1_13_adra, xt_rsc_1_13_da, xt_rsc_1_13_wea, xt_rsc_1_13_qa, xt_rsc_triosy_1_13_lz,
      xt_rsc_1_14_adra, xt_rsc_1_14_da, xt_rsc_1_14_wea, xt_rsc_1_14_qa, xt_rsc_triosy_1_14_lz,
      xt_rsc_1_15_adra, xt_rsc_1_15_da, xt_rsc_1_15_wea, xt_rsc_1_15_qa, xt_rsc_triosy_1_15_lz,
      xt_rsc_1_16_adra, xt_rsc_1_16_da, xt_rsc_1_16_wea, xt_rsc_1_16_qa, xt_rsc_triosy_1_16_lz,
      xt_rsc_1_17_adra, xt_rsc_1_17_da, xt_rsc_1_17_wea, xt_rsc_1_17_qa, xt_rsc_triosy_1_17_lz,
      xt_rsc_1_18_adra, xt_rsc_1_18_da, xt_rsc_1_18_wea, xt_rsc_1_18_qa, xt_rsc_triosy_1_18_lz,
      xt_rsc_1_19_adra, xt_rsc_1_19_da, xt_rsc_1_19_wea, xt_rsc_1_19_qa, xt_rsc_triosy_1_19_lz,
      xt_rsc_1_20_adra, xt_rsc_1_20_da, xt_rsc_1_20_wea, xt_rsc_1_20_qa, xt_rsc_triosy_1_20_lz,
      xt_rsc_1_21_adra, xt_rsc_1_21_da, xt_rsc_1_21_wea, xt_rsc_1_21_qa, xt_rsc_triosy_1_21_lz,
      xt_rsc_1_22_adra, xt_rsc_1_22_da, xt_rsc_1_22_wea, xt_rsc_1_22_qa, xt_rsc_triosy_1_22_lz,
      xt_rsc_1_23_adra, xt_rsc_1_23_da, xt_rsc_1_23_wea, xt_rsc_1_23_qa, xt_rsc_triosy_1_23_lz,
      xt_rsc_1_24_adra, xt_rsc_1_24_da, xt_rsc_1_24_wea, xt_rsc_1_24_qa, xt_rsc_triosy_1_24_lz,
      xt_rsc_1_25_adra, xt_rsc_1_25_da, xt_rsc_1_25_wea, xt_rsc_1_25_qa, xt_rsc_triosy_1_25_lz,
      xt_rsc_1_26_adra, xt_rsc_1_26_da, xt_rsc_1_26_wea, xt_rsc_1_26_qa, xt_rsc_triosy_1_26_lz,
      xt_rsc_1_27_adra, xt_rsc_1_27_da, xt_rsc_1_27_wea, xt_rsc_1_27_qa, xt_rsc_triosy_1_27_lz,
      xt_rsc_1_28_adra, xt_rsc_1_28_da, xt_rsc_1_28_wea, xt_rsc_1_28_qa, xt_rsc_triosy_1_28_lz,
      xt_rsc_1_29_adra, xt_rsc_1_29_da, xt_rsc_1_29_wea, xt_rsc_1_29_qa, xt_rsc_triosy_1_29_lz,
      xt_rsc_1_30_adra, xt_rsc_1_30_da, xt_rsc_1_30_wea, xt_rsc_1_30_qa, xt_rsc_triosy_1_30_lz,
      xt_rsc_1_31_adra, xt_rsc_1_31_da, xt_rsc_1_31_wea, xt_rsc_1_31_qa, xt_rsc_triosy_1_31_lz,
      xt_rsc_2_0_adra, xt_rsc_2_0_da, xt_rsc_2_0_wea, xt_rsc_2_0_qa, xt_rsc_triosy_2_0_lz,
      xt_rsc_2_1_adra, xt_rsc_2_1_da, xt_rsc_2_1_wea, xt_rsc_2_1_qa, xt_rsc_triosy_2_1_lz,
      xt_rsc_2_2_adra, xt_rsc_2_2_da, xt_rsc_2_2_wea, xt_rsc_2_2_qa, xt_rsc_triosy_2_2_lz,
      xt_rsc_2_3_adra, xt_rsc_2_3_da, xt_rsc_2_3_wea, xt_rsc_2_3_qa, xt_rsc_triosy_2_3_lz,
      xt_rsc_2_4_adra, xt_rsc_2_4_da, xt_rsc_2_4_wea, xt_rsc_2_4_qa, xt_rsc_triosy_2_4_lz,
      xt_rsc_2_5_adra, xt_rsc_2_5_da, xt_rsc_2_5_wea, xt_rsc_2_5_qa, xt_rsc_triosy_2_5_lz,
      xt_rsc_2_6_adra, xt_rsc_2_6_da, xt_rsc_2_6_wea, xt_rsc_2_6_qa, xt_rsc_triosy_2_6_lz,
      xt_rsc_2_7_adra, xt_rsc_2_7_da, xt_rsc_2_7_wea, xt_rsc_2_7_qa, xt_rsc_triosy_2_7_lz,
      xt_rsc_2_8_adra, xt_rsc_2_8_da, xt_rsc_2_8_wea, xt_rsc_2_8_qa, xt_rsc_triosy_2_8_lz,
      xt_rsc_2_9_adra, xt_rsc_2_9_da, xt_rsc_2_9_wea, xt_rsc_2_9_qa, xt_rsc_triosy_2_9_lz,
      xt_rsc_2_10_adra, xt_rsc_2_10_da, xt_rsc_2_10_wea, xt_rsc_2_10_qa, xt_rsc_triosy_2_10_lz,
      xt_rsc_2_11_adra, xt_rsc_2_11_da, xt_rsc_2_11_wea, xt_rsc_2_11_qa, xt_rsc_triosy_2_11_lz,
      xt_rsc_2_12_adra, xt_rsc_2_12_da, xt_rsc_2_12_wea, xt_rsc_2_12_qa, xt_rsc_triosy_2_12_lz,
      xt_rsc_2_13_adra, xt_rsc_2_13_da, xt_rsc_2_13_wea, xt_rsc_2_13_qa, xt_rsc_triosy_2_13_lz,
      xt_rsc_2_14_adra, xt_rsc_2_14_da, xt_rsc_2_14_wea, xt_rsc_2_14_qa, xt_rsc_triosy_2_14_lz,
      xt_rsc_2_15_adra, xt_rsc_2_15_da, xt_rsc_2_15_wea, xt_rsc_2_15_qa, xt_rsc_triosy_2_15_lz,
      xt_rsc_2_16_adra, xt_rsc_2_16_da, xt_rsc_2_16_wea, xt_rsc_2_16_qa, xt_rsc_triosy_2_16_lz,
      xt_rsc_2_17_adra, xt_rsc_2_17_da, xt_rsc_2_17_wea, xt_rsc_2_17_qa, xt_rsc_triosy_2_17_lz,
      xt_rsc_2_18_adra, xt_rsc_2_18_da, xt_rsc_2_18_wea, xt_rsc_2_18_qa, xt_rsc_triosy_2_18_lz,
      xt_rsc_2_19_adra, xt_rsc_2_19_da, xt_rsc_2_19_wea, xt_rsc_2_19_qa, xt_rsc_triosy_2_19_lz,
      xt_rsc_2_20_adra, xt_rsc_2_20_da, xt_rsc_2_20_wea, xt_rsc_2_20_qa, xt_rsc_triosy_2_20_lz,
      xt_rsc_2_21_adra, xt_rsc_2_21_da, xt_rsc_2_21_wea, xt_rsc_2_21_qa, xt_rsc_triosy_2_21_lz,
      xt_rsc_2_22_adra, xt_rsc_2_22_da, xt_rsc_2_22_wea, xt_rsc_2_22_qa, xt_rsc_triosy_2_22_lz,
      xt_rsc_2_23_adra, xt_rsc_2_23_da, xt_rsc_2_23_wea, xt_rsc_2_23_qa, xt_rsc_triosy_2_23_lz,
      xt_rsc_2_24_adra, xt_rsc_2_24_da, xt_rsc_2_24_wea, xt_rsc_2_24_qa, xt_rsc_triosy_2_24_lz,
      xt_rsc_2_25_adra, xt_rsc_2_25_da, xt_rsc_2_25_wea, xt_rsc_2_25_qa, xt_rsc_triosy_2_25_lz,
      xt_rsc_2_26_adra, xt_rsc_2_26_da, xt_rsc_2_26_wea, xt_rsc_2_26_qa, xt_rsc_triosy_2_26_lz,
      xt_rsc_2_27_adra, xt_rsc_2_27_da, xt_rsc_2_27_wea, xt_rsc_2_27_qa, xt_rsc_triosy_2_27_lz,
      xt_rsc_2_28_adra, xt_rsc_2_28_da, xt_rsc_2_28_wea, xt_rsc_2_28_qa, xt_rsc_triosy_2_28_lz,
      xt_rsc_2_29_adra, xt_rsc_2_29_da, xt_rsc_2_29_wea, xt_rsc_2_29_qa, xt_rsc_triosy_2_29_lz,
      xt_rsc_2_30_adra, xt_rsc_2_30_da, xt_rsc_2_30_wea, xt_rsc_2_30_qa, xt_rsc_triosy_2_30_lz,
      xt_rsc_2_31_adra, xt_rsc_2_31_da, xt_rsc_2_31_wea, xt_rsc_2_31_qa, xt_rsc_triosy_2_31_lz,
      xt_rsc_3_0_adra, xt_rsc_3_0_da, xt_rsc_3_0_wea, xt_rsc_3_0_qa, xt_rsc_triosy_3_0_lz,
      xt_rsc_3_1_adra, xt_rsc_3_1_da, xt_rsc_3_1_wea, xt_rsc_3_1_qa, xt_rsc_triosy_3_1_lz,
      xt_rsc_3_2_adra, xt_rsc_3_2_da, xt_rsc_3_2_wea, xt_rsc_3_2_qa, xt_rsc_triosy_3_2_lz,
      xt_rsc_3_3_adra, xt_rsc_3_3_da, xt_rsc_3_3_wea, xt_rsc_3_3_qa, xt_rsc_triosy_3_3_lz,
      xt_rsc_3_4_adra, xt_rsc_3_4_da, xt_rsc_3_4_wea, xt_rsc_3_4_qa, xt_rsc_triosy_3_4_lz,
      xt_rsc_3_5_adra, xt_rsc_3_5_da, xt_rsc_3_5_wea, xt_rsc_3_5_qa, xt_rsc_triosy_3_5_lz,
      xt_rsc_3_6_adra, xt_rsc_3_6_da, xt_rsc_3_6_wea, xt_rsc_3_6_qa, xt_rsc_triosy_3_6_lz,
      xt_rsc_3_7_adra, xt_rsc_3_7_da, xt_rsc_3_7_wea, xt_rsc_3_7_qa, xt_rsc_triosy_3_7_lz,
      xt_rsc_3_8_adra, xt_rsc_3_8_da, xt_rsc_3_8_wea, xt_rsc_3_8_qa, xt_rsc_triosy_3_8_lz,
      xt_rsc_3_9_adra, xt_rsc_3_9_da, xt_rsc_3_9_wea, xt_rsc_3_9_qa, xt_rsc_triosy_3_9_lz,
      xt_rsc_3_10_adra, xt_rsc_3_10_da, xt_rsc_3_10_wea, xt_rsc_3_10_qa, xt_rsc_triosy_3_10_lz,
      xt_rsc_3_11_adra, xt_rsc_3_11_da, xt_rsc_3_11_wea, xt_rsc_3_11_qa, xt_rsc_triosy_3_11_lz,
      xt_rsc_3_12_adra, xt_rsc_3_12_da, xt_rsc_3_12_wea, xt_rsc_3_12_qa, xt_rsc_triosy_3_12_lz,
      xt_rsc_3_13_adra, xt_rsc_3_13_da, xt_rsc_3_13_wea, xt_rsc_3_13_qa, xt_rsc_triosy_3_13_lz,
      xt_rsc_3_14_adra, xt_rsc_3_14_da, xt_rsc_3_14_wea, xt_rsc_3_14_qa, xt_rsc_triosy_3_14_lz,
      xt_rsc_3_15_adra, xt_rsc_3_15_da, xt_rsc_3_15_wea, xt_rsc_3_15_qa, xt_rsc_triosy_3_15_lz,
      xt_rsc_3_16_adra, xt_rsc_3_16_da, xt_rsc_3_16_wea, xt_rsc_3_16_qa, xt_rsc_triosy_3_16_lz,
      xt_rsc_3_17_adra, xt_rsc_3_17_da, xt_rsc_3_17_wea, xt_rsc_3_17_qa, xt_rsc_triosy_3_17_lz,
      xt_rsc_3_18_adra, xt_rsc_3_18_da, xt_rsc_3_18_wea, xt_rsc_3_18_qa, xt_rsc_triosy_3_18_lz,
      xt_rsc_3_19_adra, xt_rsc_3_19_da, xt_rsc_3_19_wea, xt_rsc_3_19_qa, xt_rsc_triosy_3_19_lz,
      xt_rsc_3_20_adra, xt_rsc_3_20_da, xt_rsc_3_20_wea, xt_rsc_3_20_qa, xt_rsc_triosy_3_20_lz,
      xt_rsc_3_21_adra, xt_rsc_3_21_da, xt_rsc_3_21_wea, xt_rsc_3_21_qa, xt_rsc_triosy_3_21_lz,
      xt_rsc_3_22_adra, xt_rsc_3_22_da, xt_rsc_3_22_wea, xt_rsc_3_22_qa, xt_rsc_triosy_3_22_lz,
      xt_rsc_3_23_adra, xt_rsc_3_23_da, xt_rsc_3_23_wea, xt_rsc_3_23_qa, xt_rsc_triosy_3_23_lz,
      xt_rsc_3_24_adra, xt_rsc_3_24_da, xt_rsc_3_24_wea, xt_rsc_3_24_qa, xt_rsc_triosy_3_24_lz,
      xt_rsc_3_25_adra, xt_rsc_3_25_da, xt_rsc_3_25_wea, xt_rsc_3_25_qa, xt_rsc_triosy_3_25_lz,
      xt_rsc_3_26_adra, xt_rsc_3_26_da, xt_rsc_3_26_wea, xt_rsc_3_26_qa, xt_rsc_triosy_3_26_lz,
      xt_rsc_3_27_adra, xt_rsc_3_27_da, xt_rsc_3_27_wea, xt_rsc_3_27_qa, xt_rsc_triosy_3_27_lz,
      xt_rsc_3_28_adra, xt_rsc_3_28_da, xt_rsc_3_28_wea, xt_rsc_3_28_qa, xt_rsc_triosy_3_28_lz,
      xt_rsc_3_29_adra, xt_rsc_3_29_da, xt_rsc_3_29_wea, xt_rsc_3_29_qa, xt_rsc_triosy_3_29_lz,
      xt_rsc_3_30_adra, xt_rsc_3_30_da, xt_rsc_3_30_wea, xt_rsc_3_30_qa, xt_rsc_triosy_3_30_lz,
      xt_rsc_3_31_adra, xt_rsc_3_31_da, xt_rsc_3_31_wea, xt_rsc_3_31_qa, xt_rsc_triosy_3_31_lz,
      xt_rsc_4_0_adra, xt_rsc_4_0_da, xt_rsc_4_0_wea, xt_rsc_4_0_qa, xt_rsc_triosy_4_0_lz,
      xt_rsc_4_1_adra, xt_rsc_4_1_da, xt_rsc_4_1_wea, xt_rsc_4_1_qa, xt_rsc_triosy_4_1_lz,
      xt_rsc_4_2_adra, xt_rsc_4_2_da, xt_rsc_4_2_wea, xt_rsc_4_2_qa, xt_rsc_triosy_4_2_lz,
      xt_rsc_4_3_adra, xt_rsc_4_3_da, xt_rsc_4_3_wea, xt_rsc_4_3_qa, xt_rsc_triosy_4_3_lz,
      xt_rsc_4_4_adra, xt_rsc_4_4_da, xt_rsc_4_4_wea, xt_rsc_4_4_qa, xt_rsc_triosy_4_4_lz,
      xt_rsc_4_5_adra, xt_rsc_4_5_da, xt_rsc_4_5_wea, xt_rsc_4_5_qa, xt_rsc_triosy_4_5_lz,
      xt_rsc_4_6_adra, xt_rsc_4_6_da, xt_rsc_4_6_wea, xt_rsc_4_6_qa, xt_rsc_triosy_4_6_lz,
      xt_rsc_4_7_adra, xt_rsc_4_7_da, xt_rsc_4_7_wea, xt_rsc_4_7_qa, xt_rsc_triosy_4_7_lz,
      xt_rsc_4_8_adra, xt_rsc_4_8_da, xt_rsc_4_8_wea, xt_rsc_4_8_qa, xt_rsc_triosy_4_8_lz,
      xt_rsc_4_9_adra, xt_rsc_4_9_da, xt_rsc_4_9_wea, xt_rsc_4_9_qa, xt_rsc_triosy_4_9_lz,
      xt_rsc_4_10_adra, xt_rsc_4_10_da, xt_rsc_4_10_wea, xt_rsc_4_10_qa, xt_rsc_triosy_4_10_lz,
      xt_rsc_4_11_adra, xt_rsc_4_11_da, xt_rsc_4_11_wea, xt_rsc_4_11_qa, xt_rsc_triosy_4_11_lz,
      xt_rsc_4_12_adra, xt_rsc_4_12_da, xt_rsc_4_12_wea, xt_rsc_4_12_qa, xt_rsc_triosy_4_12_lz,
      xt_rsc_4_13_adra, xt_rsc_4_13_da, xt_rsc_4_13_wea, xt_rsc_4_13_qa, xt_rsc_triosy_4_13_lz,
      xt_rsc_4_14_adra, xt_rsc_4_14_da, xt_rsc_4_14_wea, xt_rsc_4_14_qa, xt_rsc_triosy_4_14_lz,
      xt_rsc_4_15_adra, xt_rsc_4_15_da, xt_rsc_4_15_wea, xt_rsc_4_15_qa, xt_rsc_triosy_4_15_lz,
      xt_rsc_4_16_adra, xt_rsc_4_16_da, xt_rsc_4_16_wea, xt_rsc_4_16_qa, xt_rsc_triosy_4_16_lz,
      xt_rsc_4_17_adra, xt_rsc_4_17_da, xt_rsc_4_17_wea, xt_rsc_4_17_qa, xt_rsc_triosy_4_17_lz,
      xt_rsc_4_18_adra, xt_rsc_4_18_da, xt_rsc_4_18_wea, xt_rsc_4_18_qa, xt_rsc_triosy_4_18_lz,
      xt_rsc_4_19_adra, xt_rsc_4_19_da, xt_rsc_4_19_wea, xt_rsc_4_19_qa, xt_rsc_triosy_4_19_lz,
      xt_rsc_4_20_adra, xt_rsc_4_20_da, xt_rsc_4_20_wea, xt_rsc_4_20_qa, xt_rsc_triosy_4_20_lz,
      xt_rsc_4_21_adra, xt_rsc_4_21_da, xt_rsc_4_21_wea, xt_rsc_4_21_qa, xt_rsc_triosy_4_21_lz,
      xt_rsc_4_22_adra, xt_rsc_4_22_da, xt_rsc_4_22_wea, xt_rsc_4_22_qa, xt_rsc_triosy_4_22_lz,
      xt_rsc_4_23_adra, xt_rsc_4_23_da, xt_rsc_4_23_wea, xt_rsc_4_23_qa, xt_rsc_triosy_4_23_lz,
      xt_rsc_4_24_adra, xt_rsc_4_24_da, xt_rsc_4_24_wea, xt_rsc_4_24_qa, xt_rsc_triosy_4_24_lz,
      xt_rsc_4_25_adra, xt_rsc_4_25_da, xt_rsc_4_25_wea, xt_rsc_4_25_qa, xt_rsc_triosy_4_25_lz,
      xt_rsc_4_26_adra, xt_rsc_4_26_da, xt_rsc_4_26_wea, xt_rsc_4_26_qa, xt_rsc_triosy_4_26_lz,
      xt_rsc_4_27_adra, xt_rsc_4_27_da, xt_rsc_4_27_wea, xt_rsc_4_27_qa, xt_rsc_triosy_4_27_lz,
      xt_rsc_4_28_adra, xt_rsc_4_28_da, xt_rsc_4_28_wea, xt_rsc_4_28_qa, xt_rsc_triosy_4_28_lz,
      xt_rsc_4_29_adra, xt_rsc_4_29_da, xt_rsc_4_29_wea, xt_rsc_4_29_qa, xt_rsc_triosy_4_29_lz,
      xt_rsc_4_30_adra, xt_rsc_4_30_da, xt_rsc_4_30_wea, xt_rsc_4_30_qa, xt_rsc_triosy_4_30_lz,
      xt_rsc_4_31_adra, xt_rsc_4_31_da, xt_rsc_4_31_wea, xt_rsc_4_31_qa, xt_rsc_triosy_4_31_lz,
      xt_rsc_5_0_adra, xt_rsc_5_0_da, xt_rsc_5_0_wea, xt_rsc_5_0_qa, xt_rsc_triosy_5_0_lz,
      xt_rsc_5_1_adra, xt_rsc_5_1_da, xt_rsc_5_1_wea, xt_rsc_5_1_qa, xt_rsc_triosy_5_1_lz,
      xt_rsc_5_2_adra, xt_rsc_5_2_da, xt_rsc_5_2_wea, xt_rsc_5_2_qa, xt_rsc_triosy_5_2_lz,
      xt_rsc_5_3_adra, xt_rsc_5_3_da, xt_rsc_5_3_wea, xt_rsc_5_3_qa, xt_rsc_triosy_5_3_lz,
      xt_rsc_5_4_adra, xt_rsc_5_4_da, xt_rsc_5_4_wea, xt_rsc_5_4_qa, xt_rsc_triosy_5_4_lz,
      xt_rsc_5_5_adra, xt_rsc_5_5_da, xt_rsc_5_5_wea, xt_rsc_5_5_qa, xt_rsc_triosy_5_5_lz,
      xt_rsc_5_6_adra, xt_rsc_5_6_da, xt_rsc_5_6_wea, xt_rsc_5_6_qa, xt_rsc_triosy_5_6_lz,
      xt_rsc_5_7_adra, xt_rsc_5_7_da, xt_rsc_5_7_wea, xt_rsc_5_7_qa, xt_rsc_triosy_5_7_lz,
      xt_rsc_5_8_adra, xt_rsc_5_8_da, xt_rsc_5_8_wea, xt_rsc_5_8_qa, xt_rsc_triosy_5_8_lz,
      xt_rsc_5_9_adra, xt_rsc_5_9_da, xt_rsc_5_9_wea, xt_rsc_5_9_qa, xt_rsc_triosy_5_9_lz,
      xt_rsc_5_10_adra, xt_rsc_5_10_da, xt_rsc_5_10_wea, xt_rsc_5_10_qa, xt_rsc_triosy_5_10_lz,
      xt_rsc_5_11_adra, xt_rsc_5_11_da, xt_rsc_5_11_wea, xt_rsc_5_11_qa, xt_rsc_triosy_5_11_lz,
      xt_rsc_5_12_adra, xt_rsc_5_12_da, xt_rsc_5_12_wea, xt_rsc_5_12_qa, xt_rsc_triosy_5_12_lz,
      xt_rsc_5_13_adra, xt_rsc_5_13_da, xt_rsc_5_13_wea, xt_rsc_5_13_qa, xt_rsc_triosy_5_13_lz,
      xt_rsc_5_14_adra, xt_rsc_5_14_da, xt_rsc_5_14_wea, xt_rsc_5_14_qa, xt_rsc_triosy_5_14_lz,
      xt_rsc_5_15_adra, xt_rsc_5_15_da, xt_rsc_5_15_wea, xt_rsc_5_15_qa, xt_rsc_triosy_5_15_lz,
      xt_rsc_5_16_adra, xt_rsc_5_16_da, xt_rsc_5_16_wea, xt_rsc_5_16_qa, xt_rsc_triosy_5_16_lz,
      xt_rsc_5_17_adra, xt_rsc_5_17_da, xt_rsc_5_17_wea, xt_rsc_5_17_qa, xt_rsc_triosy_5_17_lz,
      xt_rsc_5_18_adra, xt_rsc_5_18_da, xt_rsc_5_18_wea, xt_rsc_5_18_qa, xt_rsc_triosy_5_18_lz,
      xt_rsc_5_19_adra, xt_rsc_5_19_da, xt_rsc_5_19_wea, xt_rsc_5_19_qa, xt_rsc_triosy_5_19_lz,
      xt_rsc_5_20_adra, xt_rsc_5_20_da, xt_rsc_5_20_wea, xt_rsc_5_20_qa, xt_rsc_triosy_5_20_lz,
      xt_rsc_5_21_adra, xt_rsc_5_21_da, xt_rsc_5_21_wea, xt_rsc_5_21_qa, xt_rsc_triosy_5_21_lz,
      xt_rsc_5_22_adra, xt_rsc_5_22_da, xt_rsc_5_22_wea, xt_rsc_5_22_qa, xt_rsc_triosy_5_22_lz,
      xt_rsc_5_23_adra, xt_rsc_5_23_da, xt_rsc_5_23_wea, xt_rsc_5_23_qa, xt_rsc_triosy_5_23_lz,
      xt_rsc_5_24_adra, xt_rsc_5_24_da, xt_rsc_5_24_wea, xt_rsc_5_24_qa, xt_rsc_triosy_5_24_lz,
      xt_rsc_5_25_adra, xt_rsc_5_25_da, xt_rsc_5_25_wea, xt_rsc_5_25_qa, xt_rsc_triosy_5_25_lz,
      xt_rsc_5_26_adra, xt_rsc_5_26_da, xt_rsc_5_26_wea, xt_rsc_5_26_qa, xt_rsc_triosy_5_26_lz,
      xt_rsc_5_27_adra, xt_rsc_5_27_da, xt_rsc_5_27_wea, xt_rsc_5_27_qa, xt_rsc_triosy_5_27_lz,
      xt_rsc_5_28_adra, xt_rsc_5_28_da, xt_rsc_5_28_wea, xt_rsc_5_28_qa, xt_rsc_triosy_5_28_lz,
      xt_rsc_5_29_adra, xt_rsc_5_29_da, xt_rsc_5_29_wea, xt_rsc_5_29_qa, xt_rsc_triosy_5_29_lz,
      xt_rsc_5_30_adra, xt_rsc_5_30_da, xt_rsc_5_30_wea, xt_rsc_5_30_qa, xt_rsc_triosy_5_30_lz,
      xt_rsc_5_31_adra, xt_rsc_5_31_da, xt_rsc_5_31_wea, xt_rsc_5_31_qa, xt_rsc_triosy_5_31_lz,
      xt_rsc_6_0_adra, xt_rsc_6_0_da, xt_rsc_6_0_wea, xt_rsc_6_0_qa, xt_rsc_triosy_6_0_lz,
      xt_rsc_6_1_adra, xt_rsc_6_1_da, xt_rsc_6_1_wea, xt_rsc_6_1_qa, xt_rsc_triosy_6_1_lz,
      xt_rsc_6_2_adra, xt_rsc_6_2_da, xt_rsc_6_2_wea, xt_rsc_6_2_qa, xt_rsc_triosy_6_2_lz,
      xt_rsc_6_3_adra, xt_rsc_6_3_da, xt_rsc_6_3_wea, xt_rsc_6_3_qa, xt_rsc_triosy_6_3_lz,
      xt_rsc_6_4_adra, xt_rsc_6_4_da, xt_rsc_6_4_wea, xt_rsc_6_4_qa, xt_rsc_triosy_6_4_lz,
      xt_rsc_6_5_adra, xt_rsc_6_5_da, xt_rsc_6_5_wea, xt_rsc_6_5_qa, xt_rsc_triosy_6_5_lz,
      xt_rsc_6_6_adra, xt_rsc_6_6_da, xt_rsc_6_6_wea, xt_rsc_6_6_qa, xt_rsc_triosy_6_6_lz,
      xt_rsc_6_7_adra, xt_rsc_6_7_da, xt_rsc_6_7_wea, xt_rsc_6_7_qa, xt_rsc_triosy_6_7_lz,
      xt_rsc_6_8_adra, xt_rsc_6_8_da, xt_rsc_6_8_wea, xt_rsc_6_8_qa, xt_rsc_triosy_6_8_lz,
      xt_rsc_6_9_adra, xt_rsc_6_9_da, xt_rsc_6_9_wea, xt_rsc_6_9_qa, xt_rsc_triosy_6_9_lz,
      xt_rsc_6_10_adra, xt_rsc_6_10_da, xt_rsc_6_10_wea, xt_rsc_6_10_qa, xt_rsc_triosy_6_10_lz,
      xt_rsc_6_11_adra, xt_rsc_6_11_da, xt_rsc_6_11_wea, xt_rsc_6_11_qa, xt_rsc_triosy_6_11_lz,
      xt_rsc_6_12_adra, xt_rsc_6_12_da, xt_rsc_6_12_wea, xt_rsc_6_12_qa, xt_rsc_triosy_6_12_lz,
      xt_rsc_6_13_adra, xt_rsc_6_13_da, xt_rsc_6_13_wea, xt_rsc_6_13_qa, xt_rsc_triosy_6_13_lz,
      xt_rsc_6_14_adra, xt_rsc_6_14_da, xt_rsc_6_14_wea, xt_rsc_6_14_qa, xt_rsc_triosy_6_14_lz,
      xt_rsc_6_15_adra, xt_rsc_6_15_da, xt_rsc_6_15_wea, xt_rsc_6_15_qa, xt_rsc_triosy_6_15_lz,
      xt_rsc_6_16_adra, xt_rsc_6_16_da, xt_rsc_6_16_wea, xt_rsc_6_16_qa, xt_rsc_triosy_6_16_lz,
      xt_rsc_6_17_adra, xt_rsc_6_17_da, xt_rsc_6_17_wea, xt_rsc_6_17_qa, xt_rsc_triosy_6_17_lz,
      xt_rsc_6_18_adra, xt_rsc_6_18_da, xt_rsc_6_18_wea, xt_rsc_6_18_qa, xt_rsc_triosy_6_18_lz,
      xt_rsc_6_19_adra, xt_rsc_6_19_da, xt_rsc_6_19_wea, xt_rsc_6_19_qa, xt_rsc_triosy_6_19_lz,
      xt_rsc_6_20_adra, xt_rsc_6_20_da, xt_rsc_6_20_wea, xt_rsc_6_20_qa, xt_rsc_triosy_6_20_lz,
      xt_rsc_6_21_adra, xt_rsc_6_21_da, xt_rsc_6_21_wea, xt_rsc_6_21_qa, xt_rsc_triosy_6_21_lz,
      xt_rsc_6_22_adra, xt_rsc_6_22_da, xt_rsc_6_22_wea, xt_rsc_6_22_qa, xt_rsc_triosy_6_22_lz,
      xt_rsc_6_23_adra, xt_rsc_6_23_da, xt_rsc_6_23_wea, xt_rsc_6_23_qa, xt_rsc_triosy_6_23_lz,
      xt_rsc_6_24_adra, xt_rsc_6_24_da, xt_rsc_6_24_wea, xt_rsc_6_24_qa, xt_rsc_triosy_6_24_lz,
      xt_rsc_6_25_adra, xt_rsc_6_25_da, xt_rsc_6_25_wea, xt_rsc_6_25_qa, xt_rsc_triosy_6_25_lz,
      xt_rsc_6_26_adra, xt_rsc_6_26_da, xt_rsc_6_26_wea, xt_rsc_6_26_qa, xt_rsc_triosy_6_26_lz,
      xt_rsc_6_27_adra, xt_rsc_6_27_da, xt_rsc_6_27_wea, xt_rsc_6_27_qa, xt_rsc_triosy_6_27_lz,
      xt_rsc_6_28_adra, xt_rsc_6_28_da, xt_rsc_6_28_wea, xt_rsc_6_28_qa, xt_rsc_triosy_6_28_lz,
      xt_rsc_6_29_adra, xt_rsc_6_29_da, xt_rsc_6_29_wea, xt_rsc_6_29_qa, xt_rsc_triosy_6_29_lz,
      xt_rsc_6_30_adra, xt_rsc_6_30_da, xt_rsc_6_30_wea, xt_rsc_6_30_qa, xt_rsc_triosy_6_30_lz,
      xt_rsc_6_31_adra, xt_rsc_6_31_da, xt_rsc_6_31_wea, xt_rsc_6_31_qa, xt_rsc_triosy_6_31_lz,
      xt_rsc_7_0_adra, xt_rsc_7_0_da, xt_rsc_7_0_wea, xt_rsc_7_0_qa, xt_rsc_triosy_7_0_lz,
      xt_rsc_7_1_adra, xt_rsc_7_1_da, xt_rsc_7_1_wea, xt_rsc_7_1_qa, xt_rsc_triosy_7_1_lz,
      xt_rsc_7_2_adra, xt_rsc_7_2_da, xt_rsc_7_2_wea, xt_rsc_7_2_qa, xt_rsc_triosy_7_2_lz,
      xt_rsc_7_3_adra, xt_rsc_7_3_da, xt_rsc_7_3_wea, xt_rsc_7_3_qa, xt_rsc_triosy_7_3_lz,
      xt_rsc_7_4_adra, xt_rsc_7_4_da, xt_rsc_7_4_wea, xt_rsc_7_4_qa, xt_rsc_triosy_7_4_lz,
      xt_rsc_7_5_adra, xt_rsc_7_5_da, xt_rsc_7_5_wea, xt_rsc_7_5_qa, xt_rsc_triosy_7_5_lz,
      xt_rsc_7_6_adra, xt_rsc_7_6_da, xt_rsc_7_6_wea, xt_rsc_7_6_qa, xt_rsc_triosy_7_6_lz,
      xt_rsc_7_7_adra, xt_rsc_7_7_da, xt_rsc_7_7_wea, xt_rsc_7_7_qa, xt_rsc_triosy_7_7_lz,
      xt_rsc_7_8_adra, xt_rsc_7_8_da, xt_rsc_7_8_wea, xt_rsc_7_8_qa, xt_rsc_triosy_7_8_lz,
      xt_rsc_7_9_adra, xt_rsc_7_9_da, xt_rsc_7_9_wea, xt_rsc_7_9_qa, xt_rsc_triosy_7_9_lz,
      xt_rsc_7_10_adra, xt_rsc_7_10_da, xt_rsc_7_10_wea, xt_rsc_7_10_qa, xt_rsc_triosy_7_10_lz,
      xt_rsc_7_11_adra, xt_rsc_7_11_da, xt_rsc_7_11_wea, xt_rsc_7_11_qa, xt_rsc_triosy_7_11_lz,
      xt_rsc_7_12_adra, xt_rsc_7_12_da, xt_rsc_7_12_wea, xt_rsc_7_12_qa, xt_rsc_triosy_7_12_lz,
      xt_rsc_7_13_adra, xt_rsc_7_13_da, xt_rsc_7_13_wea, xt_rsc_7_13_qa, xt_rsc_triosy_7_13_lz,
      xt_rsc_7_14_adra, xt_rsc_7_14_da, xt_rsc_7_14_wea, xt_rsc_7_14_qa, xt_rsc_triosy_7_14_lz,
      xt_rsc_7_15_adra, xt_rsc_7_15_da, xt_rsc_7_15_wea, xt_rsc_7_15_qa, xt_rsc_triosy_7_15_lz,
      xt_rsc_7_16_adra, xt_rsc_7_16_da, xt_rsc_7_16_wea, xt_rsc_7_16_qa, xt_rsc_triosy_7_16_lz,
      xt_rsc_7_17_adra, xt_rsc_7_17_da, xt_rsc_7_17_wea, xt_rsc_7_17_qa, xt_rsc_triosy_7_17_lz,
      xt_rsc_7_18_adra, xt_rsc_7_18_da, xt_rsc_7_18_wea, xt_rsc_7_18_qa, xt_rsc_triosy_7_18_lz,
      xt_rsc_7_19_adra, xt_rsc_7_19_da, xt_rsc_7_19_wea, xt_rsc_7_19_qa, xt_rsc_triosy_7_19_lz,
      xt_rsc_7_20_adra, xt_rsc_7_20_da, xt_rsc_7_20_wea, xt_rsc_7_20_qa, xt_rsc_triosy_7_20_lz,
      xt_rsc_7_21_adra, xt_rsc_7_21_da, xt_rsc_7_21_wea, xt_rsc_7_21_qa, xt_rsc_triosy_7_21_lz,
      xt_rsc_7_22_adra, xt_rsc_7_22_da, xt_rsc_7_22_wea, xt_rsc_7_22_qa, xt_rsc_triosy_7_22_lz,
      xt_rsc_7_23_adra, xt_rsc_7_23_da, xt_rsc_7_23_wea, xt_rsc_7_23_qa, xt_rsc_triosy_7_23_lz,
      xt_rsc_7_24_adra, xt_rsc_7_24_da, xt_rsc_7_24_wea, xt_rsc_7_24_qa, xt_rsc_triosy_7_24_lz,
      xt_rsc_7_25_adra, xt_rsc_7_25_da, xt_rsc_7_25_wea, xt_rsc_7_25_qa, xt_rsc_triosy_7_25_lz,
      xt_rsc_7_26_adra, xt_rsc_7_26_da, xt_rsc_7_26_wea, xt_rsc_7_26_qa, xt_rsc_triosy_7_26_lz,
      xt_rsc_7_27_adra, xt_rsc_7_27_da, xt_rsc_7_27_wea, xt_rsc_7_27_qa, xt_rsc_triosy_7_27_lz,
      xt_rsc_7_28_adra, xt_rsc_7_28_da, xt_rsc_7_28_wea, xt_rsc_7_28_qa, xt_rsc_triosy_7_28_lz,
      xt_rsc_7_29_adra, xt_rsc_7_29_da, xt_rsc_7_29_wea, xt_rsc_7_29_qa, xt_rsc_triosy_7_29_lz,
      xt_rsc_7_30_adra, xt_rsc_7_30_da, xt_rsc_7_30_wea, xt_rsc_7_30_qa, xt_rsc_triosy_7_30_lz,
      xt_rsc_7_31_adra, xt_rsc_7_31_da, xt_rsc_7_31_wea, xt_rsc_7_31_qa, xt_rsc_triosy_7_31_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz, twiddle_rsc_0_0_adra,
      twiddle_rsc_0_0_da, twiddle_rsc_0_0_wea, twiddle_rsc_0_0_qa, twiddle_rsc_0_0_adrb,
      twiddle_rsc_0_0_db, twiddle_rsc_0_0_web, twiddle_rsc_0_0_qb, twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_0_1_adra, twiddle_rsc_0_1_da, twiddle_rsc_0_1_wea, twiddle_rsc_0_1_qa,
      twiddle_rsc_0_1_adrb, twiddle_rsc_0_1_db, twiddle_rsc_0_1_web, twiddle_rsc_0_1_qb,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_0_2_adra, twiddle_rsc_0_2_da, twiddle_rsc_0_2_wea,
      twiddle_rsc_0_2_qa, twiddle_rsc_0_2_adrb, twiddle_rsc_0_2_db, twiddle_rsc_0_2_web,
      twiddle_rsc_0_2_qb, twiddle_rsc_triosy_0_2_lz, twiddle_rsc_0_3_adra, twiddle_rsc_0_3_da,
      twiddle_rsc_0_3_wea, twiddle_rsc_0_3_qa, twiddle_rsc_0_3_adrb, twiddle_rsc_0_3_db,
      twiddle_rsc_0_3_web, twiddle_rsc_0_3_qb, twiddle_rsc_triosy_0_3_lz, twiddle_rsc_0_4_adra,
      twiddle_rsc_0_4_da, twiddle_rsc_0_4_wea, twiddle_rsc_0_4_qa, twiddle_rsc_0_4_adrb,
      twiddle_rsc_0_4_db, twiddle_rsc_0_4_web, twiddle_rsc_0_4_qb, twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_0_5_adra, twiddle_rsc_0_5_da, twiddle_rsc_0_5_wea, twiddle_rsc_0_5_qa,
      twiddle_rsc_0_5_adrb, twiddle_rsc_0_5_db, twiddle_rsc_0_5_web, twiddle_rsc_0_5_qb,
      twiddle_rsc_triosy_0_5_lz, twiddle_rsc_0_6_adra, twiddle_rsc_0_6_da, twiddle_rsc_0_6_wea,
      twiddle_rsc_0_6_qa, twiddle_rsc_0_6_adrb, twiddle_rsc_0_6_db, twiddle_rsc_0_6_web,
      twiddle_rsc_0_6_qb, twiddle_rsc_triosy_0_6_lz, twiddle_rsc_0_7_adra, twiddle_rsc_0_7_da,
      twiddle_rsc_0_7_wea, twiddle_rsc_0_7_qa, twiddle_rsc_0_7_adrb, twiddle_rsc_0_7_db,
      twiddle_rsc_0_7_web, twiddle_rsc_0_7_qb, twiddle_rsc_triosy_0_7_lz, twiddle_rsc_0_8_adra,
      twiddle_rsc_0_8_da, twiddle_rsc_0_8_wea, twiddle_rsc_0_8_qa, twiddle_rsc_0_8_adrb,
      twiddle_rsc_0_8_db, twiddle_rsc_0_8_web, twiddle_rsc_0_8_qb, twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_0_9_adra, twiddle_rsc_0_9_da, twiddle_rsc_0_9_wea, twiddle_rsc_0_9_qa,
      twiddle_rsc_0_9_adrb, twiddle_rsc_0_9_db, twiddle_rsc_0_9_web, twiddle_rsc_0_9_qb,
      twiddle_rsc_triosy_0_9_lz, twiddle_rsc_0_10_adra, twiddle_rsc_0_10_da, twiddle_rsc_0_10_wea,
      twiddle_rsc_0_10_qa, twiddle_rsc_0_10_adrb, twiddle_rsc_0_10_db, twiddle_rsc_0_10_web,
      twiddle_rsc_0_10_qb, twiddle_rsc_triosy_0_10_lz, twiddle_rsc_0_11_adra, twiddle_rsc_0_11_da,
      twiddle_rsc_0_11_wea, twiddle_rsc_0_11_qa, twiddle_rsc_0_11_adrb, twiddle_rsc_0_11_db,
      twiddle_rsc_0_11_web, twiddle_rsc_0_11_qb, twiddle_rsc_triosy_0_11_lz, twiddle_rsc_0_12_adra,
      twiddle_rsc_0_12_da, twiddle_rsc_0_12_wea, twiddle_rsc_0_12_qa, twiddle_rsc_0_12_adrb,
      twiddle_rsc_0_12_db, twiddle_rsc_0_12_web, twiddle_rsc_0_12_qb, twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_0_13_adra, twiddle_rsc_0_13_da, twiddle_rsc_0_13_wea, twiddle_rsc_0_13_qa,
      twiddle_rsc_0_13_adrb, twiddle_rsc_0_13_db, twiddle_rsc_0_13_web, twiddle_rsc_0_13_qb,
      twiddle_rsc_triosy_0_13_lz, twiddle_rsc_0_14_adra, twiddle_rsc_0_14_da, twiddle_rsc_0_14_wea,
      twiddle_rsc_0_14_qa, twiddle_rsc_0_14_adrb, twiddle_rsc_0_14_db, twiddle_rsc_0_14_web,
      twiddle_rsc_0_14_qb, twiddle_rsc_triosy_0_14_lz, twiddle_rsc_0_15_adra, twiddle_rsc_0_15_da,
      twiddle_rsc_0_15_wea, twiddle_rsc_0_15_qa, twiddle_rsc_0_15_adrb, twiddle_rsc_0_15_db,
      twiddle_rsc_0_15_web, twiddle_rsc_0_15_qb, twiddle_rsc_triosy_0_15_lz, twiddle_h_rsc_0_0_adra,
      twiddle_h_rsc_0_0_da, twiddle_h_rsc_0_0_wea, twiddle_h_rsc_0_0_qa, twiddle_h_rsc_0_0_adrb,
      twiddle_h_rsc_0_0_db, twiddle_h_rsc_0_0_web, twiddle_h_rsc_0_0_qb, twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_0_1_adra, twiddle_h_rsc_0_1_da, twiddle_h_rsc_0_1_wea, twiddle_h_rsc_0_1_qa,
      twiddle_h_rsc_0_1_adrb, twiddle_h_rsc_0_1_db, twiddle_h_rsc_0_1_web, twiddle_h_rsc_0_1_qb,
      twiddle_h_rsc_triosy_0_1_lz, twiddle_h_rsc_0_2_adra, twiddle_h_rsc_0_2_da,
      twiddle_h_rsc_0_2_wea, twiddle_h_rsc_0_2_qa, twiddle_h_rsc_0_2_adrb, twiddle_h_rsc_0_2_db,
      twiddle_h_rsc_0_2_web, twiddle_h_rsc_0_2_qb, twiddle_h_rsc_triosy_0_2_lz, twiddle_h_rsc_0_3_adra,
      twiddle_h_rsc_0_3_da, twiddle_h_rsc_0_3_wea, twiddle_h_rsc_0_3_qa, twiddle_h_rsc_0_3_adrb,
      twiddle_h_rsc_0_3_db, twiddle_h_rsc_0_3_web, twiddle_h_rsc_0_3_qb, twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_0_4_adra, twiddle_h_rsc_0_4_da, twiddle_h_rsc_0_4_wea, twiddle_h_rsc_0_4_qa,
      twiddle_h_rsc_0_4_adrb, twiddle_h_rsc_0_4_db, twiddle_h_rsc_0_4_web, twiddle_h_rsc_0_4_qb,
      twiddle_h_rsc_triosy_0_4_lz, twiddle_h_rsc_0_5_adra, twiddle_h_rsc_0_5_da,
      twiddle_h_rsc_0_5_wea, twiddle_h_rsc_0_5_qa, twiddle_h_rsc_0_5_adrb, twiddle_h_rsc_0_5_db,
      twiddle_h_rsc_0_5_web, twiddle_h_rsc_0_5_qb, twiddle_h_rsc_triosy_0_5_lz, twiddle_h_rsc_0_6_adra,
      twiddle_h_rsc_0_6_da, twiddle_h_rsc_0_6_wea, twiddle_h_rsc_0_6_qa, twiddle_h_rsc_0_6_adrb,
      twiddle_h_rsc_0_6_db, twiddle_h_rsc_0_6_web, twiddle_h_rsc_0_6_qb, twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_0_7_adra, twiddle_h_rsc_0_7_da, twiddle_h_rsc_0_7_wea, twiddle_h_rsc_0_7_qa,
      twiddle_h_rsc_0_7_adrb, twiddle_h_rsc_0_7_db, twiddle_h_rsc_0_7_web, twiddle_h_rsc_0_7_qb,
      twiddle_h_rsc_triosy_0_7_lz, twiddle_h_rsc_0_8_adra, twiddle_h_rsc_0_8_da,
      twiddle_h_rsc_0_8_wea, twiddle_h_rsc_0_8_qa, twiddle_h_rsc_0_8_adrb, twiddle_h_rsc_0_8_db,
      twiddle_h_rsc_0_8_web, twiddle_h_rsc_0_8_qb, twiddle_h_rsc_triosy_0_8_lz, twiddle_h_rsc_0_9_adra,
      twiddle_h_rsc_0_9_da, twiddle_h_rsc_0_9_wea, twiddle_h_rsc_0_9_qa, twiddle_h_rsc_0_9_adrb,
      twiddle_h_rsc_0_9_db, twiddle_h_rsc_0_9_web, twiddle_h_rsc_0_9_qb, twiddle_h_rsc_triosy_0_9_lz,
      twiddle_h_rsc_0_10_adra, twiddle_h_rsc_0_10_da, twiddle_h_rsc_0_10_wea, twiddle_h_rsc_0_10_qa,
      twiddle_h_rsc_0_10_adrb, twiddle_h_rsc_0_10_db, twiddle_h_rsc_0_10_web, twiddle_h_rsc_0_10_qb,
      twiddle_h_rsc_triosy_0_10_lz, twiddle_h_rsc_0_11_adra, twiddle_h_rsc_0_11_da,
      twiddle_h_rsc_0_11_wea, twiddle_h_rsc_0_11_qa, twiddle_h_rsc_0_11_adrb, twiddle_h_rsc_0_11_db,
      twiddle_h_rsc_0_11_web, twiddle_h_rsc_0_11_qb, twiddle_h_rsc_triosy_0_11_lz,
      twiddle_h_rsc_0_12_adra, twiddle_h_rsc_0_12_da, twiddle_h_rsc_0_12_wea, twiddle_h_rsc_0_12_qa,
      twiddle_h_rsc_0_12_adrb, twiddle_h_rsc_0_12_db, twiddle_h_rsc_0_12_web, twiddle_h_rsc_0_12_qb,
      twiddle_h_rsc_triosy_0_12_lz, twiddle_h_rsc_0_13_adra, twiddle_h_rsc_0_13_da,
      twiddle_h_rsc_0_13_wea, twiddle_h_rsc_0_13_qa, twiddle_h_rsc_0_13_adrb, twiddle_h_rsc_0_13_db,
      twiddle_h_rsc_0_13_web, twiddle_h_rsc_0_13_qb, twiddle_h_rsc_triosy_0_13_lz,
      twiddle_h_rsc_0_14_adra, twiddle_h_rsc_0_14_da, twiddle_h_rsc_0_14_wea, twiddle_h_rsc_0_14_qa,
      twiddle_h_rsc_0_14_adrb, twiddle_h_rsc_0_14_db, twiddle_h_rsc_0_14_web, twiddle_h_rsc_0_14_qb,
      twiddle_h_rsc_triosy_0_14_lz, twiddle_h_rsc_0_15_adra, twiddle_h_rsc_0_15_da,
      twiddle_h_rsc_0_15_wea, twiddle_h_rsc_0_15_qa, twiddle_h_rsc_0_15_adrb, twiddle_h_rsc_0_15_db,
      twiddle_h_rsc_0_15_web, twiddle_h_rsc_0_15_qb, twiddle_h_rsc_triosy_0_15_lz
);
  input clk;
  input rst;
  output [3:0] xt_rsc_0_0_adra;
  output [31:0] xt_rsc_0_0_da;
  output xt_rsc_0_0_wea;
  input [31:0] xt_rsc_0_0_qa;
  output xt_rsc_triosy_0_0_lz;
  output [3:0] xt_rsc_0_1_adra;
  output [31:0] xt_rsc_0_1_da;
  output xt_rsc_0_1_wea;
  input [31:0] xt_rsc_0_1_qa;
  output xt_rsc_triosy_0_1_lz;
  output [3:0] xt_rsc_0_2_adra;
  output [31:0] xt_rsc_0_2_da;
  output xt_rsc_0_2_wea;
  input [31:0] xt_rsc_0_2_qa;
  output xt_rsc_triosy_0_2_lz;
  output [3:0] xt_rsc_0_3_adra;
  output [31:0] xt_rsc_0_3_da;
  output xt_rsc_0_3_wea;
  input [31:0] xt_rsc_0_3_qa;
  output xt_rsc_triosy_0_3_lz;
  output [3:0] xt_rsc_0_4_adra;
  output [31:0] xt_rsc_0_4_da;
  output xt_rsc_0_4_wea;
  input [31:0] xt_rsc_0_4_qa;
  output xt_rsc_triosy_0_4_lz;
  output [3:0] xt_rsc_0_5_adra;
  output [31:0] xt_rsc_0_5_da;
  output xt_rsc_0_5_wea;
  input [31:0] xt_rsc_0_5_qa;
  output xt_rsc_triosy_0_5_lz;
  output [3:0] xt_rsc_0_6_adra;
  output [31:0] xt_rsc_0_6_da;
  output xt_rsc_0_6_wea;
  input [31:0] xt_rsc_0_6_qa;
  output xt_rsc_triosy_0_6_lz;
  output [3:0] xt_rsc_0_7_adra;
  output [31:0] xt_rsc_0_7_da;
  output xt_rsc_0_7_wea;
  input [31:0] xt_rsc_0_7_qa;
  output xt_rsc_triosy_0_7_lz;
  output [3:0] xt_rsc_0_8_adra;
  output [31:0] xt_rsc_0_8_da;
  output xt_rsc_0_8_wea;
  input [31:0] xt_rsc_0_8_qa;
  output xt_rsc_triosy_0_8_lz;
  output [3:0] xt_rsc_0_9_adra;
  output [31:0] xt_rsc_0_9_da;
  output xt_rsc_0_9_wea;
  input [31:0] xt_rsc_0_9_qa;
  output xt_rsc_triosy_0_9_lz;
  output [3:0] xt_rsc_0_10_adra;
  output [31:0] xt_rsc_0_10_da;
  output xt_rsc_0_10_wea;
  input [31:0] xt_rsc_0_10_qa;
  output xt_rsc_triosy_0_10_lz;
  output [3:0] xt_rsc_0_11_adra;
  output [31:0] xt_rsc_0_11_da;
  output xt_rsc_0_11_wea;
  input [31:0] xt_rsc_0_11_qa;
  output xt_rsc_triosy_0_11_lz;
  output [3:0] xt_rsc_0_12_adra;
  output [31:0] xt_rsc_0_12_da;
  output xt_rsc_0_12_wea;
  input [31:0] xt_rsc_0_12_qa;
  output xt_rsc_triosy_0_12_lz;
  output [3:0] xt_rsc_0_13_adra;
  output [31:0] xt_rsc_0_13_da;
  output xt_rsc_0_13_wea;
  input [31:0] xt_rsc_0_13_qa;
  output xt_rsc_triosy_0_13_lz;
  output [3:0] xt_rsc_0_14_adra;
  output [31:0] xt_rsc_0_14_da;
  output xt_rsc_0_14_wea;
  input [31:0] xt_rsc_0_14_qa;
  output xt_rsc_triosy_0_14_lz;
  output [3:0] xt_rsc_0_15_adra;
  output [31:0] xt_rsc_0_15_da;
  output xt_rsc_0_15_wea;
  input [31:0] xt_rsc_0_15_qa;
  output xt_rsc_triosy_0_15_lz;
  output [3:0] xt_rsc_0_16_adra;
  output [31:0] xt_rsc_0_16_da;
  output xt_rsc_0_16_wea;
  input [31:0] xt_rsc_0_16_qa;
  output xt_rsc_triosy_0_16_lz;
  output [3:0] xt_rsc_0_17_adra;
  output [31:0] xt_rsc_0_17_da;
  output xt_rsc_0_17_wea;
  input [31:0] xt_rsc_0_17_qa;
  output xt_rsc_triosy_0_17_lz;
  output [3:0] xt_rsc_0_18_adra;
  output [31:0] xt_rsc_0_18_da;
  output xt_rsc_0_18_wea;
  input [31:0] xt_rsc_0_18_qa;
  output xt_rsc_triosy_0_18_lz;
  output [3:0] xt_rsc_0_19_adra;
  output [31:0] xt_rsc_0_19_da;
  output xt_rsc_0_19_wea;
  input [31:0] xt_rsc_0_19_qa;
  output xt_rsc_triosy_0_19_lz;
  output [3:0] xt_rsc_0_20_adra;
  output [31:0] xt_rsc_0_20_da;
  output xt_rsc_0_20_wea;
  input [31:0] xt_rsc_0_20_qa;
  output xt_rsc_triosy_0_20_lz;
  output [3:0] xt_rsc_0_21_adra;
  output [31:0] xt_rsc_0_21_da;
  output xt_rsc_0_21_wea;
  input [31:0] xt_rsc_0_21_qa;
  output xt_rsc_triosy_0_21_lz;
  output [3:0] xt_rsc_0_22_adra;
  output [31:0] xt_rsc_0_22_da;
  output xt_rsc_0_22_wea;
  input [31:0] xt_rsc_0_22_qa;
  output xt_rsc_triosy_0_22_lz;
  output [3:0] xt_rsc_0_23_adra;
  output [31:0] xt_rsc_0_23_da;
  output xt_rsc_0_23_wea;
  input [31:0] xt_rsc_0_23_qa;
  output xt_rsc_triosy_0_23_lz;
  output [3:0] xt_rsc_0_24_adra;
  output [31:0] xt_rsc_0_24_da;
  output xt_rsc_0_24_wea;
  input [31:0] xt_rsc_0_24_qa;
  output xt_rsc_triosy_0_24_lz;
  output [3:0] xt_rsc_0_25_adra;
  output [31:0] xt_rsc_0_25_da;
  output xt_rsc_0_25_wea;
  input [31:0] xt_rsc_0_25_qa;
  output xt_rsc_triosy_0_25_lz;
  output [3:0] xt_rsc_0_26_adra;
  output [31:0] xt_rsc_0_26_da;
  output xt_rsc_0_26_wea;
  input [31:0] xt_rsc_0_26_qa;
  output xt_rsc_triosy_0_26_lz;
  output [3:0] xt_rsc_0_27_adra;
  output [31:0] xt_rsc_0_27_da;
  output xt_rsc_0_27_wea;
  input [31:0] xt_rsc_0_27_qa;
  output xt_rsc_triosy_0_27_lz;
  output [3:0] xt_rsc_0_28_adra;
  output [31:0] xt_rsc_0_28_da;
  output xt_rsc_0_28_wea;
  input [31:0] xt_rsc_0_28_qa;
  output xt_rsc_triosy_0_28_lz;
  output [3:0] xt_rsc_0_29_adra;
  output [31:0] xt_rsc_0_29_da;
  output xt_rsc_0_29_wea;
  input [31:0] xt_rsc_0_29_qa;
  output xt_rsc_triosy_0_29_lz;
  output [3:0] xt_rsc_0_30_adra;
  output [31:0] xt_rsc_0_30_da;
  output xt_rsc_0_30_wea;
  input [31:0] xt_rsc_0_30_qa;
  output xt_rsc_triosy_0_30_lz;
  output [3:0] xt_rsc_0_31_adra;
  output [31:0] xt_rsc_0_31_da;
  output xt_rsc_0_31_wea;
  input [31:0] xt_rsc_0_31_qa;
  output xt_rsc_triosy_0_31_lz;
  output [3:0] xt_rsc_1_0_adra;
  output [31:0] xt_rsc_1_0_da;
  output xt_rsc_1_0_wea;
  input [31:0] xt_rsc_1_0_qa;
  output xt_rsc_triosy_1_0_lz;
  output [3:0] xt_rsc_1_1_adra;
  output [31:0] xt_rsc_1_1_da;
  output xt_rsc_1_1_wea;
  input [31:0] xt_rsc_1_1_qa;
  output xt_rsc_triosy_1_1_lz;
  output [3:0] xt_rsc_1_2_adra;
  output [31:0] xt_rsc_1_2_da;
  output xt_rsc_1_2_wea;
  input [31:0] xt_rsc_1_2_qa;
  output xt_rsc_triosy_1_2_lz;
  output [3:0] xt_rsc_1_3_adra;
  output [31:0] xt_rsc_1_3_da;
  output xt_rsc_1_3_wea;
  input [31:0] xt_rsc_1_3_qa;
  output xt_rsc_triosy_1_3_lz;
  output [3:0] xt_rsc_1_4_adra;
  output [31:0] xt_rsc_1_4_da;
  output xt_rsc_1_4_wea;
  input [31:0] xt_rsc_1_4_qa;
  output xt_rsc_triosy_1_4_lz;
  output [3:0] xt_rsc_1_5_adra;
  output [31:0] xt_rsc_1_5_da;
  output xt_rsc_1_5_wea;
  input [31:0] xt_rsc_1_5_qa;
  output xt_rsc_triosy_1_5_lz;
  output [3:0] xt_rsc_1_6_adra;
  output [31:0] xt_rsc_1_6_da;
  output xt_rsc_1_6_wea;
  input [31:0] xt_rsc_1_6_qa;
  output xt_rsc_triosy_1_6_lz;
  output [3:0] xt_rsc_1_7_adra;
  output [31:0] xt_rsc_1_7_da;
  output xt_rsc_1_7_wea;
  input [31:0] xt_rsc_1_7_qa;
  output xt_rsc_triosy_1_7_lz;
  output [3:0] xt_rsc_1_8_adra;
  output [31:0] xt_rsc_1_8_da;
  output xt_rsc_1_8_wea;
  input [31:0] xt_rsc_1_8_qa;
  output xt_rsc_triosy_1_8_lz;
  output [3:0] xt_rsc_1_9_adra;
  output [31:0] xt_rsc_1_9_da;
  output xt_rsc_1_9_wea;
  input [31:0] xt_rsc_1_9_qa;
  output xt_rsc_triosy_1_9_lz;
  output [3:0] xt_rsc_1_10_adra;
  output [31:0] xt_rsc_1_10_da;
  output xt_rsc_1_10_wea;
  input [31:0] xt_rsc_1_10_qa;
  output xt_rsc_triosy_1_10_lz;
  output [3:0] xt_rsc_1_11_adra;
  output [31:0] xt_rsc_1_11_da;
  output xt_rsc_1_11_wea;
  input [31:0] xt_rsc_1_11_qa;
  output xt_rsc_triosy_1_11_lz;
  output [3:0] xt_rsc_1_12_adra;
  output [31:0] xt_rsc_1_12_da;
  output xt_rsc_1_12_wea;
  input [31:0] xt_rsc_1_12_qa;
  output xt_rsc_triosy_1_12_lz;
  output [3:0] xt_rsc_1_13_adra;
  output [31:0] xt_rsc_1_13_da;
  output xt_rsc_1_13_wea;
  input [31:0] xt_rsc_1_13_qa;
  output xt_rsc_triosy_1_13_lz;
  output [3:0] xt_rsc_1_14_adra;
  output [31:0] xt_rsc_1_14_da;
  output xt_rsc_1_14_wea;
  input [31:0] xt_rsc_1_14_qa;
  output xt_rsc_triosy_1_14_lz;
  output [3:0] xt_rsc_1_15_adra;
  output [31:0] xt_rsc_1_15_da;
  output xt_rsc_1_15_wea;
  input [31:0] xt_rsc_1_15_qa;
  output xt_rsc_triosy_1_15_lz;
  output [3:0] xt_rsc_1_16_adra;
  output [31:0] xt_rsc_1_16_da;
  output xt_rsc_1_16_wea;
  input [31:0] xt_rsc_1_16_qa;
  output xt_rsc_triosy_1_16_lz;
  output [3:0] xt_rsc_1_17_adra;
  output [31:0] xt_rsc_1_17_da;
  output xt_rsc_1_17_wea;
  input [31:0] xt_rsc_1_17_qa;
  output xt_rsc_triosy_1_17_lz;
  output [3:0] xt_rsc_1_18_adra;
  output [31:0] xt_rsc_1_18_da;
  output xt_rsc_1_18_wea;
  input [31:0] xt_rsc_1_18_qa;
  output xt_rsc_triosy_1_18_lz;
  output [3:0] xt_rsc_1_19_adra;
  output [31:0] xt_rsc_1_19_da;
  output xt_rsc_1_19_wea;
  input [31:0] xt_rsc_1_19_qa;
  output xt_rsc_triosy_1_19_lz;
  output [3:0] xt_rsc_1_20_adra;
  output [31:0] xt_rsc_1_20_da;
  output xt_rsc_1_20_wea;
  input [31:0] xt_rsc_1_20_qa;
  output xt_rsc_triosy_1_20_lz;
  output [3:0] xt_rsc_1_21_adra;
  output [31:0] xt_rsc_1_21_da;
  output xt_rsc_1_21_wea;
  input [31:0] xt_rsc_1_21_qa;
  output xt_rsc_triosy_1_21_lz;
  output [3:0] xt_rsc_1_22_adra;
  output [31:0] xt_rsc_1_22_da;
  output xt_rsc_1_22_wea;
  input [31:0] xt_rsc_1_22_qa;
  output xt_rsc_triosy_1_22_lz;
  output [3:0] xt_rsc_1_23_adra;
  output [31:0] xt_rsc_1_23_da;
  output xt_rsc_1_23_wea;
  input [31:0] xt_rsc_1_23_qa;
  output xt_rsc_triosy_1_23_lz;
  output [3:0] xt_rsc_1_24_adra;
  output [31:0] xt_rsc_1_24_da;
  output xt_rsc_1_24_wea;
  input [31:0] xt_rsc_1_24_qa;
  output xt_rsc_triosy_1_24_lz;
  output [3:0] xt_rsc_1_25_adra;
  output [31:0] xt_rsc_1_25_da;
  output xt_rsc_1_25_wea;
  input [31:0] xt_rsc_1_25_qa;
  output xt_rsc_triosy_1_25_lz;
  output [3:0] xt_rsc_1_26_adra;
  output [31:0] xt_rsc_1_26_da;
  output xt_rsc_1_26_wea;
  input [31:0] xt_rsc_1_26_qa;
  output xt_rsc_triosy_1_26_lz;
  output [3:0] xt_rsc_1_27_adra;
  output [31:0] xt_rsc_1_27_da;
  output xt_rsc_1_27_wea;
  input [31:0] xt_rsc_1_27_qa;
  output xt_rsc_triosy_1_27_lz;
  output [3:0] xt_rsc_1_28_adra;
  output [31:0] xt_rsc_1_28_da;
  output xt_rsc_1_28_wea;
  input [31:0] xt_rsc_1_28_qa;
  output xt_rsc_triosy_1_28_lz;
  output [3:0] xt_rsc_1_29_adra;
  output [31:0] xt_rsc_1_29_da;
  output xt_rsc_1_29_wea;
  input [31:0] xt_rsc_1_29_qa;
  output xt_rsc_triosy_1_29_lz;
  output [3:0] xt_rsc_1_30_adra;
  output [31:0] xt_rsc_1_30_da;
  output xt_rsc_1_30_wea;
  input [31:0] xt_rsc_1_30_qa;
  output xt_rsc_triosy_1_30_lz;
  output [3:0] xt_rsc_1_31_adra;
  output [31:0] xt_rsc_1_31_da;
  output xt_rsc_1_31_wea;
  input [31:0] xt_rsc_1_31_qa;
  output xt_rsc_triosy_1_31_lz;
  output [3:0] xt_rsc_2_0_adra;
  output [31:0] xt_rsc_2_0_da;
  output xt_rsc_2_0_wea;
  input [31:0] xt_rsc_2_0_qa;
  output xt_rsc_triosy_2_0_lz;
  output [3:0] xt_rsc_2_1_adra;
  output [31:0] xt_rsc_2_1_da;
  output xt_rsc_2_1_wea;
  input [31:0] xt_rsc_2_1_qa;
  output xt_rsc_triosy_2_1_lz;
  output [3:0] xt_rsc_2_2_adra;
  output [31:0] xt_rsc_2_2_da;
  output xt_rsc_2_2_wea;
  input [31:0] xt_rsc_2_2_qa;
  output xt_rsc_triosy_2_2_lz;
  output [3:0] xt_rsc_2_3_adra;
  output [31:0] xt_rsc_2_3_da;
  output xt_rsc_2_3_wea;
  input [31:0] xt_rsc_2_3_qa;
  output xt_rsc_triosy_2_3_lz;
  output [3:0] xt_rsc_2_4_adra;
  output [31:0] xt_rsc_2_4_da;
  output xt_rsc_2_4_wea;
  input [31:0] xt_rsc_2_4_qa;
  output xt_rsc_triosy_2_4_lz;
  output [3:0] xt_rsc_2_5_adra;
  output [31:0] xt_rsc_2_5_da;
  output xt_rsc_2_5_wea;
  input [31:0] xt_rsc_2_5_qa;
  output xt_rsc_triosy_2_5_lz;
  output [3:0] xt_rsc_2_6_adra;
  output [31:0] xt_rsc_2_6_da;
  output xt_rsc_2_6_wea;
  input [31:0] xt_rsc_2_6_qa;
  output xt_rsc_triosy_2_6_lz;
  output [3:0] xt_rsc_2_7_adra;
  output [31:0] xt_rsc_2_7_da;
  output xt_rsc_2_7_wea;
  input [31:0] xt_rsc_2_7_qa;
  output xt_rsc_triosy_2_7_lz;
  output [3:0] xt_rsc_2_8_adra;
  output [31:0] xt_rsc_2_8_da;
  output xt_rsc_2_8_wea;
  input [31:0] xt_rsc_2_8_qa;
  output xt_rsc_triosy_2_8_lz;
  output [3:0] xt_rsc_2_9_adra;
  output [31:0] xt_rsc_2_9_da;
  output xt_rsc_2_9_wea;
  input [31:0] xt_rsc_2_9_qa;
  output xt_rsc_triosy_2_9_lz;
  output [3:0] xt_rsc_2_10_adra;
  output [31:0] xt_rsc_2_10_da;
  output xt_rsc_2_10_wea;
  input [31:0] xt_rsc_2_10_qa;
  output xt_rsc_triosy_2_10_lz;
  output [3:0] xt_rsc_2_11_adra;
  output [31:0] xt_rsc_2_11_da;
  output xt_rsc_2_11_wea;
  input [31:0] xt_rsc_2_11_qa;
  output xt_rsc_triosy_2_11_lz;
  output [3:0] xt_rsc_2_12_adra;
  output [31:0] xt_rsc_2_12_da;
  output xt_rsc_2_12_wea;
  input [31:0] xt_rsc_2_12_qa;
  output xt_rsc_triosy_2_12_lz;
  output [3:0] xt_rsc_2_13_adra;
  output [31:0] xt_rsc_2_13_da;
  output xt_rsc_2_13_wea;
  input [31:0] xt_rsc_2_13_qa;
  output xt_rsc_triosy_2_13_lz;
  output [3:0] xt_rsc_2_14_adra;
  output [31:0] xt_rsc_2_14_da;
  output xt_rsc_2_14_wea;
  input [31:0] xt_rsc_2_14_qa;
  output xt_rsc_triosy_2_14_lz;
  output [3:0] xt_rsc_2_15_adra;
  output [31:0] xt_rsc_2_15_da;
  output xt_rsc_2_15_wea;
  input [31:0] xt_rsc_2_15_qa;
  output xt_rsc_triosy_2_15_lz;
  output [3:0] xt_rsc_2_16_adra;
  output [31:0] xt_rsc_2_16_da;
  output xt_rsc_2_16_wea;
  input [31:0] xt_rsc_2_16_qa;
  output xt_rsc_triosy_2_16_lz;
  output [3:0] xt_rsc_2_17_adra;
  output [31:0] xt_rsc_2_17_da;
  output xt_rsc_2_17_wea;
  input [31:0] xt_rsc_2_17_qa;
  output xt_rsc_triosy_2_17_lz;
  output [3:0] xt_rsc_2_18_adra;
  output [31:0] xt_rsc_2_18_da;
  output xt_rsc_2_18_wea;
  input [31:0] xt_rsc_2_18_qa;
  output xt_rsc_triosy_2_18_lz;
  output [3:0] xt_rsc_2_19_adra;
  output [31:0] xt_rsc_2_19_da;
  output xt_rsc_2_19_wea;
  input [31:0] xt_rsc_2_19_qa;
  output xt_rsc_triosy_2_19_lz;
  output [3:0] xt_rsc_2_20_adra;
  output [31:0] xt_rsc_2_20_da;
  output xt_rsc_2_20_wea;
  input [31:0] xt_rsc_2_20_qa;
  output xt_rsc_triosy_2_20_lz;
  output [3:0] xt_rsc_2_21_adra;
  output [31:0] xt_rsc_2_21_da;
  output xt_rsc_2_21_wea;
  input [31:0] xt_rsc_2_21_qa;
  output xt_rsc_triosy_2_21_lz;
  output [3:0] xt_rsc_2_22_adra;
  output [31:0] xt_rsc_2_22_da;
  output xt_rsc_2_22_wea;
  input [31:0] xt_rsc_2_22_qa;
  output xt_rsc_triosy_2_22_lz;
  output [3:0] xt_rsc_2_23_adra;
  output [31:0] xt_rsc_2_23_da;
  output xt_rsc_2_23_wea;
  input [31:0] xt_rsc_2_23_qa;
  output xt_rsc_triosy_2_23_lz;
  output [3:0] xt_rsc_2_24_adra;
  output [31:0] xt_rsc_2_24_da;
  output xt_rsc_2_24_wea;
  input [31:0] xt_rsc_2_24_qa;
  output xt_rsc_triosy_2_24_lz;
  output [3:0] xt_rsc_2_25_adra;
  output [31:0] xt_rsc_2_25_da;
  output xt_rsc_2_25_wea;
  input [31:0] xt_rsc_2_25_qa;
  output xt_rsc_triosy_2_25_lz;
  output [3:0] xt_rsc_2_26_adra;
  output [31:0] xt_rsc_2_26_da;
  output xt_rsc_2_26_wea;
  input [31:0] xt_rsc_2_26_qa;
  output xt_rsc_triosy_2_26_lz;
  output [3:0] xt_rsc_2_27_adra;
  output [31:0] xt_rsc_2_27_da;
  output xt_rsc_2_27_wea;
  input [31:0] xt_rsc_2_27_qa;
  output xt_rsc_triosy_2_27_lz;
  output [3:0] xt_rsc_2_28_adra;
  output [31:0] xt_rsc_2_28_da;
  output xt_rsc_2_28_wea;
  input [31:0] xt_rsc_2_28_qa;
  output xt_rsc_triosy_2_28_lz;
  output [3:0] xt_rsc_2_29_adra;
  output [31:0] xt_rsc_2_29_da;
  output xt_rsc_2_29_wea;
  input [31:0] xt_rsc_2_29_qa;
  output xt_rsc_triosy_2_29_lz;
  output [3:0] xt_rsc_2_30_adra;
  output [31:0] xt_rsc_2_30_da;
  output xt_rsc_2_30_wea;
  input [31:0] xt_rsc_2_30_qa;
  output xt_rsc_triosy_2_30_lz;
  output [3:0] xt_rsc_2_31_adra;
  output [31:0] xt_rsc_2_31_da;
  output xt_rsc_2_31_wea;
  input [31:0] xt_rsc_2_31_qa;
  output xt_rsc_triosy_2_31_lz;
  output [3:0] xt_rsc_3_0_adra;
  output [31:0] xt_rsc_3_0_da;
  output xt_rsc_3_0_wea;
  input [31:0] xt_rsc_3_0_qa;
  output xt_rsc_triosy_3_0_lz;
  output [3:0] xt_rsc_3_1_adra;
  output [31:0] xt_rsc_3_1_da;
  output xt_rsc_3_1_wea;
  input [31:0] xt_rsc_3_1_qa;
  output xt_rsc_triosy_3_1_lz;
  output [3:0] xt_rsc_3_2_adra;
  output [31:0] xt_rsc_3_2_da;
  output xt_rsc_3_2_wea;
  input [31:0] xt_rsc_3_2_qa;
  output xt_rsc_triosy_3_2_lz;
  output [3:0] xt_rsc_3_3_adra;
  output [31:0] xt_rsc_3_3_da;
  output xt_rsc_3_3_wea;
  input [31:0] xt_rsc_3_3_qa;
  output xt_rsc_triosy_3_3_lz;
  output [3:0] xt_rsc_3_4_adra;
  output [31:0] xt_rsc_3_4_da;
  output xt_rsc_3_4_wea;
  input [31:0] xt_rsc_3_4_qa;
  output xt_rsc_triosy_3_4_lz;
  output [3:0] xt_rsc_3_5_adra;
  output [31:0] xt_rsc_3_5_da;
  output xt_rsc_3_5_wea;
  input [31:0] xt_rsc_3_5_qa;
  output xt_rsc_triosy_3_5_lz;
  output [3:0] xt_rsc_3_6_adra;
  output [31:0] xt_rsc_3_6_da;
  output xt_rsc_3_6_wea;
  input [31:0] xt_rsc_3_6_qa;
  output xt_rsc_triosy_3_6_lz;
  output [3:0] xt_rsc_3_7_adra;
  output [31:0] xt_rsc_3_7_da;
  output xt_rsc_3_7_wea;
  input [31:0] xt_rsc_3_7_qa;
  output xt_rsc_triosy_3_7_lz;
  output [3:0] xt_rsc_3_8_adra;
  output [31:0] xt_rsc_3_8_da;
  output xt_rsc_3_8_wea;
  input [31:0] xt_rsc_3_8_qa;
  output xt_rsc_triosy_3_8_lz;
  output [3:0] xt_rsc_3_9_adra;
  output [31:0] xt_rsc_3_9_da;
  output xt_rsc_3_9_wea;
  input [31:0] xt_rsc_3_9_qa;
  output xt_rsc_triosy_3_9_lz;
  output [3:0] xt_rsc_3_10_adra;
  output [31:0] xt_rsc_3_10_da;
  output xt_rsc_3_10_wea;
  input [31:0] xt_rsc_3_10_qa;
  output xt_rsc_triosy_3_10_lz;
  output [3:0] xt_rsc_3_11_adra;
  output [31:0] xt_rsc_3_11_da;
  output xt_rsc_3_11_wea;
  input [31:0] xt_rsc_3_11_qa;
  output xt_rsc_triosy_3_11_lz;
  output [3:0] xt_rsc_3_12_adra;
  output [31:0] xt_rsc_3_12_da;
  output xt_rsc_3_12_wea;
  input [31:0] xt_rsc_3_12_qa;
  output xt_rsc_triosy_3_12_lz;
  output [3:0] xt_rsc_3_13_adra;
  output [31:0] xt_rsc_3_13_da;
  output xt_rsc_3_13_wea;
  input [31:0] xt_rsc_3_13_qa;
  output xt_rsc_triosy_3_13_lz;
  output [3:0] xt_rsc_3_14_adra;
  output [31:0] xt_rsc_3_14_da;
  output xt_rsc_3_14_wea;
  input [31:0] xt_rsc_3_14_qa;
  output xt_rsc_triosy_3_14_lz;
  output [3:0] xt_rsc_3_15_adra;
  output [31:0] xt_rsc_3_15_da;
  output xt_rsc_3_15_wea;
  input [31:0] xt_rsc_3_15_qa;
  output xt_rsc_triosy_3_15_lz;
  output [3:0] xt_rsc_3_16_adra;
  output [31:0] xt_rsc_3_16_da;
  output xt_rsc_3_16_wea;
  input [31:0] xt_rsc_3_16_qa;
  output xt_rsc_triosy_3_16_lz;
  output [3:0] xt_rsc_3_17_adra;
  output [31:0] xt_rsc_3_17_da;
  output xt_rsc_3_17_wea;
  input [31:0] xt_rsc_3_17_qa;
  output xt_rsc_triosy_3_17_lz;
  output [3:0] xt_rsc_3_18_adra;
  output [31:0] xt_rsc_3_18_da;
  output xt_rsc_3_18_wea;
  input [31:0] xt_rsc_3_18_qa;
  output xt_rsc_triosy_3_18_lz;
  output [3:0] xt_rsc_3_19_adra;
  output [31:0] xt_rsc_3_19_da;
  output xt_rsc_3_19_wea;
  input [31:0] xt_rsc_3_19_qa;
  output xt_rsc_triosy_3_19_lz;
  output [3:0] xt_rsc_3_20_adra;
  output [31:0] xt_rsc_3_20_da;
  output xt_rsc_3_20_wea;
  input [31:0] xt_rsc_3_20_qa;
  output xt_rsc_triosy_3_20_lz;
  output [3:0] xt_rsc_3_21_adra;
  output [31:0] xt_rsc_3_21_da;
  output xt_rsc_3_21_wea;
  input [31:0] xt_rsc_3_21_qa;
  output xt_rsc_triosy_3_21_lz;
  output [3:0] xt_rsc_3_22_adra;
  output [31:0] xt_rsc_3_22_da;
  output xt_rsc_3_22_wea;
  input [31:0] xt_rsc_3_22_qa;
  output xt_rsc_triosy_3_22_lz;
  output [3:0] xt_rsc_3_23_adra;
  output [31:0] xt_rsc_3_23_da;
  output xt_rsc_3_23_wea;
  input [31:0] xt_rsc_3_23_qa;
  output xt_rsc_triosy_3_23_lz;
  output [3:0] xt_rsc_3_24_adra;
  output [31:0] xt_rsc_3_24_da;
  output xt_rsc_3_24_wea;
  input [31:0] xt_rsc_3_24_qa;
  output xt_rsc_triosy_3_24_lz;
  output [3:0] xt_rsc_3_25_adra;
  output [31:0] xt_rsc_3_25_da;
  output xt_rsc_3_25_wea;
  input [31:0] xt_rsc_3_25_qa;
  output xt_rsc_triosy_3_25_lz;
  output [3:0] xt_rsc_3_26_adra;
  output [31:0] xt_rsc_3_26_da;
  output xt_rsc_3_26_wea;
  input [31:0] xt_rsc_3_26_qa;
  output xt_rsc_triosy_3_26_lz;
  output [3:0] xt_rsc_3_27_adra;
  output [31:0] xt_rsc_3_27_da;
  output xt_rsc_3_27_wea;
  input [31:0] xt_rsc_3_27_qa;
  output xt_rsc_triosy_3_27_lz;
  output [3:0] xt_rsc_3_28_adra;
  output [31:0] xt_rsc_3_28_da;
  output xt_rsc_3_28_wea;
  input [31:0] xt_rsc_3_28_qa;
  output xt_rsc_triosy_3_28_lz;
  output [3:0] xt_rsc_3_29_adra;
  output [31:0] xt_rsc_3_29_da;
  output xt_rsc_3_29_wea;
  input [31:0] xt_rsc_3_29_qa;
  output xt_rsc_triosy_3_29_lz;
  output [3:0] xt_rsc_3_30_adra;
  output [31:0] xt_rsc_3_30_da;
  output xt_rsc_3_30_wea;
  input [31:0] xt_rsc_3_30_qa;
  output xt_rsc_triosy_3_30_lz;
  output [3:0] xt_rsc_3_31_adra;
  output [31:0] xt_rsc_3_31_da;
  output xt_rsc_3_31_wea;
  input [31:0] xt_rsc_3_31_qa;
  output xt_rsc_triosy_3_31_lz;
  output [3:0] xt_rsc_4_0_adra;
  output [31:0] xt_rsc_4_0_da;
  output xt_rsc_4_0_wea;
  input [31:0] xt_rsc_4_0_qa;
  output xt_rsc_triosy_4_0_lz;
  output [3:0] xt_rsc_4_1_adra;
  output [31:0] xt_rsc_4_1_da;
  output xt_rsc_4_1_wea;
  input [31:0] xt_rsc_4_1_qa;
  output xt_rsc_triosy_4_1_lz;
  output [3:0] xt_rsc_4_2_adra;
  output [31:0] xt_rsc_4_2_da;
  output xt_rsc_4_2_wea;
  input [31:0] xt_rsc_4_2_qa;
  output xt_rsc_triosy_4_2_lz;
  output [3:0] xt_rsc_4_3_adra;
  output [31:0] xt_rsc_4_3_da;
  output xt_rsc_4_3_wea;
  input [31:0] xt_rsc_4_3_qa;
  output xt_rsc_triosy_4_3_lz;
  output [3:0] xt_rsc_4_4_adra;
  output [31:0] xt_rsc_4_4_da;
  output xt_rsc_4_4_wea;
  input [31:0] xt_rsc_4_4_qa;
  output xt_rsc_triosy_4_4_lz;
  output [3:0] xt_rsc_4_5_adra;
  output [31:0] xt_rsc_4_5_da;
  output xt_rsc_4_5_wea;
  input [31:0] xt_rsc_4_5_qa;
  output xt_rsc_triosy_4_5_lz;
  output [3:0] xt_rsc_4_6_adra;
  output [31:0] xt_rsc_4_6_da;
  output xt_rsc_4_6_wea;
  input [31:0] xt_rsc_4_6_qa;
  output xt_rsc_triosy_4_6_lz;
  output [3:0] xt_rsc_4_7_adra;
  output [31:0] xt_rsc_4_7_da;
  output xt_rsc_4_7_wea;
  input [31:0] xt_rsc_4_7_qa;
  output xt_rsc_triosy_4_7_lz;
  output [3:0] xt_rsc_4_8_adra;
  output [31:0] xt_rsc_4_8_da;
  output xt_rsc_4_8_wea;
  input [31:0] xt_rsc_4_8_qa;
  output xt_rsc_triosy_4_8_lz;
  output [3:0] xt_rsc_4_9_adra;
  output [31:0] xt_rsc_4_9_da;
  output xt_rsc_4_9_wea;
  input [31:0] xt_rsc_4_9_qa;
  output xt_rsc_triosy_4_9_lz;
  output [3:0] xt_rsc_4_10_adra;
  output [31:0] xt_rsc_4_10_da;
  output xt_rsc_4_10_wea;
  input [31:0] xt_rsc_4_10_qa;
  output xt_rsc_triosy_4_10_lz;
  output [3:0] xt_rsc_4_11_adra;
  output [31:0] xt_rsc_4_11_da;
  output xt_rsc_4_11_wea;
  input [31:0] xt_rsc_4_11_qa;
  output xt_rsc_triosy_4_11_lz;
  output [3:0] xt_rsc_4_12_adra;
  output [31:0] xt_rsc_4_12_da;
  output xt_rsc_4_12_wea;
  input [31:0] xt_rsc_4_12_qa;
  output xt_rsc_triosy_4_12_lz;
  output [3:0] xt_rsc_4_13_adra;
  output [31:0] xt_rsc_4_13_da;
  output xt_rsc_4_13_wea;
  input [31:0] xt_rsc_4_13_qa;
  output xt_rsc_triosy_4_13_lz;
  output [3:0] xt_rsc_4_14_adra;
  output [31:0] xt_rsc_4_14_da;
  output xt_rsc_4_14_wea;
  input [31:0] xt_rsc_4_14_qa;
  output xt_rsc_triosy_4_14_lz;
  output [3:0] xt_rsc_4_15_adra;
  output [31:0] xt_rsc_4_15_da;
  output xt_rsc_4_15_wea;
  input [31:0] xt_rsc_4_15_qa;
  output xt_rsc_triosy_4_15_lz;
  output [3:0] xt_rsc_4_16_adra;
  output [31:0] xt_rsc_4_16_da;
  output xt_rsc_4_16_wea;
  input [31:0] xt_rsc_4_16_qa;
  output xt_rsc_triosy_4_16_lz;
  output [3:0] xt_rsc_4_17_adra;
  output [31:0] xt_rsc_4_17_da;
  output xt_rsc_4_17_wea;
  input [31:0] xt_rsc_4_17_qa;
  output xt_rsc_triosy_4_17_lz;
  output [3:0] xt_rsc_4_18_adra;
  output [31:0] xt_rsc_4_18_da;
  output xt_rsc_4_18_wea;
  input [31:0] xt_rsc_4_18_qa;
  output xt_rsc_triosy_4_18_lz;
  output [3:0] xt_rsc_4_19_adra;
  output [31:0] xt_rsc_4_19_da;
  output xt_rsc_4_19_wea;
  input [31:0] xt_rsc_4_19_qa;
  output xt_rsc_triosy_4_19_lz;
  output [3:0] xt_rsc_4_20_adra;
  output [31:0] xt_rsc_4_20_da;
  output xt_rsc_4_20_wea;
  input [31:0] xt_rsc_4_20_qa;
  output xt_rsc_triosy_4_20_lz;
  output [3:0] xt_rsc_4_21_adra;
  output [31:0] xt_rsc_4_21_da;
  output xt_rsc_4_21_wea;
  input [31:0] xt_rsc_4_21_qa;
  output xt_rsc_triosy_4_21_lz;
  output [3:0] xt_rsc_4_22_adra;
  output [31:0] xt_rsc_4_22_da;
  output xt_rsc_4_22_wea;
  input [31:0] xt_rsc_4_22_qa;
  output xt_rsc_triosy_4_22_lz;
  output [3:0] xt_rsc_4_23_adra;
  output [31:0] xt_rsc_4_23_da;
  output xt_rsc_4_23_wea;
  input [31:0] xt_rsc_4_23_qa;
  output xt_rsc_triosy_4_23_lz;
  output [3:0] xt_rsc_4_24_adra;
  output [31:0] xt_rsc_4_24_da;
  output xt_rsc_4_24_wea;
  input [31:0] xt_rsc_4_24_qa;
  output xt_rsc_triosy_4_24_lz;
  output [3:0] xt_rsc_4_25_adra;
  output [31:0] xt_rsc_4_25_da;
  output xt_rsc_4_25_wea;
  input [31:0] xt_rsc_4_25_qa;
  output xt_rsc_triosy_4_25_lz;
  output [3:0] xt_rsc_4_26_adra;
  output [31:0] xt_rsc_4_26_da;
  output xt_rsc_4_26_wea;
  input [31:0] xt_rsc_4_26_qa;
  output xt_rsc_triosy_4_26_lz;
  output [3:0] xt_rsc_4_27_adra;
  output [31:0] xt_rsc_4_27_da;
  output xt_rsc_4_27_wea;
  input [31:0] xt_rsc_4_27_qa;
  output xt_rsc_triosy_4_27_lz;
  output [3:0] xt_rsc_4_28_adra;
  output [31:0] xt_rsc_4_28_da;
  output xt_rsc_4_28_wea;
  input [31:0] xt_rsc_4_28_qa;
  output xt_rsc_triosy_4_28_lz;
  output [3:0] xt_rsc_4_29_adra;
  output [31:0] xt_rsc_4_29_da;
  output xt_rsc_4_29_wea;
  input [31:0] xt_rsc_4_29_qa;
  output xt_rsc_triosy_4_29_lz;
  output [3:0] xt_rsc_4_30_adra;
  output [31:0] xt_rsc_4_30_da;
  output xt_rsc_4_30_wea;
  input [31:0] xt_rsc_4_30_qa;
  output xt_rsc_triosy_4_30_lz;
  output [3:0] xt_rsc_4_31_adra;
  output [31:0] xt_rsc_4_31_da;
  output xt_rsc_4_31_wea;
  input [31:0] xt_rsc_4_31_qa;
  output xt_rsc_triosy_4_31_lz;
  output [3:0] xt_rsc_5_0_adra;
  output [31:0] xt_rsc_5_0_da;
  output xt_rsc_5_0_wea;
  input [31:0] xt_rsc_5_0_qa;
  output xt_rsc_triosy_5_0_lz;
  output [3:0] xt_rsc_5_1_adra;
  output [31:0] xt_rsc_5_1_da;
  output xt_rsc_5_1_wea;
  input [31:0] xt_rsc_5_1_qa;
  output xt_rsc_triosy_5_1_lz;
  output [3:0] xt_rsc_5_2_adra;
  output [31:0] xt_rsc_5_2_da;
  output xt_rsc_5_2_wea;
  input [31:0] xt_rsc_5_2_qa;
  output xt_rsc_triosy_5_2_lz;
  output [3:0] xt_rsc_5_3_adra;
  output [31:0] xt_rsc_5_3_da;
  output xt_rsc_5_3_wea;
  input [31:0] xt_rsc_5_3_qa;
  output xt_rsc_triosy_5_3_lz;
  output [3:0] xt_rsc_5_4_adra;
  output [31:0] xt_rsc_5_4_da;
  output xt_rsc_5_4_wea;
  input [31:0] xt_rsc_5_4_qa;
  output xt_rsc_triosy_5_4_lz;
  output [3:0] xt_rsc_5_5_adra;
  output [31:0] xt_rsc_5_5_da;
  output xt_rsc_5_5_wea;
  input [31:0] xt_rsc_5_5_qa;
  output xt_rsc_triosy_5_5_lz;
  output [3:0] xt_rsc_5_6_adra;
  output [31:0] xt_rsc_5_6_da;
  output xt_rsc_5_6_wea;
  input [31:0] xt_rsc_5_6_qa;
  output xt_rsc_triosy_5_6_lz;
  output [3:0] xt_rsc_5_7_adra;
  output [31:0] xt_rsc_5_7_da;
  output xt_rsc_5_7_wea;
  input [31:0] xt_rsc_5_7_qa;
  output xt_rsc_triosy_5_7_lz;
  output [3:0] xt_rsc_5_8_adra;
  output [31:0] xt_rsc_5_8_da;
  output xt_rsc_5_8_wea;
  input [31:0] xt_rsc_5_8_qa;
  output xt_rsc_triosy_5_8_lz;
  output [3:0] xt_rsc_5_9_adra;
  output [31:0] xt_rsc_5_9_da;
  output xt_rsc_5_9_wea;
  input [31:0] xt_rsc_5_9_qa;
  output xt_rsc_triosy_5_9_lz;
  output [3:0] xt_rsc_5_10_adra;
  output [31:0] xt_rsc_5_10_da;
  output xt_rsc_5_10_wea;
  input [31:0] xt_rsc_5_10_qa;
  output xt_rsc_triosy_5_10_lz;
  output [3:0] xt_rsc_5_11_adra;
  output [31:0] xt_rsc_5_11_da;
  output xt_rsc_5_11_wea;
  input [31:0] xt_rsc_5_11_qa;
  output xt_rsc_triosy_5_11_lz;
  output [3:0] xt_rsc_5_12_adra;
  output [31:0] xt_rsc_5_12_da;
  output xt_rsc_5_12_wea;
  input [31:0] xt_rsc_5_12_qa;
  output xt_rsc_triosy_5_12_lz;
  output [3:0] xt_rsc_5_13_adra;
  output [31:0] xt_rsc_5_13_da;
  output xt_rsc_5_13_wea;
  input [31:0] xt_rsc_5_13_qa;
  output xt_rsc_triosy_5_13_lz;
  output [3:0] xt_rsc_5_14_adra;
  output [31:0] xt_rsc_5_14_da;
  output xt_rsc_5_14_wea;
  input [31:0] xt_rsc_5_14_qa;
  output xt_rsc_triosy_5_14_lz;
  output [3:0] xt_rsc_5_15_adra;
  output [31:0] xt_rsc_5_15_da;
  output xt_rsc_5_15_wea;
  input [31:0] xt_rsc_5_15_qa;
  output xt_rsc_triosy_5_15_lz;
  output [3:0] xt_rsc_5_16_adra;
  output [31:0] xt_rsc_5_16_da;
  output xt_rsc_5_16_wea;
  input [31:0] xt_rsc_5_16_qa;
  output xt_rsc_triosy_5_16_lz;
  output [3:0] xt_rsc_5_17_adra;
  output [31:0] xt_rsc_5_17_da;
  output xt_rsc_5_17_wea;
  input [31:0] xt_rsc_5_17_qa;
  output xt_rsc_triosy_5_17_lz;
  output [3:0] xt_rsc_5_18_adra;
  output [31:0] xt_rsc_5_18_da;
  output xt_rsc_5_18_wea;
  input [31:0] xt_rsc_5_18_qa;
  output xt_rsc_triosy_5_18_lz;
  output [3:0] xt_rsc_5_19_adra;
  output [31:0] xt_rsc_5_19_da;
  output xt_rsc_5_19_wea;
  input [31:0] xt_rsc_5_19_qa;
  output xt_rsc_triosy_5_19_lz;
  output [3:0] xt_rsc_5_20_adra;
  output [31:0] xt_rsc_5_20_da;
  output xt_rsc_5_20_wea;
  input [31:0] xt_rsc_5_20_qa;
  output xt_rsc_triosy_5_20_lz;
  output [3:0] xt_rsc_5_21_adra;
  output [31:0] xt_rsc_5_21_da;
  output xt_rsc_5_21_wea;
  input [31:0] xt_rsc_5_21_qa;
  output xt_rsc_triosy_5_21_lz;
  output [3:0] xt_rsc_5_22_adra;
  output [31:0] xt_rsc_5_22_da;
  output xt_rsc_5_22_wea;
  input [31:0] xt_rsc_5_22_qa;
  output xt_rsc_triosy_5_22_lz;
  output [3:0] xt_rsc_5_23_adra;
  output [31:0] xt_rsc_5_23_da;
  output xt_rsc_5_23_wea;
  input [31:0] xt_rsc_5_23_qa;
  output xt_rsc_triosy_5_23_lz;
  output [3:0] xt_rsc_5_24_adra;
  output [31:0] xt_rsc_5_24_da;
  output xt_rsc_5_24_wea;
  input [31:0] xt_rsc_5_24_qa;
  output xt_rsc_triosy_5_24_lz;
  output [3:0] xt_rsc_5_25_adra;
  output [31:0] xt_rsc_5_25_da;
  output xt_rsc_5_25_wea;
  input [31:0] xt_rsc_5_25_qa;
  output xt_rsc_triosy_5_25_lz;
  output [3:0] xt_rsc_5_26_adra;
  output [31:0] xt_rsc_5_26_da;
  output xt_rsc_5_26_wea;
  input [31:0] xt_rsc_5_26_qa;
  output xt_rsc_triosy_5_26_lz;
  output [3:0] xt_rsc_5_27_adra;
  output [31:0] xt_rsc_5_27_da;
  output xt_rsc_5_27_wea;
  input [31:0] xt_rsc_5_27_qa;
  output xt_rsc_triosy_5_27_lz;
  output [3:0] xt_rsc_5_28_adra;
  output [31:0] xt_rsc_5_28_da;
  output xt_rsc_5_28_wea;
  input [31:0] xt_rsc_5_28_qa;
  output xt_rsc_triosy_5_28_lz;
  output [3:0] xt_rsc_5_29_adra;
  output [31:0] xt_rsc_5_29_da;
  output xt_rsc_5_29_wea;
  input [31:0] xt_rsc_5_29_qa;
  output xt_rsc_triosy_5_29_lz;
  output [3:0] xt_rsc_5_30_adra;
  output [31:0] xt_rsc_5_30_da;
  output xt_rsc_5_30_wea;
  input [31:0] xt_rsc_5_30_qa;
  output xt_rsc_triosy_5_30_lz;
  output [3:0] xt_rsc_5_31_adra;
  output [31:0] xt_rsc_5_31_da;
  output xt_rsc_5_31_wea;
  input [31:0] xt_rsc_5_31_qa;
  output xt_rsc_triosy_5_31_lz;
  output [3:0] xt_rsc_6_0_adra;
  output [31:0] xt_rsc_6_0_da;
  output xt_rsc_6_0_wea;
  input [31:0] xt_rsc_6_0_qa;
  output xt_rsc_triosy_6_0_lz;
  output [3:0] xt_rsc_6_1_adra;
  output [31:0] xt_rsc_6_1_da;
  output xt_rsc_6_1_wea;
  input [31:0] xt_rsc_6_1_qa;
  output xt_rsc_triosy_6_1_lz;
  output [3:0] xt_rsc_6_2_adra;
  output [31:0] xt_rsc_6_2_da;
  output xt_rsc_6_2_wea;
  input [31:0] xt_rsc_6_2_qa;
  output xt_rsc_triosy_6_2_lz;
  output [3:0] xt_rsc_6_3_adra;
  output [31:0] xt_rsc_6_3_da;
  output xt_rsc_6_3_wea;
  input [31:0] xt_rsc_6_3_qa;
  output xt_rsc_triosy_6_3_lz;
  output [3:0] xt_rsc_6_4_adra;
  output [31:0] xt_rsc_6_4_da;
  output xt_rsc_6_4_wea;
  input [31:0] xt_rsc_6_4_qa;
  output xt_rsc_triosy_6_4_lz;
  output [3:0] xt_rsc_6_5_adra;
  output [31:0] xt_rsc_6_5_da;
  output xt_rsc_6_5_wea;
  input [31:0] xt_rsc_6_5_qa;
  output xt_rsc_triosy_6_5_lz;
  output [3:0] xt_rsc_6_6_adra;
  output [31:0] xt_rsc_6_6_da;
  output xt_rsc_6_6_wea;
  input [31:0] xt_rsc_6_6_qa;
  output xt_rsc_triosy_6_6_lz;
  output [3:0] xt_rsc_6_7_adra;
  output [31:0] xt_rsc_6_7_da;
  output xt_rsc_6_7_wea;
  input [31:0] xt_rsc_6_7_qa;
  output xt_rsc_triosy_6_7_lz;
  output [3:0] xt_rsc_6_8_adra;
  output [31:0] xt_rsc_6_8_da;
  output xt_rsc_6_8_wea;
  input [31:0] xt_rsc_6_8_qa;
  output xt_rsc_triosy_6_8_lz;
  output [3:0] xt_rsc_6_9_adra;
  output [31:0] xt_rsc_6_9_da;
  output xt_rsc_6_9_wea;
  input [31:0] xt_rsc_6_9_qa;
  output xt_rsc_triosy_6_9_lz;
  output [3:0] xt_rsc_6_10_adra;
  output [31:0] xt_rsc_6_10_da;
  output xt_rsc_6_10_wea;
  input [31:0] xt_rsc_6_10_qa;
  output xt_rsc_triosy_6_10_lz;
  output [3:0] xt_rsc_6_11_adra;
  output [31:0] xt_rsc_6_11_da;
  output xt_rsc_6_11_wea;
  input [31:0] xt_rsc_6_11_qa;
  output xt_rsc_triosy_6_11_lz;
  output [3:0] xt_rsc_6_12_adra;
  output [31:0] xt_rsc_6_12_da;
  output xt_rsc_6_12_wea;
  input [31:0] xt_rsc_6_12_qa;
  output xt_rsc_triosy_6_12_lz;
  output [3:0] xt_rsc_6_13_adra;
  output [31:0] xt_rsc_6_13_da;
  output xt_rsc_6_13_wea;
  input [31:0] xt_rsc_6_13_qa;
  output xt_rsc_triosy_6_13_lz;
  output [3:0] xt_rsc_6_14_adra;
  output [31:0] xt_rsc_6_14_da;
  output xt_rsc_6_14_wea;
  input [31:0] xt_rsc_6_14_qa;
  output xt_rsc_triosy_6_14_lz;
  output [3:0] xt_rsc_6_15_adra;
  output [31:0] xt_rsc_6_15_da;
  output xt_rsc_6_15_wea;
  input [31:0] xt_rsc_6_15_qa;
  output xt_rsc_triosy_6_15_lz;
  output [3:0] xt_rsc_6_16_adra;
  output [31:0] xt_rsc_6_16_da;
  output xt_rsc_6_16_wea;
  input [31:0] xt_rsc_6_16_qa;
  output xt_rsc_triosy_6_16_lz;
  output [3:0] xt_rsc_6_17_adra;
  output [31:0] xt_rsc_6_17_da;
  output xt_rsc_6_17_wea;
  input [31:0] xt_rsc_6_17_qa;
  output xt_rsc_triosy_6_17_lz;
  output [3:0] xt_rsc_6_18_adra;
  output [31:0] xt_rsc_6_18_da;
  output xt_rsc_6_18_wea;
  input [31:0] xt_rsc_6_18_qa;
  output xt_rsc_triosy_6_18_lz;
  output [3:0] xt_rsc_6_19_adra;
  output [31:0] xt_rsc_6_19_da;
  output xt_rsc_6_19_wea;
  input [31:0] xt_rsc_6_19_qa;
  output xt_rsc_triosy_6_19_lz;
  output [3:0] xt_rsc_6_20_adra;
  output [31:0] xt_rsc_6_20_da;
  output xt_rsc_6_20_wea;
  input [31:0] xt_rsc_6_20_qa;
  output xt_rsc_triosy_6_20_lz;
  output [3:0] xt_rsc_6_21_adra;
  output [31:0] xt_rsc_6_21_da;
  output xt_rsc_6_21_wea;
  input [31:0] xt_rsc_6_21_qa;
  output xt_rsc_triosy_6_21_lz;
  output [3:0] xt_rsc_6_22_adra;
  output [31:0] xt_rsc_6_22_da;
  output xt_rsc_6_22_wea;
  input [31:0] xt_rsc_6_22_qa;
  output xt_rsc_triosy_6_22_lz;
  output [3:0] xt_rsc_6_23_adra;
  output [31:0] xt_rsc_6_23_da;
  output xt_rsc_6_23_wea;
  input [31:0] xt_rsc_6_23_qa;
  output xt_rsc_triosy_6_23_lz;
  output [3:0] xt_rsc_6_24_adra;
  output [31:0] xt_rsc_6_24_da;
  output xt_rsc_6_24_wea;
  input [31:0] xt_rsc_6_24_qa;
  output xt_rsc_triosy_6_24_lz;
  output [3:0] xt_rsc_6_25_adra;
  output [31:0] xt_rsc_6_25_da;
  output xt_rsc_6_25_wea;
  input [31:0] xt_rsc_6_25_qa;
  output xt_rsc_triosy_6_25_lz;
  output [3:0] xt_rsc_6_26_adra;
  output [31:0] xt_rsc_6_26_da;
  output xt_rsc_6_26_wea;
  input [31:0] xt_rsc_6_26_qa;
  output xt_rsc_triosy_6_26_lz;
  output [3:0] xt_rsc_6_27_adra;
  output [31:0] xt_rsc_6_27_da;
  output xt_rsc_6_27_wea;
  input [31:0] xt_rsc_6_27_qa;
  output xt_rsc_triosy_6_27_lz;
  output [3:0] xt_rsc_6_28_adra;
  output [31:0] xt_rsc_6_28_da;
  output xt_rsc_6_28_wea;
  input [31:0] xt_rsc_6_28_qa;
  output xt_rsc_triosy_6_28_lz;
  output [3:0] xt_rsc_6_29_adra;
  output [31:0] xt_rsc_6_29_da;
  output xt_rsc_6_29_wea;
  input [31:0] xt_rsc_6_29_qa;
  output xt_rsc_triosy_6_29_lz;
  output [3:0] xt_rsc_6_30_adra;
  output [31:0] xt_rsc_6_30_da;
  output xt_rsc_6_30_wea;
  input [31:0] xt_rsc_6_30_qa;
  output xt_rsc_triosy_6_30_lz;
  output [3:0] xt_rsc_6_31_adra;
  output [31:0] xt_rsc_6_31_da;
  output xt_rsc_6_31_wea;
  input [31:0] xt_rsc_6_31_qa;
  output xt_rsc_triosy_6_31_lz;
  output [3:0] xt_rsc_7_0_adra;
  output [31:0] xt_rsc_7_0_da;
  output xt_rsc_7_0_wea;
  input [31:0] xt_rsc_7_0_qa;
  output xt_rsc_triosy_7_0_lz;
  output [3:0] xt_rsc_7_1_adra;
  output [31:0] xt_rsc_7_1_da;
  output xt_rsc_7_1_wea;
  input [31:0] xt_rsc_7_1_qa;
  output xt_rsc_triosy_7_1_lz;
  output [3:0] xt_rsc_7_2_adra;
  output [31:0] xt_rsc_7_2_da;
  output xt_rsc_7_2_wea;
  input [31:0] xt_rsc_7_2_qa;
  output xt_rsc_triosy_7_2_lz;
  output [3:0] xt_rsc_7_3_adra;
  output [31:0] xt_rsc_7_3_da;
  output xt_rsc_7_3_wea;
  input [31:0] xt_rsc_7_3_qa;
  output xt_rsc_triosy_7_3_lz;
  output [3:0] xt_rsc_7_4_adra;
  output [31:0] xt_rsc_7_4_da;
  output xt_rsc_7_4_wea;
  input [31:0] xt_rsc_7_4_qa;
  output xt_rsc_triosy_7_4_lz;
  output [3:0] xt_rsc_7_5_adra;
  output [31:0] xt_rsc_7_5_da;
  output xt_rsc_7_5_wea;
  input [31:0] xt_rsc_7_5_qa;
  output xt_rsc_triosy_7_5_lz;
  output [3:0] xt_rsc_7_6_adra;
  output [31:0] xt_rsc_7_6_da;
  output xt_rsc_7_6_wea;
  input [31:0] xt_rsc_7_6_qa;
  output xt_rsc_triosy_7_6_lz;
  output [3:0] xt_rsc_7_7_adra;
  output [31:0] xt_rsc_7_7_da;
  output xt_rsc_7_7_wea;
  input [31:0] xt_rsc_7_7_qa;
  output xt_rsc_triosy_7_7_lz;
  output [3:0] xt_rsc_7_8_adra;
  output [31:0] xt_rsc_7_8_da;
  output xt_rsc_7_8_wea;
  input [31:0] xt_rsc_7_8_qa;
  output xt_rsc_triosy_7_8_lz;
  output [3:0] xt_rsc_7_9_adra;
  output [31:0] xt_rsc_7_9_da;
  output xt_rsc_7_9_wea;
  input [31:0] xt_rsc_7_9_qa;
  output xt_rsc_triosy_7_9_lz;
  output [3:0] xt_rsc_7_10_adra;
  output [31:0] xt_rsc_7_10_da;
  output xt_rsc_7_10_wea;
  input [31:0] xt_rsc_7_10_qa;
  output xt_rsc_triosy_7_10_lz;
  output [3:0] xt_rsc_7_11_adra;
  output [31:0] xt_rsc_7_11_da;
  output xt_rsc_7_11_wea;
  input [31:0] xt_rsc_7_11_qa;
  output xt_rsc_triosy_7_11_lz;
  output [3:0] xt_rsc_7_12_adra;
  output [31:0] xt_rsc_7_12_da;
  output xt_rsc_7_12_wea;
  input [31:0] xt_rsc_7_12_qa;
  output xt_rsc_triosy_7_12_lz;
  output [3:0] xt_rsc_7_13_adra;
  output [31:0] xt_rsc_7_13_da;
  output xt_rsc_7_13_wea;
  input [31:0] xt_rsc_7_13_qa;
  output xt_rsc_triosy_7_13_lz;
  output [3:0] xt_rsc_7_14_adra;
  output [31:0] xt_rsc_7_14_da;
  output xt_rsc_7_14_wea;
  input [31:0] xt_rsc_7_14_qa;
  output xt_rsc_triosy_7_14_lz;
  output [3:0] xt_rsc_7_15_adra;
  output [31:0] xt_rsc_7_15_da;
  output xt_rsc_7_15_wea;
  input [31:0] xt_rsc_7_15_qa;
  output xt_rsc_triosy_7_15_lz;
  output [3:0] xt_rsc_7_16_adra;
  output [31:0] xt_rsc_7_16_da;
  output xt_rsc_7_16_wea;
  input [31:0] xt_rsc_7_16_qa;
  output xt_rsc_triosy_7_16_lz;
  output [3:0] xt_rsc_7_17_adra;
  output [31:0] xt_rsc_7_17_da;
  output xt_rsc_7_17_wea;
  input [31:0] xt_rsc_7_17_qa;
  output xt_rsc_triosy_7_17_lz;
  output [3:0] xt_rsc_7_18_adra;
  output [31:0] xt_rsc_7_18_da;
  output xt_rsc_7_18_wea;
  input [31:0] xt_rsc_7_18_qa;
  output xt_rsc_triosy_7_18_lz;
  output [3:0] xt_rsc_7_19_adra;
  output [31:0] xt_rsc_7_19_da;
  output xt_rsc_7_19_wea;
  input [31:0] xt_rsc_7_19_qa;
  output xt_rsc_triosy_7_19_lz;
  output [3:0] xt_rsc_7_20_adra;
  output [31:0] xt_rsc_7_20_da;
  output xt_rsc_7_20_wea;
  input [31:0] xt_rsc_7_20_qa;
  output xt_rsc_triosy_7_20_lz;
  output [3:0] xt_rsc_7_21_adra;
  output [31:0] xt_rsc_7_21_da;
  output xt_rsc_7_21_wea;
  input [31:0] xt_rsc_7_21_qa;
  output xt_rsc_triosy_7_21_lz;
  output [3:0] xt_rsc_7_22_adra;
  output [31:0] xt_rsc_7_22_da;
  output xt_rsc_7_22_wea;
  input [31:0] xt_rsc_7_22_qa;
  output xt_rsc_triosy_7_22_lz;
  output [3:0] xt_rsc_7_23_adra;
  output [31:0] xt_rsc_7_23_da;
  output xt_rsc_7_23_wea;
  input [31:0] xt_rsc_7_23_qa;
  output xt_rsc_triosy_7_23_lz;
  output [3:0] xt_rsc_7_24_adra;
  output [31:0] xt_rsc_7_24_da;
  output xt_rsc_7_24_wea;
  input [31:0] xt_rsc_7_24_qa;
  output xt_rsc_triosy_7_24_lz;
  output [3:0] xt_rsc_7_25_adra;
  output [31:0] xt_rsc_7_25_da;
  output xt_rsc_7_25_wea;
  input [31:0] xt_rsc_7_25_qa;
  output xt_rsc_triosy_7_25_lz;
  output [3:0] xt_rsc_7_26_adra;
  output [31:0] xt_rsc_7_26_da;
  output xt_rsc_7_26_wea;
  input [31:0] xt_rsc_7_26_qa;
  output xt_rsc_triosy_7_26_lz;
  output [3:0] xt_rsc_7_27_adra;
  output [31:0] xt_rsc_7_27_da;
  output xt_rsc_7_27_wea;
  input [31:0] xt_rsc_7_27_qa;
  output xt_rsc_triosy_7_27_lz;
  output [3:0] xt_rsc_7_28_adra;
  output [31:0] xt_rsc_7_28_da;
  output xt_rsc_7_28_wea;
  input [31:0] xt_rsc_7_28_qa;
  output xt_rsc_triosy_7_28_lz;
  output [3:0] xt_rsc_7_29_adra;
  output [31:0] xt_rsc_7_29_da;
  output xt_rsc_7_29_wea;
  input [31:0] xt_rsc_7_29_qa;
  output xt_rsc_triosy_7_29_lz;
  output [3:0] xt_rsc_7_30_adra;
  output [31:0] xt_rsc_7_30_da;
  output xt_rsc_7_30_wea;
  input [31:0] xt_rsc_7_30_qa;
  output xt_rsc_triosy_7_30_lz;
  output [3:0] xt_rsc_7_31_adra;
  output [31:0] xt_rsc_7_31_da;
  output xt_rsc_7_31_wea;
  input [31:0] xt_rsc_7_31_qa;
  output xt_rsc_triosy_7_31_lz;
  input [31:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [31:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [7:0] twiddle_rsc_0_0_adra;
  output [31:0] twiddle_rsc_0_0_da;
  output twiddle_rsc_0_0_wea;
  input [31:0] twiddle_rsc_0_0_qa;
  output [7:0] twiddle_rsc_0_0_adrb;
  output [31:0] twiddle_rsc_0_0_db;
  output twiddle_rsc_0_0_web;
  input [31:0] twiddle_rsc_0_0_qb;
  output twiddle_rsc_triosy_0_0_lz;
  output [7:0] twiddle_rsc_0_1_adra;
  output [31:0] twiddle_rsc_0_1_da;
  output twiddle_rsc_0_1_wea;
  input [31:0] twiddle_rsc_0_1_qa;
  output [7:0] twiddle_rsc_0_1_adrb;
  output [31:0] twiddle_rsc_0_1_db;
  output twiddle_rsc_0_1_web;
  input [31:0] twiddle_rsc_0_1_qb;
  output twiddle_rsc_triosy_0_1_lz;
  output [7:0] twiddle_rsc_0_2_adra;
  output [31:0] twiddle_rsc_0_2_da;
  output twiddle_rsc_0_2_wea;
  input [31:0] twiddle_rsc_0_2_qa;
  output [7:0] twiddle_rsc_0_2_adrb;
  output [31:0] twiddle_rsc_0_2_db;
  output twiddle_rsc_0_2_web;
  input [31:0] twiddle_rsc_0_2_qb;
  output twiddle_rsc_triosy_0_2_lz;
  output [7:0] twiddle_rsc_0_3_adra;
  output [31:0] twiddle_rsc_0_3_da;
  output twiddle_rsc_0_3_wea;
  input [31:0] twiddle_rsc_0_3_qa;
  output [7:0] twiddle_rsc_0_3_adrb;
  output [31:0] twiddle_rsc_0_3_db;
  output twiddle_rsc_0_3_web;
  input [31:0] twiddle_rsc_0_3_qb;
  output twiddle_rsc_triosy_0_3_lz;
  output [7:0] twiddle_rsc_0_4_adra;
  output [31:0] twiddle_rsc_0_4_da;
  output twiddle_rsc_0_4_wea;
  input [31:0] twiddle_rsc_0_4_qa;
  output [7:0] twiddle_rsc_0_4_adrb;
  output [31:0] twiddle_rsc_0_4_db;
  output twiddle_rsc_0_4_web;
  input [31:0] twiddle_rsc_0_4_qb;
  output twiddle_rsc_triosy_0_4_lz;
  output [7:0] twiddle_rsc_0_5_adra;
  output [31:0] twiddle_rsc_0_5_da;
  output twiddle_rsc_0_5_wea;
  input [31:0] twiddle_rsc_0_5_qa;
  output [7:0] twiddle_rsc_0_5_adrb;
  output [31:0] twiddle_rsc_0_5_db;
  output twiddle_rsc_0_5_web;
  input [31:0] twiddle_rsc_0_5_qb;
  output twiddle_rsc_triosy_0_5_lz;
  output [7:0] twiddle_rsc_0_6_adra;
  output [31:0] twiddle_rsc_0_6_da;
  output twiddle_rsc_0_6_wea;
  input [31:0] twiddle_rsc_0_6_qa;
  output [7:0] twiddle_rsc_0_6_adrb;
  output [31:0] twiddle_rsc_0_6_db;
  output twiddle_rsc_0_6_web;
  input [31:0] twiddle_rsc_0_6_qb;
  output twiddle_rsc_triosy_0_6_lz;
  output [7:0] twiddle_rsc_0_7_adra;
  output [31:0] twiddle_rsc_0_7_da;
  output twiddle_rsc_0_7_wea;
  input [31:0] twiddle_rsc_0_7_qa;
  output [7:0] twiddle_rsc_0_7_adrb;
  output [31:0] twiddle_rsc_0_7_db;
  output twiddle_rsc_0_7_web;
  input [31:0] twiddle_rsc_0_7_qb;
  output twiddle_rsc_triosy_0_7_lz;
  output [7:0] twiddle_rsc_0_8_adra;
  output [31:0] twiddle_rsc_0_8_da;
  output twiddle_rsc_0_8_wea;
  input [31:0] twiddle_rsc_0_8_qa;
  output [7:0] twiddle_rsc_0_8_adrb;
  output [31:0] twiddle_rsc_0_8_db;
  output twiddle_rsc_0_8_web;
  input [31:0] twiddle_rsc_0_8_qb;
  output twiddle_rsc_triosy_0_8_lz;
  output [7:0] twiddle_rsc_0_9_adra;
  output [31:0] twiddle_rsc_0_9_da;
  output twiddle_rsc_0_9_wea;
  input [31:0] twiddle_rsc_0_9_qa;
  output [7:0] twiddle_rsc_0_9_adrb;
  output [31:0] twiddle_rsc_0_9_db;
  output twiddle_rsc_0_9_web;
  input [31:0] twiddle_rsc_0_9_qb;
  output twiddle_rsc_triosy_0_9_lz;
  output [7:0] twiddle_rsc_0_10_adra;
  output [31:0] twiddle_rsc_0_10_da;
  output twiddle_rsc_0_10_wea;
  input [31:0] twiddle_rsc_0_10_qa;
  output [7:0] twiddle_rsc_0_10_adrb;
  output [31:0] twiddle_rsc_0_10_db;
  output twiddle_rsc_0_10_web;
  input [31:0] twiddle_rsc_0_10_qb;
  output twiddle_rsc_triosy_0_10_lz;
  output [7:0] twiddle_rsc_0_11_adra;
  output [31:0] twiddle_rsc_0_11_da;
  output twiddle_rsc_0_11_wea;
  input [31:0] twiddle_rsc_0_11_qa;
  output [7:0] twiddle_rsc_0_11_adrb;
  output [31:0] twiddle_rsc_0_11_db;
  output twiddle_rsc_0_11_web;
  input [31:0] twiddle_rsc_0_11_qb;
  output twiddle_rsc_triosy_0_11_lz;
  output [7:0] twiddle_rsc_0_12_adra;
  output [31:0] twiddle_rsc_0_12_da;
  output twiddle_rsc_0_12_wea;
  input [31:0] twiddle_rsc_0_12_qa;
  output [7:0] twiddle_rsc_0_12_adrb;
  output [31:0] twiddle_rsc_0_12_db;
  output twiddle_rsc_0_12_web;
  input [31:0] twiddle_rsc_0_12_qb;
  output twiddle_rsc_triosy_0_12_lz;
  output [7:0] twiddle_rsc_0_13_adra;
  output [31:0] twiddle_rsc_0_13_da;
  output twiddle_rsc_0_13_wea;
  input [31:0] twiddle_rsc_0_13_qa;
  output [7:0] twiddle_rsc_0_13_adrb;
  output [31:0] twiddle_rsc_0_13_db;
  output twiddle_rsc_0_13_web;
  input [31:0] twiddle_rsc_0_13_qb;
  output twiddle_rsc_triosy_0_13_lz;
  output [7:0] twiddle_rsc_0_14_adra;
  output [31:0] twiddle_rsc_0_14_da;
  output twiddle_rsc_0_14_wea;
  input [31:0] twiddle_rsc_0_14_qa;
  output [7:0] twiddle_rsc_0_14_adrb;
  output [31:0] twiddle_rsc_0_14_db;
  output twiddle_rsc_0_14_web;
  input [31:0] twiddle_rsc_0_14_qb;
  output twiddle_rsc_triosy_0_14_lz;
  output [7:0] twiddle_rsc_0_15_adra;
  output [31:0] twiddle_rsc_0_15_da;
  output twiddle_rsc_0_15_wea;
  input [31:0] twiddle_rsc_0_15_qa;
  output [7:0] twiddle_rsc_0_15_adrb;
  output [31:0] twiddle_rsc_0_15_db;
  output twiddle_rsc_0_15_web;
  input [31:0] twiddle_rsc_0_15_qb;
  output twiddle_rsc_triosy_0_15_lz;
  output [7:0] twiddle_h_rsc_0_0_adra;
  output [31:0] twiddle_h_rsc_0_0_da;
  output twiddle_h_rsc_0_0_wea;
  input [31:0] twiddle_h_rsc_0_0_qa;
  output [7:0] twiddle_h_rsc_0_0_adrb;
  output [31:0] twiddle_h_rsc_0_0_db;
  output twiddle_h_rsc_0_0_web;
  input [31:0] twiddle_h_rsc_0_0_qb;
  output twiddle_h_rsc_triosy_0_0_lz;
  output [7:0] twiddle_h_rsc_0_1_adra;
  output [31:0] twiddle_h_rsc_0_1_da;
  output twiddle_h_rsc_0_1_wea;
  input [31:0] twiddle_h_rsc_0_1_qa;
  output [7:0] twiddle_h_rsc_0_1_adrb;
  output [31:0] twiddle_h_rsc_0_1_db;
  output twiddle_h_rsc_0_1_web;
  input [31:0] twiddle_h_rsc_0_1_qb;
  output twiddle_h_rsc_triosy_0_1_lz;
  output [7:0] twiddle_h_rsc_0_2_adra;
  output [31:0] twiddle_h_rsc_0_2_da;
  output twiddle_h_rsc_0_2_wea;
  input [31:0] twiddle_h_rsc_0_2_qa;
  output [7:0] twiddle_h_rsc_0_2_adrb;
  output [31:0] twiddle_h_rsc_0_2_db;
  output twiddle_h_rsc_0_2_web;
  input [31:0] twiddle_h_rsc_0_2_qb;
  output twiddle_h_rsc_triosy_0_2_lz;
  output [7:0] twiddle_h_rsc_0_3_adra;
  output [31:0] twiddle_h_rsc_0_3_da;
  output twiddle_h_rsc_0_3_wea;
  input [31:0] twiddle_h_rsc_0_3_qa;
  output [7:0] twiddle_h_rsc_0_3_adrb;
  output [31:0] twiddle_h_rsc_0_3_db;
  output twiddle_h_rsc_0_3_web;
  input [31:0] twiddle_h_rsc_0_3_qb;
  output twiddle_h_rsc_triosy_0_3_lz;
  output [7:0] twiddle_h_rsc_0_4_adra;
  output [31:0] twiddle_h_rsc_0_4_da;
  output twiddle_h_rsc_0_4_wea;
  input [31:0] twiddle_h_rsc_0_4_qa;
  output [7:0] twiddle_h_rsc_0_4_adrb;
  output [31:0] twiddle_h_rsc_0_4_db;
  output twiddle_h_rsc_0_4_web;
  input [31:0] twiddle_h_rsc_0_4_qb;
  output twiddle_h_rsc_triosy_0_4_lz;
  output [7:0] twiddle_h_rsc_0_5_adra;
  output [31:0] twiddle_h_rsc_0_5_da;
  output twiddle_h_rsc_0_5_wea;
  input [31:0] twiddle_h_rsc_0_5_qa;
  output [7:0] twiddle_h_rsc_0_5_adrb;
  output [31:0] twiddle_h_rsc_0_5_db;
  output twiddle_h_rsc_0_5_web;
  input [31:0] twiddle_h_rsc_0_5_qb;
  output twiddle_h_rsc_triosy_0_5_lz;
  output [7:0] twiddle_h_rsc_0_6_adra;
  output [31:0] twiddle_h_rsc_0_6_da;
  output twiddle_h_rsc_0_6_wea;
  input [31:0] twiddle_h_rsc_0_6_qa;
  output [7:0] twiddle_h_rsc_0_6_adrb;
  output [31:0] twiddle_h_rsc_0_6_db;
  output twiddle_h_rsc_0_6_web;
  input [31:0] twiddle_h_rsc_0_6_qb;
  output twiddle_h_rsc_triosy_0_6_lz;
  output [7:0] twiddle_h_rsc_0_7_adra;
  output [31:0] twiddle_h_rsc_0_7_da;
  output twiddle_h_rsc_0_7_wea;
  input [31:0] twiddle_h_rsc_0_7_qa;
  output [7:0] twiddle_h_rsc_0_7_adrb;
  output [31:0] twiddle_h_rsc_0_7_db;
  output twiddle_h_rsc_0_7_web;
  input [31:0] twiddle_h_rsc_0_7_qb;
  output twiddle_h_rsc_triosy_0_7_lz;
  output [7:0] twiddle_h_rsc_0_8_adra;
  output [31:0] twiddle_h_rsc_0_8_da;
  output twiddle_h_rsc_0_8_wea;
  input [31:0] twiddle_h_rsc_0_8_qa;
  output [7:0] twiddle_h_rsc_0_8_adrb;
  output [31:0] twiddle_h_rsc_0_8_db;
  output twiddle_h_rsc_0_8_web;
  input [31:0] twiddle_h_rsc_0_8_qb;
  output twiddle_h_rsc_triosy_0_8_lz;
  output [7:0] twiddle_h_rsc_0_9_adra;
  output [31:0] twiddle_h_rsc_0_9_da;
  output twiddle_h_rsc_0_9_wea;
  input [31:0] twiddle_h_rsc_0_9_qa;
  output [7:0] twiddle_h_rsc_0_9_adrb;
  output [31:0] twiddle_h_rsc_0_9_db;
  output twiddle_h_rsc_0_9_web;
  input [31:0] twiddle_h_rsc_0_9_qb;
  output twiddle_h_rsc_triosy_0_9_lz;
  output [7:0] twiddle_h_rsc_0_10_adra;
  output [31:0] twiddle_h_rsc_0_10_da;
  output twiddle_h_rsc_0_10_wea;
  input [31:0] twiddle_h_rsc_0_10_qa;
  output [7:0] twiddle_h_rsc_0_10_adrb;
  output [31:0] twiddle_h_rsc_0_10_db;
  output twiddle_h_rsc_0_10_web;
  input [31:0] twiddle_h_rsc_0_10_qb;
  output twiddle_h_rsc_triosy_0_10_lz;
  output [7:0] twiddle_h_rsc_0_11_adra;
  output [31:0] twiddle_h_rsc_0_11_da;
  output twiddle_h_rsc_0_11_wea;
  input [31:0] twiddle_h_rsc_0_11_qa;
  output [7:0] twiddle_h_rsc_0_11_adrb;
  output [31:0] twiddle_h_rsc_0_11_db;
  output twiddle_h_rsc_0_11_web;
  input [31:0] twiddle_h_rsc_0_11_qb;
  output twiddle_h_rsc_triosy_0_11_lz;
  output [7:0] twiddle_h_rsc_0_12_adra;
  output [31:0] twiddle_h_rsc_0_12_da;
  output twiddle_h_rsc_0_12_wea;
  input [31:0] twiddle_h_rsc_0_12_qa;
  output [7:0] twiddle_h_rsc_0_12_adrb;
  output [31:0] twiddle_h_rsc_0_12_db;
  output twiddle_h_rsc_0_12_web;
  input [31:0] twiddle_h_rsc_0_12_qb;
  output twiddle_h_rsc_triosy_0_12_lz;
  output [7:0] twiddle_h_rsc_0_13_adra;
  output [31:0] twiddle_h_rsc_0_13_da;
  output twiddle_h_rsc_0_13_wea;
  input [31:0] twiddle_h_rsc_0_13_qa;
  output [7:0] twiddle_h_rsc_0_13_adrb;
  output [31:0] twiddle_h_rsc_0_13_db;
  output twiddle_h_rsc_0_13_web;
  input [31:0] twiddle_h_rsc_0_13_qb;
  output twiddle_h_rsc_triosy_0_13_lz;
  output [7:0] twiddle_h_rsc_0_14_adra;
  output [31:0] twiddle_h_rsc_0_14_da;
  output twiddle_h_rsc_0_14_wea;
  input [31:0] twiddle_h_rsc_0_14_qa;
  output [7:0] twiddle_h_rsc_0_14_adrb;
  output [31:0] twiddle_h_rsc_0_14_db;
  output twiddle_h_rsc_0_14_web;
  input [31:0] twiddle_h_rsc_0_14_qb;
  output twiddle_h_rsc_triosy_0_14_lz;
  output [7:0] twiddle_h_rsc_0_15_adra;
  output [31:0] twiddle_h_rsc_0_15_da;
  output twiddle_h_rsc_0_15_wea;
  input [31:0] twiddle_h_rsc_0_15_qa;
  output [7:0] twiddle_h_rsc_0_15_adrb;
  output [31:0] twiddle_h_rsc_0_15_db;
  output twiddle_h_rsc_0_15_web;
  input [31:0] twiddle_h_rsc_0_15_qb;
  output twiddle_h_rsc_triosy_0_15_lz;


  // Interconnect Declarations
  wire yt_rsc_0_0_i_clkr_en_d;
  wire [31:0] yt_rsc_0_0_i_q_d;
  wire [31:0] yt_rsc_0_1_i_q_d;
  wire [31:0] yt_rsc_0_2_i_q_d;
  wire [31:0] yt_rsc_0_3_i_q_d;
  wire [31:0] yt_rsc_0_4_i_q_d;
  wire [31:0] yt_rsc_0_5_i_q_d;
  wire [31:0] yt_rsc_0_6_i_q_d;
  wire [31:0] yt_rsc_0_7_i_q_d;
  wire [31:0] yt_rsc_0_8_i_q_d;
  wire [31:0] yt_rsc_0_9_i_q_d;
  wire [31:0] yt_rsc_0_10_i_q_d;
  wire [31:0] yt_rsc_0_11_i_q_d;
  wire [31:0] yt_rsc_0_12_i_q_d;
  wire [31:0] yt_rsc_0_13_i_q_d;
  wire [31:0] yt_rsc_0_14_i_q_d;
  wire [31:0] yt_rsc_0_15_i_q_d;
  wire yt_rsc_0_16_i_clkr_en_d;
  wire [31:0] yt_rsc_0_16_i_q_d;
  wire [31:0] yt_rsc_0_17_i_q_d;
  wire [31:0] yt_rsc_0_18_i_q_d;
  wire [31:0] yt_rsc_0_19_i_q_d;
  wire [31:0] yt_rsc_0_20_i_q_d;
  wire [31:0] yt_rsc_0_21_i_q_d;
  wire [31:0] yt_rsc_0_22_i_q_d;
  wire [31:0] yt_rsc_0_23_i_q_d;
  wire [31:0] yt_rsc_0_24_i_q_d;
  wire [31:0] yt_rsc_0_25_i_q_d;
  wire [31:0] yt_rsc_0_26_i_q_d;
  wire [31:0] yt_rsc_0_27_i_q_d;
  wire [31:0] yt_rsc_0_28_i_q_d;
  wire [31:0] yt_rsc_0_29_i_q_d;
  wire [31:0] yt_rsc_0_30_i_q_d;
  wire [31:0] yt_rsc_0_31_i_q_d;
  wire yt_rsc_1_0_i_clkr_en_d;
  wire [31:0] yt_rsc_1_0_i_q_d;
  wire [31:0] yt_rsc_1_1_i_q_d;
  wire [31:0] yt_rsc_1_2_i_q_d;
  wire [31:0] yt_rsc_1_3_i_q_d;
  wire [31:0] yt_rsc_1_4_i_q_d;
  wire [31:0] yt_rsc_1_5_i_q_d;
  wire [31:0] yt_rsc_1_6_i_q_d;
  wire [31:0] yt_rsc_1_7_i_q_d;
  wire [31:0] yt_rsc_1_8_i_q_d;
  wire [31:0] yt_rsc_1_9_i_q_d;
  wire [31:0] yt_rsc_1_10_i_q_d;
  wire [31:0] yt_rsc_1_11_i_q_d;
  wire [31:0] yt_rsc_1_12_i_q_d;
  wire [31:0] yt_rsc_1_13_i_q_d;
  wire [31:0] yt_rsc_1_14_i_q_d;
  wire [31:0] yt_rsc_1_15_i_q_d;
  wire yt_rsc_1_16_i_clkr_en_d;
  wire [31:0] yt_rsc_1_16_i_q_d;
  wire [31:0] yt_rsc_1_17_i_q_d;
  wire [31:0] yt_rsc_1_18_i_q_d;
  wire [31:0] yt_rsc_1_19_i_q_d;
  wire [31:0] yt_rsc_1_20_i_q_d;
  wire [31:0] yt_rsc_1_21_i_q_d;
  wire [31:0] yt_rsc_1_22_i_q_d;
  wire [31:0] yt_rsc_1_23_i_q_d;
  wire [31:0] yt_rsc_1_24_i_q_d;
  wire [31:0] yt_rsc_1_25_i_q_d;
  wire [31:0] yt_rsc_1_26_i_q_d;
  wire [31:0] yt_rsc_1_27_i_q_d;
  wire [31:0] yt_rsc_1_28_i_q_d;
  wire [31:0] yt_rsc_1_29_i_q_d;
  wire [31:0] yt_rsc_1_30_i_q_d;
  wire [31:0] yt_rsc_1_31_i_q_d;
  wire yt_rsc_2_0_i_clkr_en_d;
  wire [31:0] yt_rsc_2_0_i_q_d;
  wire [31:0] yt_rsc_2_1_i_q_d;
  wire [31:0] yt_rsc_2_2_i_q_d;
  wire [31:0] yt_rsc_2_3_i_q_d;
  wire [31:0] yt_rsc_2_4_i_q_d;
  wire [31:0] yt_rsc_2_5_i_q_d;
  wire [31:0] yt_rsc_2_6_i_q_d;
  wire [31:0] yt_rsc_2_7_i_q_d;
  wire [31:0] yt_rsc_2_8_i_q_d;
  wire [31:0] yt_rsc_2_9_i_q_d;
  wire [31:0] yt_rsc_2_10_i_q_d;
  wire [31:0] yt_rsc_2_11_i_q_d;
  wire [31:0] yt_rsc_2_12_i_q_d;
  wire [31:0] yt_rsc_2_13_i_q_d;
  wire [31:0] yt_rsc_2_14_i_q_d;
  wire [31:0] yt_rsc_2_15_i_q_d;
  wire yt_rsc_2_16_i_clkr_en_d;
  wire [31:0] yt_rsc_2_16_i_q_d;
  wire [31:0] yt_rsc_2_17_i_q_d;
  wire [31:0] yt_rsc_2_18_i_q_d;
  wire [31:0] yt_rsc_2_19_i_q_d;
  wire [31:0] yt_rsc_2_20_i_q_d;
  wire [31:0] yt_rsc_2_21_i_q_d;
  wire [31:0] yt_rsc_2_22_i_q_d;
  wire [31:0] yt_rsc_2_23_i_q_d;
  wire [31:0] yt_rsc_2_24_i_q_d;
  wire [31:0] yt_rsc_2_25_i_q_d;
  wire [31:0] yt_rsc_2_26_i_q_d;
  wire [31:0] yt_rsc_2_27_i_q_d;
  wire [31:0] yt_rsc_2_28_i_q_d;
  wire [31:0] yt_rsc_2_29_i_q_d;
  wire [31:0] yt_rsc_2_30_i_q_d;
  wire [31:0] yt_rsc_2_31_i_q_d;
  wire yt_rsc_3_0_i_clkr_en_d;
  wire [31:0] yt_rsc_3_0_i_q_d;
  wire [31:0] yt_rsc_3_1_i_q_d;
  wire [31:0] yt_rsc_3_2_i_q_d;
  wire [31:0] yt_rsc_3_3_i_q_d;
  wire [31:0] yt_rsc_3_4_i_q_d;
  wire [31:0] yt_rsc_3_5_i_q_d;
  wire [31:0] yt_rsc_3_6_i_q_d;
  wire [31:0] yt_rsc_3_7_i_q_d;
  wire [31:0] yt_rsc_3_8_i_q_d;
  wire [31:0] yt_rsc_3_9_i_q_d;
  wire [31:0] yt_rsc_3_10_i_q_d;
  wire [31:0] yt_rsc_3_11_i_q_d;
  wire [31:0] yt_rsc_3_12_i_q_d;
  wire [31:0] yt_rsc_3_13_i_q_d;
  wire [31:0] yt_rsc_3_14_i_q_d;
  wire [31:0] yt_rsc_3_15_i_q_d;
  wire yt_rsc_3_16_i_clkr_en_d;
  wire [31:0] yt_rsc_3_16_i_q_d;
  wire [31:0] yt_rsc_3_17_i_q_d;
  wire [31:0] yt_rsc_3_18_i_q_d;
  wire [31:0] yt_rsc_3_19_i_q_d;
  wire [31:0] yt_rsc_3_20_i_q_d;
  wire [31:0] yt_rsc_3_21_i_q_d;
  wire [31:0] yt_rsc_3_22_i_q_d;
  wire [31:0] yt_rsc_3_23_i_q_d;
  wire [31:0] yt_rsc_3_24_i_q_d;
  wire [31:0] yt_rsc_3_25_i_q_d;
  wire [31:0] yt_rsc_3_26_i_q_d;
  wire [31:0] yt_rsc_3_27_i_q_d;
  wire [31:0] yt_rsc_3_28_i_q_d;
  wire [31:0] yt_rsc_3_29_i_q_d;
  wire [31:0] yt_rsc_3_30_i_q_d;
  wire [31:0] yt_rsc_3_31_i_q_d;
  wire yt_rsc_4_0_i_clkr_en_d;
  wire [31:0] yt_rsc_4_0_i_q_d;
  wire [31:0] yt_rsc_4_1_i_q_d;
  wire [31:0] yt_rsc_4_2_i_q_d;
  wire [31:0] yt_rsc_4_3_i_q_d;
  wire [31:0] yt_rsc_4_4_i_q_d;
  wire [31:0] yt_rsc_4_5_i_q_d;
  wire [31:0] yt_rsc_4_6_i_q_d;
  wire [31:0] yt_rsc_4_7_i_q_d;
  wire [31:0] yt_rsc_4_8_i_q_d;
  wire [31:0] yt_rsc_4_9_i_q_d;
  wire [31:0] yt_rsc_4_10_i_q_d;
  wire [31:0] yt_rsc_4_11_i_q_d;
  wire [31:0] yt_rsc_4_12_i_q_d;
  wire [31:0] yt_rsc_4_13_i_q_d;
  wire [31:0] yt_rsc_4_14_i_q_d;
  wire [31:0] yt_rsc_4_15_i_q_d;
  wire yt_rsc_4_16_i_clkr_en_d;
  wire [31:0] yt_rsc_4_16_i_q_d;
  wire [31:0] yt_rsc_4_17_i_q_d;
  wire [31:0] yt_rsc_4_18_i_q_d;
  wire [31:0] yt_rsc_4_19_i_q_d;
  wire [31:0] yt_rsc_4_20_i_q_d;
  wire [31:0] yt_rsc_4_21_i_q_d;
  wire [31:0] yt_rsc_4_22_i_q_d;
  wire [31:0] yt_rsc_4_23_i_q_d;
  wire [31:0] yt_rsc_4_24_i_q_d;
  wire [31:0] yt_rsc_4_25_i_q_d;
  wire [31:0] yt_rsc_4_26_i_q_d;
  wire [31:0] yt_rsc_4_27_i_q_d;
  wire [31:0] yt_rsc_4_28_i_q_d;
  wire [31:0] yt_rsc_4_29_i_q_d;
  wire [31:0] yt_rsc_4_30_i_q_d;
  wire [31:0] yt_rsc_4_31_i_q_d;
  wire yt_rsc_5_0_i_clkr_en_d;
  wire [31:0] yt_rsc_5_0_i_q_d;
  wire [31:0] yt_rsc_5_1_i_q_d;
  wire [31:0] yt_rsc_5_2_i_q_d;
  wire [31:0] yt_rsc_5_3_i_q_d;
  wire [31:0] yt_rsc_5_4_i_q_d;
  wire [31:0] yt_rsc_5_5_i_q_d;
  wire [31:0] yt_rsc_5_6_i_q_d;
  wire [31:0] yt_rsc_5_7_i_q_d;
  wire [31:0] yt_rsc_5_8_i_q_d;
  wire [31:0] yt_rsc_5_9_i_q_d;
  wire [31:0] yt_rsc_5_10_i_q_d;
  wire [31:0] yt_rsc_5_11_i_q_d;
  wire [31:0] yt_rsc_5_12_i_q_d;
  wire [31:0] yt_rsc_5_13_i_q_d;
  wire [31:0] yt_rsc_5_14_i_q_d;
  wire [31:0] yt_rsc_5_15_i_q_d;
  wire yt_rsc_5_16_i_clkr_en_d;
  wire [31:0] yt_rsc_5_16_i_q_d;
  wire [31:0] yt_rsc_5_17_i_q_d;
  wire [31:0] yt_rsc_5_18_i_q_d;
  wire [31:0] yt_rsc_5_19_i_q_d;
  wire [31:0] yt_rsc_5_20_i_q_d;
  wire [31:0] yt_rsc_5_21_i_q_d;
  wire [31:0] yt_rsc_5_22_i_q_d;
  wire [31:0] yt_rsc_5_23_i_q_d;
  wire [31:0] yt_rsc_5_24_i_q_d;
  wire [31:0] yt_rsc_5_25_i_q_d;
  wire [31:0] yt_rsc_5_26_i_q_d;
  wire [31:0] yt_rsc_5_27_i_q_d;
  wire [31:0] yt_rsc_5_28_i_q_d;
  wire [31:0] yt_rsc_5_29_i_q_d;
  wire [31:0] yt_rsc_5_30_i_q_d;
  wire [31:0] yt_rsc_5_31_i_q_d;
  wire yt_rsc_6_0_i_clkr_en_d;
  wire [31:0] yt_rsc_6_0_i_q_d;
  wire [31:0] yt_rsc_6_1_i_q_d;
  wire [31:0] yt_rsc_6_2_i_q_d;
  wire [31:0] yt_rsc_6_3_i_q_d;
  wire [31:0] yt_rsc_6_4_i_q_d;
  wire [31:0] yt_rsc_6_5_i_q_d;
  wire [31:0] yt_rsc_6_6_i_q_d;
  wire [31:0] yt_rsc_6_7_i_q_d;
  wire [31:0] yt_rsc_6_8_i_q_d;
  wire [31:0] yt_rsc_6_9_i_q_d;
  wire [31:0] yt_rsc_6_10_i_q_d;
  wire [31:0] yt_rsc_6_11_i_q_d;
  wire [31:0] yt_rsc_6_12_i_q_d;
  wire [31:0] yt_rsc_6_13_i_q_d;
  wire [31:0] yt_rsc_6_14_i_q_d;
  wire [31:0] yt_rsc_6_15_i_q_d;
  wire yt_rsc_6_16_i_clkr_en_d;
  wire [31:0] yt_rsc_6_16_i_q_d;
  wire [31:0] yt_rsc_6_17_i_q_d;
  wire [31:0] yt_rsc_6_18_i_q_d;
  wire [31:0] yt_rsc_6_19_i_q_d;
  wire [31:0] yt_rsc_6_20_i_q_d;
  wire [31:0] yt_rsc_6_21_i_q_d;
  wire [31:0] yt_rsc_6_22_i_q_d;
  wire [31:0] yt_rsc_6_23_i_q_d;
  wire [31:0] yt_rsc_6_24_i_q_d;
  wire [31:0] yt_rsc_6_25_i_q_d;
  wire [31:0] yt_rsc_6_26_i_q_d;
  wire [31:0] yt_rsc_6_27_i_q_d;
  wire [31:0] yt_rsc_6_28_i_q_d;
  wire [31:0] yt_rsc_6_29_i_q_d;
  wire [31:0] yt_rsc_6_30_i_q_d;
  wire [31:0] yt_rsc_6_31_i_q_d;
  wire yt_rsc_7_0_i_clkr_en_d;
  wire [31:0] yt_rsc_7_0_i_q_d;
  wire [31:0] yt_rsc_7_1_i_q_d;
  wire [31:0] yt_rsc_7_2_i_q_d;
  wire [31:0] yt_rsc_7_3_i_q_d;
  wire [31:0] yt_rsc_7_4_i_q_d;
  wire [31:0] yt_rsc_7_5_i_q_d;
  wire [31:0] yt_rsc_7_6_i_q_d;
  wire [31:0] yt_rsc_7_7_i_q_d;
  wire [31:0] yt_rsc_7_8_i_q_d;
  wire [31:0] yt_rsc_7_9_i_q_d;
  wire [31:0] yt_rsc_7_10_i_q_d;
  wire [31:0] yt_rsc_7_11_i_q_d;
  wire [31:0] yt_rsc_7_12_i_q_d;
  wire [31:0] yt_rsc_7_13_i_q_d;
  wire [31:0] yt_rsc_7_14_i_q_d;
  wire [31:0] yt_rsc_7_15_i_q_d;
  wire yt_rsc_7_16_i_clkr_en_d;
  wire [31:0] yt_rsc_7_16_i_q_d;
  wire [31:0] yt_rsc_7_17_i_q_d;
  wire [31:0] yt_rsc_7_18_i_q_d;
  wire [31:0] yt_rsc_7_19_i_q_d;
  wire [31:0] yt_rsc_7_20_i_q_d;
  wire [31:0] yt_rsc_7_21_i_q_d;
  wire [31:0] yt_rsc_7_22_i_q_d;
  wire [31:0] yt_rsc_7_23_i_q_d;
  wire [31:0] yt_rsc_7_24_i_q_d;
  wire [31:0] yt_rsc_7_25_i_q_d;
  wire [31:0] yt_rsc_7_26_i_q_d;
  wire [31:0] yt_rsc_7_27_i_q_d;
  wire [31:0] yt_rsc_7_28_i_q_d;
  wire [31:0] yt_rsc_7_29_i_q_d;
  wire [31:0] yt_rsc_7_30_i_q_d;
  wire [31:0] yt_rsc_7_31_i_q_d;
  wire [31:0] xt_rsc_0_0_i_qa_d;
  wire [31:0] xt_rsc_0_1_i_qa_d;
  wire [31:0] xt_rsc_0_2_i_qa_d;
  wire [31:0] xt_rsc_0_3_i_qa_d;
  wire [31:0] xt_rsc_0_4_i_qa_d;
  wire [31:0] xt_rsc_0_5_i_qa_d;
  wire [31:0] xt_rsc_0_6_i_qa_d;
  wire [31:0] xt_rsc_0_7_i_qa_d;
  wire [31:0] xt_rsc_0_8_i_qa_d;
  wire [31:0] xt_rsc_0_9_i_qa_d;
  wire [31:0] xt_rsc_0_10_i_qa_d;
  wire [31:0] xt_rsc_0_11_i_qa_d;
  wire [31:0] xt_rsc_0_12_i_qa_d;
  wire [31:0] xt_rsc_0_13_i_qa_d;
  wire [31:0] xt_rsc_0_14_i_qa_d;
  wire [31:0] xt_rsc_0_15_i_qa_d;
  wire [31:0] xt_rsc_0_16_i_qa_d;
  wire [31:0] xt_rsc_0_17_i_qa_d;
  wire [31:0] xt_rsc_0_18_i_qa_d;
  wire [31:0] xt_rsc_0_19_i_qa_d;
  wire [31:0] xt_rsc_0_20_i_qa_d;
  wire [31:0] xt_rsc_0_21_i_qa_d;
  wire [31:0] xt_rsc_0_22_i_qa_d;
  wire [31:0] xt_rsc_0_23_i_qa_d;
  wire [31:0] xt_rsc_0_24_i_qa_d;
  wire [31:0] xt_rsc_0_25_i_qa_d;
  wire [31:0] xt_rsc_0_26_i_qa_d;
  wire [31:0] xt_rsc_0_27_i_qa_d;
  wire [31:0] xt_rsc_0_28_i_qa_d;
  wire [31:0] xt_rsc_0_29_i_qa_d;
  wire [31:0] xt_rsc_0_30_i_qa_d;
  wire [31:0] xt_rsc_0_31_i_qa_d;
  wire [31:0] xt_rsc_1_0_i_qa_d;
  wire [31:0] xt_rsc_1_1_i_qa_d;
  wire [31:0] xt_rsc_1_2_i_qa_d;
  wire [31:0] xt_rsc_1_3_i_qa_d;
  wire [31:0] xt_rsc_1_4_i_qa_d;
  wire [31:0] xt_rsc_1_5_i_qa_d;
  wire [31:0] xt_rsc_1_6_i_qa_d;
  wire [31:0] xt_rsc_1_7_i_qa_d;
  wire [31:0] xt_rsc_1_8_i_qa_d;
  wire [31:0] xt_rsc_1_9_i_qa_d;
  wire [31:0] xt_rsc_1_10_i_qa_d;
  wire [31:0] xt_rsc_1_11_i_qa_d;
  wire [31:0] xt_rsc_1_12_i_qa_d;
  wire [31:0] xt_rsc_1_13_i_qa_d;
  wire [31:0] xt_rsc_1_14_i_qa_d;
  wire [31:0] xt_rsc_1_15_i_qa_d;
  wire [31:0] xt_rsc_1_16_i_qa_d;
  wire [31:0] xt_rsc_1_17_i_qa_d;
  wire [31:0] xt_rsc_1_18_i_qa_d;
  wire [31:0] xt_rsc_1_19_i_qa_d;
  wire [31:0] xt_rsc_1_20_i_qa_d;
  wire [31:0] xt_rsc_1_21_i_qa_d;
  wire [31:0] xt_rsc_1_22_i_qa_d;
  wire [31:0] xt_rsc_1_23_i_qa_d;
  wire [31:0] xt_rsc_1_24_i_qa_d;
  wire [31:0] xt_rsc_1_25_i_qa_d;
  wire [31:0] xt_rsc_1_26_i_qa_d;
  wire [31:0] xt_rsc_1_27_i_qa_d;
  wire [31:0] xt_rsc_1_28_i_qa_d;
  wire [31:0] xt_rsc_1_29_i_qa_d;
  wire [31:0] xt_rsc_1_30_i_qa_d;
  wire [31:0] xt_rsc_1_31_i_qa_d;
  wire [31:0] xt_rsc_2_0_i_qa_d;
  wire [31:0] xt_rsc_2_1_i_qa_d;
  wire [31:0] xt_rsc_2_2_i_qa_d;
  wire [31:0] xt_rsc_2_3_i_qa_d;
  wire [31:0] xt_rsc_2_4_i_qa_d;
  wire [31:0] xt_rsc_2_5_i_qa_d;
  wire [31:0] xt_rsc_2_6_i_qa_d;
  wire [31:0] xt_rsc_2_7_i_qa_d;
  wire [31:0] xt_rsc_2_8_i_qa_d;
  wire [31:0] xt_rsc_2_9_i_qa_d;
  wire [31:0] xt_rsc_2_10_i_qa_d;
  wire [31:0] xt_rsc_2_11_i_qa_d;
  wire [31:0] xt_rsc_2_12_i_qa_d;
  wire [31:0] xt_rsc_2_13_i_qa_d;
  wire [31:0] xt_rsc_2_14_i_qa_d;
  wire [31:0] xt_rsc_2_15_i_qa_d;
  wire [31:0] xt_rsc_2_16_i_qa_d;
  wire [31:0] xt_rsc_2_17_i_qa_d;
  wire [31:0] xt_rsc_2_18_i_qa_d;
  wire [31:0] xt_rsc_2_19_i_qa_d;
  wire [31:0] xt_rsc_2_20_i_qa_d;
  wire [31:0] xt_rsc_2_21_i_qa_d;
  wire [31:0] xt_rsc_2_22_i_qa_d;
  wire [31:0] xt_rsc_2_23_i_qa_d;
  wire [31:0] xt_rsc_2_24_i_qa_d;
  wire [31:0] xt_rsc_2_25_i_qa_d;
  wire [31:0] xt_rsc_2_26_i_qa_d;
  wire [31:0] xt_rsc_2_27_i_qa_d;
  wire [31:0] xt_rsc_2_28_i_qa_d;
  wire [31:0] xt_rsc_2_29_i_qa_d;
  wire [31:0] xt_rsc_2_30_i_qa_d;
  wire [31:0] xt_rsc_2_31_i_qa_d;
  wire [31:0] xt_rsc_3_0_i_qa_d;
  wire [31:0] xt_rsc_3_1_i_qa_d;
  wire [31:0] xt_rsc_3_2_i_qa_d;
  wire [31:0] xt_rsc_3_3_i_qa_d;
  wire [31:0] xt_rsc_3_4_i_qa_d;
  wire [31:0] xt_rsc_3_5_i_qa_d;
  wire [31:0] xt_rsc_3_6_i_qa_d;
  wire [31:0] xt_rsc_3_7_i_qa_d;
  wire [31:0] xt_rsc_3_8_i_qa_d;
  wire [31:0] xt_rsc_3_9_i_qa_d;
  wire [31:0] xt_rsc_3_10_i_qa_d;
  wire [31:0] xt_rsc_3_11_i_qa_d;
  wire [31:0] xt_rsc_3_12_i_qa_d;
  wire [31:0] xt_rsc_3_13_i_qa_d;
  wire [31:0] xt_rsc_3_14_i_qa_d;
  wire [31:0] xt_rsc_3_15_i_qa_d;
  wire [31:0] xt_rsc_3_16_i_qa_d;
  wire [31:0] xt_rsc_3_17_i_qa_d;
  wire [31:0] xt_rsc_3_18_i_qa_d;
  wire [31:0] xt_rsc_3_19_i_qa_d;
  wire [31:0] xt_rsc_3_20_i_qa_d;
  wire [31:0] xt_rsc_3_21_i_qa_d;
  wire [31:0] xt_rsc_3_22_i_qa_d;
  wire [31:0] xt_rsc_3_23_i_qa_d;
  wire [31:0] xt_rsc_3_24_i_qa_d;
  wire [31:0] xt_rsc_3_25_i_qa_d;
  wire [31:0] xt_rsc_3_26_i_qa_d;
  wire [31:0] xt_rsc_3_27_i_qa_d;
  wire [31:0] xt_rsc_3_28_i_qa_d;
  wire [31:0] xt_rsc_3_29_i_qa_d;
  wire [31:0] xt_rsc_3_30_i_qa_d;
  wire [31:0] xt_rsc_3_31_i_qa_d;
  wire [31:0] xt_rsc_4_0_i_qa_d;
  wire [31:0] xt_rsc_4_1_i_qa_d;
  wire [31:0] xt_rsc_4_2_i_qa_d;
  wire [31:0] xt_rsc_4_3_i_qa_d;
  wire [31:0] xt_rsc_4_4_i_qa_d;
  wire [31:0] xt_rsc_4_5_i_qa_d;
  wire [31:0] xt_rsc_4_6_i_qa_d;
  wire [31:0] xt_rsc_4_7_i_qa_d;
  wire [31:0] xt_rsc_4_8_i_qa_d;
  wire [31:0] xt_rsc_4_9_i_qa_d;
  wire [31:0] xt_rsc_4_10_i_qa_d;
  wire [31:0] xt_rsc_4_11_i_qa_d;
  wire [31:0] xt_rsc_4_12_i_qa_d;
  wire [31:0] xt_rsc_4_13_i_qa_d;
  wire [31:0] xt_rsc_4_14_i_qa_d;
  wire [31:0] xt_rsc_4_15_i_qa_d;
  wire [31:0] xt_rsc_4_16_i_qa_d;
  wire [31:0] xt_rsc_4_17_i_qa_d;
  wire [31:0] xt_rsc_4_18_i_qa_d;
  wire [31:0] xt_rsc_4_19_i_qa_d;
  wire [31:0] xt_rsc_4_20_i_qa_d;
  wire [31:0] xt_rsc_4_21_i_qa_d;
  wire [31:0] xt_rsc_4_22_i_qa_d;
  wire [31:0] xt_rsc_4_23_i_qa_d;
  wire [31:0] xt_rsc_4_24_i_qa_d;
  wire [31:0] xt_rsc_4_25_i_qa_d;
  wire [31:0] xt_rsc_4_26_i_qa_d;
  wire [31:0] xt_rsc_4_27_i_qa_d;
  wire [31:0] xt_rsc_4_28_i_qa_d;
  wire [31:0] xt_rsc_4_29_i_qa_d;
  wire [31:0] xt_rsc_4_30_i_qa_d;
  wire [31:0] xt_rsc_4_31_i_qa_d;
  wire [31:0] xt_rsc_5_0_i_qa_d;
  wire [31:0] xt_rsc_5_1_i_qa_d;
  wire [31:0] xt_rsc_5_2_i_qa_d;
  wire [31:0] xt_rsc_5_3_i_qa_d;
  wire [31:0] xt_rsc_5_4_i_qa_d;
  wire [31:0] xt_rsc_5_5_i_qa_d;
  wire [31:0] xt_rsc_5_6_i_qa_d;
  wire [31:0] xt_rsc_5_7_i_qa_d;
  wire [31:0] xt_rsc_5_8_i_qa_d;
  wire [31:0] xt_rsc_5_9_i_qa_d;
  wire [31:0] xt_rsc_5_10_i_qa_d;
  wire [31:0] xt_rsc_5_11_i_qa_d;
  wire [31:0] xt_rsc_5_12_i_qa_d;
  wire [31:0] xt_rsc_5_13_i_qa_d;
  wire [31:0] xt_rsc_5_14_i_qa_d;
  wire [31:0] xt_rsc_5_15_i_qa_d;
  wire [31:0] xt_rsc_5_16_i_qa_d;
  wire [31:0] xt_rsc_5_17_i_qa_d;
  wire [31:0] xt_rsc_5_18_i_qa_d;
  wire [31:0] xt_rsc_5_19_i_qa_d;
  wire [31:0] xt_rsc_5_20_i_qa_d;
  wire [31:0] xt_rsc_5_21_i_qa_d;
  wire [31:0] xt_rsc_5_22_i_qa_d;
  wire [31:0] xt_rsc_5_23_i_qa_d;
  wire [31:0] xt_rsc_5_24_i_qa_d;
  wire [31:0] xt_rsc_5_25_i_qa_d;
  wire [31:0] xt_rsc_5_26_i_qa_d;
  wire [31:0] xt_rsc_5_27_i_qa_d;
  wire [31:0] xt_rsc_5_28_i_qa_d;
  wire [31:0] xt_rsc_5_29_i_qa_d;
  wire [31:0] xt_rsc_5_30_i_qa_d;
  wire [31:0] xt_rsc_5_31_i_qa_d;
  wire [31:0] xt_rsc_6_0_i_qa_d;
  wire [31:0] xt_rsc_6_1_i_qa_d;
  wire [31:0] xt_rsc_6_2_i_qa_d;
  wire [31:0] xt_rsc_6_3_i_qa_d;
  wire [31:0] xt_rsc_6_4_i_qa_d;
  wire [31:0] xt_rsc_6_5_i_qa_d;
  wire [31:0] xt_rsc_6_6_i_qa_d;
  wire [31:0] xt_rsc_6_7_i_qa_d;
  wire [31:0] xt_rsc_6_8_i_qa_d;
  wire [31:0] xt_rsc_6_9_i_qa_d;
  wire [31:0] xt_rsc_6_10_i_qa_d;
  wire [31:0] xt_rsc_6_11_i_qa_d;
  wire [31:0] xt_rsc_6_12_i_qa_d;
  wire [31:0] xt_rsc_6_13_i_qa_d;
  wire [31:0] xt_rsc_6_14_i_qa_d;
  wire [31:0] xt_rsc_6_15_i_qa_d;
  wire [31:0] xt_rsc_6_16_i_qa_d;
  wire [31:0] xt_rsc_6_17_i_qa_d;
  wire [31:0] xt_rsc_6_18_i_qa_d;
  wire [31:0] xt_rsc_6_19_i_qa_d;
  wire [31:0] xt_rsc_6_20_i_qa_d;
  wire [31:0] xt_rsc_6_21_i_qa_d;
  wire [31:0] xt_rsc_6_22_i_qa_d;
  wire [31:0] xt_rsc_6_23_i_qa_d;
  wire [31:0] xt_rsc_6_24_i_qa_d;
  wire [31:0] xt_rsc_6_25_i_qa_d;
  wire [31:0] xt_rsc_6_26_i_qa_d;
  wire [31:0] xt_rsc_6_27_i_qa_d;
  wire [31:0] xt_rsc_6_28_i_qa_d;
  wire [31:0] xt_rsc_6_29_i_qa_d;
  wire [31:0] xt_rsc_6_30_i_qa_d;
  wire [31:0] xt_rsc_6_31_i_qa_d;
  wire [31:0] xt_rsc_7_0_i_qa_d;
  wire [31:0] xt_rsc_7_1_i_qa_d;
  wire [31:0] xt_rsc_7_2_i_qa_d;
  wire [31:0] xt_rsc_7_3_i_qa_d;
  wire [31:0] xt_rsc_7_4_i_qa_d;
  wire [31:0] xt_rsc_7_5_i_qa_d;
  wire [31:0] xt_rsc_7_6_i_qa_d;
  wire [31:0] xt_rsc_7_7_i_qa_d;
  wire [31:0] xt_rsc_7_8_i_qa_d;
  wire [31:0] xt_rsc_7_9_i_qa_d;
  wire [31:0] xt_rsc_7_10_i_qa_d;
  wire [31:0] xt_rsc_7_11_i_qa_d;
  wire [31:0] xt_rsc_7_12_i_qa_d;
  wire [31:0] xt_rsc_7_13_i_qa_d;
  wire [31:0] xt_rsc_7_14_i_qa_d;
  wire [31:0] xt_rsc_7_15_i_qa_d;
  wire [31:0] xt_rsc_7_16_i_qa_d;
  wire [31:0] xt_rsc_7_17_i_qa_d;
  wire [31:0] xt_rsc_7_18_i_qa_d;
  wire [31:0] xt_rsc_7_19_i_qa_d;
  wire [31:0] xt_rsc_7_20_i_qa_d;
  wire [31:0] xt_rsc_7_21_i_qa_d;
  wire [31:0] xt_rsc_7_22_i_qa_d;
  wire [31:0] xt_rsc_7_23_i_qa_d;
  wire [31:0] xt_rsc_7_24_i_qa_d;
  wire [31:0] xt_rsc_7_25_i_qa_d;
  wire [31:0] xt_rsc_7_26_i_qa_d;
  wire [31:0] xt_rsc_7_27_i_qa_d;
  wire [31:0] xt_rsc_7_28_i_qa_d;
  wire [31:0] xt_rsc_7_29_i_qa_d;
  wire [31:0] xt_rsc_7_30_i_qa_d;
  wire [31:0] xt_rsc_7_31_i_qa_d;
  wire [7:0] twiddle_rsc_0_0_i_adra_d;
  wire [63:0] twiddle_rsc_0_0_i_qa_d;
  wire [1:0] twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_1_i_adra_d;
  wire [63:0] twiddle_rsc_0_1_i_qa_d;
  wire [1:0] twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_2_i_adra_d;
  wire [63:0] twiddle_rsc_0_2_i_qa_d;
  wire [1:0] twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_3_i_adra_d;
  wire [63:0] twiddle_rsc_0_3_i_qa_d;
  wire [1:0] twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_4_i_adra_d;
  wire [63:0] twiddle_rsc_0_4_i_qa_d;
  wire [1:0] twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_5_i_adra_d;
  wire [63:0] twiddle_rsc_0_5_i_qa_d;
  wire [1:0] twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_6_i_adra_d;
  wire [63:0] twiddle_rsc_0_6_i_qa_d;
  wire [1:0] twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_7_i_adra_d;
  wire [63:0] twiddle_rsc_0_7_i_qa_d;
  wire [1:0] twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_8_i_adra_d;
  wire [63:0] twiddle_rsc_0_8_i_qa_d;
  wire [1:0] twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_9_i_adra_d;
  wire [63:0] twiddle_rsc_0_9_i_qa_d;
  wire [1:0] twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_10_i_adra_d;
  wire [63:0] twiddle_rsc_0_10_i_qa_d;
  wire [1:0] twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_11_i_adra_d;
  wire [63:0] twiddle_rsc_0_11_i_qa_d;
  wire [1:0] twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_12_i_adra_d;
  wire [63:0] twiddle_rsc_0_12_i_qa_d;
  wire [1:0] twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_13_i_adra_d;
  wire [63:0] twiddle_rsc_0_13_i_qa_d;
  wire [1:0] twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_14_i_adra_d;
  wire [63:0] twiddle_rsc_0_14_i_qa_d;
  wire [1:0] twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_15_i_adra_d;
  wire [63:0] twiddle_rsc_0_15_i_qa_d;
  wire [1:0] twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_0_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_0_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_1_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_1_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_2_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_2_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_3_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_3_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_4_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_4_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_5_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_5_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_6_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_6_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_7_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_7_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_8_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_8_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_9_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_9_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_10_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_10_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_11_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_11_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_12_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_12_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_13_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_13_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_14_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_14_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_15_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_15_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire yt_rsc_0_0_clkr_en;
  wire yt_rsc_0_0_clkw_en;
  wire [31:0] yt_rsc_0_0_q;
  wire [3:0] yt_rsc_0_0_radr;
  wire yt_rsc_0_0_we;
  wire [31:0] yt_rsc_0_0_d;
  wire [3:0] yt_rsc_0_0_wadr;
  wire yt_rsc_0_1_clkr_en;
  wire yt_rsc_0_1_clkw_en;
  wire [31:0] yt_rsc_0_1_q;
  wire [3:0] yt_rsc_0_1_radr;
  wire yt_rsc_0_1_we;
  wire [31:0] yt_rsc_0_1_d;
  wire [3:0] yt_rsc_0_1_wadr;
  wire yt_rsc_0_2_clkr_en;
  wire yt_rsc_0_2_clkw_en;
  wire [31:0] yt_rsc_0_2_q;
  wire [3:0] yt_rsc_0_2_radr;
  wire yt_rsc_0_2_we;
  wire [31:0] yt_rsc_0_2_d;
  wire [3:0] yt_rsc_0_2_wadr;
  wire yt_rsc_0_3_clkr_en;
  wire yt_rsc_0_3_clkw_en;
  wire [31:0] yt_rsc_0_3_q;
  wire [3:0] yt_rsc_0_3_radr;
  wire yt_rsc_0_3_we;
  wire [31:0] yt_rsc_0_3_d;
  wire [3:0] yt_rsc_0_3_wadr;
  wire yt_rsc_0_4_clkr_en;
  wire yt_rsc_0_4_clkw_en;
  wire [31:0] yt_rsc_0_4_q;
  wire [3:0] yt_rsc_0_4_radr;
  wire yt_rsc_0_4_we;
  wire [31:0] yt_rsc_0_4_d;
  wire [3:0] yt_rsc_0_4_wadr;
  wire yt_rsc_0_5_clkr_en;
  wire yt_rsc_0_5_clkw_en;
  wire [31:0] yt_rsc_0_5_q;
  wire [3:0] yt_rsc_0_5_radr;
  wire yt_rsc_0_5_we;
  wire [31:0] yt_rsc_0_5_d;
  wire [3:0] yt_rsc_0_5_wadr;
  wire yt_rsc_0_6_clkr_en;
  wire yt_rsc_0_6_clkw_en;
  wire [31:0] yt_rsc_0_6_q;
  wire [3:0] yt_rsc_0_6_radr;
  wire yt_rsc_0_6_we;
  wire [31:0] yt_rsc_0_6_d;
  wire [3:0] yt_rsc_0_6_wadr;
  wire yt_rsc_0_7_clkr_en;
  wire yt_rsc_0_7_clkw_en;
  wire [31:0] yt_rsc_0_7_q;
  wire [3:0] yt_rsc_0_7_radr;
  wire yt_rsc_0_7_we;
  wire [31:0] yt_rsc_0_7_d;
  wire [3:0] yt_rsc_0_7_wadr;
  wire yt_rsc_0_8_clkr_en;
  wire yt_rsc_0_8_clkw_en;
  wire [31:0] yt_rsc_0_8_q;
  wire [3:0] yt_rsc_0_8_radr;
  wire yt_rsc_0_8_we;
  wire [31:0] yt_rsc_0_8_d;
  wire [3:0] yt_rsc_0_8_wadr;
  wire yt_rsc_0_9_clkr_en;
  wire yt_rsc_0_9_clkw_en;
  wire [31:0] yt_rsc_0_9_q;
  wire [3:0] yt_rsc_0_9_radr;
  wire yt_rsc_0_9_we;
  wire [31:0] yt_rsc_0_9_d;
  wire [3:0] yt_rsc_0_9_wadr;
  wire yt_rsc_0_10_clkr_en;
  wire yt_rsc_0_10_clkw_en;
  wire [31:0] yt_rsc_0_10_q;
  wire [3:0] yt_rsc_0_10_radr;
  wire yt_rsc_0_10_we;
  wire [31:0] yt_rsc_0_10_d;
  wire [3:0] yt_rsc_0_10_wadr;
  wire yt_rsc_0_11_clkr_en;
  wire yt_rsc_0_11_clkw_en;
  wire [31:0] yt_rsc_0_11_q;
  wire [3:0] yt_rsc_0_11_radr;
  wire yt_rsc_0_11_we;
  wire [31:0] yt_rsc_0_11_d;
  wire [3:0] yt_rsc_0_11_wadr;
  wire yt_rsc_0_12_clkr_en;
  wire yt_rsc_0_12_clkw_en;
  wire [31:0] yt_rsc_0_12_q;
  wire [3:0] yt_rsc_0_12_radr;
  wire yt_rsc_0_12_we;
  wire [31:0] yt_rsc_0_12_d;
  wire [3:0] yt_rsc_0_12_wadr;
  wire yt_rsc_0_13_clkr_en;
  wire yt_rsc_0_13_clkw_en;
  wire [31:0] yt_rsc_0_13_q;
  wire [3:0] yt_rsc_0_13_radr;
  wire yt_rsc_0_13_we;
  wire [31:0] yt_rsc_0_13_d;
  wire [3:0] yt_rsc_0_13_wadr;
  wire yt_rsc_0_14_clkr_en;
  wire yt_rsc_0_14_clkw_en;
  wire [31:0] yt_rsc_0_14_q;
  wire [3:0] yt_rsc_0_14_radr;
  wire yt_rsc_0_14_we;
  wire [31:0] yt_rsc_0_14_d;
  wire [3:0] yt_rsc_0_14_wadr;
  wire yt_rsc_0_15_clkr_en;
  wire yt_rsc_0_15_clkw_en;
  wire [31:0] yt_rsc_0_15_q;
  wire [3:0] yt_rsc_0_15_radr;
  wire yt_rsc_0_15_we;
  wire [31:0] yt_rsc_0_15_d;
  wire [3:0] yt_rsc_0_15_wadr;
  wire yt_rsc_0_16_clkr_en;
  wire yt_rsc_0_16_clkw_en;
  wire [31:0] yt_rsc_0_16_q;
  wire [3:0] yt_rsc_0_16_radr;
  wire yt_rsc_0_16_we;
  wire [31:0] yt_rsc_0_16_d;
  wire [3:0] yt_rsc_0_16_wadr;
  wire yt_rsc_0_17_clkr_en;
  wire yt_rsc_0_17_clkw_en;
  wire [31:0] yt_rsc_0_17_q;
  wire [3:0] yt_rsc_0_17_radr;
  wire yt_rsc_0_17_we;
  wire [31:0] yt_rsc_0_17_d;
  wire [3:0] yt_rsc_0_17_wadr;
  wire yt_rsc_0_18_clkr_en;
  wire yt_rsc_0_18_clkw_en;
  wire [31:0] yt_rsc_0_18_q;
  wire [3:0] yt_rsc_0_18_radr;
  wire yt_rsc_0_18_we;
  wire [31:0] yt_rsc_0_18_d;
  wire [3:0] yt_rsc_0_18_wadr;
  wire yt_rsc_0_19_clkr_en;
  wire yt_rsc_0_19_clkw_en;
  wire [31:0] yt_rsc_0_19_q;
  wire [3:0] yt_rsc_0_19_radr;
  wire yt_rsc_0_19_we;
  wire [31:0] yt_rsc_0_19_d;
  wire [3:0] yt_rsc_0_19_wadr;
  wire yt_rsc_0_20_clkr_en;
  wire yt_rsc_0_20_clkw_en;
  wire [31:0] yt_rsc_0_20_q;
  wire [3:0] yt_rsc_0_20_radr;
  wire yt_rsc_0_20_we;
  wire [31:0] yt_rsc_0_20_d;
  wire [3:0] yt_rsc_0_20_wadr;
  wire yt_rsc_0_21_clkr_en;
  wire yt_rsc_0_21_clkw_en;
  wire [31:0] yt_rsc_0_21_q;
  wire [3:0] yt_rsc_0_21_radr;
  wire yt_rsc_0_21_we;
  wire [31:0] yt_rsc_0_21_d;
  wire [3:0] yt_rsc_0_21_wadr;
  wire yt_rsc_0_22_clkr_en;
  wire yt_rsc_0_22_clkw_en;
  wire [31:0] yt_rsc_0_22_q;
  wire [3:0] yt_rsc_0_22_radr;
  wire yt_rsc_0_22_we;
  wire [31:0] yt_rsc_0_22_d;
  wire [3:0] yt_rsc_0_22_wadr;
  wire yt_rsc_0_23_clkr_en;
  wire yt_rsc_0_23_clkw_en;
  wire [31:0] yt_rsc_0_23_q;
  wire [3:0] yt_rsc_0_23_radr;
  wire yt_rsc_0_23_we;
  wire [31:0] yt_rsc_0_23_d;
  wire [3:0] yt_rsc_0_23_wadr;
  wire yt_rsc_0_24_clkr_en;
  wire yt_rsc_0_24_clkw_en;
  wire [31:0] yt_rsc_0_24_q;
  wire [3:0] yt_rsc_0_24_radr;
  wire yt_rsc_0_24_we;
  wire [31:0] yt_rsc_0_24_d;
  wire [3:0] yt_rsc_0_24_wadr;
  wire yt_rsc_0_25_clkr_en;
  wire yt_rsc_0_25_clkw_en;
  wire [31:0] yt_rsc_0_25_q;
  wire [3:0] yt_rsc_0_25_radr;
  wire yt_rsc_0_25_we;
  wire [31:0] yt_rsc_0_25_d;
  wire [3:0] yt_rsc_0_25_wadr;
  wire yt_rsc_0_26_clkr_en;
  wire yt_rsc_0_26_clkw_en;
  wire [31:0] yt_rsc_0_26_q;
  wire [3:0] yt_rsc_0_26_radr;
  wire yt_rsc_0_26_we;
  wire [31:0] yt_rsc_0_26_d;
  wire [3:0] yt_rsc_0_26_wadr;
  wire yt_rsc_0_27_clkr_en;
  wire yt_rsc_0_27_clkw_en;
  wire [31:0] yt_rsc_0_27_q;
  wire [3:0] yt_rsc_0_27_radr;
  wire yt_rsc_0_27_we;
  wire [31:0] yt_rsc_0_27_d;
  wire [3:0] yt_rsc_0_27_wadr;
  wire yt_rsc_0_28_clkr_en;
  wire yt_rsc_0_28_clkw_en;
  wire [31:0] yt_rsc_0_28_q;
  wire [3:0] yt_rsc_0_28_radr;
  wire yt_rsc_0_28_we;
  wire [31:0] yt_rsc_0_28_d;
  wire [3:0] yt_rsc_0_28_wadr;
  wire yt_rsc_0_29_clkr_en;
  wire yt_rsc_0_29_clkw_en;
  wire [31:0] yt_rsc_0_29_q;
  wire [3:0] yt_rsc_0_29_radr;
  wire yt_rsc_0_29_we;
  wire [31:0] yt_rsc_0_29_d;
  wire [3:0] yt_rsc_0_29_wadr;
  wire yt_rsc_0_30_clkr_en;
  wire yt_rsc_0_30_clkw_en;
  wire [31:0] yt_rsc_0_30_q;
  wire [3:0] yt_rsc_0_30_radr;
  wire yt_rsc_0_30_we;
  wire [31:0] yt_rsc_0_30_d;
  wire [3:0] yt_rsc_0_30_wadr;
  wire yt_rsc_0_31_clkr_en;
  wire yt_rsc_0_31_clkw_en;
  wire [31:0] yt_rsc_0_31_q;
  wire [3:0] yt_rsc_0_31_radr;
  wire yt_rsc_0_31_we;
  wire [31:0] yt_rsc_0_31_d;
  wire [3:0] yt_rsc_0_31_wadr;
  wire yt_rsc_1_0_clkr_en;
  wire yt_rsc_1_0_clkw_en;
  wire [31:0] yt_rsc_1_0_q;
  wire [3:0] yt_rsc_1_0_radr;
  wire yt_rsc_1_0_we;
  wire [31:0] yt_rsc_1_0_d;
  wire [3:0] yt_rsc_1_0_wadr;
  wire yt_rsc_1_1_clkr_en;
  wire yt_rsc_1_1_clkw_en;
  wire [31:0] yt_rsc_1_1_q;
  wire [3:0] yt_rsc_1_1_radr;
  wire yt_rsc_1_1_we;
  wire [31:0] yt_rsc_1_1_d;
  wire [3:0] yt_rsc_1_1_wadr;
  wire yt_rsc_1_2_clkr_en;
  wire yt_rsc_1_2_clkw_en;
  wire [31:0] yt_rsc_1_2_q;
  wire [3:0] yt_rsc_1_2_radr;
  wire yt_rsc_1_2_we;
  wire [31:0] yt_rsc_1_2_d;
  wire [3:0] yt_rsc_1_2_wadr;
  wire yt_rsc_1_3_clkr_en;
  wire yt_rsc_1_3_clkw_en;
  wire [31:0] yt_rsc_1_3_q;
  wire [3:0] yt_rsc_1_3_radr;
  wire yt_rsc_1_3_we;
  wire [31:0] yt_rsc_1_3_d;
  wire [3:0] yt_rsc_1_3_wadr;
  wire yt_rsc_1_4_clkr_en;
  wire yt_rsc_1_4_clkw_en;
  wire [31:0] yt_rsc_1_4_q;
  wire [3:0] yt_rsc_1_4_radr;
  wire yt_rsc_1_4_we;
  wire [31:0] yt_rsc_1_4_d;
  wire [3:0] yt_rsc_1_4_wadr;
  wire yt_rsc_1_5_clkr_en;
  wire yt_rsc_1_5_clkw_en;
  wire [31:0] yt_rsc_1_5_q;
  wire [3:0] yt_rsc_1_5_radr;
  wire yt_rsc_1_5_we;
  wire [31:0] yt_rsc_1_5_d;
  wire [3:0] yt_rsc_1_5_wadr;
  wire yt_rsc_1_6_clkr_en;
  wire yt_rsc_1_6_clkw_en;
  wire [31:0] yt_rsc_1_6_q;
  wire [3:0] yt_rsc_1_6_radr;
  wire yt_rsc_1_6_we;
  wire [31:0] yt_rsc_1_6_d;
  wire [3:0] yt_rsc_1_6_wadr;
  wire yt_rsc_1_7_clkr_en;
  wire yt_rsc_1_7_clkw_en;
  wire [31:0] yt_rsc_1_7_q;
  wire [3:0] yt_rsc_1_7_radr;
  wire yt_rsc_1_7_we;
  wire [31:0] yt_rsc_1_7_d;
  wire [3:0] yt_rsc_1_7_wadr;
  wire yt_rsc_1_8_clkr_en;
  wire yt_rsc_1_8_clkw_en;
  wire [31:0] yt_rsc_1_8_q;
  wire [3:0] yt_rsc_1_8_radr;
  wire yt_rsc_1_8_we;
  wire [31:0] yt_rsc_1_8_d;
  wire [3:0] yt_rsc_1_8_wadr;
  wire yt_rsc_1_9_clkr_en;
  wire yt_rsc_1_9_clkw_en;
  wire [31:0] yt_rsc_1_9_q;
  wire [3:0] yt_rsc_1_9_radr;
  wire yt_rsc_1_9_we;
  wire [31:0] yt_rsc_1_9_d;
  wire [3:0] yt_rsc_1_9_wadr;
  wire yt_rsc_1_10_clkr_en;
  wire yt_rsc_1_10_clkw_en;
  wire [31:0] yt_rsc_1_10_q;
  wire [3:0] yt_rsc_1_10_radr;
  wire yt_rsc_1_10_we;
  wire [31:0] yt_rsc_1_10_d;
  wire [3:0] yt_rsc_1_10_wadr;
  wire yt_rsc_1_11_clkr_en;
  wire yt_rsc_1_11_clkw_en;
  wire [31:0] yt_rsc_1_11_q;
  wire [3:0] yt_rsc_1_11_radr;
  wire yt_rsc_1_11_we;
  wire [31:0] yt_rsc_1_11_d;
  wire [3:0] yt_rsc_1_11_wadr;
  wire yt_rsc_1_12_clkr_en;
  wire yt_rsc_1_12_clkw_en;
  wire [31:0] yt_rsc_1_12_q;
  wire [3:0] yt_rsc_1_12_radr;
  wire yt_rsc_1_12_we;
  wire [31:0] yt_rsc_1_12_d;
  wire [3:0] yt_rsc_1_12_wadr;
  wire yt_rsc_1_13_clkr_en;
  wire yt_rsc_1_13_clkw_en;
  wire [31:0] yt_rsc_1_13_q;
  wire [3:0] yt_rsc_1_13_radr;
  wire yt_rsc_1_13_we;
  wire [31:0] yt_rsc_1_13_d;
  wire [3:0] yt_rsc_1_13_wadr;
  wire yt_rsc_1_14_clkr_en;
  wire yt_rsc_1_14_clkw_en;
  wire [31:0] yt_rsc_1_14_q;
  wire [3:0] yt_rsc_1_14_radr;
  wire yt_rsc_1_14_we;
  wire [31:0] yt_rsc_1_14_d;
  wire [3:0] yt_rsc_1_14_wadr;
  wire yt_rsc_1_15_clkr_en;
  wire yt_rsc_1_15_clkw_en;
  wire [31:0] yt_rsc_1_15_q;
  wire [3:0] yt_rsc_1_15_radr;
  wire yt_rsc_1_15_we;
  wire [31:0] yt_rsc_1_15_d;
  wire [3:0] yt_rsc_1_15_wadr;
  wire yt_rsc_1_16_clkr_en;
  wire yt_rsc_1_16_clkw_en;
  wire [31:0] yt_rsc_1_16_q;
  wire [3:0] yt_rsc_1_16_radr;
  wire yt_rsc_1_16_we;
  wire [31:0] yt_rsc_1_16_d;
  wire [3:0] yt_rsc_1_16_wadr;
  wire yt_rsc_1_17_clkr_en;
  wire yt_rsc_1_17_clkw_en;
  wire [31:0] yt_rsc_1_17_q;
  wire [3:0] yt_rsc_1_17_radr;
  wire yt_rsc_1_17_we;
  wire [31:0] yt_rsc_1_17_d;
  wire [3:0] yt_rsc_1_17_wadr;
  wire yt_rsc_1_18_clkr_en;
  wire yt_rsc_1_18_clkw_en;
  wire [31:0] yt_rsc_1_18_q;
  wire [3:0] yt_rsc_1_18_radr;
  wire yt_rsc_1_18_we;
  wire [31:0] yt_rsc_1_18_d;
  wire [3:0] yt_rsc_1_18_wadr;
  wire yt_rsc_1_19_clkr_en;
  wire yt_rsc_1_19_clkw_en;
  wire [31:0] yt_rsc_1_19_q;
  wire [3:0] yt_rsc_1_19_radr;
  wire yt_rsc_1_19_we;
  wire [31:0] yt_rsc_1_19_d;
  wire [3:0] yt_rsc_1_19_wadr;
  wire yt_rsc_1_20_clkr_en;
  wire yt_rsc_1_20_clkw_en;
  wire [31:0] yt_rsc_1_20_q;
  wire [3:0] yt_rsc_1_20_radr;
  wire yt_rsc_1_20_we;
  wire [31:0] yt_rsc_1_20_d;
  wire [3:0] yt_rsc_1_20_wadr;
  wire yt_rsc_1_21_clkr_en;
  wire yt_rsc_1_21_clkw_en;
  wire [31:0] yt_rsc_1_21_q;
  wire [3:0] yt_rsc_1_21_radr;
  wire yt_rsc_1_21_we;
  wire [31:0] yt_rsc_1_21_d;
  wire [3:0] yt_rsc_1_21_wadr;
  wire yt_rsc_1_22_clkr_en;
  wire yt_rsc_1_22_clkw_en;
  wire [31:0] yt_rsc_1_22_q;
  wire [3:0] yt_rsc_1_22_radr;
  wire yt_rsc_1_22_we;
  wire [31:0] yt_rsc_1_22_d;
  wire [3:0] yt_rsc_1_22_wadr;
  wire yt_rsc_1_23_clkr_en;
  wire yt_rsc_1_23_clkw_en;
  wire [31:0] yt_rsc_1_23_q;
  wire [3:0] yt_rsc_1_23_radr;
  wire yt_rsc_1_23_we;
  wire [31:0] yt_rsc_1_23_d;
  wire [3:0] yt_rsc_1_23_wadr;
  wire yt_rsc_1_24_clkr_en;
  wire yt_rsc_1_24_clkw_en;
  wire [31:0] yt_rsc_1_24_q;
  wire [3:0] yt_rsc_1_24_radr;
  wire yt_rsc_1_24_we;
  wire [31:0] yt_rsc_1_24_d;
  wire [3:0] yt_rsc_1_24_wadr;
  wire yt_rsc_1_25_clkr_en;
  wire yt_rsc_1_25_clkw_en;
  wire [31:0] yt_rsc_1_25_q;
  wire [3:0] yt_rsc_1_25_radr;
  wire yt_rsc_1_25_we;
  wire [31:0] yt_rsc_1_25_d;
  wire [3:0] yt_rsc_1_25_wadr;
  wire yt_rsc_1_26_clkr_en;
  wire yt_rsc_1_26_clkw_en;
  wire [31:0] yt_rsc_1_26_q;
  wire [3:0] yt_rsc_1_26_radr;
  wire yt_rsc_1_26_we;
  wire [31:0] yt_rsc_1_26_d;
  wire [3:0] yt_rsc_1_26_wadr;
  wire yt_rsc_1_27_clkr_en;
  wire yt_rsc_1_27_clkw_en;
  wire [31:0] yt_rsc_1_27_q;
  wire [3:0] yt_rsc_1_27_radr;
  wire yt_rsc_1_27_we;
  wire [31:0] yt_rsc_1_27_d;
  wire [3:0] yt_rsc_1_27_wadr;
  wire yt_rsc_1_28_clkr_en;
  wire yt_rsc_1_28_clkw_en;
  wire [31:0] yt_rsc_1_28_q;
  wire [3:0] yt_rsc_1_28_radr;
  wire yt_rsc_1_28_we;
  wire [31:0] yt_rsc_1_28_d;
  wire [3:0] yt_rsc_1_28_wadr;
  wire yt_rsc_1_29_clkr_en;
  wire yt_rsc_1_29_clkw_en;
  wire [31:0] yt_rsc_1_29_q;
  wire [3:0] yt_rsc_1_29_radr;
  wire yt_rsc_1_29_we;
  wire [31:0] yt_rsc_1_29_d;
  wire [3:0] yt_rsc_1_29_wadr;
  wire yt_rsc_1_30_clkr_en;
  wire yt_rsc_1_30_clkw_en;
  wire [31:0] yt_rsc_1_30_q;
  wire [3:0] yt_rsc_1_30_radr;
  wire yt_rsc_1_30_we;
  wire [31:0] yt_rsc_1_30_d;
  wire [3:0] yt_rsc_1_30_wadr;
  wire yt_rsc_1_31_clkr_en;
  wire yt_rsc_1_31_clkw_en;
  wire [31:0] yt_rsc_1_31_q;
  wire [3:0] yt_rsc_1_31_radr;
  wire yt_rsc_1_31_we;
  wire [31:0] yt_rsc_1_31_d;
  wire [3:0] yt_rsc_1_31_wadr;
  wire yt_rsc_2_0_clkr_en;
  wire yt_rsc_2_0_clkw_en;
  wire [31:0] yt_rsc_2_0_q;
  wire [3:0] yt_rsc_2_0_radr;
  wire yt_rsc_2_0_we;
  wire [31:0] yt_rsc_2_0_d;
  wire [3:0] yt_rsc_2_0_wadr;
  wire yt_rsc_2_1_clkr_en;
  wire yt_rsc_2_1_clkw_en;
  wire [31:0] yt_rsc_2_1_q;
  wire [3:0] yt_rsc_2_1_radr;
  wire yt_rsc_2_1_we;
  wire [31:0] yt_rsc_2_1_d;
  wire [3:0] yt_rsc_2_1_wadr;
  wire yt_rsc_2_2_clkr_en;
  wire yt_rsc_2_2_clkw_en;
  wire [31:0] yt_rsc_2_2_q;
  wire [3:0] yt_rsc_2_2_radr;
  wire yt_rsc_2_2_we;
  wire [31:0] yt_rsc_2_2_d;
  wire [3:0] yt_rsc_2_2_wadr;
  wire yt_rsc_2_3_clkr_en;
  wire yt_rsc_2_3_clkw_en;
  wire [31:0] yt_rsc_2_3_q;
  wire [3:0] yt_rsc_2_3_radr;
  wire yt_rsc_2_3_we;
  wire [31:0] yt_rsc_2_3_d;
  wire [3:0] yt_rsc_2_3_wadr;
  wire yt_rsc_2_4_clkr_en;
  wire yt_rsc_2_4_clkw_en;
  wire [31:0] yt_rsc_2_4_q;
  wire [3:0] yt_rsc_2_4_radr;
  wire yt_rsc_2_4_we;
  wire [31:0] yt_rsc_2_4_d;
  wire [3:0] yt_rsc_2_4_wadr;
  wire yt_rsc_2_5_clkr_en;
  wire yt_rsc_2_5_clkw_en;
  wire [31:0] yt_rsc_2_5_q;
  wire [3:0] yt_rsc_2_5_radr;
  wire yt_rsc_2_5_we;
  wire [31:0] yt_rsc_2_5_d;
  wire [3:0] yt_rsc_2_5_wadr;
  wire yt_rsc_2_6_clkr_en;
  wire yt_rsc_2_6_clkw_en;
  wire [31:0] yt_rsc_2_6_q;
  wire [3:0] yt_rsc_2_6_radr;
  wire yt_rsc_2_6_we;
  wire [31:0] yt_rsc_2_6_d;
  wire [3:0] yt_rsc_2_6_wadr;
  wire yt_rsc_2_7_clkr_en;
  wire yt_rsc_2_7_clkw_en;
  wire [31:0] yt_rsc_2_7_q;
  wire [3:0] yt_rsc_2_7_radr;
  wire yt_rsc_2_7_we;
  wire [31:0] yt_rsc_2_7_d;
  wire [3:0] yt_rsc_2_7_wadr;
  wire yt_rsc_2_8_clkr_en;
  wire yt_rsc_2_8_clkw_en;
  wire [31:0] yt_rsc_2_8_q;
  wire [3:0] yt_rsc_2_8_radr;
  wire yt_rsc_2_8_we;
  wire [31:0] yt_rsc_2_8_d;
  wire [3:0] yt_rsc_2_8_wadr;
  wire yt_rsc_2_9_clkr_en;
  wire yt_rsc_2_9_clkw_en;
  wire [31:0] yt_rsc_2_9_q;
  wire [3:0] yt_rsc_2_9_radr;
  wire yt_rsc_2_9_we;
  wire [31:0] yt_rsc_2_9_d;
  wire [3:0] yt_rsc_2_9_wadr;
  wire yt_rsc_2_10_clkr_en;
  wire yt_rsc_2_10_clkw_en;
  wire [31:0] yt_rsc_2_10_q;
  wire [3:0] yt_rsc_2_10_radr;
  wire yt_rsc_2_10_we;
  wire [31:0] yt_rsc_2_10_d;
  wire [3:0] yt_rsc_2_10_wadr;
  wire yt_rsc_2_11_clkr_en;
  wire yt_rsc_2_11_clkw_en;
  wire [31:0] yt_rsc_2_11_q;
  wire [3:0] yt_rsc_2_11_radr;
  wire yt_rsc_2_11_we;
  wire [31:0] yt_rsc_2_11_d;
  wire [3:0] yt_rsc_2_11_wadr;
  wire yt_rsc_2_12_clkr_en;
  wire yt_rsc_2_12_clkw_en;
  wire [31:0] yt_rsc_2_12_q;
  wire [3:0] yt_rsc_2_12_radr;
  wire yt_rsc_2_12_we;
  wire [31:0] yt_rsc_2_12_d;
  wire [3:0] yt_rsc_2_12_wadr;
  wire yt_rsc_2_13_clkr_en;
  wire yt_rsc_2_13_clkw_en;
  wire [31:0] yt_rsc_2_13_q;
  wire [3:0] yt_rsc_2_13_radr;
  wire yt_rsc_2_13_we;
  wire [31:0] yt_rsc_2_13_d;
  wire [3:0] yt_rsc_2_13_wadr;
  wire yt_rsc_2_14_clkr_en;
  wire yt_rsc_2_14_clkw_en;
  wire [31:0] yt_rsc_2_14_q;
  wire [3:0] yt_rsc_2_14_radr;
  wire yt_rsc_2_14_we;
  wire [31:0] yt_rsc_2_14_d;
  wire [3:0] yt_rsc_2_14_wadr;
  wire yt_rsc_2_15_clkr_en;
  wire yt_rsc_2_15_clkw_en;
  wire [31:0] yt_rsc_2_15_q;
  wire [3:0] yt_rsc_2_15_radr;
  wire yt_rsc_2_15_we;
  wire [31:0] yt_rsc_2_15_d;
  wire [3:0] yt_rsc_2_15_wadr;
  wire yt_rsc_2_16_clkr_en;
  wire yt_rsc_2_16_clkw_en;
  wire [31:0] yt_rsc_2_16_q;
  wire [3:0] yt_rsc_2_16_radr;
  wire yt_rsc_2_16_we;
  wire [31:0] yt_rsc_2_16_d;
  wire [3:0] yt_rsc_2_16_wadr;
  wire yt_rsc_2_17_clkr_en;
  wire yt_rsc_2_17_clkw_en;
  wire [31:0] yt_rsc_2_17_q;
  wire [3:0] yt_rsc_2_17_radr;
  wire yt_rsc_2_17_we;
  wire [31:0] yt_rsc_2_17_d;
  wire [3:0] yt_rsc_2_17_wadr;
  wire yt_rsc_2_18_clkr_en;
  wire yt_rsc_2_18_clkw_en;
  wire [31:0] yt_rsc_2_18_q;
  wire [3:0] yt_rsc_2_18_radr;
  wire yt_rsc_2_18_we;
  wire [31:0] yt_rsc_2_18_d;
  wire [3:0] yt_rsc_2_18_wadr;
  wire yt_rsc_2_19_clkr_en;
  wire yt_rsc_2_19_clkw_en;
  wire [31:0] yt_rsc_2_19_q;
  wire [3:0] yt_rsc_2_19_radr;
  wire yt_rsc_2_19_we;
  wire [31:0] yt_rsc_2_19_d;
  wire [3:0] yt_rsc_2_19_wadr;
  wire yt_rsc_2_20_clkr_en;
  wire yt_rsc_2_20_clkw_en;
  wire [31:0] yt_rsc_2_20_q;
  wire [3:0] yt_rsc_2_20_radr;
  wire yt_rsc_2_20_we;
  wire [31:0] yt_rsc_2_20_d;
  wire [3:0] yt_rsc_2_20_wadr;
  wire yt_rsc_2_21_clkr_en;
  wire yt_rsc_2_21_clkw_en;
  wire [31:0] yt_rsc_2_21_q;
  wire [3:0] yt_rsc_2_21_radr;
  wire yt_rsc_2_21_we;
  wire [31:0] yt_rsc_2_21_d;
  wire [3:0] yt_rsc_2_21_wadr;
  wire yt_rsc_2_22_clkr_en;
  wire yt_rsc_2_22_clkw_en;
  wire [31:0] yt_rsc_2_22_q;
  wire [3:0] yt_rsc_2_22_radr;
  wire yt_rsc_2_22_we;
  wire [31:0] yt_rsc_2_22_d;
  wire [3:0] yt_rsc_2_22_wadr;
  wire yt_rsc_2_23_clkr_en;
  wire yt_rsc_2_23_clkw_en;
  wire [31:0] yt_rsc_2_23_q;
  wire [3:0] yt_rsc_2_23_radr;
  wire yt_rsc_2_23_we;
  wire [31:0] yt_rsc_2_23_d;
  wire [3:0] yt_rsc_2_23_wadr;
  wire yt_rsc_2_24_clkr_en;
  wire yt_rsc_2_24_clkw_en;
  wire [31:0] yt_rsc_2_24_q;
  wire [3:0] yt_rsc_2_24_radr;
  wire yt_rsc_2_24_we;
  wire [31:0] yt_rsc_2_24_d;
  wire [3:0] yt_rsc_2_24_wadr;
  wire yt_rsc_2_25_clkr_en;
  wire yt_rsc_2_25_clkw_en;
  wire [31:0] yt_rsc_2_25_q;
  wire [3:0] yt_rsc_2_25_radr;
  wire yt_rsc_2_25_we;
  wire [31:0] yt_rsc_2_25_d;
  wire [3:0] yt_rsc_2_25_wadr;
  wire yt_rsc_2_26_clkr_en;
  wire yt_rsc_2_26_clkw_en;
  wire [31:0] yt_rsc_2_26_q;
  wire [3:0] yt_rsc_2_26_radr;
  wire yt_rsc_2_26_we;
  wire [31:0] yt_rsc_2_26_d;
  wire [3:0] yt_rsc_2_26_wadr;
  wire yt_rsc_2_27_clkr_en;
  wire yt_rsc_2_27_clkw_en;
  wire [31:0] yt_rsc_2_27_q;
  wire [3:0] yt_rsc_2_27_radr;
  wire yt_rsc_2_27_we;
  wire [31:0] yt_rsc_2_27_d;
  wire [3:0] yt_rsc_2_27_wadr;
  wire yt_rsc_2_28_clkr_en;
  wire yt_rsc_2_28_clkw_en;
  wire [31:0] yt_rsc_2_28_q;
  wire [3:0] yt_rsc_2_28_radr;
  wire yt_rsc_2_28_we;
  wire [31:0] yt_rsc_2_28_d;
  wire [3:0] yt_rsc_2_28_wadr;
  wire yt_rsc_2_29_clkr_en;
  wire yt_rsc_2_29_clkw_en;
  wire [31:0] yt_rsc_2_29_q;
  wire [3:0] yt_rsc_2_29_radr;
  wire yt_rsc_2_29_we;
  wire [31:0] yt_rsc_2_29_d;
  wire [3:0] yt_rsc_2_29_wadr;
  wire yt_rsc_2_30_clkr_en;
  wire yt_rsc_2_30_clkw_en;
  wire [31:0] yt_rsc_2_30_q;
  wire [3:0] yt_rsc_2_30_radr;
  wire yt_rsc_2_30_we;
  wire [31:0] yt_rsc_2_30_d;
  wire [3:0] yt_rsc_2_30_wadr;
  wire yt_rsc_2_31_clkr_en;
  wire yt_rsc_2_31_clkw_en;
  wire [31:0] yt_rsc_2_31_q;
  wire [3:0] yt_rsc_2_31_radr;
  wire yt_rsc_2_31_we;
  wire [31:0] yt_rsc_2_31_d;
  wire [3:0] yt_rsc_2_31_wadr;
  wire yt_rsc_3_0_clkr_en;
  wire yt_rsc_3_0_clkw_en;
  wire [31:0] yt_rsc_3_0_q;
  wire [3:0] yt_rsc_3_0_radr;
  wire yt_rsc_3_0_we;
  wire [31:0] yt_rsc_3_0_d;
  wire [3:0] yt_rsc_3_0_wadr;
  wire yt_rsc_3_1_clkr_en;
  wire yt_rsc_3_1_clkw_en;
  wire [31:0] yt_rsc_3_1_q;
  wire [3:0] yt_rsc_3_1_radr;
  wire yt_rsc_3_1_we;
  wire [31:0] yt_rsc_3_1_d;
  wire [3:0] yt_rsc_3_1_wadr;
  wire yt_rsc_3_2_clkr_en;
  wire yt_rsc_3_2_clkw_en;
  wire [31:0] yt_rsc_3_2_q;
  wire [3:0] yt_rsc_3_2_radr;
  wire yt_rsc_3_2_we;
  wire [31:0] yt_rsc_3_2_d;
  wire [3:0] yt_rsc_3_2_wadr;
  wire yt_rsc_3_3_clkr_en;
  wire yt_rsc_3_3_clkw_en;
  wire [31:0] yt_rsc_3_3_q;
  wire [3:0] yt_rsc_3_3_radr;
  wire yt_rsc_3_3_we;
  wire [31:0] yt_rsc_3_3_d;
  wire [3:0] yt_rsc_3_3_wadr;
  wire yt_rsc_3_4_clkr_en;
  wire yt_rsc_3_4_clkw_en;
  wire [31:0] yt_rsc_3_4_q;
  wire [3:0] yt_rsc_3_4_radr;
  wire yt_rsc_3_4_we;
  wire [31:0] yt_rsc_3_4_d;
  wire [3:0] yt_rsc_3_4_wadr;
  wire yt_rsc_3_5_clkr_en;
  wire yt_rsc_3_5_clkw_en;
  wire [31:0] yt_rsc_3_5_q;
  wire [3:0] yt_rsc_3_5_radr;
  wire yt_rsc_3_5_we;
  wire [31:0] yt_rsc_3_5_d;
  wire [3:0] yt_rsc_3_5_wadr;
  wire yt_rsc_3_6_clkr_en;
  wire yt_rsc_3_6_clkw_en;
  wire [31:0] yt_rsc_3_6_q;
  wire [3:0] yt_rsc_3_6_radr;
  wire yt_rsc_3_6_we;
  wire [31:0] yt_rsc_3_6_d;
  wire [3:0] yt_rsc_3_6_wadr;
  wire yt_rsc_3_7_clkr_en;
  wire yt_rsc_3_7_clkw_en;
  wire [31:0] yt_rsc_3_7_q;
  wire [3:0] yt_rsc_3_7_radr;
  wire yt_rsc_3_7_we;
  wire [31:0] yt_rsc_3_7_d;
  wire [3:0] yt_rsc_3_7_wadr;
  wire yt_rsc_3_8_clkr_en;
  wire yt_rsc_3_8_clkw_en;
  wire [31:0] yt_rsc_3_8_q;
  wire [3:0] yt_rsc_3_8_radr;
  wire yt_rsc_3_8_we;
  wire [31:0] yt_rsc_3_8_d;
  wire [3:0] yt_rsc_3_8_wadr;
  wire yt_rsc_3_9_clkr_en;
  wire yt_rsc_3_9_clkw_en;
  wire [31:0] yt_rsc_3_9_q;
  wire [3:0] yt_rsc_3_9_radr;
  wire yt_rsc_3_9_we;
  wire [31:0] yt_rsc_3_9_d;
  wire [3:0] yt_rsc_3_9_wadr;
  wire yt_rsc_3_10_clkr_en;
  wire yt_rsc_3_10_clkw_en;
  wire [31:0] yt_rsc_3_10_q;
  wire [3:0] yt_rsc_3_10_radr;
  wire yt_rsc_3_10_we;
  wire [31:0] yt_rsc_3_10_d;
  wire [3:0] yt_rsc_3_10_wadr;
  wire yt_rsc_3_11_clkr_en;
  wire yt_rsc_3_11_clkw_en;
  wire [31:0] yt_rsc_3_11_q;
  wire [3:0] yt_rsc_3_11_radr;
  wire yt_rsc_3_11_we;
  wire [31:0] yt_rsc_3_11_d;
  wire [3:0] yt_rsc_3_11_wadr;
  wire yt_rsc_3_12_clkr_en;
  wire yt_rsc_3_12_clkw_en;
  wire [31:0] yt_rsc_3_12_q;
  wire [3:0] yt_rsc_3_12_radr;
  wire yt_rsc_3_12_we;
  wire [31:0] yt_rsc_3_12_d;
  wire [3:0] yt_rsc_3_12_wadr;
  wire yt_rsc_3_13_clkr_en;
  wire yt_rsc_3_13_clkw_en;
  wire [31:0] yt_rsc_3_13_q;
  wire [3:0] yt_rsc_3_13_radr;
  wire yt_rsc_3_13_we;
  wire [31:0] yt_rsc_3_13_d;
  wire [3:0] yt_rsc_3_13_wadr;
  wire yt_rsc_3_14_clkr_en;
  wire yt_rsc_3_14_clkw_en;
  wire [31:0] yt_rsc_3_14_q;
  wire [3:0] yt_rsc_3_14_radr;
  wire yt_rsc_3_14_we;
  wire [31:0] yt_rsc_3_14_d;
  wire [3:0] yt_rsc_3_14_wadr;
  wire yt_rsc_3_15_clkr_en;
  wire yt_rsc_3_15_clkw_en;
  wire [31:0] yt_rsc_3_15_q;
  wire [3:0] yt_rsc_3_15_radr;
  wire yt_rsc_3_15_we;
  wire [31:0] yt_rsc_3_15_d;
  wire [3:0] yt_rsc_3_15_wadr;
  wire yt_rsc_3_16_clkr_en;
  wire yt_rsc_3_16_clkw_en;
  wire [31:0] yt_rsc_3_16_q;
  wire [3:0] yt_rsc_3_16_radr;
  wire yt_rsc_3_16_we;
  wire [31:0] yt_rsc_3_16_d;
  wire [3:0] yt_rsc_3_16_wadr;
  wire yt_rsc_3_17_clkr_en;
  wire yt_rsc_3_17_clkw_en;
  wire [31:0] yt_rsc_3_17_q;
  wire [3:0] yt_rsc_3_17_radr;
  wire yt_rsc_3_17_we;
  wire [31:0] yt_rsc_3_17_d;
  wire [3:0] yt_rsc_3_17_wadr;
  wire yt_rsc_3_18_clkr_en;
  wire yt_rsc_3_18_clkw_en;
  wire [31:0] yt_rsc_3_18_q;
  wire [3:0] yt_rsc_3_18_radr;
  wire yt_rsc_3_18_we;
  wire [31:0] yt_rsc_3_18_d;
  wire [3:0] yt_rsc_3_18_wadr;
  wire yt_rsc_3_19_clkr_en;
  wire yt_rsc_3_19_clkw_en;
  wire [31:0] yt_rsc_3_19_q;
  wire [3:0] yt_rsc_3_19_radr;
  wire yt_rsc_3_19_we;
  wire [31:0] yt_rsc_3_19_d;
  wire [3:0] yt_rsc_3_19_wadr;
  wire yt_rsc_3_20_clkr_en;
  wire yt_rsc_3_20_clkw_en;
  wire [31:0] yt_rsc_3_20_q;
  wire [3:0] yt_rsc_3_20_radr;
  wire yt_rsc_3_20_we;
  wire [31:0] yt_rsc_3_20_d;
  wire [3:0] yt_rsc_3_20_wadr;
  wire yt_rsc_3_21_clkr_en;
  wire yt_rsc_3_21_clkw_en;
  wire [31:0] yt_rsc_3_21_q;
  wire [3:0] yt_rsc_3_21_radr;
  wire yt_rsc_3_21_we;
  wire [31:0] yt_rsc_3_21_d;
  wire [3:0] yt_rsc_3_21_wadr;
  wire yt_rsc_3_22_clkr_en;
  wire yt_rsc_3_22_clkw_en;
  wire [31:0] yt_rsc_3_22_q;
  wire [3:0] yt_rsc_3_22_radr;
  wire yt_rsc_3_22_we;
  wire [31:0] yt_rsc_3_22_d;
  wire [3:0] yt_rsc_3_22_wadr;
  wire yt_rsc_3_23_clkr_en;
  wire yt_rsc_3_23_clkw_en;
  wire [31:0] yt_rsc_3_23_q;
  wire [3:0] yt_rsc_3_23_radr;
  wire yt_rsc_3_23_we;
  wire [31:0] yt_rsc_3_23_d;
  wire [3:0] yt_rsc_3_23_wadr;
  wire yt_rsc_3_24_clkr_en;
  wire yt_rsc_3_24_clkw_en;
  wire [31:0] yt_rsc_3_24_q;
  wire [3:0] yt_rsc_3_24_radr;
  wire yt_rsc_3_24_we;
  wire [31:0] yt_rsc_3_24_d;
  wire [3:0] yt_rsc_3_24_wadr;
  wire yt_rsc_3_25_clkr_en;
  wire yt_rsc_3_25_clkw_en;
  wire [31:0] yt_rsc_3_25_q;
  wire [3:0] yt_rsc_3_25_radr;
  wire yt_rsc_3_25_we;
  wire [31:0] yt_rsc_3_25_d;
  wire [3:0] yt_rsc_3_25_wadr;
  wire yt_rsc_3_26_clkr_en;
  wire yt_rsc_3_26_clkw_en;
  wire [31:0] yt_rsc_3_26_q;
  wire [3:0] yt_rsc_3_26_radr;
  wire yt_rsc_3_26_we;
  wire [31:0] yt_rsc_3_26_d;
  wire [3:0] yt_rsc_3_26_wadr;
  wire yt_rsc_3_27_clkr_en;
  wire yt_rsc_3_27_clkw_en;
  wire [31:0] yt_rsc_3_27_q;
  wire [3:0] yt_rsc_3_27_radr;
  wire yt_rsc_3_27_we;
  wire [31:0] yt_rsc_3_27_d;
  wire [3:0] yt_rsc_3_27_wadr;
  wire yt_rsc_3_28_clkr_en;
  wire yt_rsc_3_28_clkw_en;
  wire [31:0] yt_rsc_3_28_q;
  wire [3:0] yt_rsc_3_28_radr;
  wire yt_rsc_3_28_we;
  wire [31:0] yt_rsc_3_28_d;
  wire [3:0] yt_rsc_3_28_wadr;
  wire yt_rsc_3_29_clkr_en;
  wire yt_rsc_3_29_clkw_en;
  wire [31:0] yt_rsc_3_29_q;
  wire [3:0] yt_rsc_3_29_radr;
  wire yt_rsc_3_29_we;
  wire [31:0] yt_rsc_3_29_d;
  wire [3:0] yt_rsc_3_29_wadr;
  wire yt_rsc_3_30_clkr_en;
  wire yt_rsc_3_30_clkw_en;
  wire [31:0] yt_rsc_3_30_q;
  wire [3:0] yt_rsc_3_30_radr;
  wire yt_rsc_3_30_we;
  wire [31:0] yt_rsc_3_30_d;
  wire [3:0] yt_rsc_3_30_wadr;
  wire yt_rsc_3_31_clkr_en;
  wire yt_rsc_3_31_clkw_en;
  wire [31:0] yt_rsc_3_31_q;
  wire [3:0] yt_rsc_3_31_radr;
  wire yt_rsc_3_31_we;
  wire [31:0] yt_rsc_3_31_d;
  wire [3:0] yt_rsc_3_31_wadr;
  wire yt_rsc_4_0_clkr_en;
  wire yt_rsc_4_0_clkw_en;
  wire [31:0] yt_rsc_4_0_q;
  wire [3:0] yt_rsc_4_0_radr;
  wire yt_rsc_4_0_we;
  wire [31:0] yt_rsc_4_0_d;
  wire [3:0] yt_rsc_4_0_wadr;
  wire yt_rsc_4_1_clkr_en;
  wire yt_rsc_4_1_clkw_en;
  wire [31:0] yt_rsc_4_1_q;
  wire [3:0] yt_rsc_4_1_radr;
  wire yt_rsc_4_1_we;
  wire [31:0] yt_rsc_4_1_d;
  wire [3:0] yt_rsc_4_1_wadr;
  wire yt_rsc_4_2_clkr_en;
  wire yt_rsc_4_2_clkw_en;
  wire [31:0] yt_rsc_4_2_q;
  wire [3:0] yt_rsc_4_2_radr;
  wire yt_rsc_4_2_we;
  wire [31:0] yt_rsc_4_2_d;
  wire [3:0] yt_rsc_4_2_wadr;
  wire yt_rsc_4_3_clkr_en;
  wire yt_rsc_4_3_clkw_en;
  wire [31:0] yt_rsc_4_3_q;
  wire [3:0] yt_rsc_4_3_radr;
  wire yt_rsc_4_3_we;
  wire [31:0] yt_rsc_4_3_d;
  wire [3:0] yt_rsc_4_3_wadr;
  wire yt_rsc_4_4_clkr_en;
  wire yt_rsc_4_4_clkw_en;
  wire [31:0] yt_rsc_4_4_q;
  wire [3:0] yt_rsc_4_4_radr;
  wire yt_rsc_4_4_we;
  wire [31:0] yt_rsc_4_4_d;
  wire [3:0] yt_rsc_4_4_wadr;
  wire yt_rsc_4_5_clkr_en;
  wire yt_rsc_4_5_clkw_en;
  wire [31:0] yt_rsc_4_5_q;
  wire [3:0] yt_rsc_4_5_radr;
  wire yt_rsc_4_5_we;
  wire [31:0] yt_rsc_4_5_d;
  wire [3:0] yt_rsc_4_5_wadr;
  wire yt_rsc_4_6_clkr_en;
  wire yt_rsc_4_6_clkw_en;
  wire [31:0] yt_rsc_4_6_q;
  wire [3:0] yt_rsc_4_6_radr;
  wire yt_rsc_4_6_we;
  wire [31:0] yt_rsc_4_6_d;
  wire [3:0] yt_rsc_4_6_wadr;
  wire yt_rsc_4_7_clkr_en;
  wire yt_rsc_4_7_clkw_en;
  wire [31:0] yt_rsc_4_7_q;
  wire [3:0] yt_rsc_4_7_radr;
  wire yt_rsc_4_7_we;
  wire [31:0] yt_rsc_4_7_d;
  wire [3:0] yt_rsc_4_7_wadr;
  wire yt_rsc_4_8_clkr_en;
  wire yt_rsc_4_8_clkw_en;
  wire [31:0] yt_rsc_4_8_q;
  wire [3:0] yt_rsc_4_8_radr;
  wire yt_rsc_4_8_we;
  wire [31:0] yt_rsc_4_8_d;
  wire [3:0] yt_rsc_4_8_wadr;
  wire yt_rsc_4_9_clkr_en;
  wire yt_rsc_4_9_clkw_en;
  wire [31:0] yt_rsc_4_9_q;
  wire [3:0] yt_rsc_4_9_radr;
  wire yt_rsc_4_9_we;
  wire [31:0] yt_rsc_4_9_d;
  wire [3:0] yt_rsc_4_9_wadr;
  wire yt_rsc_4_10_clkr_en;
  wire yt_rsc_4_10_clkw_en;
  wire [31:0] yt_rsc_4_10_q;
  wire [3:0] yt_rsc_4_10_radr;
  wire yt_rsc_4_10_we;
  wire [31:0] yt_rsc_4_10_d;
  wire [3:0] yt_rsc_4_10_wadr;
  wire yt_rsc_4_11_clkr_en;
  wire yt_rsc_4_11_clkw_en;
  wire [31:0] yt_rsc_4_11_q;
  wire [3:0] yt_rsc_4_11_radr;
  wire yt_rsc_4_11_we;
  wire [31:0] yt_rsc_4_11_d;
  wire [3:0] yt_rsc_4_11_wadr;
  wire yt_rsc_4_12_clkr_en;
  wire yt_rsc_4_12_clkw_en;
  wire [31:0] yt_rsc_4_12_q;
  wire [3:0] yt_rsc_4_12_radr;
  wire yt_rsc_4_12_we;
  wire [31:0] yt_rsc_4_12_d;
  wire [3:0] yt_rsc_4_12_wadr;
  wire yt_rsc_4_13_clkr_en;
  wire yt_rsc_4_13_clkw_en;
  wire [31:0] yt_rsc_4_13_q;
  wire [3:0] yt_rsc_4_13_radr;
  wire yt_rsc_4_13_we;
  wire [31:0] yt_rsc_4_13_d;
  wire [3:0] yt_rsc_4_13_wadr;
  wire yt_rsc_4_14_clkr_en;
  wire yt_rsc_4_14_clkw_en;
  wire [31:0] yt_rsc_4_14_q;
  wire [3:0] yt_rsc_4_14_radr;
  wire yt_rsc_4_14_we;
  wire [31:0] yt_rsc_4_14_d;
  wire [3:0] yt_rsc_4_14_wadr;
  wire yt_rsc_4_15_clkr_en;
  wire yt_rsc_4_15_clkw_en;
  wire [31:0] yt_rsc_4_15_q;
  wire [3:0] yt_rsc_4_15_radr;
  wire yt_rsc_4_15_we;
  wire [31:0] yt_rsc_4_15_d;
  wire [3:0] yt_rsc_4_15_wadr;
  wire yt_rsc_4_16_clkr_en;
  wire yt_rsc_4_16_clkw_en;
  wire [31:0] yt_rsc_4_16_q;
  wire [3:0] yt_rsc_4_16_radr;
  wire yt_rsc_4_16_we;
  wire [31:0] yt_rsc_4_16_d;
  wire [3:0] yt_rsc_4_16_wadr;
  wire yt_rsc_4_17_clkr_en;
  wire yt_rsc_4_17_clkw_en;
  wire [31:0] yt_rsc_4_17_q;
  wire [3:0] yt_rsc_4_17_radr;
  wire yt_rsc_4_17_we;
  wire [31:0] yt_rsc_4_17_d;
  wire [3:0] yt_rsc_4_17_wadr;
  wire yt_rsc_4_18_clkr_en;
  wire yt_rsc_4_18_clkw_en;
  wire [31:0] yt_rsc_4_18_q;
  wire [3:0] yt_rsc_4_18_radr;
  wire yt_rsc_4_18_we;
  wire [31:0] yt_rsc_4_18_d;
  wire [3:0] yt_rsc_4_18_wadr;
  wire yt_rsc_4_19_clkr_en;
  wire yt_rsc_4_19_clkw_en;
  wire [31:0] yt_rsc_4_19_q;
  wire [3:0] yt_rsc_4_19_radr;
  wire yt_rsc_4_19_we;
  wire [31:0] yt_rsc_4_19_d;
  wire [3:0] yt_rsc_4_19_wadr;
  wire yt_rsc_4_20_clkr_en;
  wire yt_rsc_4_20_clkw_en;
  wire [31:0] yt_rsc_4_20_q;
  wire [3:0] yt_rsc_4_20_radr;
  wire yt_rsc_4_20_we;
  wire [31:0] yt_rsc_4_20_d;
  wire [3:0] yt_rsc_4_20_wadr;
  wire yt_rsc_4_21_clkr_en;
  wire yt_rsc_4_21_clkw_en;
  wire [31:0] yt_rsc_4_21_q;
  wire [3:0] yt_rsc_4_21_radr;
  wire yt_rsc_4_21_we;
  wire [31:0] yt_rsc_4_21_d;
  wire [3:0] yt_rsc_4_21_wadr;
  wire yt_rsc_4_22_clkr_en;
  wire yt_rsc_4_22_clkw_en;
  wire [31:0] yt_rsc_4_22_q;
  wire [3:0] yt_rsc_4_22_radr;
  wire yt_rsc_4_22_we;
  wire [31:0] yt_rsc_4_22_d;
  wire [3:0] yt_rsc_4_22_wadr;
  wire yt_rsc_4_23_clkr_en;
  wire yt_rsc_4_23_clkw_en;
  wire [31:0] yt_rsc_4_23_q;
  wire [3:0] yt_rsc_4_23_radr;
  wire yt_rsc_4_23_we;
  wire [31:0] yt_rsc_4_23_d;
  wire [3:0] yt_rsc_4_23_wadr;
  wire yt_rsc_4_24_clkr_en;
  wire yt_rsc_4_24_clkw_en;
  wire [31:0] yt_rsc_4_24_q;
  wire [3:0] yt_rsc_4_24_radr;
  wire yt_rsc_4_24_we;
  wire [31:0] yt_rsc_4_24_d;
  wire [3:0] yt_rsc_4_24_wadr;
  wire yt_rsc_4_25_clkr_en;
  wire yt_rsc_4_25_clkw_en;
  wire [31:0] yt_rsc_4_25_q;
  wire [3:0] yt_rsc_4_25_radr;
  wire yt_rsc_4_25_we;
  wire [31:0] yt_rsc_4_25_d;
  wire [3:0] yt_rsc_4_25_wadr;
  wire yt_rsc_4_26_clkr_en;
  wire yt_rsc_4_26_clkw_en;
  wire [31:0] yt_rsc_4_26_q;
  wire [3:0] yt_rsc_4_26_radr;
  wire yt_rsc_4_26_we;
  wire [31:0] yt_rsc_4_26_d;
  wire [3:0] yt_rsc_4_26_wadr;
  wire yt_rsc_4_27_clkr_en;
  wire yt_rsc_4_27_clkw_en;
  wire [31:0] yt_rsc_4_27_q;
  wire [3:0] yt_rsc_4_27_radr;
  wire yt_rsc_4_27_we;
  wire [31:0] yt_rsc_4_27_d;
  wire [3:0] yt_rsc_4_27_wadr;
  wire yt_rsc_4_28_clkr_en;
  wire yt_rsc_4_28_clkw_en;
  wire [31:0] yt_rsc_4_28_q;
  wire [3:0] yt_rsc_4_28_radr;
  wire yt_rsc_4_28_we;
  wire [31:0] yt_rsc_4_28_d;
  wire [3:0] yt_rsc_4_28_wadr;
  wire yt_rsc_4_29_clkr_en;
  wire yt_rsc_4_29_clkw_en;
  wire [31:0] yt_rsc_4_29_q;
  wire [3:0] yt_rsc_4_29_radr;
  wire yt_rsc_4_29_we;
  wire [31:0] yt_rsc_4_29_d;
  wire [3:0] yt_rsc_4_29_wadr;
  wire yt_rsc_4_30_clkr_en;
  wire yt_rsc_4_30_clkw_en;
  wire [31:0] yt_rsc_4_30_q;
  wire [3:0] yt_rsc_4_30_radr;
  wire yt_rsc_4_30_we;
  wire [31:0] yt_rsc_4_30_d;
  wire [3:0] yt_rsc_4_30_wadr;
  wire yt_rsc_4_31_clkr_en;
  wire yt_rsc_4_31_clkw_en;
  wire [31:0] yt_rsc_4_31_q;
  wire [3:0] yt_rsc_4_31_radr;
  wire yt_rsc_4_31_we;
  wire [31:0] yt_rsc_4_31_d;
  wire [3:0] yt_rsc_4_31_wadr;
  wire yt_rsc_5_0_clkr_en;
  wire yt_rsc_5_0_clkw_en;
  wire [31:0] yt_rsc_5_0_q;
  wire [3:0] yt_rsc_5_0_radr;
  wire yt_rsc_5_0_we;
  wire [31:0] yt_rsc_5_0_d;
  wire [3:0] yt_rsc_5_0_wadr;
  wire yt_rsc_5_1_clkr_en;
  wire yt_rsc_5_1_clkw_en;
  wire [31:0] yt_rsc_5_1_q;
  wire [3:0] yt_rsc_5_1_radr;
  wire yt_rsc_5_1_we;
  wire [31:0] yt_rsc_5_1_d;
  wire [3:0] yt_rsc_5_1_wadr;
  wire yt_rsc_5_2_clkr_en;
  wire yt_rsc_5_2_clkw_en;
  wire [31:0] yt_rsc_5_2_q;
  wire [3:0] yt_rsc_5_2_radr;
  wire yt_rsc_5_2_we;
  wire [31:0] yt_rsc_5_2_d;
  wire [3:0] yt_rsc_5_2_wadr;
  wire yt_rsc_5_3_clkr_en;
  wire yt_rsc_5_3_clkw_en;
  wire [31:0] yt_rsc_5_3_q;
  wire [3:0] yt_rsc_5_3_radr;
  wire yt_rsc_5_3_we;
  wire [31:0] yt_rsc_5_3_d;
  wire [3:0] yt_rsc_5_3_wadr;
  wire yt_rsc_5_4_clkr_en;
  wire yt_rsc_5_4_clkw_en;
  wire [31:0] yt_rsc_5_4_q;
  wire [3:0] yt_rsc_5_4_radr;
  wire yt_rsc_5_4_we;
  wire [31:0] yt_rsc_5_4_d;
  wire [3:0] yt_rsc_5_4_wadr;
  wire yt_rsc_5_5_clkr_en;
  wire yt_rsc_5_5_clkw_en;
  wire [31:0] yt_rsc_5_5_q;
  wire [3:0] yt_rsc_5_5_radr;
  wire yt_rsc_5_5_we;
  wire [31:0] yt_rsc_5_5_d;
  wire [3:0] yt_rsc_5_5_wadr;
  wire yt_rsc_5_6_clkr_en;
  wire yt_rsc_5_6_clkw_en;
  wire [31:0] yt_rsc_5_6_q;
  wire [3:0] yt_rsc_5_6_radr;
  wire yt_rsc_5_6_we;
  wire [31:0] yt_rsc_5_6_d;
  wire [3:0] yt_rsc_5_6_wadr;
  wire yt_rsc_5_7_clkr_en;
  wire yt_rsc_5_7_clkw_en;
  wire [31:0] yt_rsc_5_7_q;
  wire [3:0] yt_rsc_5_7_radr;
  wire yt_rsc_5_7_we;
  wire [31:0] yt_rsc_5_7_d;
  wire [3:0] yt_rsc_5_7_wadr;
  wire yt_rsc_5_8_clkr_en;
  wire yt_rsc_5_8_clkw_en;
  wire [31:0] yt_rsc_5_8_q;
  wire [3:0] yt_rsc_5_8_radr;
  wire yt_rsc_5_8_we;
  wire [31:0] yt_rsc_5_8_d;
  wire [3:0] yt_rsc_5_8_wadr;
  wire yt_rsc_5_9_clkr_en;
  wire yt_rsc_5_9_clkw_en;
  wire [31:0] yt_rsc_5_9_q;
  wire [3:0] yt_rsc_5_9_radr;
  wire yt_rsc_5_9_we;
  wire [31:0] yt_rsc_5_9_d;
  wire [3:0] yt_rsc_5_9_wadr;
  wire yt_rsc_5_10_clkr_en;
  wire yt_rsc_5_10_clkw_en;
  wire [31:0] yt_rsc_5_10_q;
  wire [3:0] yt_rsc_5_10_radr;
  wire yt_rsc_5_10_we;
  wire [31:0] yt_rsc_5_10_d;
  wire [3:0] yt_rsc_5_10_wadr;
  wire yt_rsc_5_11_clkr_en;
  wire yt_rsc_5_11_clkw_en;
  wire [31:0] yt_rsc_5_11_q;
  wire [3:0] yt_rsc_5_11_radr;
  wire yt_rsc_5_11_we;
  wire [31:0] yt_rsc_5_11_d;
  wire [3:0] yt_rsc_5_11_wadr;
  wire yt_rsc_5_12_clkr_en;
  wire yt_rsc_5_12_clkw_en;
  wire [31:0] yt_rsc_5_12_q;
  wire [3:0] yt_rsc_5_12_radr;
  wire yt_rsc_5_12_we;
  wire [31:0] yt_rsc_5_12_d;
  wire [3:0] yt_rsc_5_12_wadr;
  wire yt_rsc_5_13_clkr_en;
  wire yt_rsc_5_13_clkw_en;
  wire [31:0] yt_rsc_5_13_q;
  wire [3:0] yt_rsc_5_13_radr;
  wire yt_rsc_5_13_we;
  wire [31:0] yt_rsc_5_13_d;
  wire [3:0] yt_rsc_5_13_wadr;
  wire yt_rsc_5_14_clkr_en;
  wire yt_rsc_5_14_clkw_en;
  wire [31:0] yt_rsc_5_14_q;
  wire [3:0] yt_rsc_5_14_radr;
  wire yt_rsc_5_14_we;
  wire [31:0] yt_rsc_5_14_d;
  wire [3:0] yt_rsc_5_14_wadr;
  wire yt_rsc_5_15_clkr_en;
  wire yt_rsc_5_15_clkw_en;
  wire [31:0] yt_rsc_5_15_q;
  wire [3:0] yt_rsc_5_15_radr;
  wire yt_rsc_5_15_we;
  wire [31:0] yt_rsc_5_15_d;
  wire [3:0] yt_rsc_5_15_wadr;
  wire yt_rsc_5_16_clkr_en;
  wire yt_rsc_5_16_clkw_en;
  wire [31:0] yt_rsc_5_16_q;
  wire [3:0] yt_rsc_5_16_radr;
  wire yt_rsc_5_16_we;
  wire [31:0] yt_rsc_5_16_d;
  wire [3:0] yt_rsc_5_16_wadr;
  wire yt_rsc_5_17_clkr_en;
  wire yt_rsc_5_17_clkw_en;
  wire [31:0] yt_rsc_5_17_q;
  wire [3:0] yt_rsc_5_17_radr;
  wire yt_rsc_5_17_we;
  wire [31:0] yt_rsc_5_17_d;
  wire [3:0] yt_rsc_5_17_wadr;
  wire yt_rsc_5_18_clkr_en;
  wire yt_rsc_5_18_clkw_en;
  wire [31:0] yt_rsc_5_18_q;
  wire [3:0] yt_rsc_5_18_radr;
  wire yt_rsc_5_18_we;
  wire [31:0] yt_rsc_5_18_d;
  wire [3:0] yt_rsc_5_18_wadr;
  wire yt_rsc_5_19_clkr_en;
  wire yt_rsc_5_19_clkw_en;
  wire [31:0] yt_rsc_5_19_q;
  wire [3:0] yt_rsc_5_19_radr;
  wire yt_rsc_5_19_we;
  wire [31:0] yt_rsc_5_19_d;
  wire [3:0] yt_rsc_5_19_wadr;
  wire yt_rsc_5_20_clkr_en;
  wire yt_rsc_5_20_clkw_en;
  wire [31:0] yt_rsc_5_20_q;
  wire [3:0] yt_rsc_5_20_radr;
  wire yt_rsc_5_20_we;
  wire [31:0] yt_rsc_5_20_d;
  wire [3:0] yt_rsc_5_20_wadr;
  wire yt_rsc_5_21_clkr_en;
  wire yt_rsc_5_21_clkw_en;
  wire [31:0] yt_rsc_5_21_q;
  wire [3:0] yt_rsc_5_21_radr;
  wire yt_rsc_5_21_we;
  wire [31:0] yt_rsc_5_21_d;
  wire [3:0] yt_rsc_5_21_wadr;
  wire yt_rsc_5_22_clkr_en;
  wire yt_rsc_5_22_clkw_en;
  wire [31:0] yt_rsc_5_22_q;
  wire [3:0] yt_rsc_5_22_radr;
  wire yt_rsc_5_22_we;
  wire [31:0] yt_rsc_5_22_d;
  wire [3:0] yt_rsc_5_22_wadr;
  wire yt_rsc_5_23_clkr_en;
  wire yt_rsc_5_23_clkw_en;
  wire [31:0] yt_rsc_5_23_q;
  wire [3:0] yt_rsc_5_23_radr;
  wire yt_rsc_5_23_we;
  wire [31:0] yt_rsc_5_23_d;
  wire [3:0] yt_rsc_5_23_wadr;
  wire yt_rsc_5_24_clkr_en;
  wire yt_rsc_5_24_clkw_en;
  wire [31:0] yt_rsc_5_24_q;
  wire [3:0] yt_rsc_5_24_radr;
  wire yt_rsc_5_24_we;
  wire [31:0] yt_rsc_5_24_d;
  wire [3:0] yt_rsc_5_24_wadr;
  wire yt_rsc_5_25_clkr_en;
  wire yt_rsc_5_25_clkw_en;
  wire [31:0] yt_rsc_5_25_q;
  wire [3:0] yt_rsc_5_25_radr;
  wire yt_rsc_5_25_we;
  wire [31:0] yt_rsc_5_25_d;
  wire [3:0] yt_rsc_5_25_wadr;
  wire yt_rsc_5_26_clkr_en;
  wire yt_rsc_5_26_clkw_en;
  wire [31:0] yt_rsc_5_26_q;
  wire [3:0] yt_rsc_5_26_radr;
  wire yt_rsc_5_26_we;
  wire [31:0] yt_rsc_5_26_d;
  wire [3:0] yt_rsc_5_26_wadr;
  wire yt_rsc_5_27_clkr_en;
  wire yt_rsc_5_27_clkw_en;
  wire [31:0] yt_rsc_5_27_q;
  wire [3:0] yt_rsc_5_27_radr;
  wire yt_rsc_5_27_we;
  wire [31:0] yt_rsc_5_27_d;
  wire [3:0] yt_rsc_5_27_wadr;
  wire yt_rsc_5_28_clkr_en;
  wire yt_rsc_5_28_clkw_en;
  wire [31:0] yt_rsc_5_28_q;
  wire [3:0] yt_rsc_5_28_radr;
  wire yt_rsc_5_28_we;
  wire [31:0] yt_rsc_5_28_d;
  wire [3:0] yt_rsc_5_28_wadr;
  wire yt_rsc_5_29_clkr_en;
  wire yt_rsc_5_29_clkw_en;
  wire [31:0] yt_rsc_5_29_q;
  wire [3:0] yt_rsc_5_29_radr;
  wire yt_rsc_5_29_we;
  wire [31:0] yt_rsc_5_29_d;
  wire [3:0] yt_rsc_5_29_wadr;
  wire yt_rsc_5_30_clkr_en;
  wire yt_rsc_5_30_clkw_en;
  wire [31:0] yt_rsc_5_30_q;
  wire [3:0] yt_rsc_5_30_radr;
  wire yt_rsc_5_30_we;
  wire [31:0] yt_rsc_5_30_d;
  wire [3:0] yt_rsc_5_30_wadr;
  wire yt_rsc_5_31_clkr_en;
  wire yt_rsc_5_31_clkw_en;
  wire [31:0] yt_rsc_5_31_q;
  wire [3:0] yt_rsc_5_31_radr;
  wire yt_rsc_5_31_we;
  wire [31:0] yt_rsc_5_31_d;
  wire [3:0] yt_rsc_5_31_wadr;
  wire yt_rsc_6_0_clkr_en;
  wire yt_rsc_6_0_clkw_en;
  wire [31:0] yt_rsc_6_0_q;
  wire [3:0] yt_rsc_6_0_radr;
  wire yt_rsc_6_0_we;
  wire [31:0] yt_rsc_6_0_d;
  wire [3:0] yt_rsc_6_0_wadr;
  wire yt_rsc_6_1_clkr_en;
  wire yt_rsc_6_1_clkw_en;
  wire [31:0] yt_rsc_6_1_q;
  wire [3:0] yt_rsc_6_1_radr;
  wire yt_rsc_6_1_we;
  wire [31:0] yt_rsc_6_1_d;
  wire [3:0] yt_rsc_6_1_wadr;
  wire yt_rsc_6_2_clkr_en;
  wire yt_rsc_6_2_clkw_en;
  wire [31:0] yt_rsc_6_2_q;
  wire [3:0] yt_rsc_6_2_radr;
  wire yt_rsc_6_2_we;
  wire [31:0] yt_rsc_6_2_d;
  wire [3:0] yt_rsc_6_2_wadr;
  wire yt_rsc_6_3_clkr_en;
  wire yt_rsc_6_3_clkw_en;
  wire [31:0] yt_rsc_6_3_q;
  wire [3:0] yt_rsc_6_3_radr;
  wire yt_rsc_6_3_we;
  wire [31:0] yt_rsc_6_3_d;
  wire [3:0] yt_rsc_6_3_wadr;
  wire yt_rsc_6_4_clkr_en;
  wire yt_rsc_6_4_clkw_en;
  wire [31:0] yt_rsc_6_4_q;
  wire [3:0] yt_rsc_6_4_radr;
  wire yt_rsc_6_4_we;
  wire [31:0] yt_rsc_6_4_d;
  wire [3:0] yt_rsc_6_4_wadr;
  wire yt_rsc_6_5_clkr_en;
  wire yt_rsc_6_5_clkw_en;
  wire [31:0] yt_rsc_6_5_q;
  wire [3:0] yt_rsc_6_5_radr;
  wire yt_rsc_6_5_we;
  wire [31:0] yt_rsc_6_5_d;
  wire [3:0] yt_rsc_6_5_wadr;
  wire yt_rsc_6_6_clkr_en;
  wire yt_rsc_6_6_clkw_en;
  wire [31:0] yt_rsc_6_6_q;
  wire [3:0] yt_rsc_6_6_radr;
  wire yt_rsc_6_6_we;
  wire [31:0] yt_rsc_6_6_d;
  wire [3:0] yt_rsc_6_6_wadr;
  wire yt_rsc_6_7_clkr_en;
  wire yt_rsc_6_7_clkw_en;
  wire [31:0] yt_rsc_6_7_q;
  wire [3:0] yt_rsc_6_7_radr;
  wire yt_rsc_6_7_we;
  wire [31:0] yt_rsc_6_7_d;
  wire [3:0] yt_rsc_6_7_wadr;
  wire yt_rsc_6_8_clkr_en;
  wire yt_rsc_6_8_clkw_en;
  wire [31:0] yt_rsc_6_8_q;
  wire [3:0] yt_rsc_6_8_radr;
  wire yt_rsc_6_8_we;
  wire [31:0] yt_rsc_6_8_d;
  wire [3:0] yt_rsc_6_8_wadr;
  wire yt_rsc_6_9_clkr_en;
  wire yt_rsc_6_9_clkw_en;
  wire [31:0] yt_rsc_6_9_q;
  wire [3:0] yt_rsc_6_9_radr;
  wire yt_rsc_6_9_we;
  wire [31:0] yt_rsc_6_9_d;
  wire [3:0] yt_rsc_6_9_wadr;
  wire yt_rsc_6_10_clkr_en;
  wire yt_rsc_6_10_clkw_en;
  wire [31:0] yt_rsc_6_10_q;
  wire [3:0] yt_rsc_6_10_radr;
  wire yt_rsc_6_10_we;
  wire [31:0] yt_rsc_6_10_d;
  wire [3:0] yt_rsc_6_10_wadr;
  wire yt_rsc_6_11_clkr_en;
  wire yt_rsc_6_11_clkw_en;
  wire [31:0] yt_rsc_6_11_q;
  wire [3:0] yt_rsc_6_11_radr;
  wire yt_rsc_6_11_we;
  wire [31:0] yt_rsc_6_11_d;
  wire [3:0] yt_rsc_6_11_wadr;
  wire yt_rsc_6_12_clkr_en;
  wire yt_rsc_6_12_clkw_en;
  wire [31:0] yt_rsc_6_12_q;
  wire [3:0] yt_rsc_6_12_radr;
  wire yt_rsc_6_12_we;
  wire [31:0] yt_rsc_6_12_d;
  wire [3:0] yt_rsc_6_12_wadr;
  wire yt_rsc_6_13_clkr_en;
  wire yt_rsc_6_13_clkw_en;
  wire [31:0] yt_rsc_6_13_q;
  wire [3:0] yt_rsc_6_13_radr;
  wire yt_rsc_6_13_we;
  wire [31:0] yt_rsc_6_13_d;
  wire [3:0] yt_rsc_6_13_wadr;
  wire yt_rsc_6_14_clkr_en;
  wire yt_rsc_6_14_clkw_en;
  wire [31:0] yt_rsc_6_14_q;
  wire [3:0] yt_rsc_6_14_radr;
  wire yt_rsc_6_14_we;
  wire [31:0] yt_rsc_6_14_d;
  wire [3:0] yt_rsc_6_14_wadr;
  wire yt_rsc_6_15_clkr_en;
  wire yt_rsc_6_15_clkw_en;
  wire [31:0] yt_rsc_6_15_q;
  wire [3:0] yt_rsc_6_15_radr;
  wire yt_rsc_6_15_we;
  wire [31:0] yt_rsc_6_15_d;
  wire [3:0] yt_rsc_6_15_wadr;
  wire yt_rsc_6_16_clkr_en;
  wire yt_rsc_6_16_clkw_en;
  wire [31:0] yt_rsc_6_16_q;
  wire [3:0] yt_rsc_6_16_radr;
  wire yt_rsc_6_16_we;
  wire [31:0] yt_rsc_6_16_d;
  wire [3:0] yt_rsc_6_16_wadr;
  wire yt_rsc_6_17_clkr_en;
  wire yt_rsc_6_17_clkw_en;
  wire [31:0] yt_rsc_6_17_q;
  wire [3:0] yt_rsc_6_17_radr;
  wire yt_rsc_6_17_we;
  wire [31:0] yt_rsc_6_17_d;
  wire [3:0] yt_rsc_6_17_wadr;
  wire yt_rsc_6_18_clkr_en;
  wire yt_rsc_6_18_clkw_en;
  wire [31:0] yt_rsc_6_18_q;
  wire [3:0] yt_rsc_6_18_radr;
  wire yt_rsc_6_18_we;
  wire [31:0] yt_rsc_6_18_d;
  wire [3:0] yt_rsc_6_18_wadr;
  wire yt_rsc_6_19_clkr_en;
  wire yt_rsc_6_19_clkw_en;
  wire [31:0] yt_rsc_6_19_q;
  wire [3:0] yt_rsc_6_19_radr;
  wire yt_rsc_6_19_we;
  wire [31:0] yt_rsc_6_19_d;
  wire [3:0] yt_rsc_6_19_wadr;
  wire yt_rsc_6_20_clkr_en;
  wire yt_rsc_6_20_clkw_en;
  wire [31:0] yt_rsc_6_20_q;
  wire [3:0] yt_rsc_6_20_radr;
  wire yt_rsc_6_20_we;
  wire [31:0] yt_rsc_6_20_d;
  wire [3:0] yt_rsc_6_20_wadr;
  wire yt_rsc_6_21_clkr_en;
  wire yt_rsc_6_21_clkw_en;
  wire [31:0] yt_rsc_6_21_q;
  wire [3:0] yt_rsc_6_21_radr;
  wire yt_rsc_6_21_we;
  wire [31:0] yt_rsc_6_21_d;
  wire [3:0] yt_rsc_6_21_wadr;
  wire yt_rsc_6_22_clkr_en;
  wire yt_rsc_6_22_clkw_en;
  wire [31:0] yt_rsc_6_22_q;
  wire [3:0] yt_rsc_6_22_radr;
  wire yt_rsc_6_22_we;
  wire [31:0] yt_rsc_6_22_d;
  wire [3:0] yt_rsc_6_22_wadr;
  wire yt_rsc_6_23_clkr_en;
  wire yt_rsc_6_23_clkw_en;
  wire [31:0] yt_rsc_6_23_q;
  wire [3:0] yt_rsc_6_23_radr;
  wire yt_rsc_6_23_we;
  wire [31:0] yt_rsc_6_23_d;
  wire [3:0] yt_rsc_6_23_wadr;
  wire yt_rsc_6_24_clkr_en;
  wire yt_rsc_6_24_clkw_en;
  wire [31:0] yt_rsc_6_24_q;
  wire [3:0] yt_rsc_6_24_radr;
  wire yt_rsc_6_24_we;
  wire [31:0] yt_rsc_6_24_d;
  wire [3:0] yt_rsc_6_24_wadr;
  wire yt_rsc_6_25_clkr_en;
  wire yt_rsc_6_25_clkw_en;
  wire [31:0] yt_rsc_6_25_q;
  wire [3:0] yt_rsc_6_25_radr;
  wire yt_rsc_6_25_we;
  wire [31:0] yt_rsc_6_25_d;
  wire [3:0] yt_rsc_6_25_wadr;
  wire yt_rsc_6_26_clkr_en;
  wire yt_rsc_6_26_clkw_en;
  wire [31:0] yt_rsc_6_26_q;
  wire [3:0] yt_rsc_6_26_radr;
  wire yt_rsc_6_26_we;
  wire [31:0] yt_rsc_6_26_d;
  wire [3:0] yt_rsc_6_26_wadr;
  wire yt_rsc_6_27_clkr_en;
  wire yt_rsc_6_27_clkw_en;
  wire [31:0] yt_rsc_6_27_q;
  wire [3:0] yt_rsc_6_27_radr;
  wire yt_rsc_6_27_we;
  wire [31:0] yt_rsc_6_27_d;
  wire [3:0] yt_rsc_6_27_wadr;
  wire yt_rsc_6_28_clkr_en;
  wire yt_rsc_6_28_clkw_en;
  wire [31:0] yt_rsc_6_28_q;
  wire [3:0] yt_rsc_6_28_radr;
  wire yt_rsc_6_28_we;
  wire [31:0] yt_rsc_6_28_d;
  wire [3:0] yt_rsc_6_28_wadr;
  wire yt_rsc_6_29_clkr_en;
  wire yt_rsc_6_29_clkw_en;
  wire [31:0] yt_rsc_6_29_q;
  wire [3:0] yt_rsc_6_29_radr;
  wire yt_rsc_6_29_we;
  wire [31:0] yt_rsc_6_29_d;
  wire [3:0] yt_rsc_6_29_wadr;
  wire yt_rsc_6_30_clkr_en;
  wire yt_rsc_6_30_clkw_en;
  wire [31:0] yt_rsc_6_30_q;
  wire [3:0] yt_rsc_6_30_radr;
  wire yt_rsc_6_30_we;
  wire [31:0] yt_rsc_6_30_d;
  wire [3:0] yt_rsc_6_30_wadr;
  wire yt_rsc_6_31_clkr_en;
  wire yt_rsc_6_31_clkw_en;
  wire [31:0] yt_rsc_6_31_q;
  wire [3:0] yt_rsc_6_31_radr;
  wire yt_rsc_6_31_we;
  wire [31:0] yt_rsc_6_31_d;
  wire [3:0] yt_rsc_6_31_wadr;
  wire yt_rsc_7_0_clkr_en;
  wire yt_rsc_7_0_clkw_en;
  wire [31:0] yt_rsc_7_0_q;
  wire [3:0] yt_rsc_7_0_radr;
  wire yt_rsc_7_0_we;
  wire [31:0] yt_rsc_7_0_d;
  wire [3:0] yt_rsc_7_0_wadr;
  wire yt_rsc_7_1_clkr_en;
  wire yt_rsc_7_1_clkw_en;
  wire [31:0] yt_rsc_7_1_q;
  wire [3:0] yt_rsc_7_1_radr;
  wire yt_rsc_7_1_we;
  wire [31:0] yt_rsc_7_1_d;
  wire [3:0] yt_rsc_7_1_wadr;
  wire yt_rsc_7_2_clkr_en;
  wire yt_rsc_7_2_clkw_en;
  wire [31:0] yt_rsc_7_2_q;
  wire [3:0] yt_rsc_7_2_radr;
  wire yt_rsc_7_2_we;
  wire [31:0] yt_rsc_7_2_d;
  wire [3:0] yt_rsc_7_2_wadr;
  wire yt_rsc_7_3_clkr_en;
  wire yt_rsc_7_3_clkw_en;
  wire [31:0] yt_rsc_7_3_q;
  wire [3:0] yt_rsc_7_3_radr;
  wire yt_rsc_7_3_we;
  wire [31:0] yt_rsc_7_3_d;
  wire [3:0] yt_rsc_7_3_wadr;
  wire yt_rsc_7_4_clkr_en;
  wire yt_rsc_7_4_clkw_en;
  wire [31:0] yt_rsc_7_4_q;
  wire [3:0] yt_rsc_7_4_radr;
  wire yt_rsc_7_4_we;
  wire [31:0] yt_rsc_7_4_d;
  wire [3:0] yt_rsc_7_4_wadr;
  wire yt_rsc_7_5_clkr_en;
  wire yt_rsc_7_5_clkw_en;
  wire [31:0] yt_rsc_7_5_q;
  wire [3:0] yt_rsc_7_5_radr;
  wire yt_rsc_7_5_we;
  wire [31:0] yt_rsc_7_5_d;
  wire [3:0] yt_rsc_7_5_wadr;
  wire yt_rsc_7_6_clkr_en;
  wire yt_rsc_7_6_clkw_en;
  wire [31:0] yt_rsc_7_6_q;
  wire [3:0] yt_rsc_7_6_radr;
  wire yt_rsc_7_6_we;
  wire [31:0] yt_rsc_7_6_d;
  wire [3:0] yt_rsc_7_6_wadr;
  wire yt_rsc_7_7_clkr_en;
  wire yt_rsc_7_7_clkw_en;
  wire [31:0] yt_rsc_7_7_q;
  wire [3:0] yt_rsc_7_7_radr;
  wire yt_rsc_7_7_we;
  wire [31:0] yt_rsc_7_7_d;
  wire [3:0] yt_rsc_7_7_wadr;
  wire yt_rsc_7_8_clkr_en;
  wire yt_rsc_7_8_clkw_en;
  wire [31:0] yt_rsc_7_8_q;
  wire [3:0] yt_rsc_7_8_radr;
  wire yt_rsc_7_8_we;
  wire [31:0] yt_rsc_7_8_d;
  wire [3:0] yt_rsc_7_8_wadr;
  wire yt_rsc_7_9_clkr_en;
  wire yt_rsc_7_9_clkw_en;
  wire [31:0] yt_rsc_7_9_q;
  wire [3:0] yt_rsc_7_9_radr;
  wire yt_rsc_7_9_we;
  wire [31:0] yt_rsc_7_9_d;
  wire [3:0] yt_rsc_7_9_wadr;
  wire yt_rsc_7_10_clkr_en;
  wire yt_rsc_7_10_clkw_en;
  wire [31:0] yt_rsc_7_10_q;
  wire [3:0] yt_rsc_7_10_radr;
  wire yt_rsc_7_10_we;
  wire [31:0] yt_rsc_7_10_d;
  wire [3:0] yt_rsc_7_10_wadr;
  wire yt_rsc_7_11_clkr_en;
  wire yt_rsc_7_11_clkw_en;
  wire [31:0] yt_rsc_7_11_q;
  wire [3:0] yt_rsc_7_11_radr;
  wire yt_rsc_7_11_we;
  wire [31:0] yt_rsc_7_11_d;
  wire [3:0] yt_rsc_7_11_wadr;
  wire yt_rsc_7_12_clkr_en;
  wire yt_rsc_7_12_clkw_en;
  wire [31:0] yt_rsc_7_12_q;
  wire [3:0] yt_rsc_7_12_radr;
  wire yt_rsc_7_12_we;
  wire [31:0] yt_rsc_7_12_d;
  wire [3:0] yt_rsc_7_12_wadr;
  wire yt_rsc_7_13_clkr_en;
  wire yt_rsc_7_13_clkw_en;
  wire [31:0] yt_rsc_7_13_q;
  wire [3:0] yt_rsc_7_13_radr;
  wire yt_rsc_7_13_we;
  wire [31:0] yt_rsc_7_13_d;
  wire [3:0] yt_rsc_7_13_wadr;
  wire yt_rsc_7_14_clkr_en;
  wire yt_rsc_7_14_clkw_en;
  wire [31:0] yt_rsc_7_14_q;
  wire [3:0] yt_rsc_7_14_radr;
  wire yt_rsc_7_14_we;
  wire [31:0] yt_rsc_7_14_d;
  wire [3:0] yt_rsc_7_14_wadr;
  wire yt_rsc_7_15_clkr_en;
  wire yt_rsc_7_15_clkw_en;
  wire [31:0] yt_rsc_7_15_q;
  wire [3:0] yt_rsc_7_15_radr;
  wire yt_rsc_7_15_we;
  wire [31:0] yt_rsc_7_15_d;
  wire [3:0] yt_rsc_7_15_wadr;
  wire yt_rsc_7_16_clkr_en;
  wire yt_rsc_7_16_clkw_en;
  wire [31:0] yt_rsc_7_16_q;
  wire [3:0] yt_rsc_7_16_radr;
  wire yt_rsc_7_16_we;
  wire [31:0] yt_rsc_7_16_d;
  wire [3:0] yt_rsc_7_16_wadr;
  wire yt_rsc_7_17_clkr_en;
  wire yt_rsc_7_17_clkw_en;
  wire [31:0] yt_rsc_7_17_q;
  wire [3:0] yt_rsc_7_17_radr;
  wire yt_rsc_7_17_we;
  wire [31:0] yt_rsc_7_17_d;
  wire [3:0] yt_rsc_7_17_wadr;
  wire yt_rsc_7_18_clkr_en;
  wire yt_rsc_7_18_clkw_en;
  wire [31:0] yt_rsc_7_18_q;
  wire [3:0] yt_rsc_7_18_radr;
  wire yt_rsc_7_18_we;
  wire [31:0] yt_rsc_7_18_d;
  wire [3:0] yt_rsc_7_18_wadr;
  wire yt_rsc_7_19_clkr_en;
  wire yt_rsc_7_19_clkw_en;
  wire [31:0] yt_rsc_7_19_q;
  wire [3:0] yt_rsc_7_19_radr;
  wire yt_rsc_7_19_we;
  wire [31:0] yt_rsc_7_19_d;
  wire [3:0] yt_rsc_7_19_wadr;
  wire yt_rsc_7_20_clkr_en;
  wire yt_rsc_7_20_clkw_en;
  wire [31:0] yt_rsc_7_20_q;
  wire [3:0] yt_rsc_7_20_radr;
  wire yt_rsc_7_20_we;
  wire [31:0] yt_rsc_7_20_d;
  wire [3:0] yt_rsc_7_20_wadr;
  wire yt_rsc_7_21_clkr_en;
  wire yt_rsc_7_21_clkw_en;
  wire [31:0] yt_rsc_7_21_q;
  wire [3:0] yt_rsc_7_21_radr;
  wire yt_rsc_7_21_we;
  wire [31:0] yt_rsc_7_21_d;
  wire [3:0] yt_rsc_7_21_wadr;
  wire yt_rsc_7_22_clkr_en;
  wire yt_rsc_7_22_clkw_en;
  wire [31:0] yt_rsc_7_22_q;
  wire [3:0] yt_rsc_7_22_radr;
  wire yt_rsc_7_22_we;
  wire [31:0] yt_rsc_7_22_d;
  wire [3:0] yt_rsc_7_22_wadr;
  wire yt_rsc_7_23_clkr_en;
  wire yt_rsc_7_23_clkw_en;
  wire [31:0] yt_rsc_7_23_q;
  wire [3:0] yt_rsc_7_23_radr;
  wire yt_rsc_7_23_we;
  wire [31:0] yt_rsc_7_23_d;
  wire [3:0] yt_rsc_7_23_wadr;
  wire yt_rsc_7_24_clkr_en;
  wire yt_rsc_7_24_clkw_en;
  wire [31:0] yt_rsc_7_24_q;
  wire [3:0] yt_rsc_7_24_radr;
  wire yt_rsc_7_24_we;
  wire [31:0] yt_rsc_7_24_d;
  wire [3:0] yt_rsc_7_24_wadr;
  wire yt_rsc_7_25_clkr_en;
  wire yt_rsc_7_25_clkw_en;
  wire [31:0] yt_rsc_7_25_q;
  wire [3:0] yt_rsc_7_25_radr;
  wire yt_rsc_7_25_we;
  wire [31:0] yt_rsc_7_25_d;
  wire [3:0] yt_rsc_7_25_wadr;
  wire yt_rsc_7_26_clkr_en;
  wire yt_rsc_7_26_clkw_en;
  wire [31:0] yt_rsc_7_26_q;
  wire [3:0] yt_rsc_7_26_radr;
  wire yt_rsc_7_26_we;
  wire [31:0] yt_rsc_7_26_d;
  wire [3:0] yt_rsc_7_26_wadr;
  wire yt_rsc_7_27_clkr_en;
  wire yt_rsc_7_27_clkw_en;
  wire [31:0] yt_rsc_7_27_q;
  wire [3:0] yt_rsc_7_27_radr;
  wire yt_rsc_7_27_we;
  wire [31:0] yt_rsc_7_27_d;
  wire [3:0] yt_rsc_7_27_wadr;
  wire yt_rsc_7_28_clkr_en;
  wire yt_rsc_7_28_clkw_en;
  wire [31:0] yt_rsc_7_28_q;
  wire [3:0] yt_rsc_7_28_radr;
  wire yt_rsc_7_28_we;
  wire [31:0] yt_rsc_7_28_d;
  wire [3:0] yt_rsc_7_28_wadr;
  wire yt_rsc_7_29_clkr_en;
  wire yt_rsc_7_29_clkw_en;
  wire [31:0] yt_rsc_7_29_q;
  wire [3:0] yt_rsc_7_29_radr;
  wire yt_rsc_7_29_we;
  wire [31:0] yt_rsc_7_29_d;
  wire [3:0] yt_rsc_7_29_wadr;
  wire yt_rsc_7_30_clkr_en;
  wire yt_rsc_7_30_clkw_en;
  wire [31:0] yt_rsc_7_30_q;
  wire [3:0] yt_rsc_7_30_radr;
  wire yt_rsc_7_30_we;
  wire [31:0] yt_rsc_7_30_d;
  wire [3:0] yt_rsc_7_30_wadr;
  wire yt_rsc_7_31_clkr_en;
  wire yt_rsc_7_31_clkw_en;
  wire [31:0] yt_rsc_7_31_q;
  wire [3:0] yt_rsc_7_31_radr;
  wire yt_rsc_7_31_we;
  wire [31:0] yt_rsc_7_31_d;
  wire [3:0] yt_rsc_7_31_wadr;
  wire [31:0] yt_rsc_0_0_i_d_d_iff;
  wire [3:0] yt_rsc_0_0_i_radr_d_iff;
  wire [3:0] yt_rsc_0_0_i_wadr_d_iff;
  wire yt_rsc_0_0_i_we_d_iff;
  wire yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire [31:0] yt_rsc_0_1_i_d_d_iff;
  wire [3:0] yt_rsc_0_1_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_2_i_d_d_iff;
  wire [3:0] yt_rsc_0_2_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_3_i_d_d_iff;
  wire [3:0] yt_rsc_0_3_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_4_i_d_d_iff;
  wire [3:0] yt_rsc_0_4_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_5_i_d_d_iff;
  wire [3:0] yt_rsc_0_5_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_6_i_d_d_iff;
  wire [3:0] yt_rsc_0_6_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_7_i_d_d_iff;
  wire [31:0] yt_rsc_0_8_i_d_d_iff;
  wire [31:0] yt_rsc_0_9_i_d_d_iff;
  wire [31:0] yt_rsc_0_10_i_d_d_iff;
  wire [3:0] yt_rsc_0_10_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_11_i_d_d_iff;
  wire [3:0] yt_rsc_0_11_i_wadr_d_iff;
  wire [31:0] yt_rsc_0_12_i_d_d_iff;
  wire [31:0] yt_rsc_0_13_i_d_d_iff;
  wire [31:0] yt_rsc_0_14_i_d_d_iff;
  wire [31:0] yt_rsc_0_15_i_d_d_iff;
  wire yt_rsc_0_16_i_we_d_iff;
  wire yt_rsc_1_0_i_we_d_iff;
  wire yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire yt_rsc_1_16_i_we_d_iff;
  wire yt_rsc_2_0_i_we_d_iff;
  wire yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire yt_rsc_2_16_i_we_d_iff;
  wire yt_rsc_3_0_i_we_d_iff;
  wire yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire yt_rsc_3_16_i_we_d_iff;
  wire [31:0] yt_rsc_4_0_i_d_d_iff;
  wire [3:0] yt_rsc_4_0_i_wadr_d_iff;
  wire yt_rsc_4_0_i_we_d_iff;
  wire yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire [31:0] yt_rsc_4_1_i_d_d_iff;
  wire [3:0] yt_rsc_4_1_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_2_i_d_d_iff;
  wire [3:0] yt_rsc_4_2_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_3_i_d_d_iff;
  wire [3:0] yt_rsc_4_3_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_4_i_d_d_iff;
  wire [3:0] yt_rsc_4_4_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_5_i_d_d_iff;
  wire [3:0] yt_rsc_4_5_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_6_i_d_d_iff;
  wire [3:0] yt_rsc_4_6_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_7_i_d_d_iff;
  wire [31:0] yt_rsc_4_8_i_d_d_iff;
  wire [31:0] yt_rsc_4_9_i_d_d_iff;
  wire [3:0] yt_rsc_4_9_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_10_i_d_d_iff;
  wire [3:0] yt_rsc_4_10_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_11_i_d_d_iff;
  wire [3:0] yt_rsc_4_11_i_wadr_d_iff;
  wire [31:0] yt_rsc_4_12_i_d_d_iff;
  wire [31:0] yt_rsc_4_13_i_d_d_iff;
  wire [31:0] yt_rsc_4_14_i_d_d_iff;
  wire [31:0] yt_rsc_4_15_i_d_d_iff;
  wire yt_rsc_4_16_i_we_d_iff;
  wire yt_rsc_5_0_i_we_d_iff;
  wire yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire yt_rsc_5_16_i_we_d_iff;
  wire yt_rsc_6_0_i_we_d_iff;
  wire yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire yt_rsc_6_16_i_we_d_iff;
  wire yt_rsc_7_0_i_we_d_iff;
  wire yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff;
  wire yt_rsc_7_16_i_we_d_iff;
  wire [3:0] xt_rsc_0_0_i_adra_d_iff;
  wire [31:0] xt_rsc_0_0_i_da_d_iff;
  wire xt_rsc_0_0_i_wea_d_iff;
  wire xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire [3:0] xt_rsc_0_1_i_adra_d_iff;
  wire [31:0] xt_rsc_0_1_i_da_d_iff;
  wire [3:0] xt_rsc_0_2_i_adra_d_iff;
  wire [31:0] xt_rsc_0_2_i_da_d_iff;
  wire [3:0] xt_rsc_0_3_i_adra_d_iff;
  wire [31:0] xt_rsc_0_3_i_da_d_iff;
  wire [3:0] xt_rsc_0_4_i_adra_d_iff;
  wire [31:0] xt_rsc_0_4_i_da_d_iff;
  wire [3:0] xt_rsc_0_5_i_adra_d_iff;
  wire [31:0] xt_rsc_0_5_i_da_d_iff;
  wire [3:0] xt_rsc_0_6_i_adra_d_iff;
  wire [31:0] xt_rsc_0_6_i_da_d_iff;
  wire [3:0] xt_rsc_0_7_i_adra_d_iff;
  wire [31:0] xt_rsc_0_7_i_da_d_iff;
  wire [3:0] xt_rsc_0_8_i_adra_d_iff;
  wire [31:0] xt_rsc_0_8_i_da_d_iff;
  wire [3:0] xt_rsc_0_9_i_adra_d_iff;
  wire [31:0] xt_rsc_0_9_i_da_d_iff;
  wire [3:0] xt_rsc_0_10_i_adra_d_iff;
  wire [31:0] xt_rsc_0_10_i_da_d_iff;
  wire [3:0] xt_rsc_0_11_i_adra_d_iff;
  wire [31:0] xt_rsc_0_11_i_da_d_iff;
  wire [3:0] xt_rsc_0_12_i_adra_d_iff;
  wire [31:0] xt_rsc_0_12_i_da_d_iff;
  wire [3:0] xt_rsc_0_13_i_adra_d_iff;
  wire [31:0] xt_rsc_0_13_i_da_d_iff;
  wire [3:0] xt_rsc_0_14_i_adra_d_iff;
  wire [31:0] xt_rsc_0_14_i_da_d_iff;
  wire [3:0] xt_rsc_0_15_i_adra_d_iff;
  wire [31:0] xt_rsc_0_15_i_da_d_iff;
  wire xt_rsc_0_16_i_wea_d_iff;
  wire xt_rsc_1_0_i_wea_d_iff;
  wire xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire xt_rsc_1_16_i_wea_d_iff;
  wire xt_rsc_2_0_i_wea_d_iff;
  wire xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire xt_rsc_2_16_i_wea_d_iff;
  wire xt_rsc_3_0_i_wea_d_iff;
  wire xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire xt_rsc_3_16_i_wea_d_iff;
  wire [31:0] xt_rsc_4_0_i_da_d_iff;
  wire xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire [3:0] xt_rsc_4_1_i_adra_d_iff;
  wire [31:0] xt_rsc_4_1_i_da_d_iff;
  wire [3:0] xt_rsc_4_2_i_adra_d_iff;
  wire [31:0] xt_rsc_4_2_i_da_d_iff;
  wire [31:0] xt_rsc_4_3_i_da_d_iff;
  wire [31:0] xt_rsc_4_4_i_da_d_iff;
  wire [31:0] xt_rsc_4_5_i_da_d_iff;
  wire [31:0] xt_rsc_4_6_i_da_d_iff;
  wire [31:0] xt_rsc_4_7_i_da_d_iff;
  wire [31:0] xt_rsc_4_8_i_da_d_iff;
  wire [3:0] xt_rsc_4_9_i_adra_d_iff;
  wire [31:0] xt_rsc_4_9_i_da_d_iff;
  wire [3:0] xt_rsc_4_10_i_adra_d_iff;
  wire [31:0] xt_rsc_4_10_i_da_d_iff;
  wire [31:0] xt_rsc_4_11_i_da_d_iff;
  wire [31:0] xt_rsc_4_12_i_da_d_iff;
  wire [31:0] xt_rsc_4_13_i_da_d_iff;
  wire [31:0] xt_rsc_4_14_i_da_d_iff;
  wire [31:0] xt_rsc_4_15_i_da_d_iff;
  wire xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;
  wire xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_twiddle_rsc_0_0_i_adra_d;
  assign nl_twiddle_rsc_0_0_i_adra_d = {8'b00000000 , twiddle_rsc_0_0_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_1_i_adra_d;
  assign nl_twiddle_rsc_0_1_i_adra_d = {8'b00000000 , twiddle_rsc_0_1_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_2_i_adra_d;
  assign nl_twiddle_rsc_0_2_i_adra_d = {8'b00000000 , twiddle_rsc_0_2_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_3_i_adra_d;
  assign nl_twiddle_rsc_0_3_i_adra_d = {8'b00000000 , twiddle_rsc_0_3_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_4_i_adra_d;
  assign nl_twiddle_rsc_0_4_i_adra_d = {8'b00000000 , twiddle_rsc_0_4_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_5_i_adra_d;
  assign nl_twiddle_rsc_0_5_i_adra_d = {8'b00000000 , twiddle_rsc_0_5_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_6_i_adra_d;
  assign nl_twiddle_rsc_0_6_i_adra_d = {8'b00000000 , twiddle_rsc_0_6_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_7_i_adra_d;
  assign nl_twiddle_rsc_0_7_i_adra_d = {8'b00000000 , twiddle_rsc_0_7_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_8_i_adra_d;
  assign nl_twiddle_rsc_0_8_i_adra_d = {8'b00000000 , twiddle_rsc_0_8_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_9_i_adra_d;
  assign nl_twiddle_rsc_0_9_i_adra_d = {8'b00000000 , twiddle_rsc_0_9_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_10_i_adra_d;
  assign nl_twiddle_rsc_0_10_i_adra_d = {8'b00000000 , twiddle_rsc_0_10_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_11_i_adra_d;
  assign nl_twiddle_rsc_0_11_i_adra_d = {8'b00000000 , twiddle_rsc_0_11_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_12_i_adra_d;
  assign nl_twiddle_rsc_0_12_i_adra_d = {8'b00000000 , twiddle_rsc_0_12_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_13_i_adra_d;
  assign nl_twiddle_rsc_0_13_i_adra_d = {8'b00000000 , twiddle_rsc_0_13_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_14_i_adra_d;
  assign nl_twiddle_rsc_0_14_i_adra_d = {8'b00000000 , twiddle_rsc_0_14_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_15_i_adra_d;
  assign nl_twiddle_rsc_0_15_i_adra_d = {8'b00000000 , twiddle_rsc_0_15_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_0_i_adra_d;
  assign nl_twiddle_h_rsc_0_0_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_0_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_1_i_adra_d;
  assign nl_twiddle_h_rsc_0_1_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_1_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_2_i_adra_d;
  assign nl_twiddle_h_rsc_0_2_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_2_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_3_i_adra_d;
  assign nl_twiddle_h_rsc_0_3_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_3_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_4_i_adra_d;
  assign nl_twiddle_h_rsc_0_4_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_4_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_5_i_adra_d;
  assign nl_twiddle_h_rsc_0_5_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_5_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_6_i_adra_d;
  assign nl_twiddle_h_rsc_0_6_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_6_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_7_i_adra_d;
  assign nl_twiddle_h_rsc_0_7_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_7_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_8_i_adra_d;
  assign nl_twiddle_h_rsc_0_8_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_8_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_9_i_adra_d;
  assign nl_twiddle_h_rsc_0_9_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_9_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_10_i_adra_d;
  assign nl_twiddle_h_rsc_0_10_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_10_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_11_i_adra_d;
  assign nl_twiddle_h_rsc_0_11_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_11_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_12_i_adra_d;
  assign nl_twiddle_h_rsc_0_12_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_12_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_13_i_adra_d;
  assign nl_twiddle_h_rsc_0_13_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_13_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_14_i_adra_d;
  assign nl_twiddle_h_rsc_0_14_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_14_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_15_i_adra_d;
  assign nl_twiddle_h_rsc_0_15_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_15_i_adra_d};
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_0_clkr_en),
      .d(yt_rsc_0_0_d),
      .q(yt_rsc_0_0_q),
      .radr(yt_rsc_0_0_radr),
      .wadr(yt_rsc_0_0_wadr),
      .we(yt_rsc_0_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_1_clkr_en),
      .d(yt_rsc_0_1_d),
      .q(yt_rsc_0_1_q),
      .radr(yt_rsc_0_1_radr),
      .wadr(yt_rsc_0_1_wadr),
      .we(yt_rsc_0_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_2_clkr_en),
      .d(yt_rsc_0_2_d),
      .q(yt_rsc_0_2_q),
      .radr(yt_rsc_0_2_radr),
      .wadr(yt_rsc_0_2_wadr),
      .we(yt_rsc_0_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_3_clkr_en),
      .d(yt_rsc_0_3_d),
      .q(yt_rsc_0_3_q),
      .radr(yt_rsc_0_3_radr),
      .wadr(yt_rsc_0_3_wadr),
      .we(yt_rsc_0_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_4_clkr_en),
      .d(yt_rsc_0_4_d),
      .q(yt_rsc_0_4_q),
      .radr(yt_rsc_0_4_radr),
      .wadr(yt_rsc_0_4_wadr),
      .we(yt_rsc_0_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_5_clkr_en),
      .d(yt_rsc_0_5_d),
      .q(yt_rsc_0_5_q),
      .radr(yt_rsc_0_5_radr),
      .wadr(yt_rsc_0_5_wadr),
      .we(yt_rsc_0_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_6_clkr_en),
      .d(yt_rsc_0_6_d),
      .q(yt_rsc_0_6_q),
      .radr(yt_rsc_0_6_radr),
      .wadr(yt_rsc_0_6_wadr),
      .we(yt_rsc_0_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_7_clkr_en),
      .d(yt_rsc_0_7_d),
      .q(yt_rsc_0_7_q),
      .radr(yt_rsc_0_7_radr),
      .wadr(yt_rsc_0_7_wadr),
      .we(yt_rsc_0_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_8_clkr_en),
      .d(yt_rsc_0_8_d),
      .q(yt_rsc_0_8_q),
      .radr(yt_rsc_0_8_radr),
      .wadr(yt_rsc_0_8_wadr),
      .we(yt_rsc_0_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_9_clkr_en),
      .d(yt_rsc_0_9_d),
      .q(yt_rsc_0_9_q),
      .radr(yt_rsc_0_9_radr),
      .wadr(yt_rsc_0_9_wadr),
      .we(yt_rsc_0_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_10_clkr_en),
      .d(yt_rsc_0_10_d),
      .q(yt_rsc_0_10_q),
      .radr(yt_rsc_0_10_radr),
      .wadr(yt_rsc_0_10_wadr),
      .we(yt_rsc_0_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_11_clkr_en),
      .d(yt_rsc_0_11_d),
      .q(yt_rsc_0_11_q),
      .radr(yt_rsc_0_11_radr),
      .wadr(yt_rsc_0_11_wadr),
      .we(yt_rsc_0_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_12_clkr_en),
      .d(yt_rsc_0_12_d),
      .q(yt_rsc_0_12_q),
      .radr(yt_rsc_0_12_radr),
      .wadr(yt_rsc_0_12_wadr),
      .we(yt_rsc_0_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_13_clkr_en),
      .d(yt_rsc_0_13_d),
      .q(yt_rsc_0_13_q),
      .radr(yt_rsc_0_13_radr),
      .wadr(yt_rsc_0_13_wadr),
      .we(yt_rsc_0_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_14_clkr_en),
      .d(yt_rsc_0_14_d),
      .q(yt_rsc_0_14_q),
      .radr(yt_rsc_0_14_radr),
      .wadr(yt_rsc_0_14_wadr),
      .we(yt_rsc_0_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_15_clkr_en),
      .d(yt_rsc_0_15_d),
      .q(yt_rsc_0_15_q),
      .radr(yt_rsc_0_15_radr),
      .wadr(yt_rsc_0_15_wadr),
      .we(yt_rsc_0_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_16_clkr_en),
      .d(yt_rsc_0_16_d),
      .q(yt_rsc_0_16_q),
      .radr(yt_rsc_0_16_radr),
      .wadr(yt_rsc_0_16_wadr),
      .we(yt_rsc_0_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_17_clkr_en),
      .d(yt_rsc_0_17_d),
      .q(yt_rsc_0_17_q),
      .radr(yt_rsc_0_17_radr),
      .wadr(yt_rsc_0_17_wadr),
      .we(yt_rsc_0_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_18_clkr_en),
      .d(yt_rsc_0_18_d),
      .q(yt_rsc_0_18_q),
      .radr(yt_rsc_0_18_radr),
      .wadr(yt_rsc_0_18_wadr),
      .we(yt_rsc_0_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_19_clkr_en),
      .d(yt_rsc_0_19_d),
      .q(yt_rsc_0_19_q),
      .radr(yt_rsc_0_19_radr),
      .wadr(yt_rsc_0_19_wadr),
      .we(yt_rsc_0_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_20_clkr_en),
      .d(yt_rsc_0_20_d),
      .q(yt_rsc_0_20_q),
      .radr(yt_rsc_0_20_radr),
      .wadr(yt_rsc_0_20_wadr),
      .we(yt_rsc_0_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_21_clkr_en),
      .d(yt_rsc_0_21_d),
      .q(yt_rsc_0_21_q),
      .radr(yt_rsc_0_21_radr),
      .wadr(yt_rsc_0_21_wadr),
      .we(yt_rsc_0_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_22_clkr_en),
      .d(yt_rsc_0_22_d),
      .q(yt_rsc_0_22_q),
      .radr(yt_rsc_0_22_radr),
      .wadr(yt_rsc_0_22_wadr),
      .we(yt_rsc_0_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_23_clkr_en),
      .d(yt_rsc_0_23_d),
      .q(yt_rsc_0_23_q),
      .radr(yt_rsc_0_23_radr),
      .wadr(yt_rsc_0_23_wadr),
      .we(yt_rsc_0_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_24_clkr_en),
      .d(yt_rsc_0_24_d),
      .q(yt_rsc_0_24_q),
      .radr(yt_rsc_0_24_radr),
      .wadr(yt_rsc_0_24_wadr),
      .we(yt_rsc_0_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_25_clkr_en),
      .d(yt_rsc_0_25_d),
      .q(yt_rsc_0_25_q),
      .radr(yt_rsc_0_25_radr),
      .wadr(yt_rsc_0_25_wadr),
      .we(yt_rsc_0_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_26_clkr_en),
      .d(yt_rsc_0_26_d),
      .q(yt_rsc_0_26_q),
      .radr(yt_rsc_0_26_radr),
      .wadr(yt_rsc_0_26_wadr),
      .we(yt_rsc_0_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_27_clkr_en),
      .d(yt_rsc_0_27_d),
      .q(yt_rsc_0_27_q),
      .radr(yt_rsc_0_27_radr),
      .wadr(yt_rsc_0_27_wadr),
      .we(yt_rsc_0_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_28_clkr_en),
      .d(yt_rsc_0_28_d),
      .q(yt_rsc_0_28_q),
      .radr(yt_rsc_0_28_radr),
      .wadr(yt_rsc_0_28_wadr),
      .we(yt_rsc_0_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_29_clkr_en),
      .d(yt_rsc_0_29_d),
      .q(yt_rsc_0_29_q),
      .radr(yt_rsc_0_29_radr),
      .wadr(yt_rsc_0_29_wadr),
      .we(yt_rsc_0_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_30_clkr_en),
      .d(yt_rsc_0_30_d),
      .q(yt_rsc_0_30_q),
      .radr(yt_rsc_0_30_radr),
      .wadr(yt_rsc_0_30_wadr),
      .we(yt_rsc_0_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_0_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_0_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_0_31_clkr_en),
      .d(yt_rsc_0_31_d),
      .q(yt_rsc_0_31_q),
      .radr(yt_rsc_0_31_radr),
      .wadr(yt_rsc_0_31_wadr),
      .we(yt_rsc_0_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_0_clkr_en),
      .d(yt_rsc_1_0_d),
      .q(yt_rsc_1_0_q),
      .radr(yt_rsc_1_0_radr),
      .wadr(yt_rsc_1_0_wadr),
      .we(yt_rsc_1_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_1_clkr_en),
      .d(yt_rsc_1_1_d),
      .q(yt_rsc_1_1_q),
      .radr(yt_rsc_1_1_radr),
      .wadr(yt_rsc_1_1_wadr),
      .we(yt_rsc_1_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_2_clkr_en),
      .d(yt_rsc_1_2_d),
      .q(yt_rsc_1_2_q),
      .radr(yt_rsc_1_2_radr),
      .wadr(yt_rsc_1_2_wadr),
      .we(yt_rsc_1_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_3_clkr_en),
      .d(yt_rsc_1_3_d),
      .q(yt_rsc_1_3_q),
      .radr(yt_rsc_1_3_radr),
      .wadr(yt_rsc_1_3_wadr),
      .we(yt_rsc_1_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_4_clkr_en),
      .d(yt_rsc_1_4_d),
      .q(yt_rsc_1_4_q),
      .radr(yt_rsc_1_4_radr),
      .wadr(yt_rsc_1_4_wadr),
      .we(yt_rsc_1_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_5_clkr_en),
      .d(yt_rsc_1_5_d),
      .q(yt_rsc_1_5_q),
      .radr(yt_rsc_1_5_radr),
      .wadr(yt_rsc_1_5_wadr),
      .we(yt_rsc_1_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_6_clkr_en),
      .d(yt_rsc_1_6_d),
      .q(yt_rsc_1_6_q),
      .radr(yt_rsc_1_6_radr),
      .wadr(yt_rsc_1_6_wadr),
      .we(yt_rsc_1_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_7_clkr_en),
      .d(yt_rsc_1_7_d),
      .q(yt_rsc_1_7_q),
      .radr(yt_rsc_1_7_radr),
      .wadr(yt_rsc_1_7_wadr),
      .we(yt_rsc_1_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_8_clkr_en),
      .d(yt_rsc_1_8_d),
      .q(yt_rsc_1_8_q),
      .radr(yt_rsc_1_8_radr),
      .wadr(yt_rsc_1_8_wadr),
      .we(yt_rsc_1_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_9_clkr_en),
      .d(yt_rsc_1_9_d),
      .q(yt_rsc_1_9_q),
      .radr(yt_rsc_1_9_radr),
      .wadr(yt_rsc_1_9_wadr),
      .we(yt_rsc_1_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_10_clkr_en),
      .d(yt_rsc_1_10_d),
      .q(yt_rsc_1_10_q),
      .radr(yt_rsc_1_10_radr),
      .wadr(yt_rsc_1_10_wadr),
      .we(yt_rsc_1_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_11_clkr_en),
      .d(yt_rsc_1_11_d),
      .q(yt_rsc_1_11_q),
      .radr(yt_rsc_1_11_radr),
      .wadr(yt_rsc_1_11_wadr),
      .we(yt_rsc_1_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_12_clkr_en),
      .d(yt_rsc_1_12_d),
      .q(yt_rsc_1_12_q),
      .radr(yt_rsc_1_12_radr),
      .wadr(yt_rsc_1_12_wadr),
      .we(yt_rsc_1_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_13_clkr_en),
      .d(yt_rsc_1_13_d),
      .q(yt_rsc_1_13_q),
      .radr(yt_rsc_1_13_radr),
      .wadr(yt_rsc_1_13_wadr),
      .we(yt_rsc_1_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_14_clkr_en),
      .d(yt_rsc_1_14_d),
      .q(yt_rsc_1_14_q),
      .radr(yt_rsc_1_14_radr),
      .wadr(yt_rsc_1_14_wadr),
      .we(yt_rsc_1_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_15_clkr_en),
      .d(yt_rsc_1_15_d),
      .q(yt_rsc_1_15_q),
      .radr(yt_rsc_1_15_radr),
      .wadr(yt_rsc_1_15_wadr),
      .we(yt_rsc_1_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_16_clkr_en),
      .d(yt_rsc_1_16_d),
      .q(yt_rsc_1_16_q),
      .radr(yt_rsc_1_16_radr),
      .wadr(yt_rsc_1_16_wadr),
      .we(yt_rsc_1_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_17_clkr_en),
      .d(yt_rsc_1_17_d),
      .q(yt_rsc_1_17_q),
      .radr(yt_rsc_1_17_radr),
      .wadr(yt_rsc_1_17_wadr),
      .we(yt_rsc_1_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_18_clkr_en),
      .d(yt_rsc_1_18_d),
      .q(yt_rsc_1_18_q),
      .radr(yt_rsc_1_18_radr),
      .wadr(yt_rsc_1_18_wadr),
      .we(yt_rsc_1_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_19_clkr_en),
      .d(yt_rsc_1_19_d),
      .q(yt_rsc_1_19_q),
      .radr(yt_rsc_1_19_radr),
      .wadr(yt_rsc_1_19_wadr),
      .we(yt_rsc_1_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_20_clkr_en),
      .d(yt_rsc_1_20_d),
      .q(yt_rsc_1_20_q),
      .radr(yt_rsc_1_20_radr),
      .wadr(yt_rsc_1_20_wadr),
      .we(yt_rsc_1_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_21_clkr_en),
      .d(yt_rsc_1_21_d),
      .q(yt_rsc_1_21_q),
      .radr(yt_rsc_1_21_radr),
      .wadr(yt_rsc_1_21_wadr),
      .we(yt_rsc_1_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_22_clkr_en),
      .d(yt_rsc_1_22_d),
      .q(yt_rsc_1_22_q),
      .radr(yt_rsc_1_22_radr),
      .wadr(yt_rsc_1_22_wadr),
      .we(yt_rsc_1_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_23_clkr_en),
      .d(yt_rsc_1_23_d),
      .q(yt_rsc_1_23_q),
      .radr(yt_rsc_1_23_radr),
      .wadr(yt_rsc_1_23_wadr),
      .we(yt_rsc_1_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_24_clkr_en),
      .d(yt_rsc_1_24_d),
      .q(yt_rsc_1_24_q),
      .radr(yt_rsc_1_24_radr),
      .wadr(yt_rsc_1_24_wadr),
      .we(yt_rsc_1_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_25_clkr_en),
      .d(yt_rsc_1_25_d),
      .q(yt_rsc_1_25_q),
      .radr(yt_rsc_1_25_radr),
      .wadr(yt_rsc_1_25_wadr),
      .we(yt_rsc_1_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_26_clkr_en),
      .d(yt_rsc_1_26_d),
      .q(yt_rsc_1_26_q),
      .radr(yt_rsc_1_26_radr),
      .wadr(yt_rsc_1_26_wadr),
      .we(yt_rsc_1_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_27_clkr_en),
      .d(yt_rsc_1_27_d),
      .q(yt_rsc_1_27_q),
      .radr(yt_rsc_1_27_radr),
      .wadr(yt_rsc_1_27_wadr),
      .we(yt_rsc_1_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_28_clkr_en),
      .d(yt_rsc_1_28_d),
      .q(yt_rsc_1_28_q),
      .radr(yt_rsc_1_28_radr),
      .wadr(yt_rsc_1_28_wadr),
      .we(yt_rsc_1_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_29_clkr_en),
      .d(yt_rsc_1_29_d),
      .q(yt_rsc_1_29_q),
      .radr(yt_rsc_1_29_radr),
      .wadr(yt_rsc_1_29_wadr),
      .we(yt_rsc_1_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_30_clkr_en),
      .d(yt_rsc_1_30_d),
      .q(yt_rsc_1_30_q),
      .radr(yt_rsc_1_30_radr),
      .wadr(yt_rsc_1_30_wadr),
      .we(yt_rsc_1_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_1_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_1_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_1_31_clkr_en),
      .d(yt_rsc_1_31_d),
      .q(yt_rsc_1_31_q),
      .radr(yt_rsc_1_31_radr),
      .wadr(yt_rsc_1_31_wadr),
      .we(yt_rsc_1_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_0_clkr_en),
      .d(yt_rsc_2_0_d),
      .q(yt_rsc_2_0_q),
      .radr(yt_rsc_2_0_radr),
      .wadr(yt_rsc_2_0_wadr),
      .we(yt_rsc_2_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_1_clkr_en),
      .d(yt_rsc_2_1_d),
      .q(yt_rsc_2_1_q),
      .radr(yt_rsc_2_1_radr),
      .wadr(yt_rsc_2_1_wadr),
      .we(yt_rsc_2_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_2_clkr_en),
      .d(yt_rsc_2_2_d),
      .q(yt_rsc_2_2_q),
      .radr(yt_rsc_2_2_radr),
      .wadr(yt_rsc_2_2_wadr),
      .we(yt_rsc_2_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_3_clkr_en),
      .d(yt_rsc_2_3_d),
      .q(yt_rsc_2_3_q),
      .radr(yt_rsc_2_3_radr),
      .wadr(yt_rsc_2_3_wadr),
      .we(yt_rsc_2_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_4_clkr_en),
      .d(yt_rsc_2_4_d),
      .q(yt_rsc_2_4_q),
      .radr(yt_rsc_2_4_radr),
      .wadr(yt_rsc_2_4_wadr),
      .we(yt_rsc_2_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_5_clkr_en),
      .d(yt_rsc_2_5_d),
      .q(yt_rsc_2_5_q),
      .radr(yt_rsc_2_5_radr),
      .wadr(yt_rsc_2_5_wadr),
      .we(yt_rsc_2_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_6_clkr_en),
      .d(yt_rsc_2_6_d),
      .q(yt_rsc_2_6_q),
      .radr(yt_rsc_2_6_radr),
      .wadr(yt_rsc_2_6_wadr),
      .we(yt_rsc_2_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_7_clkr_en),
      .d(yt_rsc_2_7_d),
      .q(yt_rsc_2_7_q),
      .radr(yt_rsc_2_7_radr),
      .wadr(yt_rsc_2_7_wadr),
      .we(yt_rsc_2_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_8_clkr_en),
      .d(yt_rsc_2_8_d),
      .q(yt_rsc_2_8_q),
      .radr(yt_rsc_2_8_radr),
      .wadr(yt_rsc_2_8_wadr),
      .we(yt_rsc_2_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_9_clkr_en),
      .d(yt_rsc_2_9_d),
      .q(yt_rsc_2_9_q),
      .radr(yt_rsc_2_9_radr),
      .wadr(yt_rsc_2_9_wadr),
      .we(yt_rsc_2_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_10_clkr_en),
      .d(yt_rsc_2_10_d),
      .q(yt_rsc_2_10_q),
      .radr(yt_rsc_2_10_radr),
      .wadr(yt_rsc_2_10_wadr),
      .we(yt_rsc_2_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_11_clkr_en),
      .d(yt_rsc_2_11_d),
      .q(yt_rsc_2_11_q),
      .radr(yt_rsc_2_11_radr),
      .wadr(yt_rsc_2_11_wadr),
      .we(yt_rsc_2_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_12_clkr_en),
      .d(yt_rsc_2_12_d),
      .q(yt_rsc_2_12_q),
      .radr(yt_rsc_2_12_radr),
      .wadr(yt_rsc_2_12_wadr),
      .we(yt_rsc_2_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_13_clkr_en),
      .d(yt_rsc_2_13_d),
      .q(yt_rsc_2_13_q),
      .radr(yt_rsc_2_13_radr),
      .wadr(yt_rsc_2_13_wadr),
      .we(yt_rsc_2_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_14_clkr_en),
      .d(yt_rsc_2_14_d),
      .q(yt_rsc_2_14_q),
      .radr(yt_rsc_2_14_radr),
      .wadr(yt_rsc_2_14_wadr),
      .we(yt_rsc_2_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_15_clkr_en),
      .d(yt_rsc_2_15_d),
      .q(yt_rsc_2_15_q),
      .radr(yt_rsc_2_15_radr),
      .wadr(yt_rsc_2_15_wadr),
      .we(yt_rsc_2_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_16_clkr_en),
      .d(yt_rsc_2_16_d),
      .q(yt_rsc_2_16_q),
      .radr(yt_rsc_2_16_radr),
      .wadr(yt_rsc_2_16_wadr),
      .we(yt_rsc_2_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_17_clkr_en),
      .d(yt_rsc_2_17_d),
      .q(yt_rsc_2_17_q),
      .radr(yt_rsc_2_17_radr),
      .wadr(yt_rsc_2_17_wadr),
      .we(yt_rsc_2_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_18_clkr_en),
      .d(yt_rsc_2_18_d),
      .q(yt_rsc_2_18_q),
      .radr(yt_rsc_2_18_radr),
      .wadr(yt_rsc_2_18_wadr),
      .we(yt_rsc_2_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_19_clkr_en),
      .d(yt_rsc_2_19_d),
      .q(yt_rsc_2_19_q),
      .radr(yt_rsc_2_19_radr),
      .wadr(yt_rsc_2_19_wadr),
      .we(yt_rsc_2_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_20_clkr_en),
      .d(yt_rsc_2_20_d),
      .q(yt_rsc_2_20_q),
      .radr(yt_rsc_2_20_radr),
      .wadr(yt_rsc_2_20_wadr),
      .we(yt_rsc_2_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_21_clkr_en),
      .d(yt_rsc_2_21_d),
      .q(yt_rsc_2_21_q),
      .radr(yt_rsc_2_21_radr),
      .wadr(yt_rsc_2_21_wadr),
      .we(yt_rsc_2_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_22_clkr_en),
      .d(yt_rsc_2_22_d),
      .q(yt_rsc_2_22_q),
      .radr(yt_rsc_2_22_radr),
      .wadr(yt_rsc_2_22_wadr),
      .we(yt_rsc_2_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_23_clkr_en),
      .d(yt_rsc_2_23_d),
      .q(yt_rsc_2_23_q),
      .radr(yt_rsc_2_23_radr),
      .wadr(yt_rsc_2_23_wadr),
      .we(yt_rsc_2_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_24_clkr_en),
      .d(yt_rsc_2_24_d),
      .q(yt_rsc_2_24_q),
      .radr(yt_rsc_2_24_radr),
      .wadr(yt_rsc_2_24_wadr),
      .we(yt_rsc_2_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_25_clkr_en),
      .d(yt_rsc_2_25_d),
      .q(yt_rsc_2_25_q),
      .radr(yt_rsc_2_25_radr),
      .wadr(yt_rsc_2_25_wadr),
      .we(yt_rsc_2_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_26_clkr_en),
      .d(yt_rsc_2_26_d),
      .q(yt_rsc_2_26_q),
      .radr(yt_rsc_2_26_radr),
      .wadr(yt_rsc_2_26_wadr),
      .we(yt_rsc_2_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_27_clkr_en),
      .d(yt_rsc_2_27_d),
      .q(yt_rsc_2_27_q),
      .radr(yt_rsc_2_27_radr),
      .wadr(yt_rsc_2_27_wadr),
      .we(yt_rsc_2_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_28_clkr_en),
      .d(yt_rsc_2_28_d),
      .q(yt_rsc_2_28_q),
      .radr(yt_rsc_2_28_radr),
      .wadr(yt_rsc_2_28_wadr),
      .we(yt_rsc_2_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_29_clkr_en),
      .d(yt_rsc_2_29_d),
      .q(yt_rsc_2_29_q),
      .radr(yt_rsc_2_29_radr),
      .wadr(yt_rsc_2_29_wadr),
      .we(yt_rsc_2_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_30_clkr_en),
      .d(yt_rsc_2_30_d),
      .q(yt_rsc_2_30_q),
      .radr(yt_rsc_2_30_radr),
      .wadr(yt_rsc_2_30_wadr),
      .we(yt_rsc_2_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_2_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_2_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_2_31_clkr_en),
      .d(yt_rsc_2_31_d),
      .q(yt_rsc_2_31_q),
      .radr(yt_rsc_2_31_radr),
      .wadr(yt_rsc_2_31_wadr),
      .we(yt_rsc_2_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_0_clkr_en),
      .d(yt_rsc_3_0_d),
      .q(yt_rsc_3_0_q),
      .radr(yt_rsc_3_0_radr),
      .wadr(yt_rsc_3_0_wadr),
      .we(yt_rsc_3_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_1_clkr_en),
      .d(yt_rsc_3_1_d),
      .q(yt_rsc_3_1_q),
      .radr(yt_rsc_3_1_radr),
      .wadr(yt_rsc_3_1_wadr),
      .we(yt_rsc_3_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_2_clkr_en),
      .d(yt_rsc_3_2_d),
      .q(yt_rsc_3_2_q),
      .radr(yt_rsc_3_2_radr),
      .wadr(yt_rsc_3_2_wadr),
      .we(yt_rsc_3_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_3_clkr_en),
      .d(yt_rsc_3_3_d),
      .q(yt_rsc_3_3_q),
      .radr(yt_rsc_3_3_radr),
      .wadr(yt_rsc_3_3_wadr),
      .we(yt_rsc_3_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_4_clkr_en),
      .d(yt_rsc_3_4_d),
      .q(yt_rsc_3_4_q),
      .radr(yt_rsc_3_4_radr),
      .wadr(yt_rsc_3_4_wadr),
      .we(yt_rsc_3_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_5_clkr_en),
      .d(yt_rsc_3_5_d),
      .q(yt_rsc_3_5_q),
      .radr(yt_rsc_3_5_radr),
      .wadr(yt_rsc_3_5_wadr),
      .we(yt_rsc_3_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_6_clkr_en),
      .d(yt_rsc_3_6_d),
      .q(yt_rsc_3_6_q),
      .radr(yt_rsc_3_6_radr),
      .wadr(yt_rsc_3_6_wadr),
      .we(yt_rsc_3_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_7_clkr_en),
      .d(yt_rsc_3_7_d),
      .q(yt_rsc_3_7_q),
      .radr(yt_rsc_3_7_radr),
      .wadr(yt_rsc_3_7_wadr),
      .we(yt_rsc_3_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_8_clkr_en),
      .d(yt_rsc_3_8_d),
      .q(yt_rsc_3_8_q),
      .radr(yt_rsc_3_8_radr),
      .wadr(yt_rsc_3_8_wadr),
      .we(yt_rsc_3_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_9_clkr_en),
      .d(yt_rsc_3_9_d),
      .q(yt_rsc_3_9_q),
      .radr(yt_rsc_3_9_radr),
      .wadr(yt_rsc_3_9_wadr),
      .we(yt_rsc_3_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_10_clkr_en),
      .d(yt_rsc_3_10_d),
      .q(yt_rsc_3_10_q),
      .radr(yt_rsc_3_10_radr),
      .wadr(yt_rsc_3_10_wadr),
      .we(yt_rsc_3_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_11_clkr_en),
      .d(yt_rsc_3_11_d),
      .q(yt_rsc_3_11_q),
      .radr(yt_rsc_3_11_radr),
      .wadr(yt_rsc_3_11_wadr),
      .we(yt_rsc_3_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_12_clkr_en),
      .d(yt_rsc_3_12_d),
      .q(yt_rsc_3_12_q),
      .radr(yt_rsc_3_12_radr),
      .wadr(yt_rsc_3_12_wadr),
      .we(yt_rsc_3_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_13_clkr_en),
      .d(yt_rsc_3_13_d),
      .q(yt_rsc_3_13_q),
      .radr(yt_rsc_3_13_radr),
      .wadr(yt_rsc_3_13_wadr),
      .we(yt_rsc_3_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_14_clkr_en),
      .d(yt_rsc_3_14_d),
      .q(yt_rsc_3_14_q),
      .radr(yt_rsc_3_14_radr),
      .wadr(yt_rsc_3_14_wadr),
      .we(yt_rsc_3_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_15_clkr_en),
      .d(yt_rsc_3_15_d),
      .q(yt_rsc_3_15_q),
      .radr(yt_rsc_3_15_radr),
      .wadr(yt_rsc_3_15_wadr),
      .we(yt_rsc_3_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_16_clkr_en),
      .d(yt_rsc_3_16_d),
      .q(yt_rsc_3_16_q),
      .radr(yt_rsc_3_16_radr),
      .wadr(yt_rsc_3_16_wadr),
      .we(yt_rsc_3_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_17_clkr_en),
      .d(yt_rsc_3_17_d),
      .q(yt_rsc_3_17_q),
      .radr(yt_rsc_3_17_radr),
      .wadr(yt_rsc_3_17_wadr),
      .we(yt_rsc_3_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_18_clkr_en),
      .d(yt_rsc_3_18_d),
      .q(yt_rsc_3_18_q),
      .radr(yt_rsc_3_18_radr),
      .wadr(yt_rsc_3_18_wadr),
      .we(yt_rsc_3_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_19_clkr_en),
      .d(yt_rsc_3_19_d),
      .q(yt_rsc_3_19_q),
      .radr(yt_rsc_3_19_radr),
      .wadr(yt_rsc_3_19_wadr),
      .we(yt_rsc_3_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_20_clkr_en),
      .d(yt_rsc_3_20_d),
      .q(yt_rsc_3_20_q),
      .radr(yt_rsc_3_20_radr),
      .wadr(yt_rsc_3_20_wadr),
      .we(yt_rsc_3_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_21_clkr_en),
      .d(yt_rsc_3_21_d),
      .q(yt_rsc_3_21_q),
      .radr(yt_rsc_3_21_radr),
      .wadr(yt_rsc_3_21_wadr),
      .we(yt_rsc_3_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_22_clkr_en),
      .d(yt_rsc_3_22_d),
      .q(yt_rsc_3_22_q),
      .radr(yt_rsc_3_22_radr),
      .wadr(yt_rsc_3_22_wadr),
      .we(yt_rsc_3_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_23_clkr_en),
      .d(yt_rsc_3_23_d),
      .q(yt_rsc_3_23_q),
      .radr(yt_rsc_3_23_radr),
      .wadr(yt_rsc_3_23_wadr),
      .we(yt_rsc_3_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_24_clkr_en),
      .d(yt_rsc_3_24_d),
      .q(yt_rsc_3_24_q),
      .radr(yt_rsc_3_24_radr),
      .wadr(yt_rsc_3_24_wadr),
      .we(yt_rsc_3_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_25_clkr_en),
      .d(yt_rsc_3_25_d),
      .q(yt_rsc_3_25_q),
      .radr(yt_rsc_3_25_radr),
      .wadr(yt_rsc_3_25_wadr),
      .we(yt_rsc_3_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_26_clkr_en),
      .d(yt_rsc_3_26_d),
      .q(yt_rsc_3_26_q),
      .radr(yt_rsc_3_26_radr),
      .wadr(yt_rsc_3_26_wadr),
      .we(yt_rsc_3_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_27_clkr_en),
      .d(yt_rsc_3_27_d),
      .q(yt_rsc_3_27_q),
      .radr(yt_rsc_3_27_radr),
      .wadr(yt_rsc_3_27_wadr),
      .we(yt_rsc_3_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_28_clkr_en),
      .d(yt_rsc_3_28_d),
      .q(yt_rsc_3_28_q),
      .radr(yt_rsc_3_28_radr),
      .wadr(yt_rsc_3_28_wadr),
      .we(yt_rsc_3_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_29_clkr_en),
      .d(yt_rsc_3_29_d),
      .q(yt_rsc_3_29_q),
      .radr(yt_rsc_3_29_radr),
      .wadr(yt_rsc_3_29_wadr),
      .we(yt_rsc_3_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_30_clkr_en),
      .d(yt_rsc_3_30_d),
      .q(yt_rsc_3_30_q),
      .radr(yt_rsc_3_30_radr),
      .wadr(yt_rsc_3_30_wadr),
      .we(yt_rsc_3_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_3_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_3_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_3_31_clkr_en),
      .d(yt_rsc_3_31_d),
      .q(yt_rsc_3_31_q),
      .radr(yt_rsc_3_31_radr),
      .wadr(yt_rsc_3_31_wadr),
      .we(yt_rsc_3_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_0_clkr_en),
      .d(yt_rsc_4_0_d),
      .q(yt_rsc_4_0_q),
      .radr(yt_rsc_4_0_radr),
      .wadr(yt_rsc_4_0_wadr),
      .we(yt_rsc_4_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_1_clkr_en),
      .d(yt_rsc_4_1_d),
      .q(yt_rsc_4_1_q),
      .radr(yt_rsc_4_1_radr),
      .wadr(yt_rsc_4_1_wadr),
      .we(yt_rsc_4_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_2_clkr_en),
      .d(yt_rsc_4_2_d),
      .q(yt_rsc_4_2_q),
      .radr(yt_rsc_4_2_radr),
      .wadr(yt_rsc_4_2_wadr),
      .we(yt_rsc_4_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_3_clkr_en),
      .d(yt_rsc_4_3_d),
      .q(yt_rsc_4_3_q),
      .radr(yt_rsc_4_3_radr),
      .wadr(yt_rsc_4_3_wadr),
      .we(yt_rsc_4_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_4_clkr_en),
      .d(yt_rsc_4_4_d),
      .q(yt_rsc_4_4_q),
      .radr(yt_rsc_4_4_radr),
      .wadr(yt_rsc_4_4_wadr),
      .we(yt_rsc_4_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_5_clkr_en),
      .d(yt_rsc_4_5_d),
      .q(yt_rsc_4_5_q),
      .radr(yt_rsc_4_5_radr),
      .wadr(yt_rsc_4_5_wadr),
      .we(yt_rsc_4_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_6_clkr_en),
      .d(yt_rsc_4_6_d),
      .q(yt_rsc_4_6_q),
      .radr(yt_rsc_4_6_radr),
      .wadr(yt_rsc_4_6_wadr),
      .we(yt_rsc_4_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_7_clkr_en),
      .d(yt_rsc_4_7_d),
      .q(yt_rsc_4_7_q),
      .radr(yt_rsc_4_7_radr),
      .wadr(yt_rsc_4_7_wadr),
      .we(yt_rsc_4_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_8_clkr_en),
      .d(yt_rsc_4_8_d),
      .q(yt_rsc_4_8_q),
      .radr(yt_rsc_4_8_radr),
      .wadr(yt_rsc_4_8_wadr),
      .we(yt_rsc_4_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_9_clkr_en),
      .d(yt_rsc_4_9_d),
      .q(yt_rsc_4_9_q),
      .radr(yt_rsc_4_9_radr),
      .wadr(yt_rsc_4_9_wadr),
      .we(yt_rsc_4_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_10_clkr_en),
      .d(yt_rsc_4_10_d),
      .q(yt_rsc_4_10_q),
      .radr(yt_rsc_4_10_radr),
      .wadr(yt_rsc_4_10_wadr),
      .we(yt_rsc_4_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_11_clkr_en),
      .d(yt_rsc_4_11_d),
      .q(yt_rsc_4_11_q),
      .radr(yt_rsc_4_11_radr),
      .wadr(yt_rsc_4_11_wadr),
      .we(yt_rsc_4_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_12_clkr_en),
      .d(yt_rsc_4_12_d),
      .q(yt_rsc_4_12_q),
      .radr(yt_rsc_4_12_radr),
      .wadr(yt_rsc_4_12_wadr),
      .we(yt_rsc_4_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_13_clkr_en),
      .d(yt_rsc_4_13_d),
      .q(yt_rsc_4_13_q),
      .radr(yt_rsc_4_13_radr),
      .wadr(yt_rsc_4_13_wadr),
      .we(yt_rsc_4_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_14_clkr_en),
      .d(yt_rsc_4_14_d),
      .q(yt_rsc_4_14_q),
      .radr(yt_rsc_4_14_radr),
      .wadr(yt_rsc_4_14_wadr),
      .we(yt_rsc_4_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_15_clkr_en),
      .d(yt_rsc_4_15_d),
      .q(yt_rsc_4_15_q),
      .radr(yt_rsc_4_15_radr),
      .wadr(yt_rsc_4_15_wadr),
      .we(yt_rsc_4_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_16_clkr_en),
      .d(yt_rsc_4_16_d),
      .q(yt_rsc_4_16_q),
      .radr(yt_rsc_4_16_radr),
      .wadr(yt_rsc_4_16_wadr),
      .we(yt_rsc_4_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_17_clkr_en),
      .d(yt_rsc_4_17_d),
      .q(yt_rsc_4_17_q),
      .radr(yt_rsc_4_17_radr),
      .wadr(yt_rsc_4_17_wadr),
      .we(yt_rsc_4_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_18_clkr_en),
      .d(yt_rsc_4_18_d),
      .q(yt_rsc_4_18_q),
      .radr(yt_rsc_4_18_radr),
      .wadr(yt_rsc_4_18_wadr),
      .we(yt_rsc_4_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_19_clkr_en),
      .d(yt_rsc_4_19_d),
      .q(yt_rsc_4_19_q),
      .radr(yt_rsc_4_19_radr),
      .wadr(yt_rsc_4_19_wadr),
      .we(yt_rsc_4_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_20_clkr_en),
      .d(yt_rsc_4_20_d),
      .q(yt_rsc_4_20_q),
      .radr(yt_rsc_4_20_radr),
      .wadr(yt_rsc_4_20_wadr),
      .we(yt_rsc_4_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_21_clkr_en),
      .d(yt_rsc_4_21_d),
      .q(yt_rsc_4_21_q),
      .radr(yt_rsc_4_21_radr),
      .wadr(yt_rsc_4_21_wadr),
      .we(yt_rsc_4_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_22_clkr_en),
      .d(yt_rsc_4_22_d),
      .q(yt_rsc_4_22_q),
      .radr(yt_rsc_4_22_radr),
      .wadr(yt_rsc_4_22_wadr),
      .we(yt_rsc_4_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_23_clkr_en),
      .d(yt_rsc_4_23_d),
      .q(yt_rsc_4_23_q),
      .radr(yt_rsc_4_23_radr),
      .wadr(yt_rsc_4_23_wadr),
      .we(yt_rsc_4_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_24_clkr_en),
      .d(yt_rsc_4_24_d),
      .q(yt_rsc_4_24_q),
      .radr(yt_rsc_4_24_radr),
      .wadr(yt_rsc_4_24_wadr),
      .we(yt_rsc_4_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_25_clkr_en),
      .d(yt_rsc_4_25_d),
      .q(yt_rsc_4_25_q),
      .radr(yt_rsc_4_25_radr),
      .wadr(yt_rsc_4_25_wadr),
      .we(yt_rsc_4_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_26_clkr_en),
      .d(yt_rsc_4_26_d),
      .q(yt_rsc_4_26_q),
      .radr(yt_rsc_4_26_radr),
      .wadr(yt_rsc_4_26_wadr),
      .we(yt_rsc_4_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_27_clkr_en),
      .d(yt_rsc_4_27_d),
      .q(yt_rsc_4_27_q),
      .radr(yt_rsc_4_27_radr),
      .wadr(yt_rsc_4_27_wadr),
      .we(yt_rsc_4_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_28_clkr_en),
      .d(yt_rsc_4_28_d),
      .q(yt_rsc_4_28_q),
      .radr(yt_rsc_4_28_radr),
      .wadr(yt_rsc_4_28_wadr),
      .we(yt_rsc_4_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_29_clkr_en),
      .d(yt_rsc_4_29_d),
      .q(yt_rsc_4_29_q),
      .radr(yt_rsc_4_29_radr),
      .wadr(yt_rsc_4_29_wadr),
      .we(yt_rsc_4_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_30_clkr_en),
      .d(yt_rsc_4_30_d),
      .q(yt_rsc_4_30_q),
      .radr(yt_rsc_4_30_radr),
      .wadr(yt_rsc_4_30_wadr),
      .we(yt_rsc_4_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_4_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_4_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_4_31_clkr_en),
      .d(yt_rsc_4_31_d),
      .q(yt_rsc_4_31_q),
      .radr(yt_rsc_4_31_radr),
      .wadr(yt_rsc_4_31_wadr),
      .we(yt_rsc_4_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_0_clkr_en),
      .d(yt_rsc_5_0_d),
      .q(yt_rsc_5_0_q),
      .radr(yt_rsc_5_0_radr),
      .wadr(yt_rsc_5_0_wadr),
      .we(yt_rsc_5_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_1_clkr_en),
      .d(yt_rsc_5_1_d),
      .q(yt_rsc_5_1_q),
      .radr(yt_rsc_5_1_radr),
      .wadr(yt_rsc_5_1_wadr),
      .we(yt_rsc_5_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_2_clkr_en),
      .d(yt_rsc_5_2_d),
      .q(yt_rsc_5_2_q),
      .radr(yt_rsc_5_2_radr),
      .wadr(yt_rsc_5_2_wadr),
      .we(yt_rsc_5_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_3_clkr_en),
      .d(yt_rsc_5_3_d),
      .q(yt_rsc_5_3_q),
      .radr(yt_rsc_5_3_radr),
      .wadr(yt_rsc_5_3_wadr),
      .we(yt_rsc_5_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_4_clkr_en),
      .d(yt_rsc_5_4_d),
      .q(yt_rsc_5_4_q),
      .radr(yt_rsc_5_4_radr),
      .wadr(yt_rsc_5_4_wadr),
      .we(yt_rsc_5_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_5_clkr_en),
      .d(yt_rsc_5_5_d),
      .q(yt_rsc_5_5_q),
      .radr(yt_rsc_5_5_radr),
      .wadr(yt_rsc_5_5_wadr),
      .we(yt_rsc_5_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_6_clkr_en),
      .d(yt_rsc_5_6_d),
      .q(yt_rsc_5_6_q),
      .radr(yt_rsc_5_6_radr),
      .wadr(yt_rsc_5_6_wadr),
      .we(yt_rsc_5_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_7_clkr_en),
      .d(yt_rsc_5_7_d),
      .q(yt_rsc_5_7_q),
      .radr(yt_rsc_5_7_radr),
      .wadr(yt_rsc_5_7_wadr),
      .we(yt_rsc_5_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_8_clkr_en),
      .d(yt_rsc_5_8_d),
      .q(yt_rsc_5_8_q),
      .radr(yt_rsc_5_8_radr),
      .wadr(yt_rsc_5_8_wadr),
      .we(yt_rsc_5_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_9_clkr_en),
      .d(yt_rsc_5_9_d),
      .q(yt_rsc_5_9_q),
      .radr(yt_rsc_5_9_radr),
      .wadr(yt_rsc_5_9_wadr),
      .we(yt_rsc_5_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_10_clkr_en),
      .d(yt_rsc_5_10_d),
      .q(yt_rsc_5_10_q),
      .radr(yt_rsc_5_10_radr),
      .wadr(yt_rsc_5_10_wadr),
      .we(yt_rsc_5_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_11_clkr_en),
      .d(yt_rsc_5_11_d),
      .q(yt_rsc_5_11_q),
      .radr(yt_rsc_5_11_radr),
      .wadr(yt_rsc_5_11_wadr),
      .we(yt_rsc_5_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_12_clkr_en),
      .d(yt_rsc_5_12_d),
      .q(yt_rsc_5_12_q),
      .radr(yt_rsc_5_12_radr),
      .wadr(yt_rsc_5_12_wadr),
      .we(yt_rsc_5_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_13_clkr_en),
      .d(yt_rsc_5_13_d),
      .q(yt_rsc_5_13_q),
      .radr(yt_rsc_5_13_radr),
      .wadr(yt_rsc_5_13_wadr),
      .we(yt_rsc_5_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_14_clkr_en),
      .d(yt_rsc_5_14_d),
      .q(yt_rsc_5_14_q),
      .radr(yt_rsc_5_14_radr),
      .wadr(yt_rsc_5_14_wadr),
      .we(yt_rsc_5_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_15_clkr_en),
      .d(yt_rsc_5_15_d),
      .q(yt_rsc_5_15_q),
      .radr(yt_rsc_5_15_radr),
      .wadr(yt_rsc_5_15_wadr),
      .we(yt_rsc_5_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_16_clkr_en),
      .d(yt_rsc_5_16_d),
      .q(yt_rsc_5_16_q),
      .radr(yt_rsc_5_16_radr),
      .wadr(yt_rsc_5_16_wadr),
      .we(yt_rsc_5_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_17_clkr_en),
      .d(yt_rsc_5_17_d),
      .q(yt_rsc_5_17_q),
      .radr(yt_rsc_5_17_radr),
      .wadr(yt_rsc_5_17_wadr),
      .we(yt_rsc_5_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_18_clkr_en),
      .d(yt_rsc_5_18_d),
      .q(yt_rsc_5_18_q),
      .radr(yt_rsc_5_18_radr),
      .wadr(yt_rsc_5_18_wadr),
      .we(yt_rsc_5_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_19_clkr_en),
      .d(yt_rsc_5_19_d),
      .q(yt_rsc_5_19_q),
      .radr(yt_rsc_5_19_radr),
      .wadr(yt_rsc_5_19_wadr),
      .we(yt_rsc_5_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_20_clkr_en),
      .d(yt_rsc_5_20_d),
      .q(yt_rsc_5_20_q),
      .radr(yt_rsc_5_20_radr),
      .wadr(yt_rsc_5_20_wadr),
      .we(yt_rsc_5_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_21_clkr_en),
      .d(yt_rsc_5_21_d),
      .q(yt_rsc_5_21_q),
      .radr(yt_rsc_5_21_radr),
      .wadr(yt_rsc_5_21_wadr),
      .we(yt_rsc_5_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_22_clkr_en),
      .d(yt_rsc_5_22_d),
      .q(yt_rsc_5_22_q),
      .radr(yt_rsc_5_22_radr),
      .wadr(yt_rsc_5_22_wadr),
      .we(yt_rsc_5_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_23_clkr_en),
      .d(yt_rsc_5_23_d),
      .q(yt_rsc_5_23_q),
      .radr(yt_rsc_5_23_radr),
      .wadr(yt_rsc_5_23_wadr),
      .we(yt_rsc_5_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_24_clkr_en),
      .d(yt_rsc_5_24_d),
      .q(yt_rsc_5_24_q),
      .radr(yt_rsc_5_24_radr),
      .wadr(yt_rsc_5_24_wadr),
      .we(yt_rsc_5_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_25_clkr_en),
      .d(yt_rsc_5_25_d),
      .q(yt_rsc_5_25_q),
      .radr(yt_rsc_5_25_radr),
      .wadr(yt_rsc_5_25_wadr),
      .we(yt_rsc_5_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_26_clkr_en),
      .d(yt_rsc_5_26_d),
      .q(yt_rsc_5_26_q),
      .radr(yt_rsc_5_26_radr),
      .wadr(yt_rsc_5_26_wadr),
      .we(yt_rsc_5_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_27_clkr_en),
      .d(yt_rsc_5_27_d),
      .q(yt_rsc_5_27_q),
      .radr(yt_rsc_5_27_radr),
      .wadr(yt_rsc_5_27_wadr),
      .we(yt_rsc_5_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_28_clkr_en),
      .d(yt_rsc_5_28_d),
      .q(yt_rsc_5_28_q),
      .radr(yt_rsc_5_28_radr),
      .wadr(yt_rsc_5_28_wadr),
      .we(yt_rsc_5_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_29_clkr_en),
      .d(yt_rsc_5_29_d),
      .q(yt_rsc_5_29_q),
      .radr(yt_rsc_5_29_radr),
      .wadr(yt_rsc_5_29_wadr),
      .we(yt_rsc_5_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_30_clkr_en),
      .d(yt_rsc_5_30_d),
      .q(yt_rsc_5_30_q),
      .radr(yt_rsc_5_30_radr),
      .wadr(yt_rsc_5_30_wadr),
      .we(yt_rsc_5_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_5_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_5_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_5_31_clkr_en),
      .d(yt_rsc_5_31_d),
      .q(yt_rsc_5_31_q),
      .radr(yt_rsc_5_31_radr),
      .wadr(yt_rsc_5_31_wadr),
      .we(yt_rsc_5_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_0_clkr_en),
      .d(yt_rsc_6_0_d),
      .q(yt_rsc_6_0_q),
      .radr(yt_rsc_6_0_radr),
      .wadr(yt_rsc_6_0_wadr),
      .we(yt_rsc_6_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_1_clkr_en),
      .d(yt_rsc_6_1_d),
      .q(yt_rsc_6_1_q),
      .radr(yt_rsc_6_1_radr),
      .wadr(yt_rsc_6_1_wadr),
      .we(yt_rsc_6_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_2_clkr_en),
      .d(yt_rsc_6_2_d),
      .q(yt_rsc_6_2_q),
      .radr(yt_rsc_6_2_radr),
      .wadr(yt_rsc_6_2_wadr),
      .we(yt_rsc_6_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_3_clkr_en),
      .d(yt_rsc_6_3_d),
      .q(yt_rsc_6_3_q),
      .radr(yt_rsc_6_3_radr),
      .wadr(yt_rsc_6_3_wadr),
      .we(yt_rsc_6_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_4_clkr_en),
      .d(yt_rsc_6_4_d),
      .q(yt_rsc_6_4_q),
      .radr(yt_rsc_6_4_radr),
      .wadr(yt_rsc_6_4_wadr),
      .we(yt_rsc_6_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_5_clkr_en),
      .d(yt_rsc_6_5_d),
      .q(yt_rsc_6_5_q),
      .radr(yt_rsc_6_5_radr),
      .wadr(yt_rsc_6_5_wadr),
      .we(yt_rsc_6_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_6_clkr_en),
      .d(yt_rsc_6_6_d),
      .q(yt_rsc_6_6_q),
      .radr(yt_rsc_6_6_radr),
      .wadr(yt_rsc_6_6_wadr),
      .we(yt_rsc_6_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_7_clkr_en),
      .d(yt_rsc_6_7_d),
      .q(yt_rsc_6_7_q),
      .radr(yt_rsc_6_7_radr),
      .wadr(yt_rsc_6_7_wadr),
      .we(yt_rsc_6_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_8_clkr_en),
      .d(yt_rsc_6_8_d),
      .q(yt_rsc_6_8_q),
      .radr(yt_rsc_6_8_radr),
      .wadr(yt_rsc_6_8_wadr),
      .we(yt_rsc_6_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_9_clkr_en),
      .d(yt_rsc_6_9_d),
      .q(yt_rsc_6_9_q),
      .radr(yt_rsc_6_9_radr),
      .wadr(yt_rsc_6_9_wadr),
      .we(yt_rsc_6_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_10_clkr_en),
      .d(yt_rsc_6_10_d),
      .q(yt_rsc_6_10_q),
      .radr(yt_rsc_6_10_radr),
      .wadr(yt_rsc_6_10_wadr),
      .we(yt_rsc_6_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_11_clkr_en),
      .d(yt_rsc_6_11_d),
      .q(yt_rsc_6_11_q),
      .radr(yt_rsc_6_11_radr),
      .wadr(yt_rsc_6_11_wadr),
      .we(yt_rsc_6_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_12_clkr_en),
      .d(yt_rsc_6_12_d),
      .q(yt_rsc_6_12_q),
      .radr(yt_rsc_6_12_radr),
      .wadr(yt_rsc_6_12_wadr),
      .we(yt_rsc_6_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_13_clkr_en),
      .d(yt_rsc_6_13_d),
      .q(yt_rsc_6_13_q),
      .radr(yt_rsc_6_13_radr),
      .wadr(yt_rsc_6_13_wadr),
      .we(yt_rsc_6_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_14_clkr_en),
      .d(yt_rsc_6_14_d),
      .q(yt_rsc_6_14_q),
      .radr(yt_rsc_6_14_radr),
      .wadr(yt_rsc_6_14_wadr),
      .we(yt_rsc_6_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_15_clkr_en),
      .d(yt_rsc_6_15_d),
      .q(yt_rsc_6_15_q),
      .radr(yt_rsc_6_15_radr),
      .wadr(yt_rsc_6_15_wadr),
      .we(yt_rsc_6_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_16_clkr_en),
      .d(yt_rsc_6_16_d),
      .q(yt_rsc_6_16_q),
      .radr(yt_rsc_6_16_radr),
      .wadr(yt_rsc_6_16_wadr),
      .we(yt_rsc_6_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_17_clkr_en),
      .d(yt_rsc_6_17_d),
      .q(yt_rsc_6_17_q),
      .radr(yt_rsc_6_17_radr),
      .wadr(yt_rsc_6_17_wadr),
      .we(yt_rsc_6_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_18_clkr_en),
      .d(yt_rsc_6_18_d),
      .q(yt_rsc_6_18_q),
      .radr(yt_rsc_6_18_radr),
      .wadr(yt_rsc_6_18_wadr),
      .we(yt_rsc_6_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_19_clkr_en),
      .d(yt_rsc_6_19_d),
      .q(yt_rsc_6_19_q),
      .radr(yt_rsc_6_19_radr),
      .wadr(yt_rsc_6_19_wadr),
      .we(yt_rsc_6_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_20_clkr_en),
      .d(yt_rsc_6_20_d),
      .q(yt_rsc_6_20_q),
      .radr(yt_rsc_6_20_radr),
      .wadr(yt_rsc_6_20_wadr),
      .we(yt_rsc_6_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_21_clkr_en),
      .d(yt_rsc_6_21_d),
      .q(yt_rsc_6_21_q),
      .radr(yt_rsc_6_21_radr),
      .wadr(yt_rsc_6_21_wadr),
      .we(yt_rsc_6_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_22_clkr_en),
      .d(yt_rsc_6_22_d),
      .q(yt_rsc_6_22_q),
      .radr(yt_rsc_6_22_radr),
      .wadr(yt_rsc_6_22_wadr),
      .we(yt_rsc_6_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_23_clkr_en),
      .d(yt_rsc_6_23_d),
      .q(yt_rsc_6_23_q),
      .radr(yt_rsc_6_23_radr),
      .wadr(yt_rsc_6_23_wadr),
      .we(yt_rsc_6_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_24_clkr_en),
      .d(yt_rsc_6_24_d),
      .q(yt_rsc_6_24_q),
      .radr(yt_rsc_6_24_radr),
      .wadr(yt_rsc_6_24_wadr),
      .we(yt_rsc_6_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_25_clkr_en),
      .d(yt_rsc_6_25_d),
      .q(yt_rsc_6_25_q),
      .radr(yt_rsc_6_25_radr),
      .wadr(yt_rsc_6_25_wadr),
      .we(yt_rsc_6_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_26_clkr_en),
      .d(yt_rsc_6_26_d),
      .q(yt_rsc_6_26_q),
      .radr(yt_rsc_6_26_radr),
      .wadr(yt_rsc_6_26_wadr),
      .we(yt_rsc_6_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_27_clkr_en),
      .d(yt_rsc_6_27_d),
      .q(yt_rsc_6_27_q),
      .radr(yt_rsc_6_27_radr),
      .wadr(yt_rsc_6_27_wadr),
      .we(yt_rsc_6_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_28_clkr_en),
      .d(yt_rsc_6_28_d),
      .q(yt_rsc_6_28_q),
      .radr(yt_rsc_6_28_radr),
      .wadr(yt_rsc_6_28_wadr),
      .we(yt_rsc_6_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_29_clkr_en),
      .d(yt_rsc_6_29_d),
      .q(yt_rsc_6_29_q),
      .radr(yt_rsc_6_29_radr),
      .wadr(yt_rsc_6_29_wadr),
      .we(yt_rsc_6_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_30_clkr_en),
      .d(yt_rsc_6_30_d),
      .q(yt_rsc_6_30_q),
      .radr(yt_rsc_6_30_radr),
      .wadr(yt_rsc_6_30_wadr),
      .we(yt_rsc_6_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_6_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_6_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_6_31_clkr_en),
      .d(yt_rsc_6_31_d),
      .q(yt_rsc_6_31_q),
      .radr(yt_rsc_6_31_radr),
      .wadr(yt_rsc_6_31_wadr),
      .we(yt_rsc_6_31_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_0_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_0_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_0_clkr_en),
      .d(yt_rsc_7_0_d),
      .q(yt_rsc_7_0_q),
      .radr(yt_rsc_7_0_radr),
      .wadr(yt_rsc_7_0_wadr),
      .we(yt_rsc_7_0_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_1_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_1_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_1_clkr_en),
      .d(yt_rsc_7_1_d),
      .q(yt_rsc_7_1_q),
      .radr(yt_rsc_7_1_radr),
      .wadr(yt_rsc_7_1_wadr),
      .we(yt_rsc_7_1_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_2_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_2_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_2_clkr_en),
      .d(yt_rsc_7_2_d),
      .q(yt_rsc_7_2_q),
      .radr(yt_rsc_7_2_radr),
      .wadr(yt_rsc_7_2_wadr),
      .we(yt_rsc_7_2_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_3_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_3_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_3_clkr_en),
      .d(yt_rsc_7_3_d),
      .q(yt_rsc_7_3_q),
      .radr(yt_rsc_7_3_radr),
      .wadr(yt_rsc_7_3_wadr),
      .we(yt_rsc_7_3_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_4_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_4_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_4_clkr_en),
      .d(yt_rsc_7_4_d),
      .q(yt_rsc_7_4_q),
      .radr(yt_rsc_7_4_radr),
      .wadr(yt_rsc_7_4_wadr),
      .we(yt_rsc_7_4_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_5_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_5_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_5_clkr_en),
      .d(yt_rsc_7_5_d),
      .q(yt_rsc_7_5_q),
      .radr(yt_rsc_7_5_radr),
      .wadr(yt_rsc_7_5_wadr),
      .we(yt_rsc_7_5_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_6_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_6_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_6_clkr_en),
      .d(yt_rsc_7_6_d),
      .q(yt_rsc_7_6_q),
      .radr(yt_rsc_7_6_radr),
      .wadr(yt_rsc_7_6_wadr),
      .we(yt_rsc_7_6_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_7_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_7_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_7_clkr_en),
      .d(yt_rsc_7_7_d),
      .q(yt_rsc_7_7_q),
      .radr(yt_rsc_7_7_radr),
      .wadr(yt_rsc_7_7_wadr),
      .we(yt_rsc_7_7_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_8_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_8_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_8_clkr_en),
      .d(yt_rsc_7_8_d),
      .q(yt_rsc_7_8_q),
      .radr(yt_rsc_7_8_radr),
      .wadr(yt_rsc_7_8_wadr),
      .we(yt_rsc_7_8_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_9_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_9_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_9_clkr_en),
      .d(yt_rsc_7_9_d),
      .q(yt_rsc_7_9_q),
      .radr(yt_rsc_7_9_radr),
      .wadr(yt_rsc_7_9_wadr),
      .we(yt_rsc_7_9_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_10_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_10_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_10_clkr_en),
      .d(yt_rsc_7_10_d),
      .q(yt_rsc_7_10_q),
      .radr(yt_rsc_7_10_radr),
      .wadr(yt_rsc_7_10_wadr),
      .we(yt_rsc_7_10_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_11_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_11_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_11_clkr_en),
      .d(yt_rsc_7_11_d),
      .q(yt_rsc_7_11_q),
      .radr(yt_rsc_7_11_radr),
      .wadr(yt_rsc_7_11_wadr),
      .we(yt_rsc_7_11_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_12_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_12_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_12_clkr_en),
      .d(yt_rsc_7_12_d),
      .q(yt_rsc_7_12_q),
      .radr(yt_rsc_7_12_radr),
      .wadr(yt_rsc_7_12_wadr),
      .we(yt_rsc_7_12_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_13_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_13_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_13_clkr_en),
      .d(yt_rsc_7_13_d),
      .q(yt_rsc_7_13_q),
      .radr(yt_rsc_7_13_radr),
      .wadr(yt_rsc_7_13_wadr),
      .we(yt_rsc_7_13_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_14_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_14_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_14_clkr_en),
      .d(yt_rsc_7_14_d),
      .q(yt_rsc_7_14_q),
      .radr(yt_rsc_7_14_radr),
      .wadr(yt_rsc_7_14_wadr),
      .we(yt_rsc_7_14_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_15_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_15_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_15_clkr_en),
      .d(yt_rsc_7_15_d),
      .q(yt_rsc_7_15_q),
      .radr(yt_rsc_7_15_radr),
      .wadr(yt_rsc_7_15_wadr),
      .we(yt_rsc_7_15_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_16_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_16_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_16_clkr_en),
      .d(yt_rsc_7_16_d),
      .q(yt_rsc_7_16_q),
      .radr(yt_rsc_7_16_radr),
      .wadr(yt_rsc_7_16_wadr),
      .we(yt_rsc_7_16_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_17_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_17_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_17_clkr_en),
      .d(yt_rsc_7_17_d),
      .q(yt_rsc_7_17_q),
      .radr(yt_rsc_7_17_radr),
      .wadr(yt_rsc_7_17_wadr),
      .we(yt_rsc_7_17_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_18_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_18_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_18_clkr_en),
      .d(yt_rsc_7_18_d),
      .q(yt_rsc_7_18_q),
      .radr(yt_rsc_7_18_radr),
      .wadr(yt_rsc_7_18_wadr),
      .we(yt_rsc_7_18_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_19_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_19_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_19_clkr_en),
      .d(yt_rsc_7_19_d),
      .q(yt_rsc_7_19_q),
      .radr(yt_rsc_7_19_radr),
      .wadr(yt_rsc_7_19_wadr),
      .we(yt_rsc_7_19_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_20_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_20_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_20_clkr_en),
      .d(yt_rsc_7_20_d),
      .q(yt_rsc_7_20_q),
      .radr(yt_rsc_7_20_radr),
      .wadr(yt_rsc_7_20_wadr),
      .we(yt_rsc_7_20_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_21_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_21_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_21_clkr_en),
      .d(yt_rsc_7_21_d),
      .q(yt_rsc_7_21_q),
      .radr(yt_rsc_7_21_radr),
      .wadr(yt_rsc_7_21_wadr),
      .we(yt_rsc_7_21_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_22_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_22_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_22_clkr_en),
      .d(yt_rsc_7_22_d),
      .q(yt_rsc_7_22_q),
      .radr(yt_rsc_7_22_radr),
      .wadr(yt_rsc_7_22_wadr),
      .we(yt_rsc_7_22_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_23_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_23_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_23_clkr_en),
      .d(yt_rsc_7_23_d),
      .q(yt_rsc_7_23_q),
      .radr(yt_rsc_7_23_radr),
      .wadr(yt_rsc_7_23_wadr),
      .we(yt_rsc_7_23_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_24_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_24_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_24_clkr_en),
      .d(yt_rsc_7_24_d),
      .q(yt_rsc_7_24_q),
      .radr(yt_rsc_7_24_radr),
      .wadr(yt_rsc_7_24_wadr),
      .we(yt_rsc_7_24_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_25_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_25_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_25_clkr_en),
      .d(yt_rsc_7_25_d),
      .q(yt_rsc_7_25_q),
      .radr(yt_rsc_7_25_radr),
      .wadr(yt_rsc_7_25_wadr),
      .we(yt_rsc_7_25_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_26_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_26_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_26_clkr_en),
      .d(yt_rsc_7_26_d),
      .q(yt_rsc_7_26_q),
      .radr(yt_rsc_7_26_radr),
      .wadr(yt_rsc_7_26_wadr),
      .we(yt_rsc_7_26_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_27_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_27_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_27_clkr_en),
      .d(yt_rsc_7_27_d),
      .q(yt_rsc_7_27_q),
      .radr(yt_rsc_7_27_radr),
      .wadr(yt_rsc_7_27_wadr),
      .we(yt_rsc_7_27_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_28_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_28_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_28_clkr_en),
      .d(yt_rsc_7_28_d),
      .q(yt_rsc_7_28_q),
      .radr(yt_rsc_7_28_radr),
      .wadr(yt_rsc_7_28_wadr),
      .we(yt_rsc_7_28_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_29_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_29_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_29_clkr_en),
      .d(yt_rsc_7_29_d),
      .q(yt_rsc_7_29_q),
      .radr(yt_rsc_7_29_radr),
      .wadr(yt_rsc_7_29_wadr),
      .we(yt_rsc_7_29_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_30_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_30_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_30_clkr_en),
      .d(yt_rsc_7_30_d),
      .q(yt_rsc_7_30_q),
      .radr(yt_rsc_7_30_radr),
      .wadr(yt_rsc_7_30_wadr),
      .we(yt_rsc_7_30_we)
    );
  BLOCK_1R1W_RBW_DUAL #(.addr_width(32'sd4),
  .data_width(32'sd32),
  .depth(32'sd16),
  .latency(32'sd1)) yt_rsc_7_31_comp (
      .clkr(clk),
      .clkr_en(yt_rsc_7_31_clkr_en),
      .clkw(clk),
      .clkw_en(yt_rsc_7_31_clkr_en),
      .d(yt_rsc_7_31_d),
      .q(yt_rsc_7_31_q),
      .radr(yt_rsc_7_31_radr),
      .wadr(yt_rsc_7_31_wadr),
      .we(yt_rsc_7_31_we)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_7_4_32_16_16_32_1_gen yt_rsc_0_0_i
      (
      .clkr_en(yt_rsc_0_0_clkr_en),
      .clkw_en(yt_rsc_0_0_clkw_en),
      .q(yt_rsc_0_0_q),
      .radr(yt_rsc_0_0_radr),
      .we(yt_rsc_0_0_we),
      .d(yt_rsc_0_0_d),
      .wadr(yt_rsc_0_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_0_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_8_4_32_16_16_32_1_gen yt_rsc_0_1_i
      (
      .clkr_en(yt_rsc_0_1_clkr_en),
      .clkw_en(yt_rsc_0_1_clkw_en),
      .q(yt_rsc_0_1_q),
      .radr(yt_rsc_0_1_radr),
      .we(yt_rsc_0_1_we),
      .d(yt_rsc_0_1_d),
      .wadr(yt_rsc_0_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_0_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_9_4_32_16_16_32_1_gen yt_rsc_0_2_i
      (
      .clkr_en(yt_rsc_0_2_clkr_en),
      .clkw_en(yt_rsc_0_2_clkw_en),
      .q(yt_rsc_0_2_q),
      .radr(yt_rsc_0_2_radr),
      .we(yt_rsc_0_2_we),
      .d(yt_rsc_0_2_d),
      .wadr(yt_rsc_0_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_0_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_10_4_32_16_16_32_1_gen yt_rsc_0_3_i
      (
      .clkr_en(yt_rsc_0_3_clkr_en),
      .clkw_en(yt_rsc_0_3_clkw_en),
      .q(yt_rsc_0_3_q),
      .radr(yt_rsc_0_3_radr),
      .we(yt_rsc_0_3_we),
      .d(yt_rsc_0_3_d),
      .wadr(yt_rsc_0_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_0_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_11_4_32_16_16_32_1_gen yt_rsc_0_4_i
      (
      .clkr_en(yt_rsc_0_4_clkr_en),
      .clkw_en(yt_rsc_0_4_clkw_en),
      .q(yt_rsc_0_4_q),
      .radr(yt_rsc_0_4_radr),
      .we(yt_rsc_0_4_we),
      .d(yt_rsc_0_4_d),
      .wadr(yt_rsc_0_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_0_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_12_4_32_16_16_32_1_gen yt_rsc_0_5_i
      (
      .clkr_en(yt_rsc_0_5_clkr_en),
      .clkw_en(yt_rsc_0_5_clkw_en),
      .q(yt_rsc_0_5_q),
      .radr(yt_rsc_0_5_radr),
      .we(yt_rsc_0_5_we),
      .d(yt_rsc_0_5_d),
      .wadr(yt_rsc_0_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_0_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_13_4_32_16_16_32_1_gen yt_rsc_0_6_i
      (
      .clkr_en(yt_rsc_0_6_clkr_en),
      .clkw_en(yt_rsc_0_6_clkw_en),
      .q(yt_rsc_0_6_q),
      .radr(yt_rsc_0_6_radr),
      .we(yt_rsc_0_6_we),
      .d(yt_rsc_0_6_d),
      .wadr(yt_rsc_0_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_0_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_14_4_32_16_16_32_1_gen yt_rsc_0_7_i
      (
      .clkr_en(yt_rsc_0_7_clkr_en),
      .clkw_en(yt_rsc_0_7_clkw_en),
      .q(yt_rsc_0_7_q),
      .radr(yt_rsc_0_7_radr),
      .we(yt_rsc_0_7_we),
      .d(yt_rsc_0_7_d),
      .wadr(yt_rsc_0_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_0_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_15_4_32_16_16_32_1_gen yt_rsc_0_8_i
      (
      .clkr_en(yt_rsc_0_8_clkr_en),
      .clkw_en(yt_rsc_0_8_clkw_en),
      .q(yt_rsc_0_8_q),
      .radr(yt_rsc_0_8_radr),
      .we(yt_rsc_0_8_we),
      .d(yt_rsc_0_8_d),
      .wadr(yt_rsc_0_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_0_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_16_4_32_16_16_32_1_gen yt_rsc_0_9_i
      (
      .clkr_en(yt_rsc_0_9_clkr_en),
      .clkw_en(yt_rsc_0_9_clkw_en),
      .q(yt_rsc_0_9_q),
      .radr(yt_rsc_0_9_radr),
      .we(yt_rsc_0_9_we),
      .d(yt_rsc_0_9_d),
      .wadr(yt_rsc_0_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_0_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_17_4_32_16_16_32_1_gen yt_rsc_0_10_i
      (
      .clkr_en(yt_rsc_0_10_clkr_en),
      .clkw_en(yt_rsc_0_10_clkw_en),
      .q(yt_rsc_0_10_q),
      .radr(yt_rsc_0_10_radr),
      .we(yt_rsc_0_10_we),
      .d(yt_rsc_0_10_d),
      .wadr(yt_rsc_0_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_0_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_18_4_32_16_16_32_1_gen yt_rsc_0_11_i
      (
      .clkr_en(yt_rsc_0_11_clkr_en),
      .clkw_en(yt_rsc_0_11_clkw_en),
      .q(yt_rsc_0_11_q),
      .radr(yt_rsc_0_11_radr),
      .we(yt_rsc_0_11_we),
      .d(yt_rsc_0_11_d),
      .wadr(yt_rsc_0_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_0_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_19_4_32_16_16_32_1_gen yt_rsc_0_12_i
      (
      .clkr_en(yt_rsc_0_12_clkr_en),
      .clkw_en(yt_rsc_0_12_clkw_en),
      .q(yt_rsc_0_12_q),
      .radr(yt_rsc_0_12_radr),
      .we(yt_rsc_0_12_we),
      .d(yt_rsc_0_12_d),
      .wadr(yt_rsc_0_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_0_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_20_4_32_16_16_32_1_gen yt_rsc_0_13_i
      (
      .clkr_en(yt_rsc_0_13_clkr_en),
      .clkw_en(yt_rsc_0_13_clkw_en),
      .q(yt_rsc_0_13_q),
      .radr(yt_rsc_0_13_radr),
      .we(yt_rsc_0_13_we),
      .d(yt_rsc_0_13_d),
      .wadr(yt_rsc_0_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_0_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_21_4_32_16_16_32_1_gen yt_rsc_0_14_i
      (
      .clkr_en(yt_rsc_0_14_clkr_en),
      .clkw_en(yt_rsc_0_14_clkw_en),
      .q(yt_rsc_0_14_q),
      .radr(yt_rsc_0_14_radr),
      .we(yt_rsc_0_14_we),
      .d(yt_rsc_0_14_d),
      .wadr(yt_rsc_0_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_0_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_22_4_32_16_16_32_1_gen yt_rsc_0_15_i
      (
      .clkr_en(yt_rsc_0_15_clkr_en),
      .clkw_en(yt_rsc_0_15_clkw_en),
      .q(yt_rsc_0_15_q),
      .radr(yt_rsc_0_15_radr),
      .we(yt_rsc_0_15_we),
      .d(yt_rsc_0_15_d),
      .wadr(yt_rsc_0_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_0_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_0_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_23_4_32_16_16_32_1_gen yt_rsc_0_16_i
      (
      .clkr_en(yt_rsc_0_16_clkr_en),
      .clkw_en(yt_rsc_0_16_clkw_en),
      .q(yt_rsc_0_16_q),
      .radr(yt_rsc_0_16_radr),
      .we(yt_rsc_0_16_we),
      .d(yt_rsc_0_16_d),
      .wadr(yt_rsc_0_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_0_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_24_4_32_16_16_32_1_gen yt_rsc_0_17_i
      (
      .clkr_en(yt_rsc_0_17_clkr_en),
      .clkw_en(yt_rsc_0_17_clkw_en),
      .q(yt_rsc_0_17_q),
      .radr(yt_rsc_0_17_radr),
      .we(yt_rsc_0_17_we),
      .d(yt_rsc_0_17_d),
      .wadr(yt_rsc_0_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_0_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_25_4_32_16_16_32_1_gen yt_rsc_0_18_i
      (
      .clkr_en(yt_rsc_0_18_clkr_en),
      .clkw_en(yt_rsc_0_18_clkw_en),
      .q(yt_rsc_0_18_q),
      .radr(yt_rsc_0_18_radr),
      .we(yt_rsc_0_18_we),
      .d(yt_rsc_0_18_d),
      .wadr(yt_rsc_0_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_0_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_26_4_32_16_16_32_1_gen yt_rsc_0_19_i
      (
      .clkr_en(yt_rsc_0_19_clkr_en),
      .clkw_en(yt_rsc_0_19_clkw_en),
      .q(yt_rsc_0_19_q),
      .radr(yt_rsc_0_19_radr),
      .we(yt_rsc_0_19_we),
      .d(yt_rsc_0_19_d),
      .wadr(yt_rsc_0_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_0_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_27_4_32_16_16_32_1_gen yt_rsc_0_20_i
      (
      .clkr_en(yt_rsc_0_20_clkr_en),
      .clkw_en(yt_rsc_0_20_clkw_en),
      .q(yt_rsc_0_20_q),
      .radr(yt_rsc_0_20_radr),
      .we(yt_rsc_0_20_we),
      .d(yt_rsc_0_20_d),
      .wadr(yt_rsc_0_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_0_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_28_4_32_16_16_32_1_gen yt_rsc_0_21_i
      (
      .clkr_en(yt_rsc_0_21_clkr_en),
      .clkw_en(yt_rsc_0_21_clkw_en),
      .q(yt_rsc_0_21_q),
      .radr(yt_rsc_0_21_radr),
      .we(yt_rsc_0_21_we),
      .d(yt_rsc_0_21_d),
      .wadr(yt_rsc_0_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_0_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_29_4_32_16_16_32_1_gen yt_rsc_0_22_i
      (
      .clkr_en(yt_rsc_0_22_clkr_en),
      .clkw_en(yt_rsc_0_22_clkw_en),
      .q(yt_rsc_0_22_q),
      .radr(yt_rsc_0_22_radr),
      .we(yt_rsc_0_22_we),
      .d(yt_rsc_0_22_d),
      .wadr(yt_rsc_0_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_0_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_30_4_32_16_16_32_1_gen yt_rsc_0_23_i
      (
      .clkr_en(yt_rsc_0_23_clkr_en),
      .clkw_en(yt_rsc_0_23_clkw_en),
      .q(yt_rsc_0_23_q),
      .radr(yt_rsc_0_23_radr),
      .we(yt_rsc_0_23_we),
      .d(yt_rsc_0_23_d),
      .wadr(yt_rsc_0_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_0_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_31_4_32_16_16_32_1_gen yt_rsc_0_24_i
      (
      .clkr_en(yt_rsc_0_24_clkr_en),
      .clkw_en(yt_rsc_0_24_clkw_en),
      .q(yt_rsc_0_24_q),
      .radr(yt_rsc_0_24_radr),
      .we(yt_rsc_0_24_we),
      .d(yt_rsc_0_24_d),
      .wadr(yt_rsc_0_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_0_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_32_4_32_16_16_32_1_gen yt_rsc_0_25_i
      (
      .clkr_en(yt_rsc_0_25_clkr_en),
      .clkw_en(yt_rsc_0_25_clkw_en),
      .q(yt_rsc_0_25_q),
      .radr(yt_rsc_0_25_radr),
      .we(yt_rsc_0_25_we),
      .d(yt_rsc_0_25_d),
      .wadr(yt_rsc_0_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_0_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_33_4_32_16_16_32_1_gen yt_rsc_0_26_i
      (
      .clkr_en(yt_rsc_0_26_clkr_en),
      .clkw_en(yt_rsc_0_26_clkw_en),
      .q(yt_rsc_0_26_q),
      .radr(yt_rsc_0_26_radr),
      .we(yt_rsc_0_26_we),
      .d(yt_rsc_0_26_d),
      .wadr(yt_rsc_0_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_0_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_34_4_32_16_16_32_1_gen yt_rsc_0_27_i
      (
      .clkr_en(yt_rsc_0_27_clkr_en),
      .clkw_en(yt_rsc_0_27_clkw_en),
      .q(yt_rsc_0_27_q),
      .radr(yt_rsc_0_27_radr),
      .we(yt_rsc_0_27_we),
      .d(yt_rsc_0_27_d),
      .wadr(yt_rsc_0_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_0_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_35_4_32_16_16_32_1_gen yt_rsc_0_28_i
      (
      .clkr_en(yt_rsc_0_28_clkr_en),
      .clkw_en(yt_rsc_0_28_clkw_en),
      .q(yt_rsc_0_28_q),
      .radr(yt_rsc_0_28_radr),
      .we(yt_rsc_0_28_we),
      .d(yt_rsc_0_28_d),
      .wadr(yt_rsc_0_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_0_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_36_4_32_16_16_32_1_gen yt_rsc_0_29_i
      (
      .clkr_en(yt_rsc_0_29_clkr_en),
      .clkw_en(yt_rsc_0_29_clkw_en),
      .q(yt_rsc_0_29_q),
      .radr(yt_rsc_0_29_radr),
      .we(yt_rsc_0_29_we),
      .d(yt_rsc_0_29_d),
      .wadr(yt_rsc_0_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_0_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_37_4_32_16_16_32_1_gen yt_rsc_0_30_i
      (
      .clkr_en(yt_rsc_0_30_clkr_en),
      .clkw_en(yt_rsc_0_30_clkw_en),
      .q(yt_rsc_0_30_q),
      .radr(yt_rsc_0_30_radr),
      .we(yt_rsc_0_30_we),
      .d(yt_rsc_0_30_d),
      .wadr(yt_rsc_0_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_0_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_38_4_32_16_16_32_1_gen yt_rsc_0_31_i
      (
      .clkr_en(yt_rsc_0_31_clkr_en),
      .clkw_en(yt_rsc_0_31_clkw_en),
      .q(yt_rsc_0_31_q),
      .radr(yt_rsc_0_31_radr),
      .we(yt_rsc_0_31_we),
      .d(yt_rsc_0_31_d),
      .wadr(yt_rsc_0_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_0_16_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_0_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_39_4_32_16_16_32_1_gen yt_rsc_1_0_i
      (
      .clkr_en(yt_rsc_1_0_clkr_en),
      .clkw_en(yt_rsc_1_0_clkw_en),
      .q(yt_rsc_1_0_q),
      .radr(yt_rsc_1_0_radr),
      .we(yt_rsc_1_0_we),
      .d(yt_rsc_1_0_d),
      .wadr(yt_rsc_1_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_1_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_40_4_32_16_16_32_1_gen yt_rsc_1_1_i
      (
      .clkr_en(yt_rsc_1_1_clkr_en),
      .clkw_en(yt_rsc_1_1_clkw_en),
      .q(yt_rsc_1_1_q),
      .radr(yt_rsc_1_1_radr),
      .we(yt_rsc_1_1_we),
      .d(yt_rsc_1_1_d),
      .wadr(yt_rsc_1_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_1_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_41_4_32_16_16_32_1_gen yt_rsc_1_2_i
      (
      .clkr_en(yt_rsc_1_2_clkr_en),
      .clkw_en(yt_rsc_1_2_clkw_en),
      .q(yt_rsc_1_2_q),
      .radr(yt_rsc_1_2_radr),
      .we(yt_rsc_1_2_we),
      .d(yt_rsc_1_2_d),
      .wadr(yt_rsc_1_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_1_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_42_4_32_16_16_32_1_gen yt_rsc_1_3_i
      (
      .clkr_en(yt_rsc_1_3_clkr_en),
      .clkw_en(yt_rsc_1_3_clkw_en),
      .q(yt_rsc_1_3_q),
      .radr(yt_rsc_1_3_radr),
      .we(yt_rsc_1_3_we),
      .d(yt_rsc_1_3_d),
      .wadr(yt_rsc_1_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_1_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_43_4_32_16_16_32_1_gen yt_rsc_1_4_i
      (
      .clkr_en(yt_rsc_1_4_clkr_en),
      .clkw_en(yt_rsc_1_4_clkw_en),
      .q(yt_rsc_1_4_q),
      .radr(yt_rsc_1_4_radr),
      .we(yt_rsc_1_4_we),
      .d(yt_rsc_1_4_d),
      .wadr(yt_rsc_1_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_1_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_44_4_32_16_16_32_1_gen yt_rsc_1_5_i
      (
      .clkr_en(yt_rsc_1_5_clkr_en),
      .clkw_en(yt_rsc_1_5_clkw_en),
      .q(yt_rsc_1_5_q),
      .radr(yt_rsc_1_5_radr),
      .we(yt_rsc_1_5_we),
      .d(yt_rsc_1_5_d),
      .wadr(yt_rsc_1_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_1_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_45_4_32_16_16_32_1_gen yt_rsc_1_6_i
      (
      .clkr_en(yt_rsc_1_6_clkr_en),
      .clkw_en(yt_rsc_1_6_clkw_en),
      .q(yt_rsc_1_6_q),
      .radr(yt_rsc_1_6_radr),
      .we(yt_rsc_1_6_we),
      .d(yt_rsc_1_6_d),
      .wadr(yt_rsc_1_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_1_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_46_4_32_16_16_32_1_gen yt_rsc_1_7_i
      (
      .clkr_en(yt_rsc_1_7_clkr_en),
      .clkw_en(yt_rsc_1_7_clkw_en),
      .q(yt_rsc_1_7_q),
      .radr(yt_rsc_1_7_radr),
      .we(yt_rsc_1_7_we),
      .d(yt_rsc_1_7_d),
      .wadr(yt_rsc_1_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_1_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_47_4_32_16_16_32_1_gen yt_rsc_1_8_i
      (
      .clkr_en(yt_rsc_1_8_clkr_en),
      .clkw_en(yt_rsc_1_8_clkw_en),
      .q(yt_rsc_1_8_q),
      .radr(yt_rsc_1_8_radr),
      .we(yt_rsc_1_8_we),
      .d(yt_rsc_1_8_d),
      .wadr(yt_rsc_1_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_1_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_48_4_32_16_16_32_1_gen yt_rsc_1_9_i
      (
      .clkr_en(yt_rsc_1_9_clkr_en),
      .clkw_en(yt_rsc_1_9_clkw_en),
      .q(yt_rsc_1_9_q),
      .radr(yt_rsc_1_9_radr),
      .we(yt_rsc_1_9_we),
      .d(yt_rsc_1_9_d),
      .wadr(yt_rsc_1_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_1_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_49_4_32_16_16_32_1_gen yt_rsc_1_10_i
      (
      .clkr_en(yt_rsc_1_10_clkr_en),
      .clkw_en(yt_rsc_1_10_clkw_en),
      .q(yt_rsc_1_10_q),
      .radr(yt_rsc_1_10_radr),
      .we(yt_rsc_1_10_we),
      .d(yt_rsc_1_10_d),
      .wadr(yt_rsc_1_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_1_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_50_4_32_16_16_32_1_gen yt_rsc_1_11_i
      (
      .clkr_en(yt_rsc_1_11_clkr_en),
      .clkw_en(yt_rsc_1_11_clkw_en),
      .q(yt_rsc_1_11_q),
      .radr(yt_rsc_1_11_radr),
      .we(yt_rsc_1_11_we),
      .d(yt_rsc_1_11_d),
      .wadr(yt_rsc_1_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_1_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_51_4_32_16_16_32_1_gen yt_rsc_1_12_i
      (
      .clkr_en(yt_rsc_1_12_clkr_en),
      .clkw_en(yt_rsc_1_12_clkw_en),
      .q(yt_rsc_1_12_q),
      .radr(yt_rsc_1_12_radr),
      .we(yt_rsc_1_12_we),
      .d(yt_rsc_1_12_d),
      .wadr(yt_rsc_1_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_1_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_52_4_32_16_16_32_1_gen yt_rsc_1_13_i
      (
      .clkr_en(yt_rsc_1_13_clkr_en),
      .clkw_en(yt_rsc_1_13_clkw_en),
      .q(yt_rsc_1_13_q),
      .radr(yt_rsc_1_13_radr),
      .we(yt_rsc_1_13_we),
      .d(yt_rsc_1_13_d),
      .wadr(yt_rsc_1_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_1_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_53_4_32_16_16_32_1_gen yt_rsc_1_14_i
      (
      .clkr_en(yt_rsc_1_14_clkr_en),
      .clkw_en(yt_rsc_1_14_clkw_en),
      .q(yt_rsc_1_14_q),
      .radr(yt_rsc_1_14_radr),
      .we(yt_rsc_1_14_we),
      .d(yt_rsc_1_14_d),
      .wadr(yt_rsc_1_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_1_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_54_4_32_16_16_32_1_gen yt_rsc_1_15_i
      (
      .clkr_en(yt_rsc_1_15_clkr_en),
      .clkw_en(yt_rsc_1_15_clkw_en),
      .q(yt_rsc_1_15_q),
      .radr(yt_rsc_1_15_radr),
      .we(yt_rsc_1_15_we),
      .d(yt_rsc_1_15_d),
      .wadr(yt_rsc_1_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_0_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_1_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_1_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_55_4_32_16_16_32_1_gen yt_rsc_1_16_i
      (
      .clkr_en(yt_rsc_1_16_clkr_en),
      .clkw_en(yt_rsc_1_16_clkw_en),
      .q(yt_rsc_1_16_q),
      .radr(yt_rsc_1_16_radr),
      .we(yt_rsc_1_16_we),
      .d(yt_rsc_1_16_d),
      .wadr(yt_rsc_1_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_1_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_56_4_32_16_16_32_1_gen yt_rsc_1_17_i
      (
      .clkr_en(yt_rsc_1_17_clkr_en),
      .clkw_en(yt_rsc_1_17_clkw_en),
      .q(yt_rsc_1_17_q),
      .radr(yt_rsc_1_17_radr),
      .we(yt_rsc_1_17_we),
      .d(yt_rsc_1_17_d),
      .wadr(yt_rsc_1_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_1_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_57_4_32_16_16_32_1_gen yt_rsc_1_18_i
      (
      .clkr_en(yt_rsc_1_18_clkr_en),
      .clkw_en(yt_rsc_1_18_clkw_en),
      .q(yt_rsc_1_18_q),
      .radr(yt_rsc_1_18_radr),
      .we(yt_rsc_1_18_we),
      .d(yt_rsc_1_18_d),
      .wadr(yt_rsc_1_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_1_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_58_4_32_16_16_32_1_gen yt_rsc_1_19_i
      (
      .clkr_en(yt_rsc_1_19_clkr_en),
      .clkw_en(yt_rsc_1_19_clkw_en),
      .q(yt_rsc_1_19_q),
      .radr(yt_rsc_1_19_radr),
      .we(yt_rsc_1_19_we),
      .d(yt_rsc_1_19_d),
      .wadr(yt_rsc_1_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_1_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_59_4_32_16_16_32_1_gen yt_rsc_1_20_i
      (
      .clkr_en(yt_rsc_1_20_clkr_en),
      .clkw_en(yt_rsc_1_20_clkw_en),
      .q(yt_rsc_1_20_q),
      .radr(yt_rsc_1_20_radr),
      .we(yt_rsc_1_20_we),
      .d(yt_rsc_1_20_d),
      .wadr(yt_rsc_1_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_1_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_60_4_32_16_16_32_1_gen yt_rsc_1_21_i
      (
      .clkr_en(yt_rsc_1_21_clkr_en),
      .clkw_en(yt_rsc_1_21_clkw_en),
      .q(yt_rsc_1_21_q),
      .radr(yt_rsc_1_21_radr),
      .we(yt_rsc_1_21_we),
      .d(yt_rsc_1_21_d),
      .wadr(yt_rsc_1_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_1_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_61_4_32_16_16_32_1_gen yt_rsc_1_22_i
      (
      .clkr_en(yt_rsc_1_22_clkr_en),
      .clkw_en(yt_rsc_1_22_clkw_en),
      .q(yt_rsc_1_22_q),
      .radr(yt_rsc_1_22_radr),
      .we(yt_rsc_1_22_we),
      .d(yt_rsc_1_22_d),
      .wadr(yt_rsc_1_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_1_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_62_4_32_16_16_32_1_gen yt_rsc_1_23_i
      (
      .clkr_en(yt_rsc_1_23_clkr_en),
      .clkw_en(yt_rsc_1_23_clkw_en),
      .q(yt_rsc_1_23_q),
      .radr(yt_rsc_1_23_radr),
      .we(yt_rsc_1_23_we),
      .d(yt_rsc_1_23_d),
      .wadr(yt_rsc_1_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_1_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_63_4_32_16_16_32_1_gen yt_rsc_1_24_i
      (
      .clkr_en(yt_rsc_1_24_clkr_en),
      .clkw_en(yt_rsc_1_24_clkw_en),
      .q(yt_rsc_1_24_q),
      .radr(yt_rsc_1_24_radr),
      .we(yt_rsc_1_24_we),
      .d(yt_rsc_1_24_d),
      .wadr(yt_rsc_1_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_1_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_64_4_32_16_16_32_1_gen yt_rsc_1_25_i
      (
      .clkr_en(yt_rsc_1_25_clkr_en),
      .clkw_en(yt_rsc_1_25_clkw_en),
      .q(yt_rsc_1_25_q),
      .radr(yt_rsc_1_25_radr),
      .we(yt_rsc_1_25_we),
      .d(yt_rsc_1_25_d),
      .wadr(yt_rsc_1_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_1_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_65_4_32_16_16_32_1_gen yt_rsc_1_26_i
      (
      .clkr_en(yt_rsc_1_26_clkr_en),
      .clkw_en(yt_rsc_1_26_clkw_en),
      .q(yt_rsc_1_26_q),
      .radr(yt_rsc_1_26_radr),
      .we(yt_rsc_1_26_we),
      .d(yt_rsc_1_26_d),
      .wadr(yt_rsc_1_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_1_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_66_4_32_16_16_32_1_gen yt_rsc_1_27_i
      (
      .clkr_en(yt_rsc_1_27_clkr_en),
      .clkw_en(yt_rsc_1_27_clkw_en),
      .q(yt_rsc_1_27_q),
      .radr(yt_rsc_1_27_radr),
      .we(yt_rsc_1_27_we),
      .d(yt_rsc_1_27_d),
      .wadr(yt_rsc_1_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_1_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_67_4_32_16_16_32_1_gen yt_rsc_1_28_i
      (
      .clkr_en(yt_rsc_1_28_clkr_en),
      .clkw_en(yt_rsc_1_28_clkw_en),
      .q(yt_rsc_1_28_q),
      .radr(yt_rsc_1_28_radr),
      .we(yt_rsc_1_28_we),
      .d(yt_rsc_1_28_d),
      .wadr(yt_rsc_1_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_1_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_68_4_32_16_16_32_1_gen yt_rsc_1_29_i
      (
      .clkr_en(yt_rsc_1_29_clkr_en),
      .clkw_en(yt_rsc_1_29_clkw_en),
      .q(yt_rsc_1_29_q),
      .radr(yt_rsc_1_29_radr),
      .we(yt_rsc_1_29_we),
      .d(yt_rsc_1_29_d),
      .wadr(yt_rsc_1_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_1_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_69_4_32_16_16_32_1_gen yt_rsc_1_30_i
      (
      .clkr_en(yt_rsc_1_30_clkr_en),
      .clkw_en(yt_rsc_1_30_clkw_en),
      .q(yt_rsc_1_30_q),
      .radr(yt_rsc_1_30_radr),
      .we(yt_rsc_1_30_we),
      .d(yt_rsc_1_30_d),
      .wadr(yt_rsc_1_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_1_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_70_4_32_16_16_32_1_gen yt_rsc_1_31_i
      (
      .clkr_en(yt_rsc_1_31_clkr_en),
      .clkw_en(yt_rsc_1_31_clkw_en),
      .q(yt_rsc_1_31_q),
      .radr(yt_rsc_1_31_radr),
      .we(yt_rsc_1_31_we),
      .d(yt_rsc_1_31_d),
      .wadr(yt_rsc_1_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_1_16_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_1_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_1_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_1_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_71_4_32_16_16_32_1_gen yt_rsc_2_0_i
      (
      .clkr_en(yt_rsc_2_0_clkr_en),
      .clkw_en(yt_rsc_2_0_clkw_en),
      .q(yt_rsc_2_0_q),
      .radr(yt_rsc_2_0_radr),
      .we(yt_rsc_2_0_we),
      .d(yt_rsc_2_0_d),
      .wadr(yt_rsc_2_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_2_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_72_4_32_16_16_32_1_gen yt_rsc_2_1_i
      (
      .clkr_en(yt_rsc_2_1_clkr_en),
      .clkw_en(yt_rsc_2_1_clkw_en),
      .q(yt_rsc_2_1_q),
      .radr(yt_rsc_2_1_radr),
      .we(yt_rsc_2_1_we),
      .d(yt_rsc_2_1_d),
      .wadr(yt_rsc_2_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_2_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_73_4_32_16_16_32_1_gen yt_rsc_2_2_i
      (
      .clkr_en(yt_rsc_2_2_clkr_en),
      .clkw_en(yt_rsc_2_2_clkw_en),
      .q(yt_rsc_2_2_q),
      .radr(yt_rsc_2_2_radr),
      .we(yt_rsc_2_2_we),
      .d(yt_rsc_2_2_d),
      .wadr(yt_rsc_2_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_2_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_74_4_32_16_16_32_1_gen yt_rsc_2_3_i
      (
      .clkr_en(yt_rsc_2_3_clkr_en),
      .clkw_en(yt_rsc_2_3_clkw_en),
      .q(yt_rsc_2_3_q),
      .radr(yt_rsc_2_3_radr),
      .we(yt_rsc_2_3_we),
      .d(yt_rsc_2_3_d),
      .wadr(yt_rsc_2_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_2_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_75_4_32_16_16_32_1_gen yt_rsc_2_4_i
      (
      .clkr_en(yt_rsc_2_4_clkr_en),
      .clkw_en(yt_rsc_2_4_clkw_en),
      .q(yt_rsc_2_4_q),
      .radr(yt_rsc_2_4_radr),
      .we(yt_rsc_2_4_we),
      .d(yt_rsc_2_4_d),
      .wadr(yt_rsc_2_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_2_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_76_4_32_16_16_32_1_gen yt_rsc_2_5_i
      (
      .clkr_en(yt_rsc_2_5_clkr_en),
      .clkw_en(yt_rsc_2_5_clkw_en),
      .q(yt_rsc_2_5_q),
      .radr(yt_rsc_2_5_radr),
      .we(yt_rsc_2_5_we),
      .d(yt_rsc_2_5_d),
      .wadr(yt_rsc_2_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_2_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_77_4_32_16_16_32_1_gen yt_rsc_2_6_i
      (
      .clkr_en(yt_rsc_2_6_clkr_en),
      .clkw_en(yt_rsc_2_6_clkw_en),
      .q(yt_rsc_2_6_q),
      .radr(yt_rsc_2_6_radr),
      .we(yt_rsc_2_6_we),
      .d(yt_rsc_2_6_d),
      .wadr(yt_rsc_2_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_2_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_78_4_32_16_16_32_1_gen yt_rsc_2_7_i
      (
      .clkr_en(yt_rsc_2_7_clkr_en),
      .clkw_en(yt_rsc_2_7_clkw_en),
      .q(yt_rsc_2_7_q),
      .radr(yt_rsc_2_7_radr),
      .we(yt_rsc_2_7_we),
      .d(yt_rsc_2_7_d),
      .wadr(yt_rsc_2_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_2_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_79_4_32_16_16_32_1_gen yt_rsc_2_8_i
      (
      .clkr_en(yt_rsc_2_8_clkr_en),
      .clkw_en(yt_rsc_2_8_clkw_en),
      .q(yt_rsc_2_8_q),
      .radr(yt_rsc_2_8_radr),
      .we(yt_rsc_2_8_we),
      .d(yt_rsc_2_8_d),
      .wadr(yt_rsc_2_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_2_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_80_4_32_16_16_32_1_gen yt_rsc_2_9_i
      (
      .clkr_en(yt_rsc_2_9_clkr_en),
      .clkw_en(yt_rsc_2_9_clkw_en),
      .q(yt_rsc_2_9_q),
      .radr(yt_rsc_2_9_radr),
      .we(yt_rsc_2_9_we),
      .d(yt_rsc_2_9_d),
      .wadr(yt_rsc_2_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_2_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_81_4_32_16_16_32_1_gen yt_rsc_2_10_i
      (
      .clkr_en(yt_rsc_2_10_clkr_en),
      .clkw_en(yt_rsc_2_10_clkw_en),
      .q(yt_rsc_2_10_q),
      .radr(yt_rsc_2_10_radr),
      .we(yt_rsc_2_10_we),
      .d(yt_rsc_2_10_d),
      .wadr(yt_rsc_2_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_2_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_82_4_32_16_16_32_1_gen yt_rsc_2_11_i
      (
      .clkr_en(yt_rsc_2_11_clkr_en),
      .clkw_en(yt_rsc_2_11_clkw_en),
      .q(yt_rsc_2_11_q),
      .radr(yt_rsc_2_11_radr),
      .we(yt_rsc_2_11_we),
      .d(yt_rsc_2_11_d),
      .wadr(yt_rsc_2_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_2_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_83_4_32_16_16_32_1_gen yt_rsc_2_12_i
      (
      .clkr_en(yt_rsc_2_12_clkr_en),
      .clkw_en(yt_rsc_2_12_clkw_en),
      .q(yt_rsc_2_12_q),
      .radr(yt_rsc_2_12_radr),
      .we(yt_rsc_2_12_we),
      .d(yt_rsc_2_12_d),
      .wadr(yt_rsc_2_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_2_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_84_4_32_16_16_32_1_gen yt_rsc_2_13_i
      (
      .clkr_en(yt_rsc_2_13_clkr_en),
      .clkw_en(yt_rsc_2_13_clkw_en),
      .q(yt_rsc_2_13_q),
      .radr(yt_rsc_2_13_radr),
      .we(yt_rsc_2_13_we),
      .d(yt_rsc_2_13_d),
      .wadr(yt_rsc_2_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_2_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_85_4_32_16_16_32_1_gen yt_rsc_2_14_i
      (
      .clkr_en(yt_rsc_2_14_clkr_en),
      .clkw_en(yt_rsc_2_14_clkw_en),
      .q(yt_rsc_2_14_q),
      .radr(yt_rsc_2_14_radr),
      .we(yt_rsc_2_14_we),
      .d(yt_rsc_2_14_d),
      .wadr(yt_rsc_2_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_2_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_86_4_32_16_16_32_1_gen yt_rsc_2_15_i
      (
      .clkr_en(yt_rsc_2_15_clkr_en),
      .clkw_en(yt_rsc_2_15_clkw_en),
      .q(yt_rsc_2_15_q),
      .radr(yt_rsc_2_15_radr),
      .we(yt_rsc_2_15_we),
      .d(yt_rsc_2_15_d),
      .wadr(yt_rsc_2_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_0_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_2_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_2_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_87_4_32_16_16_32_1_gen yt_rsc_2_16_i
      (
      .clkr_en(yt_rsc_2_16_clkr_en),
      .clkw_en(yt_rsc_2_16_clkw_en),
      .q(yt_rsc_2_16_q),
      .radr(yt_rsc_2_16_radr),
      .we(yt_rsc_2_16_we),
      .d(yt_rsc_2_16_d),
      .wadr(yt_rsc_2_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_2_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_88_4_32_16_16_32_1_gen yt_rsc_2_17_i
      (
      .clkr_en(yt_rsc_2_17_clkr_en),
      .clkw_en(yt_rsc_2_17_clkw_en),
      .q(yt_rsc_2_17_q),
      .radr(yt_rsc_2_17_radr),
      .we(yt_rsc_2_17_we),
      .d(yt_rsc_2_17_d),
      .wadr(yt_rsc_2_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_2_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_89_4_32_16_16_32_1_gen yt_rsc_2_18_i
      (
      .clkr_en(yt_rsc_2_18_clkr_en),
      .clkw_en(yt_rsc_2_18_clkw_en),
      .q(yt_rsc_2_18_q),
      .radr(yt_rsc_2_18_radr),
      .we(yt_rsc_2_18_we),
      .d(yt_rsc_2_18_d),
      .wadr(yt_rsc_2_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_2_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_90_4_32_16_16_32_1_gen yt_rsc_2_19_i
      (
      .clkr_en(yt_rsc_2_19_clkr_en),
      .clkw_en(yt_rsc_2_19_clkw_en),
      .q(yt_rsc_2_19_q),
      .radr(yt_rsc_2_19_radr),
      .we(yt_rsc_2_19_we),
      .d(yt_rsc_2_19_d),
      .wadr(yt_rsc_2_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_2_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_91_4_32_16_16_32_1_gen yt_rsc_2_20_i
      (
      .clkr_en(yt_rsc_2_20_clkr_en),
      .clkw_en(yt_rsc_2_20_clkw_en),
      .q(yt_rsc_2_20_q),
      .radr(yt_rsc_2_20_radr),
      .we(yt_rsc_2_20_we),
      .d(yt_rsc_2_20_d),
      .wadr(yt_rsc_2_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_2_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_92_4_32_16_16_32_1_gen yt_rsc_2_21_i
      (
      .clkr_en(yt_rsc_2_21_clkr_en),
      .clkw_en(yt_rsc_2_21_clkw_en),
      .q(yt_rsc_2_21_q),
      .radr(yt_rsc_2_21_radr),
      .we(yt_rsc_2_21_we),
      .d(yt_rsc_2_21_d),
      .wadr(yt_rsc_2_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_2_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_93_4_32_16_16_32_1_gen yt_rsc_2_22_i
      (
      .clkr_en(yt_rsc_2_22_clkr_en),
      .clkw_en(yt_rsc_2_22_clkw_en),
      .q(yt_rsc_2_22_q),
      .radr(yt_rsc_2_22_radr),
      .we(yt_rsc_2_22_we),
      .d(yt_rsc_2_22_d),
      .wadr(yt_rsc_2_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_2_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_94_4_32_16_16_32_1_gen yt_rsc_2_23_i
      (
      .clkr_en(yt_rsc_2_23_clkr_en),
      .clkw_en(yt_rsc_2_23_clkw_en),
      .q(yt_rsc_2_23_q),
      .radr(yt_rsc_2_23_radr),
      .we(yt_rsc_2_23_we),
      .d(yt_rsc_2_23_d),
      .wadr(yt_rsc_2_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_2_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_95_4_32_16_16_32_1_gen yt_rsc_2_24_i
      (
      .clkr_en(yt_rsc_2_24_clkr_en),
      .clkw_en(yt_rsc_2_24_clkw_en),
      .q(yt_rsc_2_24_q),
      .radr(yt_rsc_2_24_radr),
      .we(yt_rsc_2_24_we),
      .d(yt_rsc_2_24_d),
      .wadr(yt_rsc_2_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_2_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_96_4_32_16_16_32_1_gen yt_rsc_2_25_i
      (
      .clkr_en(yt_rsc_2_25_clkr_en),
      .clkw_en(yt_rsc_2_25_clkw_en),
      .q(yt_rsc_2_25_q),
      .radr(yt_rsc_2_25_radr),
      .we(yt_rsc_2_25_we),
      .d(yt_rsc_2_25_d),
      .wadr(yt_rsc_2_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_2_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_97_4_32_16_16_32_1_gen yt_rsc_2_26_i
      (
      .clkr_en(yt_rsc_2_26_clkr_en),
      .clkw_en(yt_rsc_2_26_clkw_en),
      .q(yt_rsc_2_26_q),
      .radr(yt_rsc_2_26_radr),
      .we(yt_rsc_2_26_we),
      .d(yt_rsc_2_26_d),
      .wadr(yt_rsc_2_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_2_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_98_4_32_16_16_32_1_gen yt_rsc_2_27_i
      (
      .clkr_en(yt_rsc_2_27_clkr_en),
      .clkw_en(yt_rsc_2_27_clkw_en),
      .q(yt_rsc_2_27_q),
      .radr(yt_rsc_2_27_radr),
      .we(yt_rsc_2_27_we),
      .d(yt_rsc_2_27_d),
      .wadr(yt_rsc_2_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_2_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_99_4_32_16_16_32_1_gen yt_rsc_2_28_i
      (
      .clkr_en(yt_rsc_2_28_clkr_en),
      .clkw_en(yt_rsc_2_28_clkw_en),
      .q(yt_rsc_2_28_q),
      .radr(yt_rsc_2_28_radr),
      .we(yt_rsc_2_28_we),
      .d(yt_rsc_2_28_d),
      .wadr(yt_rsc_2_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_2_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_100_4_32_16_16_32_1_gen yt_rsc_2_29_i
      (
      .clkr_en(yt_rsc_2_29_clkr_en),
      .clkw_en(yt_rsc_2_29_clkw_en),
      .q(yt_rsc_2_29_q),
      .radr(yt_rsc_2_29_radr),
      .we(yt_rsc_2_29_we),
      .d(yt_rsc_2_29_d),
      .wadr(yt_rsc_2_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_2_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_101_4_32_16_16_32_1_gen yt_rsc_2_30_i
      (
      .clkr_en(yt_rsc_2_30_clkr_en),
      .clkw_en(yt_rsc_2_30_clkw_en),
      .q(yt_rsc_2_30_q),
      .radr(yt_rsc_2_30_radr),
      .we(yt_rsc_2_30_we),
      .d(yt_rsc_2_30_d),
      .wadr(yt_rsc_2_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_2_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_102_4_32_16_16_32_1_gen yt_rsc_2_31_i
      (
      .clkr_en(yt_rsc_2_31_clkr_en),
      .clkw_en(yt_rsc_2_31_clkw_en),
      .q(yt_rsc_2_31_q),
      .radr(yt_rsc_2_31_radr),
      .we(yt_rsc_2_31_we),
      .d(yt_rsc_2_31_d),
      .wadr(yt_rsc_2_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_2_16_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_2_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_2_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_2_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_103_4_32_16_16_32_1_gen yt_rsc_3_0_i
      (
      .clkr_en(yt_rsc_3_0_clkr_en),
      .clkw_en(yt_rsc_3_0_clkw_en),
      .q(yt_rsc_3_0_q),
      .radr(yt_rsc_3_0_radr),
      .we(yt_rsc_3_0_we),
      .d(yt_rsc_3_0_d),
      .wadr(yt_rsc_3_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_3_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_104_4_32_16_16_32_1_gen yt_rsc_3_1_i
      (
      .clkr_en(yt_rsc_3_1_clkr_en),
      .clkw_en(yt_rsc_3_1_clkw_en),
      .q(yt_rsc_3_1_q),
      .radr(yt_rsc_3_1_radr),
      .we(yt_rsc_3_1_we),
      .d(yt_rsc_3_1_d),
      .wadr(yt_rsc_3_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_3_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_105_4_32_16_16_32_1_gen yt_rsc_3_2_i
      (
      .clkr_en(yt_rsc_3_2_clkr_en),
      .clkw_en(yt_rsc_3_2_clkw_en),
      .q(yt_rsc_3_2_q),
      .radr(yt_rsc_3_2_radr),
      .we(yt_rsc_3_2_we),
      .d(yt_rsc_3_2_d),
      .wadr(yt_rsc_3_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_3_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_106_4_32_16_16_32_1_gen yt_rsc_3_3_i
      (
      .clkr_en(yt_rsc_3_3_clkr_en),
      .clkw_en(yt_rsc_3_3_clkw_en),
      .q(yt_rsc_3_3_q),
      .radr(yt_rsc_3_3_radr),
      .we(yt_rsc_3_3_we),
      .d(yt_rsc_3_3_d),
      .wadr(yt_rsc_3_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_3_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_107_4_32_16_16_32_1_gen yt_rsc_3_4_i
      (
      .clkr_en(yt_rsc_3_4_clkr_en),
      .clkw_en(yt_rsc_3_4_clkw_en),
      .q(yt_rsc_3_4_q),
      .radr(yt_rsc_3_4_radr),
      .we(yt_rsc_3_4_we),
      .d(yt_rsc_3_4_d),
      .wadr(yt_rsc_3_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_3_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_108_4_32_16_16_32_1_gen yt_rsc_3_5_i
      (
      .clkr_en(yt_rsc_3_5_clkr_en),
      .clkw_en(yt_rsc_3_5_clkw_en),
      .q(yt_rsc_3_5_q),
      .radr(yt_rsc_3_5_radr),
      .we(yt_rsc_3_5_we),
      .d(yt_rsc_3_5_d),
      .wadr(yt_rsc_3_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_3_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_109_4_32_16_16_32_1_gen yt_rsc_3_6_i
      (
      .clkr_en(yt_rsc_3_6_clkr_en),
      .clkw_en(yt_rsc_3_6_clkw_en),
      .q(yt_rsc_3_6_q),
      .radr(yt_rsc_3_6_radr),
      .we(yt_rsc_3_6_we),
      .d(yt_rsc_3_6_d),
      .wadr(yt_rsc_3_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_3_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_110_4_32_16_16_32_1_gen yt_rsc_3_7_i
      (
      .clkr_en(yt_rsc_3_7_clkr_en),
      .clkw_en(yt_rsc_3_7_clkw_en),
      .q(yt_rsc_3_7_q),
      .radr(yt_rsc_3_7_radr),
      .we(yt_rsc_3_7_we),
      .d(yt_rsc_3_7_d),
      .wadr(yt_rsc_3_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_3_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_111_4_32_16_16_32_1_gen yt_rsc_3_8_i
      (
      .clkr_en(yt_rsc_3_8_clkr_en),
      .clkw_en(yt_rsc_3_8_clkw_en),
      .q(yt_rsc_3_8_q),
      .radr(yt_rsc_3_8_radr),
      .we(yt_rsc_3_8_we),
      .d(yt_rsc_3_8_d),
      .wadr(yt_rsc_3_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_3_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_112_4_32_16_16_32_1_gen yt_rsc_3_9_i
      (
      .clkr_en(yt_rsc_3_9_clkr_en),
      .clkw_en(yt_rsc_3_9_clkw_en),
      .q(yt_rsc_3_9_q),
      .radr(yt_rsc_3_9_radr),
      .we(yt_rsc_3_9_we),
      .d(yt_rsc_3_9_d),
      .wadr(yt_rsc_3_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_3_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_113_4_32_16_16_32_1_gen yt_rsc_3_10_i
      (
      .clkr_en(yt_rsc_3_10_clkr_en),
      .clkw_en(yt_rsc_3_10_clkw_en),
      .q(yt_rsc_3_10_q),
      .radr(yt_rsc_3_10_radr),
      .we(yt_rsc_3_10_we),
      .d(yt_rsc_3_10_d),
      .wadr(yt_rsc_3_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_3_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_114_4_32_16_16_32_1_gen yt_rsc_3_11_i
      (
      .clkr_en(yt_rsc_3_11_clkr_en),
      .clkw_en(yt_rsc_3_11_clkw_en),
      .q(yt_rsc_3_11_q),
      .radr(yt_rsc_3_11_radr),
      .we(yt_rsc_3_11_we),
      .d(yt_rsc_3_11_d),
      .wadr(yt_rsc_3_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_3_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_115_4_32_16_16_32_1_gen yt_rsc_3_12_i
      (
      .clkr_en(yt_rsc_3_12_clkr_en),
      .clkw_en(yt_rsc_3_12_clkw_en),
      .q(yt_rsc_3_12_q),
      .radr(yt_rsc_3_12_radr),
      .we(yt_rsc_3_12_we),
      .d(yt_rsc_3_12_d),
      .wadr(yt_rsc_3_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_3_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_116_4_32_16_16_32_1_gen yt_rsc_3_13_i
      (
      .clkr_en(yt_rsc_3_13_clkr_en),
      .clkw_en(yt_rsc_3_13_clkw_en),
      .q(yt_rsc_3_13_q),
      .radr(yt_rsc_3_13_radr),
      .we(yt_rsc_3_13_we),
      .d(yt_rsc_3_13_d),
      .wadr(yt_rsc_3_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_3_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_117_4_32_16_16_32_1_gen yt_rsc_3_14_i
      (
      .clkr_en(yt_rsc_3_14_clkr_en),
      .clkw_en(yt_rsc_3_14_clkw_en),
      .q(yt_rsc_3_14_q),
      .radr(yt_rsc_3_14_radr),
      .we(yt_rsc_3_14_we),
      .d(yt_rsc_3_14_d),
      .wadr(yt_rsc_3_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_3_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_118_4_32_16_16_32_1_gen yt_rsc_3_15_i
      (
      .clkr_en(yt_rsc_3_15_clkr_en),
      .clkw_en(yt_rsc_3_15_clkw_en),
      .q(yt_rsc_3_15_q),
      .radr(yt_rsc_3_15_radr),
      .we(yt_rsc_3_15_we),
      .d(yt_rsc_3_15_d),
      .wadr(yt_rsc_3_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_0_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_3_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_3_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_119_4_32_16_16_32_1_gen yt_rsc_3_16_i
      (
      .clkr_en(yt_rsc_3_16_clkr_en),
      .clkw_en(yt_rsc_3_16_clkw_en),
      .q(yt_rsc_3_16_q),
      .radr(yt_rsc_3_16_radr),
      .we(yt_rsc_3_16_we),
      .d(yt_rsc_3_16_d),
      .wadr(yt_rsc_3_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_0_i_d_d_iff),
      .q_d(yt_rsc_3_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_120_4_32_16_16_32_1_gen yt_rsc_3_17_i
      (
      .clkr_en(yt_rsc_3_17_clkr_en),
      .clkw_en(yt_rsc_3_17_clkw_en),
      .q(yt_rsc_3_17_q),
      .radr(yt_rsc_3_17_radr),
      .we(yt_rsc_3_17_we),
      .d(yt_rsc_3_17_d),
      .wadr(yt_rsc_3_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_1_i_d_d_iff),
      .q_d(yt_rsc_3_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_121_4_32_16_16_32_1_gen yt_rsc_3_18_i
      (
      .clkr_en(yt_rsc_3_18_clkr_en),
      .clkw_en(yt_rsc_3_18_clkw_en),
      .q(yt_rsc_3_18_q),
      .radr(yt_rsc_3_18_radr),
      .we(yt_rsc_3_18_we),
      .d(yt_rsc_3_18_d),
      .wadr(yt_rsc_3_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_2_i_d_d_iff),
      .q_d(yt_rsc_3_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_122_4_32_16_16_32_1_gen yt_rsc_3_19_i
      (
      .clkr_en(yt_rsc_3_19_clkr_en),
      .clkw_en(yt_rsc_3_19_clkw_en),
      .q(yt_rsc_3_19_q),
      .radr(yt_rsc_3_19_radr),
      .we(yt_rsc_3_19_we),
      .d(yt_rsc_3_19_d),
      .wadr(yt_rsc_3_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_3_i_d_d_iff),
      .q_d(yt_rsc_3_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_123_4_32_16_16_32_1_gen yt_rsc_3_20_i
      (
      .clkr_en(yt_rsc_3_20_clkr_en),
      .clkw_en(yt_rsc_3_20_clkw_en),
      .q(yt_rsc_3_20_q),
      .radr(yt_rsc_3_20_radr),
      .we(yt_rsc_3_20_we),
      .d(yt_rsc_3_20_d),
      .wadr(yt_rsc_3_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_4_i_d_d_iff),
      .q_d(yt_rsc_3_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_124_4_32_16_16_32_1_gen yt_rsc_3_21_i
      (
      .clkr_en(yt_rsc_3_21_clkr_en),
      .clkw_en(yt_rsc_3_21_clkw_en),
      .q(yt_rsc_3_21_q),
      .radr(yt_rsc_3_21_radr),
      .we(yt_rsc_3_21_we),
      .d(yt_rsc_3_21_d),
      .wadr(yt_rsc_3_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_5_i_d_d_iff),
      .q_d(yt_rsc_3_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_125_4_32_16_16_32_1_gen yt_rsc_3_22_i
      (
      .clkr_en(yt_rsc_3_22_clkr_en),
      .clkw_en(yt_rsc_3_22_clkw_en),
      .q(yt_rsc_3_22_q),
      .radr(yt_rsc_3_22_radr),
      .we(yt_rsc_3_22_we),
      .d(yt_rsc_3_22_d),
      .wadr(yt_rsc_3_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_6_i_d_d_iff),
      .q_d(yt_rsc_3_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_126_4_32_16_16_32_1_gen yt_rsc_3_23_i
      (
      .clkr_en(yt_rsc_3_23_clkr_en),
      .clkw_en(yt_rsc_3_23_clkw_en),
      .q(yt_rsc_3_23_q),
      .radr(yt_rsc_3_23_radr),
      .we(yt_rsc_3_23_we),
      .d(yt_rsc_3_23_d),
      .wadr(yt_rsc_3_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_7_i_d_d_iff),
      .q_d(yt_rsc_3_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_0_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_127_4_32_16_16_32_1_gen yt_rsc_3_24_i
      (
      .clkr_en(yt_rsc_3_24_clkr_en),
      .clkw_en(yt_rsc_3_24_clkw_en),
      .q(yt_rsc_3_24_q),
      .radr(yt_rsc_3_24_radr),
      .we(yt_rsc_3_24_we),
      .d(yt_rsc_3_24_d),
      .wadr(yt_rsc_3_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_8_i_d_d_iff),
      .q_d(yt_rsc_3_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_1_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_128_4_32_16_16_32_1_gen yt_rsc_3_25_i
      (
      .clkr_en(yt_rsc_3_25_clkr_en),
      .clkw_en(yt_rsc_3_25_clkw_en),
      .q(yt_rsc_3_25_q),
      .radr(yt_rsc_3_25_radr),
      .we(yt_rsc_3_25_we),
      .d(yt_rsc_3_25_d),
      .wadr(yt_rsc_3_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_9_i_d_d_iff),
      .q_d(yt_rsc_3_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_2_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_129_4_32_16_16_32_1_gen yt_rsc_3_26_i
      (
      .clkr_en(yt_rsc_3_26_clkr_en),
      .clkw_en(yt_rsc_3_26_clkw_en),
      .q(yt_rsc_3_26_q),
      .radr(yt_rsc_3_26_radr),
      .we(yt_rsc_3_26_we),
      .d(yt_rsc_3_26_d),
      .wadr(yt_rsc_3_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_10_i_d_d_iff),
      .q_d(yt_rsc_3_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_10_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_130_4_32_16_16_32_1_gen yt_rsc_3_27_i
      (
      .clkr_en(yt_rsc_3_27_clkr_en),
      .clkw_en(yt_rsc_3_27_clkw_en),
      .q(yt_rsc_3_27_q),
      .radr(yt_rsc_3_27_radr),
      .we(yt_rsc_3_27_we),
      .d(yt_rsc_3_27_d),
      .wadr(yt_rsc_3_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_11_i_d_d_iff),
      .q_d(yt_rsc_3_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_11_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_131_4_32_16_16_32_1_gen yt_rsc_3_28_i
      (
      .clkr_en(yt_rsc_3_28_clkr_en),
      .clkw_en(yt_rsc_3_28_clkw_en),
      .q(yt_rsc_3_28_q),
      .radr(yt_rsc_3_28_radr),
      .we(yt_rsc_3_28_we),
      .d(yt_rsc_3_28_d),
      .wadr(yt_rsc_3_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_12_i_d_d_iff),
      .q_d(yt_rsc_3_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_3_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_132_4_32_16_16_32_1_gen yt_rsc_3_29_i
      (
      .clkr_en(yt_rsc_3_29_clkr_en),
      .clkw_en(yt_rsc_3_29_clkw_en),
      .q(yt_rsc_3_29_q),
      .radr(yt_rsc_3_29_radr),
      .we(yt_rsc_3_29_we),
      .d(yt_rsc_3_29_d),
      .wadr(yt_rsc_3_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_13_i_d_d_iff),
      .q_d(yt_rsc_3_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_4_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_133_4_32_16_16_32_1_gen yt_rsc_3_30_i
      (
      .clkr_en(yt_rsc_3_30_clkr_en),
      .clkw_en(yt_rsc_3_30_clkw_en),
      .q(yt_rsc_3_30_q),
      .radr(yt_rsc_3_30_radr),
      .we(yt_rsc_3_30_we),
      .d(yt_rsc_3_30_d),
      .wadr(yt_rsc_3_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_14_i_d_d_iff),
      .q_d(yt_rsc_3_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_5_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_134_4_32_16_16_32_1_gen yt_rsc_3_31_i
      (
      .clkr_en(yt_rsc_3_31_clkr_en),
      .clkw_en(yt_rsc_3_31_clkw_en),
      .q(yt_rsc_3_31_q),
      .radr(yt_rsc_3_31_radr),
      .we(yt_rsc_3_31_we),
      .d(yt_rsc_3_31_d),
      .wadr(yt_rsc_3_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_3_16_i_clkr_en_d),
      .d_d(yt_rsc_0_15_i_d_d_iff),
      .q_d(yt_rsc_3_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_0_6_i_wadr_d_iff),
      .we_d(yt_rsc_3_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_3_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_135_4_32_16_16_32_1_gen yt_rsc_4_0_i
      (
      .clkr_en(yt_rsc_4_0_clkr_en),
      .clkw_en(yt_rsc_4_0_clkw_en),
      .q(yt_rsc_4_0_q),
      .radr(yt_rsc_4_0_radr),
      .we(yt_rsc_4_0_we),
      .d(yt_rsc_4_0_d),
      .wadr(yt_rsc_4_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_4_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_136_4_32_16_16_32_1_gen yt_rsc_4_1_i
      (
      .clkr_en(yt_rsc_4_1_clkr_en),
      .clkw_en(yt_rsc_4_1_clkw_en),
      .q(yt_rsc_4_1_q),
      .radr(yt_rsc_4_1_radr),
      .we(yt_rsc_4_1_we),
      .d(yt_rsc_4_1_d),
      .wadr(yt_rsc_4_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_4_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_137_4_32_16_16_32_1_gen yt_rsc_4_2_i
      (
      .clkr_en(yt_rsc_4_2_clkr_en),
      .clkw_en(yt_rsc_4_2_clkw_en),
      .q(yt_rsc_4_2_q),
      .radr(yt_rsc_4_2_radr),
      .we(yt_rsc_4_2_we),
      .d(yt_rsc_4_2_d),
      .wadr(yt_rsc_4_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_4_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_138_4_32_16_16_32_1_gen yt_rsc_4_3_i
      (
      .clkr_en(yt_rsc_4_3_clkr_en),
      .clkw_en(yt_rsc_4_3_clkw_en),
      .q(yt_rsc_4_3_q),
      .radr(yt_rsc_4_3_radr),
      .we(yt_rsc_4_3_we),
      .d(yt_rsc_4_3_d),
      .wadr(yt_rsc_4_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_4_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_139_4_32_16_16_32_1_gen yt_rsc_4_4_i
      (
      .clkr_en(yt_rsc_4_4_clkr_en),
      .clkw_en(yt_rsc_4_4_clkw_en),
      .q(yt_rsc_4_4_q),
      .radr(yt_rsc_4_4_radr),
      .we(yt_rsc_4_4_we),
      .d(yt_rsc_4_4_d),
      .wadr(yt_rsc_4_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_4_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_140_4_32_16_16_32_1_gen yt_rsc_4_5_i
      (
      .clkr_en(yt_rsc_4_5_clkr_en),
      .clkw_en(yt_rsc_4_5_clkw_en),
      .q(yt_rsc_4_5_q),
      .radr(yt_rsc_4_5_radr),
      .we(yt_rsc_4_5_we),
      .d(yt_rsc_4_5_d),
      .wadr(yt_rsc_4_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_4_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_141_4_32_16_16_32_1_gen yt_rsc_4_6_i
      (
      .clkr_en(yt_rsc_4_6_clkr_en),
      .clkw_en(yt_rsc_4_6_clkw_en),
      .q(yt_rsc_4_6_q),
      .radr(yt_rsc_4_6_radr),
      .we(yt_rsc_4_6_we),
      .d(yt_rsc_4_6_d),
      .wadr(yt_rsc_4_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_4_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_142_4_32_16_16_32_1_gen yt_rsc_4_7_i
      (
      .clkr_en(yt_rsc_4_7_clkr_en),
      .clkw_en(yt_rsc_4_7_clkw_en),
      .q(yt_rsc_4_7_q),
      .radr(yt_rsc_4_7_radr),
      .we(yt_rsc_4_7_we),
      .d(yt_rsc_4_7_d),
      .wadr(yt_rsc_4_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_4_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_143_4_32_16_16_32_1_gen yt_rsc_4_8_i
      (
      .clkr_en(yt_rsc_4_8_clkr_en),
      .clkw_en(yt_rsc_4_8_clkw_en),
      .q(yt_rsc_4_8_q),
      .radr(yt_rsc_4_8_radr),
      .we(yt_rsc_4_8_we),
      .d(yt_rsc_4_8_d),
      .wadr(yt_rsc_4_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_4_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_144_4_32_16_16_32_1_gen yt_rsc_4_9_i
      (
      .clkr_en(yt_rsc_4_9_clkr_en),
      .clkw_en(yt_rsc_4_9_clkw_en),
      .q(yt_rsc_4_9_q),
      .radr(yt_rsc_4_9_radr),
      .we(yt_rsc_4_9_we),
      .d(yt_rsc_4_9_d),
      .wadr(yt_rsc_4_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_4_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_145_4_32_16_16_32_1_gen yt_rsc_4_10_i
      (
      .clkr_en(yt_rsc_4_10_clkr_en),
      .clkw_en(yt_rsc_4_10_clkw_en),
      .q(yt_rsc_4_10_q),
      .radr(yt_rsc_4_10_radr),
      .we(yt_rsc_4_10_we),
      .d(yt_rsc_4_10_d),
      .wadr(yt_rsc_4_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_4_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_146_4_32_16_16_32_1_gen yt_rsc_4_11_i
      (
      .clkr_en(yt_rsc_4_11_clkr_en),
      .clkw_en(yt_rsc_4_11_clkw_en),
      .q(yt_rsc_4_11_q),
      .radr(yt_rsc_4_11_radr),
      .we(yt_rsc_4_11_we),
      .d(yt_rsc_4_11_d),
      .wadr(yt_rsc_4_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_4_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_147_4_32_16_16_32_1_gen yt_rsc_4_12_i
      (
      .clkr_en(yt_rsc_4_12_clkr_en),
      .clkw_en(yt_rsc_4_12_clkw_en),
      .q(yt_rsc_4_12_q),
      .radr(yt_rsc_4_12_radr),
      .we(yt_rsc_4_12_we),
      .d(yt_rsc_4_12_d),
      .wadr(yt_rsc_4_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_4_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_148_4_32_16_16_32_1_gen yt_rsc_4_13_i
      (
      .clkr_en(yt_rsc_4_13_clkr_en),
      .clkw_en(yt_rsc_4_13_clkw_en),
      .q(yt_rsc_4_13_q),
      .radr(yt_rsc_4_13_radr),
      .we(yt_rsc_4_13_we),
      .d(yt_rsc_4_13_d),
      .wadr(yt_rsc_4_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_4_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_149_4_32_16_16_32_1_gen yt_rsc_4_14_i
      (
      .clkr_en(yt_rsc_4_14_clkr_en),
      .clkw_en(yt_rsc_4_14_clkw_en),
      .q(yt_rsc_4_14_q),
      .radr(yt_rsc_4_14_radr),
      .we(yt_rsc_4_14_we),
      .d(yt_rsc_4_14_d),
      .wadr(yt_rsc_4_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_4_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_150_4_32_16_16_32_1_gen yt_rsc_4_15_i
      (
      .clkr_en(yt_rsc_4_15_clkr_en),
      .clkw_en(yt_rsc_4_15_clkw_en),
      .q(yt_rsc_4_15_q),
      .radr(yt_rsc_4_15_radr),
      .we(yt_rsc_4_15_we),
      .d(yt_rsc_4_15_d),
      .wadr(yt_rsc_4_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_0_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_4_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_4_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_151_4_32_16_16_32_1_gen yt_rsc_4_16_i
      (
      .clkr_en(yt_rsc_4_16_clkr_en),
      .clkw_en(yt_rsc_4_16_clkw_en),
      .q(yt_rsc_4_16_q),
      .radr(yt_rsc_4_16_radr),
      .we(yt_rsc_4_16_we),
      .d(yt_rsc_4_16_d),
      .wadr(yt_rsc_4_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_4_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_152_4_32_16_16_32_1_gen yt_rsc_4_17_i
      (
      .clkr_en(yt_rsc_4_17_clkr_en),
      .clkw_en(yt_rsc_4_17_clkw_en),
      .q(yt_rsc_4_17_q),
      .radr(yt_rsc_4_17_radr),
      .we(yt_rsc_4_17_we),
      .d(yt_rsc_4_17_d),
      .wadr(yt_rsc_4_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_4_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_153_4_32_16_16_32_1_gen yt_rsc_4_18_i
      (
      .clkr_en(yt_rsc_4_18_clkr_en),
      .clkw_en(yt_rsc_4_18_clkw_en),
      .q(yt_rsc_4_18_q),
      .radr(yt_rsc_4_18_radr),
      .we(yt_rsc_4_18_we),
      .d(yt_rsc_4_18_d),
      .wadr(yt_rsc_4_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_4_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_154_4_32_16_16_32_1_gen yt_rsc_4_19_i
      (
      .clkr_en(yt_rsc_4_19_clkr_en),
      .clkw_en(yt_rsc_4_19_clkw_en),
      .q(yt_rsc_4_19_q),
      .radr(yt_rsc_4_19_radr),
      .we(yt_rsc_4_19_we),
      .d(yt_rsc_4_19_d),
      .wadr(yt_rsc_4_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_4_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_155_4_32_16_16_32_1_gen yt_rsc_4_20_i
      (
      .clkr_en(yt_rsc_4_20_clkr_en),
      .clkw_en(yt_rsc_4_20_clkw_en),
      .q(yt_rsc_4_20_q),
      .radr(yt_rsc_4_20_radr),
      .we(yt_rsc_4_20_we),
      .d(yt_rsc_4_20_d),
      .wadr(yt_rsc_4_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_4_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_156_4_32_16_16_32_1_gen yt_rsc_4_21_i
      (
      .clkr_en(yt_rsc_4_21_clkr_en),
      .clkw_en(yt_rsc_4_21_clkw_en),
      .q(yt_rsc_4_21_q),
      .radr(yt_rsc_4_21_radr),
      .we(yt_rsc_4_21_we),
      .d(yt_rsc_4_21_d),
      .wadr(yt_rsc_4_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_4_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_157_4_32_16_16_32_1_gen yt_rsc_4_22_i
      (
      .clkr_en(yt_rsc_4_22_clkr_en),
      .clkw_en(yt_rsc_4_22_clkw_en),
      .q(yt_rsc_4_22_q),
      .radr(yt_rsc_4_22_radr),
      .we(yt_rsc_4_22_we),
      .d(yt_rsc_4_22_d),
      .wadr(yt_rsc_4_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_4_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_158_4_32_16_16_32_1_gen yt_rsc_4_23_i
      (
      .clkr_en(yt_rsc_4_23_clkr_en),
      .clkw_en(yt_rsc_4_23_clkw_en),
      .q(yt_rsc_4_23_q),
      .radr(yt_rsc_4_23_radr),
      .we(yt_rsc_4_23_we),
      .d(yt_rsc_4_23_d),
      .wadr(yt_rsc_4_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_4_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_159_4_32_16_16_32_1_gen yt_rsc_4_24_i
      (
      .clkr_en(yt_rsc_4_24_clkr_en),
      .clkw_en(yt_rsc_4_24_clkw_en),
      .q(yt_rsc_4_24_q),
      .radr(yt_rsc_4_24_radr),
      .we(yt_rsc_4_24_we),
      .d(yt_rsc_4_24_d),
      .wadr(yt_rsc_4_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_4_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_160_4_32_16_16_32_1_gen yt_rsc_4_25_i
      (
      .clkr_en(yt_rsc_4_25_clkr_en),
      .clkw_en(yt_rsc_4_25_clkw_en),
      .q(yt_rsc_4_25_q),
      .radr(yt_rsc_4_25_radr),
      .we(yt_rsc_4_25_we),
      .d(yt_rsc_4_25_d),
      .wadr(yt_rsc_4_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_4_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_161_4_32_16_16_32_1_gen yt_rsc_4_26_i
      (
      .clkr_en(yt_rsc_4_26_clkr_en),
      .clkw_en(yt_rsc_4_26_clkw_en),
      .q(yt_rsc_4_26_q),
      .radr(yt_rsc_4_26_radr),
      .we(yt_rsc_4_26_we),
      .d(yt_rsc_4_26_d),
      .wadr(yt_rsc_4_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_4_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_162_4_32_16_16_32_1_gen yt_rsc_4_27_i
      (
      .clkr_en(yt_rsc_4_27_clkr_en),
      .clkw_en(yt_rsc_4_27_clkw_en),
      .q(yt_rsc_4_27_q),
      .radr(yt_rsc_4_27_radr),
      .we(yt_rsc_4_27_we),
      .d(yt_rsc_4_27_d),
      .wadr(yt_rsc_4_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_4_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_163_4_32_16_16_32_1_gen yt_rsc_4_28_i
      (
      .clkr_en(yt_rsc_4_28_clkr_en),
      .clkw_en(yt_rsc_4_28_clkw_en),
      .q(yt_rsc_4_28_q),
      .radr(yt_rsc_4_28_radr),
      .we(yt_rsc_4_28_we),
      .d(yt_rsc_4_28_d),
      .wadr(yt_rsc_4_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_4_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_164_4_32_16_16_32_1_gen yt_rsc_4_29_i
      (
      .clkr_en(yt_rsc_4_29_clkr_en),
      .clkw_en(yt_rsc_4_29_clkw_en),
      .q(yt_rsc_4_29_q),
      .radr(yt_rsc_4_29_radr),
      .we(yt_rsc_4_29_we),
      .d(yt_rsc_4_29_d),
      .wadr(yt_rsc_4_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_4_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_165_4_32_16_16_32_1_gen yt_rsc_4_30_i
      (
      .clkr_en(yt_rsc_4_30_clkr_en),
      .clkw_en(yt_rsc_4_30_clkw_en),
      .q(yt_rsc_4_30_q),
      .radr(yt_rsc_4_30_radr),
      .we(yt_rsc_4_30_we),
      .d(yt_rsc_4_30_d),
      .wadr(yt_rsc_4_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_4_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_166_4_32_16_16_32_1_gen yt_rsc_4_31_i
      (
      .clkr_en(yt_rsc_4_31_clkr_en),
      .clkw_en(yt_rsc_4_31_clkw_en),
      .q(yt_rsc_4_31_q),
      .radr(yt_rsc_4_31_radr),
      .we(yt_rsc_4_31_we),
      .d(yt_rsc_4_31_d),
      .wadr(yt_rsc_4_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_4_16_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_4_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_4_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_4_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_167_4_32_16_16_32_1_gen yt_rsc_5_0_i
      (
      .clkr_en(yt_rsc_5_0_clkr_en),
      .clkw_en(yt_rsc_5_0_clkw_en),
      .q(yt_rsc_5_0_q),
      .radr(yt_rsc_5_0_radr),
      .we(yt_rsc_5_0_we),
      .d(yt_rsc_5_0_d),
      .wadr(yt_rsc_5_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_5_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_168_4_32_16_16_32_1_gen yt_rsc_5_1_i
      (
      .clkr_en(yt_rsc_5_1_clkr_en),
      .clkw_en(yt_rsc_5_1_clkw_en),
      .q(yt_rsc_5_1_q),
      .radr(yt_rsc_5_1_radr),
      .we(yt_rsc_5_1_we),
      .d(yt_rsc_5_1_d),
      .wadr(yt_rsc_5_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_5_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_169_4_32_16_16_32_1_gen yt_rsc_5_2_i
      (
      .clkr_en(yt_rsc_5_2_clkr_en),
      .clkw_en(yt_rsc_5_2_clkw_en),
      .q(yt_rsc_5_2_q),
      .radr(yt_rsc_5_2_radr),
      .we(yt_rsc_5_2_we),
      .d(yt_rsc_5_2_d),
      .wadr(yt_rsc_5_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_5_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_170_4_32_16_16_32_1_gen yt_rsc_5_3_i
      (
      .clkr_en(yt_rsc_5_3_clkr_en),
      .clkw_en(yt_rsc_5_3_clkw_en),
      .q(yt_rsc_5_3_q),
      .radr(yt_rsc_5_3_radr),
      .we(yt_rsc_5_3_we),
      .d(yt_rsc_5_3_d),
      .wadr(yt_rsc_5_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_5_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_171_4_32_16_16_32_1_gen yt_rsc_5_4_i
      (
      .clkr_en(yt_rsc_5_4_clkr_en),
      .clkw_en(yt_rsc_5_4_clkw_en),
      .q(yt_rsc_5_4_q),
      .radr(yt_rsc_5_4_radr),
      .we(yt_rsc_5_4_we),
      .d(yt_rsc_5_4_d),
      .wadr(yt_rsc_5_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_5_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_172_4_32_16_16_32_1_gen yt_rsc_5_5_i
      (
      .clkr_en(yt_rsc_5_5_clkr_en),
      .clkw_en(yt_rsc_5_5_clkw_en),
      .q(yt_rsc_5_5_q),
      .radr(yt_rsc_5_5_radr),
      .we(yt_rsc_5_5_we),
      .d(yt_rsc_5_5_d),
      .wadr(yt_rsc_5_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_5_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_173_4_32_16_16_32_1_gen yt_rsc_5_6_i
      (
      .clkr_en(yt_rsc_5_6_clkr_en),
      .clkw_en(yt_rsc_5_6_clkw_en),
      .q(yt_rsc_5_6_q),
      .radr(yt_rsc_5_6_radr),
      .we(yt_rsc_5_6_we),
      .d(yt_rsc_5_6_d),
      .wadr(yt_rsc_5_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_5_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_174_4_32_16_16_32_1_gen yt_rsc_5_7_i
      (
      .clkr_en(yt_rsc_5_7_clkr_en),
      .clkw_en(yt_rsc_5_7_clkw_en),
      .q(yt_rsc_5_7_q),
      .radr(yt_rsc_5_7_radr),
      .we(yt_rsc_5_7_we),
      .d(yt_rsc_5_7_d),
      .wadr(yt_rsc_5_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_5_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_175_4_32_16_16_32_1_gen yt_rsc_5_8_i
      (
      .clkr_en(yt_rsc_5_8_clkr_en),
      .clkw_en(yt_rsc_5_8_clkw_en),
      .q(yt_rsc_5_8_q),
      .radr(yt_rsc_5_8_radr),
      .we(yt_rsc_5_8_we),
      .d(yt_rsc_5_8_d),
      .wadr(yt_rsc_5_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_5_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_176_4_32_16_16_32_1_gen yt_rsc_5_9_i
      (
      .clkr_en(yt_rsc_5_9_clkr_en),
      .clkw_en(yt_rsc_5_9_clkw_en),
      .q(yt_rsc_5_9_q),
      .radr(yt_rsc_5_9_radr),
      .we(yt_rsc_5_9_we),
      .d(yt_rsc_5_9_d),
      .wadr(yt_rsc_5_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_5_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_177_4_32_16_16_32_1_gen yt_rsc_5_10_i
      (
      .clkr_en(yt_rsc_5_10_clkr_en),
      .clkw_en(yt_rsc_5_10_clkw_en),
      .q(yt_rsc_5_10_q),
      .radr(yt_rsc_5_10_radr),
      .we(yt_rsc_5_10_we),
      .d(yt_rsc_5_10_d),
      .wadr(yt_rsc_5_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_5_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_178_4_32_16_16_32_1_gen yt_rsc_5_11_i
      (
      .clkr_en(yt_rsc_5_11_clkr_en),
      .clkw_en(yt_rsc_5_11_clkw_en),
      .q(yt_rsc_5_11_q),
      .radr(yt_rsc_5_11_radr),
      .we(yt_rsc_5_11_we),
      .d(yt_rsc_5_11_d),
      .wadr(yt_rsc_5_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_5_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_179_4_32_16_16_32_1_gen yt_rsc_5_12_i
      (
      .clkr_en(yt_rsc_5_12_clkr_en),
      .clkw_en(yt_rsc_5_12_clkw_en),
      .q(yt_rsc_5_12_q),
      .radr(yt_rsc_5_12_radr),
      .we(yt_rsc_5_12_we),
      .d(yt_rsc_5_12_d),
      .wadr(yt_rsc_5_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_5_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_180_4_32_16_16_32_1_gen yt_rsc_5_13_i
      (
      .clkr_en(yt_rsc_5_13_clkr_en),
      .clkw_en(yt_rsc_5_13_clkw_en),
      .q(yt_rsc_5_13_q),
      .radr(yt_rsc_5_13_radr),
      .we(yt_rsc_5_13_we),
      .d(yt_rsc_5_13_d),
      .wadr(yt_rsc_5_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_5_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_181_4_32_16_16_32_1_gen yt_rsc_5_14_i
      (
      .clkr_en(yt_rsc_5_14_clkr_en),
      .clkw_en(yt_rsc_5_14_clkw_en),
      .q(yt_rsc_5_14_q),
      .radr(yt_rsc_5_14_radr),
      .we(yt_rsc_5_14_we),
      .d(yt_rsc_5_14_d),
      .wadr(yt_rsc_5_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_5_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_182_4_32_16_16_32_1_gen yt_rsc_5_15_i
      (
      .clkr_en(yt_rsc_5_15_clkr_en),
      .clkw_en(yt_rsc_5_15_clkw_en),
      .q(yt_rsc_5_15_q),
      .radr(yt_rsc_5_15_radr),
      .we(yt_rsc_5_15_we),
      .d(yt_rsc_5_15_d),
      .wadr(yt_rsc_5_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_0_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_5_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_5_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_183_4_32_16_16_32_1_gen yt_rsc_5_16_i
      (
      .clkr_en(yt_rsc_5_16_clkr_en),
      .clkw_en(yt_rsc_5_16_clkw_en),
      .q(yt_rsc_5_16_q),
      .radr(yt_rsc_5_16_radr),
      .we(yt_rsc_5_16_we),
      .d(yt_rsc_5_16_d),
      .wadr(yt_rsc_5_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_5_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_184_4_32_16_16_32_1_gen yt_rsc_5_17_i
      (
      .clkr_en(yt_rsc_5_17_clkr_en),
      .clkw_en(yt_rsc_5_17_clkw_en),
      .q(yt_rsc_5_17_q),
      .radr(yt_rsc_5_17_radr),
      .we(yt_rsc_5_17_we),
      .d(yt_rsc_5_17_d),
      .wadr(yt_rsc_5_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_5_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_185_4_32_16_16_32_1_gen yt_rsc_5_18_i
      (
      .clkr_en(yt_rsc_5_18_clkr_en),
      .clkw_en(yt_rsc_5_18_clkw_en),
      .q(yt_rsc_5_18_q),
      .radr(yt_rsc_5_18_radr),
      .we(yt_rsc_5_18_we),
      .d(yt_rsc_5_18_d),
      .wadr(yt_rsc_5_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_5_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_186_4_32_16_16_32_1_gen yt_rsc_5_19_i
      (
      .clkr_en(yt_rsc_5_19_clkr_en),
      .clkw_en(yt_rsc_5_19_clkw_en),
      .q(yt_rsc_5_19_q),
      .radr(yt_rsc_5_19_radr),
      .we(yt_rsc_5_19_we),
      .d(yt_rsc_5_19_d),
      .wadr(yt_rsc_5_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_5_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_187_4_32_16_16_32_1_gen yt_rsc_5_20_i
      (
      .clkr_en(yt_rsc_5_20_clkr_en),
      .clkw_en(yt_rsc_5_20_clkw_en),
      .q(yt_rsc_5_20_q),
      .radr(yt_rsc_5_20_radr),
      .we(yt_rsc_5_20_we),
      .d(yt_rsc_5_20_d),
      .wadr(yt_rsc_5_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_5_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_188_4_32_16_16_32_1_gen yt_rsc_5_21_i
      (
      .clkr_en(yt_rsc_5_21_clkr_en),
      .clkw_en(yt_rsc_5_21_clkw_en),
      .q(yt_rsc_5_21_q),
      .radr(yt_rsc_5_21_radr),
      .we(yt_rsc_5_21_we),
      .d(yt_rsc_5_21_d),
      .wadr(yt_rsc_5_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_5_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_189_4_32_16_16_32_1_gen yt_rsc_5_22_i
      (
      .clkr_en(yt_rsc_5_22_clkr_en),
      .clkw_en(yt_rsc_5_22_clkw_en),
      .q(yt_rsc_5_22_q),
      .radr(yt_rsc_5_22_radr),
      .we(yt_rsc_5_22_we),
      .d(yt_rsc_5_22_d),
      .wadr(yt_rsc_5_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_5_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_190_4_32_16_16_32_1_gen yt_rsc_5_23_i
      (
      .clkr_en(yt_rsc_5_23_clkr_en),
      .clkw_en(yt_rsc_5_23_clkw_en),
      .q(yt_rsc_5_23_q),
      .radr(yt_rsc_5_23_radr),
      .we(yt_rsc_5_23_we),
      .d(yt_rsc_5_23_d),
      .wadr(yt_rsc_5_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_5_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_191_4_32_16_16_32_1_gen yt_rsc_5_24_i
      (
      .clkr_en(yt_rsc_5_24_clkr_en),
      .clkw_en(yt_rsc_5_24_clkw_en),
      .q(yt_rsc_5_24_q),
      .radr(yt_rsc_5_24_radr),
      .we(yt_rsc_5_24_we),
      .d(yt_rsc_5_24_d),
      .wadr(yt_rsc_5_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_5_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_192_4_32_16_16_32_1_gen yt_rsc_5_25_i
      (
      .clkr_en(yt_rsc_5_25_clkr_en),
      .clkw_en(yt_rsc_5_25_clkw_en),
      .q(yt_rsc_5_25_q),
      .radr(yt_rsc_5_25_radr),
      .we(yt_rsc_5_25_we),
      .d(yt_rsc_5_25_d),
      .wadr(yt_rsc_5_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_5_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_193_4_32_16_16_32_1_gen yt_rsc_5_26_i
      (
      .clkr_en(yt_rsc_5_26_clkr_en),
      .clkw_en(yt_rsc_5_26_clkw_en),
      .q(yt_rsc_5_26_q),
      .radr(yt_rsc_5_26_radr),
      .we(yt_rsc_5_26_we),
      .d(yt_rsc_5_26_d),
      .wadr(yt_rsc_5_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_5_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_194_4_32_16_16_32_1_gen yt_rsc_5_27_i
      (
      .clkr_en(yt_rsc_5_27_clkr_en),
      .clkw_en(yt_rsc_5_27_clkw_en),
      .q(yt_rsc_5_27_q),
      .radr(yt_rsc_5_27_radr),
      .we(yt_rsc_5_27_we),
      .d(yt_rsc_5_27_d),
      .wadr(yt_rsc_5_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_5_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_195_4_32_16_16_32_1_gen yt_rsc_5_28_i
      (
      .clkr_en(yt_rsc_5_28_clkr_en),
      .clkw_en(yt_rsc_5_28_clkw_en),
      .q(yt_rsc_5_28_q),
      .radr(yt_rsc_5_28_radr),
      .we(yt_rsc_5_28_we),
      .d(yt_rsc_5_28_d),
      .wadr(yt_rsc_5_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_5_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_196_4_32_16_16_32_1_gen yt_rsc_5_29_i
      (
      .clkr_en(yt_rsc_5_29_clkr_en),
      .clkw_en(yt_rsc_5_29_clkw_en),
      .q(yt_rsc_5_29_q),
      .radr(yt_rsc_5_29_radr),
      .we(yt_rsc_5_29_we),
      .d(yt_rsc_5_29_d),
      .wadr(yt_rsc_5_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_5_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_197_4_32_16_16_32_1_gen yt_rsc_5_30_i
      (
      .clkr_en(yt_rsc_5_30_clkr_en),
      .clkw_en(yt_rsc_5_30_clkw_en),
      .q(yt_rsc_5_30_q),
      .radr(yt_rsc_5_30_radr),
      .we(yt_rsc_5_30_we),
      .d(yt_rsc_5_30_d),
      .wadr(yt_rsc_5_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_5_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_198_4_32_16_16_32_1_gen yt_rsc_5_31_i
      (
      .clkr_en(yt_rsc_5_31_clkr_en),
      .clkw_en(yt_rsc_5_31_clkw_en),
      .q(yt_rsc_5_31_q),
      .radr(yt_rsc_5_31_radr),
      .we(yt_rsc_5_31_we),
      .d(yt_rsc_5_31_d),
      .wadr(yt_rsc_5_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_5_16_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_5_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_5_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_5_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_199_4_32_16_16_32_1_gen yt_rsc_6_0_i
      (
      .clkr_en(yt_rsc_6_0_clkr_en),
      .clkw_en(yt_rsc_6_0_clkw_en),
      .q(yt_rsc_6_0_q),
      .radr(yt_rsc_6_0_radr),
      .we(yt_rsc_6_0_we),
      .d(yt_rsc_6_0_d),
      .wadr(yt_rsc_6_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_6_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_200_4_32_16_16_32_1_gen yt_rsc_6_1_i
      (
      .clkr_en(yt_rsc_6_1_clkr_en),
      .clkw_en(yt_rsc_6_1_clkw_en),
      .q(yt_rsc_6_1_q),
      .radr(yt_rsc_6_1_radr),
      .we(yt_rsc_6_1_we),
      .d(yt_rsc_6_1_d),
      .wadr(yt_rsc_6_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_6_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_201_4_32_16_16_32_1_gen yt_rsc_6_2_i
      (
      .clkr_en(yt_rsc_6_2_clkr_en),
      .clkw_en(yt_rsc_6_2_clkw_en),
      .q(yt_rsc_6_2_q),
      .radr(yt_rsc_6_2_radr),
      .we(yt_rsc_6_2_we),
      .d(yt_rsc_6_2_d),
      .wadr(yt_rsc_6_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_6_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_202_4_32_16_16_32_1_gen yt_rsc_6_3_i
      (
      .clkr_en(yt_rsc_6_3_clkr_en),
      .clkw_en(yt_rsc_6_3_clkw_en),
      .q(yt_rsc_6_3_q),
      .radr(yt_rsc_6_3_radr),
      .we(yt_rsc_6_3_we),
      .d(yt_rsc_6_3_d),
      .wadr(yt_rsc_6_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_6_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_203_4_32_16_16_32_1_gen yt_rsc_6_4_i
      (
      .clkr_en(yt_rsc_6_4_clkr_en),
      .clkw_en(yt_rsc_6_4_clkw_en),
      .q(yt_rsc_6_4_q),
      .radr(yt_rsc_6_4_radr),
      .we(yt_rsc_6_4_we),
      .d(yt_rsc_6_4_d),
      .wadr(yt_rsc_6_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_6_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_204_4_32_16_16_32_1_gen yt_rsc_6_5_i
      (
      .clkr_en(yt_rsc_6_5_clkr_en),
      .clkw_en(yt_rsc_6_5_clkw_en),
      .q(yt_rsc_6_5_q),
      .radr(yt_rsc_6_5_radr),
      .we(yt_rsc_6_5_we),
      .d(yt_rsc_6_5_d),
      .wadr(yt_rsc_6_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_6_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_205_4_32_16_16_32_1_gen yt_rsc_6_6_i
      (
      .clkr_en(yt_rsc_6_6_clkr_en),
      .clkw_en(yt_rsc_6_6_clkw_en),
      .q(yt_rsc_6_6_q),
      .radr(yt_rsc_6_6_radr),
      .we(yt_rsc_6_6_we),
      .d(yt_rsc_6_6_d),
      .wadr(yt_rsc_6_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_6_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_206_4_32_16_16_32_1_gen yt_rsc_6_7_i
      (
      .clkr_en(yt_rsc_6_7_clkr_en),
      .clkw_en(yt_rsc_6_7_clkw_en),
      .q(yt_rsc_6_7_q),
      .radr(yt_rsc_6_7_radr),
      .we(yt_rsc_6_7_we),
      .d(yt_rsc_6_7_d),
      .wadr(yt_rsc_6_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_6_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_207_4_32_16_16_32_1_gen yt_rsc_6_8_i
      (
      .clkr_en(yt_rsc_6_8_clkr_en),
      .clkw_en(yt_rsc_6_8_clkw_en),
      .q(yt_rsc_6_8_q),
      .radr(yt_rsc_6_8_radr),
      .we(yt_rsc_6_8_we),
      .d(yt_rsc_6_8_d),
      .wadr(yt_rsc_6_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_6_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_208_4_32_16_16_32_1_gen yt_rsc_6_9_i
      (
      .clkr_en(yt_rsc_6_9_clkr_en),
      .clkw_en(yt_rsc_6_9_clkw_en),
      .q(yt_rsc_6_9_q),
      .radr(yt_rsc_6_9_radr),
      .we(yt_rsc_6_9_we),
      .d(yt_rsc_6_9_d),
      .wadr(yt_rsc_6_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_6_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_209_4_32_16_16_32_1_gen yt_rsc_6_10_i
      (
      .clkr_en(yt_rsc_6_10_clkr_en),
      .clkw_en(yt_rsc_6_10_clkw_en),
      .q(yt_rsc_6_10_q),
      .radr(yt_rsc_6_10_radr),
      .we(yt_rsc_6_10_we),
      .d(yt_rsc_6_10_d),
      .wadr(yt_rsc_6_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_6_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_210_4_32_16_16_32_1_gen yt_rsc_6_11_i
      (
      .clkr_en(yt_rsc_6_11_clkr_en),
      .clkw_en(yt_rsc_6_11_clkw_en),
      .q(yt_rsc_6_11_q),
      .radr(yt_rsc_6_11_radr),
      .we(yt_rsc_6_11_we),
      .d(yt_rsc_6_11_d),
      .wadr(yt_rsc_6_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_6_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_211_4_32_16_16_32_1_gen yt_rsc_6_12_i
      (
      .clkr_en(yt_rsc_6_12_clkr_en),
      .clkw_en(yt_rsc_6_12_clkw_en),
      .q(yt_rsc_6_12_q),
      .radr(yt_rsc_6_12_radr),
      .we(yt_rsc_6_12_we),
      .d(yt_rsc_6_12_d),
      .wadr(yt_rsc_6_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_6_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_212_4_32_16_16_32_1_gen yt_rsc_6_13_i
      (
      .clkr_en(yt_rsc_6_13_clkr_en),
      .clkw_en(yt_rsc_6_13_clkw_en),
      .q(yt_rsc_6_13_q),
      .radr(yt_rsc_6_13_radr),
      .we(yt_rsc_6_13_we),
      .d(yt_rsc_6_13_d),
      .wadr(yt_rsc_6_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_6_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_213_4_32_16_16_32_1_gen yt_rsc_6_14_i
      (
      .clkr_en(yt_rsc_6_14_clkr_en),
      .clkw_en(yt_rsc_6_14_clkw_en),
      .q(yt_rsc_6_14_q),
      .radr(yt_rsc_6_14_radr),
      .we(yt_rsc_6_14_we),
      .d(yt_rsc_6_14_d),
      .wadr(yt_rsc_6_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_6_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_214_4_32_16_16_32_1_gen yt_rsc_6_15_i
      (
      .clkr_en(yt_rsc_6_15_clkr_en),
      .clkw_en(yt_rsc_6_15_clkw_en),
      .q(yt_rsc_6_15_q),
      .radr(yt_rsc_6_15_radr),
      .we(yt_rsc_6_15_we),
      .d(yt_rsc_6_15_d),
      .wadr(yt_rsc_6_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_0_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_6_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_6_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_215_4_32_16_16_32_1_gen yt_rsc_6_16_i
      (
      .clkr_en(yt_rsc_6_16_clkr_en),
      .clkw_en(yt_rsc_6_16_clkw_en),
      .q(yt_rsc_6_16_q),
      .radr(yt_rsc_6_16_radr),
      .we(yt_rsc_6_16_we),
      .d(yt_rsc_6_16_d),
      .wadr(yt_rsc_6_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_6_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_216_4_32_16_16_32_1_gen yt_rsc_6_17_i
      (
      .clkr_en(yt_rsc_6_17_clkr_en),
      .clkw_en(yt_rsc_6_17_clkw_en),
      .q(yt_rsc_6_17_q),
      .radr(yt_rsc_6_17_radr),
      .we(yt_rsc_6_17_we),
      .d(yt_rsc_6_17_d),
      .wadr(yt_rsc_6_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_6_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_217_4_32_16_16_32_1_gen yt_rsc_6_18_i
      (
      .clkr_en(yt_rsc_6_18_clkr_en),
      .clkw_en(yt_rsc_6_18_clkw_en),
      .q(yt_rsc_6_18_q),
      .radr(yt_rsc_6_18_radr),
      .we(yt_rsc_6_18_we),
      .d(yt_rsc_6_18_d),
      .wadr(yt_rsc_6_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_6_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_218_4_32_16_16_32_1_gen yt_rsc_6_19_i
      (
      .clkr_en(yt_rsc_6_19_clkr_en),
      .clkw_en(yt_rsc_6_19_clkw_en),
      .q(yt_rsc_6_19_q),
      .radr(yt_rsc_6_19_radr),
      .we(yt_rsc_6_19_we),
      .d(yt_rsc_6_19_d),
      .wadr(yt_rsc_6_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_6_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_219_4_32_16_16_32_1_gen yt_rsc_6_20_i
      (
      .clkr_en(yt_rsc_6_20_clkr_en),
      .clkw_en(yt_rsc_6_20_clkw_en),
      .q(yt_rsc_6_20_q),
      .radr(yt_rsc_6_20_radr),
      .we(yt_rsc_6_20_we),
      .d(yt_rsc_6_20_d),
      .wadr(yt_rsc_6_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_6_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_220_4_32_16_16_32_1_gen yt_rsc_6_21_i
      (
      .clkr_en(yt_rsc_6_21_clkr_en),
      .clkw_en(yt_rsc_6_21_clkw_en),
      .q(yt_rsc_6_21_q),
      .radr(yt_rsc_6_21_radr),
      .we(yt_rsc_6_21_we),
      .d(yt_rsc_6_21_d),
      .wadr(yt_rsc_6_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_6_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_221_4_32_16_16_32_1_gen yt_rsc_6_22_i
      (
      .clkr_en(yt_rsc_6_22_clkr_en),
      .clkw_en(yt_rsc_6_22_clkw_en),
      .q(yt_rsc_6_22_q),
      .radr(yt_rsc_6_22_radr),
      .we(yt_rsc_6_22_we),
      .d(yt_rsc_6_22_d),
      .wadr(yt_rsc_6_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_6_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_222_4_32_16_16_32_1_gen yt_rsc_6_23_i
      (
      .clkr_en(yt_rsc_6_23_clkr_en),
      .clkw_en(yt_rsc_6_23_clkw_en),
      .q(yt_rsc_6_23_q),
      .radr(yt_rsc_6_23_radr),
      .we(yt_rsc_6_23_we),
      .d(yt_rsc_6_23_d),
      .wadr(yt_rsc_6_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_6_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_223_4_32_16_16_32_1_gen yt_rsc_6_24_i
      (
      .clkr_en(yt_rsc_6_24_clkr_en),
      .clkw_en(yt_rsc_6_24_clkw_en),
      .q(yt_rsc_6_24_q),
      .radr(yt_rsc_6_24_radr),
      .we(yt_rsc_6_24_we),
      .d(yt_rsc_6_24_d),
      .wadr(yt_rsc_6_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_6_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_224_4_32_16_16_32_1_gen yt_rsc_6_25_i
      (
      .clkr_en(yt_rsc_6_25_clkr_en),
      .clkw_en(yt_rsc_6_25_clkw_en),
      .q(yt_rsc_6_25_q),
      .radr(yt_rsc_6_25_radr),
      .we(yt_rsc_6_25_we),
      .d(yt_rsc_6_25_d),
      .wadr(yt_rsc_6_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_6_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_225_4_32_16_16_32_1_gen yt_rsc_6_26_i
      (
      .clkr_en(yt_rsc_6_26_clkr_en),
      .clkw_en(yt_rsc_6_26_clkw_en),
      .q(yt_rsc_6_26_q),
      .radr(yt_rsc_6_26_radr),
      .we(yt_rsc_6_26_we),
      .d(yt_rsc_6_26_d),
      .wadr(yt_rsc_6_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_6_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_226_4_32_16_16_32_1_gen yt_rsc_6_27_i
      (
      .clkr_en(yt_rsc_6_27_clkr_en),
      .clkw_en(yt_rsc_6_27_clkw_en),
      .q(yt_rsc_6_27_q),
      .radr(yt_rsc_6_27_radr),
      .we(yt_rsc_6_27_we),
      .d(yt_rsc_6_27_d),
      .wadr(yt_rsc_6_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_6_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_227_4_32_16_16_32_1_gen yt_rsc_6_28_i
      (
      .clkr_en(yt_rsc_6_28_clkr_en),
      .clkw_en(yt_rsc_6_28_clkw_en),
      .q(yt_rsc_6_28_q),
      .radr(yt_rsc_6_28_radr),
      .we(yt_rsc_6_28_we),
      .d(yt_rsc_6_28_d),
      .wadr(yt_rsc_6_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_6_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_228_4_32_16_16_32_1_gen yt_rsc_6_29_i
      (
      .clkr_en(yt_rsc_6_29_clkr_en),
      .clkw_en(yt_rsc_6_29_clkw_en),
      .q(yt_rsc_6_29_q),
      .radr(yt_rsc_6_29_radr),
      .we(yt_rsc_6_29_we),
      .d(yt_rsc_6_29_d),
      .wadr(yt_rsc_6_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_6_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_229_4_32_16_16_32_1_gen yt_rsc_6_30_i
      (
      .clkr_en(yt_rsc_6_30_clkr_en),
      .clkw_en(yt_rsc_6_30_clkw_en),
      .q(yt_rsc_6_30_q),
      .radr(yt_rsc_6_30_radr),
      .we(yt_rsc_6_30_we),
      .d(yt_rsc_6_30_d),
      .wadr(yt_rsc_6_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_6_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_230_4_32_16_16_32_1_gen yt_rsc_6_31_i
      (
      .clkr_en(yt_rsc_6_31_clkr_en),
      .clkw_en(yt_rsc_6_31_clkw_en),
      .q(yt_rsc_6_31_q),
      .radr(yt_rsc_6_31_radr),
      .we(yt_rsc_6_31_we),
      .d(yt_rsc_6_31_d),
      .wadr(yt_rsc_6_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_6_16_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_6_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_6_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_6_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_231_4_32_16_16_32_1_gen yt_rsc_7_0_i
      (
      .clkr_en(yt_rsc_7_0_clkr_en),
      .clkw_en(yt_rsc_7_0_clkw_en),
      .q(yt_rsc_7_0_q),
      .radr(yt_rsc_7_0_radr),
      .we(yt_rsc_7_0_we),
      .d(yt_rsc_7_0_d),
      .wadr(yt_rsc_7_0_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_7_0_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_232_4_32_16_16_32_1_gen yt_rsc_7_1_i
      (
      .clkr_en(yt_rsc_7_1_clkr_en),
      .clkw_en(yt_rsc_7_1_clkw_en),
      .q(yt_rsc_7_1_q),
      .radr(yt_rsc_7_1_radr),
      .we(yt_rsc_7_1_we),
      .d(yt_rsc_7_1_d),
      .wadr(yt_rsc_7_1_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_7_1_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_233_4_32_16_16_32_1_gen yt_rsc_7_2_i
      (
      .clkr_en(yt_rsc_7_2_clkr_en),
      .clkw_en(yt_rsc_7_2_clkw_en),
      .q(yt_rsc_7_2_q),
      .radr(yt_rsc_7_2_radr),
      .we(yt_rsc_7_2_we),
      .d(yt_rsc_7_2_d),
      .wadr(yt_rsc_7_2_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_7_2_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_234_4_32_16_16_32_1_gen yt_rsc_7_3_i
      (
      .clkr_en(yt_rsc_7_3_clkr_en),
      .clkw_en(yt_rsc_7_3_clkw_en),
      .q(yt_rsc_7_3_q),
      .radr(yt_rsc_7_3_radr),
      .we(yt_rsc_7_3_we),
      .d(yt_rsc_7_3_d),
      .wadr(yt_rsc_7_3_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_7_3_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_235_4_32_16_16_32_1_gen yt_rsc_7_4_i
      (
      .clkr_en(yt_rsc_7_4_clkr_en),
      .clkw_en(yt_rsc_7_4_clkw_en),
      .q(yt_rsc_7_4_q),
      .radr(yt_rsc_7_4_radr),
      .we(yt_rsc_7_4_we),
      .d(yt_rsc_7_4_d),
      .wadr(yt_rsc_7_4_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_7_4_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_236_4_32_16_16_32_1_gen yt_rsc_7_5_i
      (
      .clkr_en(yt_rsc_7_5_clkr_en),
      .clkw_en(yt_rsc_7_5_clkw_en),
      .q(yt_rsc_7_5_q),
      .radr(yt_rsc_7_5_radr),
      .we(yt_rsc_7_5_we),
      .d(yt_rsc_7_5_d),
      .wadr(yt_rsc_7_5_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_7_5_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_237_4_32_16_16_32_1_gen yt_rsc_7_6_i
      (
      .clkr_en(yt_rsc_7_6_clkr_en),
      .clkw_en(yt_rsc_7_6_clkw_en),
      .q(yt_rsc_7_6_q),
      .radr(yt_rsc_7_6_radr),
      .we(yt_rsc_7_6_we),
      .d(yt_rsc_7_6_d),
      .wadr(yt_rsc_7_6_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_7_6_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_238_4_32_16_16_32_1_gen yt_rsc_7_7_i
      (
      .clkr_en(yt_rsc_7_7_clkr_en),
      .clkw_en(yt_rsc_7_7_clkw_en),
      .q(yt_rsc_7_7_q),
      .radr(yt_rsc_7_7_radr),
      .we(yt_rsc_7_7_we),
      .d(yt_rsc_7_7_d),
      .wadr(yt_rsc_7_7_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_7_7_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_239_4_32_16_16_32_1_gen yt_rsc_7_8_i
      (
      .clkr_en(yt_rsc_7_8_clkr_en),
      .clkw_en(yt_rsc_7_8_clkw_en),
      .q(yt_rsc_7_8_q),
      .radr(yt_rsc_7_8_radr),
      .we(yt_rsc_7_8_we),
      .d(yt_rsc_7_8_d),
      .wadr(yt_rsc_7_8_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_7_8_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_240_4_32_16_16_32_1_gen yt_rsc_7_9_i
      (
      .clkr_en(yt_rsc_7_9_clkr_en),
      .clkw_en(yt_rsc_7_9_clkw_en),
      .q(yt_rsc_7_9_q),
      .radr(yt_rsc_7_9_radr),
      .we(yt_rsc_7_9_we),
      .d(yt_rsc_7_9_d),
      .wadr(yt_rsc_7_9_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_7_9_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_241_4_32_16_16_32_1_gen yt_rsc_7_10_i
      (
      .clkr_en(yt_rsc_7_10_clkr_en),
      .clkw_en(yt_rsc_7_10_clkw_en),
      .q(yt_rsc_7_10_q),
      .radr(yt_rsc_7_10_radr),
      .we(yt_rsc_7_10_we),
      .d(yt_rsc_7_10_d),
      .wadr(yt_rsc_7_10_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_7_10_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_242_4_32_16_16_32_1_gen yt_rsc_7_11_i
      (
      .clkr_en(yt_rsc_7_11_clkr_en),
      .clkw_en(yt_rsc_7_11_clkw_en),
      .q(yt_rsc_7_11_q),
      .radr(yt_rsc_7_11_radr),
      .we(yt_rsc_7_11_we),
      .d(yt_rsc_7_11_d),
      .wadr(yt_rsc_7_11_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_7_11_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_243_4_32_16_16_32_1_gen yt_rsc_7_12_i
      (
      .clkr_en(yt_rsc_7_12_clkr_en),
      .clkw_en(yt_rsc_7_12_clkw_en),
      .q(yt_rsc_7_12_q),
      .radr(yt_rsc_7_12_radr),
      .we(yt_rsc_7_12_we),
      .d(yt_rsc_7_12_d),
      .wadr(yt_rsc_7_12_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_7_12_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_244_4_32_16_16_32_1_gen yt_rsc_7_13_i
      (
      .clkr_en(yt_rsc_7_13_clkr_en),
      .clkw_en(yt_rsc_7_13_clkw_en),
      .q(yt_rsc_7_13_q),
      .radr(yt_rsc_7_13_radr),
      .we(yt_rsc_7_13_we),
      .d(yt_rsc_7_13_d),
      .wadr(yt_rsc_7_13_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_7_13_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_245_4_32_16_16_32_1_gen yt_rsc_7_14_i
      (
      .clkr_en(yt_rsc_7_14_clkr_en),
      .clkw_en(yt_rsc_7_14_clkw_en),
      .q(yt_rsc_7_14_q),
      .radr(yt_rsc_7_14_radr),
      .we(yt_rsc_7_14_we),
      .d(yt_rsc_7_14_d),
      .wadr(yt_rsc_7_14_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_7_14_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_246_4_32_16_16_32_1_gen yt_rsc_7_15_i
      (
      .clkr_en(yt_rsc_7_15_clkr_en),
      .clkw_en(yt_rsc_7_15_clkw_en),
      .q(yt_rsc_7_15_q),
      .radr(yt_rsc_7_15_radr),
      .we(yt_rsc_7_15_we),
      .d(yt_rsc_7_15_d),
      .wadr(yt_rsc_7_15_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_0_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_7_15_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_7_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_247_4_32_16_16_32_1_gen yt_rsc_7_16_i
      (
      .clkr_en(yt_rsc_7_16_clkr_en),
      .clkw_en(yt_rsc_7_16_clkw_en),
      .q(yt_rsc_7_16_q),
      .radr(yt_rsc_7_16_radr),
      .we(yt_rsc_7_16_we),
      .d(yt_rsc_7_16_d),
      .wadr(yt_rsc_7_16_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_0_i_d_d_iff),
      .q_d(yt_rsc_7_16_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_248_4_32_16_16_32_1_gen yt_rsc_7_17_i
      (
      .clkr_en(yt_rsc_7_17_clkr_en),
      .clkw_en(yt_rsc_7_17_clkw_en),
      .q(yt_rsc_7_17_q),
      .radr(yt_rsc_7_17_radr),
      .we(yt_rsc_7_17_we),
      .d(yt_rsc_7_17_d),
      .wadr(yt_rsc_7_17_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_1_i_d_d_iff),
      .q_d(yt_rsc_7_17_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_249_4_32_16_16_32_1_gen yt_rsc_7_18_i
      (
      .clkr_en(yt_rsc_7_18_clkr_en),
      .clkw_en(yt_rsc_7_18_clkw_en),
      .q(yt_rsc_7_18_q),
      .radr(yt_rsc_7_18_radr),
      .we(yt_rsc_7_18_we),
      .d(yt_rsc_7_18_d),
      .wadr(yt_rsc_7_18_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_2_i_d_d_iff),
      .q_d(yt_rsc_7_18_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_2_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_250_4_32_16_16_32_1_gen yt_rsc_7_19_i
      (
      .clkr_en(yt_rsc_7_19_clkr_en),
      .clkw_en(yt_rsc_7_19_clkw_en),
      .q(yt_rsc_7_19_q),
      .radr(yt_rsc_7_19_radr),
      .we(yt_rsc_7_19_we),
      .d(yt_rsc_7_19_d),
      .wadr(yt_rsc_7_19_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_3_i_d_d_iff),
      .q_d(yt_rsc_7_19_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_251_4_32_16_16_32_1_gen yt_rsc_7_20_i
      (
      .clkr_en(yt_rsc_7_20_clkr_en),
      .clkw_en(yt_rsc_7_20_clkw_en),
      .q(yt_rsc_7_20_q),
      .radr(yt_rsc_7_20_radr),
      .we(yt_rsc_7_20_we),
      .d(yt_rsc_7_20_d),
      .wadr(yt_rsc_7_20_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_4_i_d_d_iff),
      .q_d(yt_rsc_7_20_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_252_4_32_16_16_32_1_gen yt_rsc_7_21_i
      (
      .clkr_en(yt_rsc_7_21_clkr_en),
      .clkw_en(yt_rsc_7_21_clkw_en),
      .q(yt_rsc_7_21_q),
      .radr(yt_rsc_7_21_radr),
      .we(yt_rsc_7_21_we),
      .d(yt_rsc_7_21_d),
      .wadr(yt_rsc_7_21_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_5_i_d_d_iff),
      .q_d(yt_rsc_7_21_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_253_4_32_16_16_32_1_gen yt_rsc_7_22_i
      (
      .clkr_en(yt_rsc_7_22_clkr_en),
      .clkw_en(yt_rsc_7_22_clkw_en),
      .q(yt_rsc_7_22_q),
      .radr(yt_rsc_7_22_radr),
      .we(yt_rsc_7_22_we),
      .d(yt_rsc_7_22_d),
      .wadr(yt_rsc_7_22_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_6_i_d_d_iff),
      .q_d(yt_rsc_7_22_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_254_4_32_16_16_32_1_gen yt_rsc_7_23_i
      (
      .clkr_en(yt_rsc_7_23_clkr_en),
      .clkw_en(yt_rsc_7_23_clkw_en),
      .q(yt_rsc_7_23_q),
      .radr(yt_rsc_7_23_radr),
      .we(yt_rsc_7_23_we),
      .d(yt_rsc_7_23_d),
      .wadr(yt_rsc_7_23_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_7_i_d_d_iff),
      .q_d(yt_rsc_7_23_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_0_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_255_4_32_16_16_32_1_gen yt_rsc_7_24_i
      (
      .clkr_en(yt_rsc_7_24_clkr_en),
      .clkw_en(yt_rsc_7_24_clkw_en),
      .q(yt_rsc_7_24_q),
      .radr(yt_rsc_7_24_radr),
      .we(yt_rsc_7_24_we),
      .d(yt_rsc_7_24_d),
      .wadr(yt_rsc_7_24_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_8_i_d_d_iff),
      .q_d(yt_rsc_7_24_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_1_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_256_4_32_16_16_32_1_gen yt_rsc_7_25_i
      (
      .clkr_en(yt_rsc_7_25_clkr_en),
      .clkw_en(yt_rsc_7_25_clkw_en),
      .q(yt_rsc_7_25_q),
      .radr(yt_rsc_7_25_radr),
      .we(yt_rsc_7_25_we),
      .d(yt_rsc_7_25_d),
      .wadr(yt_rsc_7_25_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_9_i_d_d_iff),
      .q_d(yt_rsc_7_25_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_9_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_257_4_32_16_16_32_1_gen yt_rsc_7_26_i
      (
      .clkr_en(yt_rsc_7_26_clkr_en),
      .clkw_en(yt_rsc_7_26_clkw_en),
      .q(yt_rsc_7_26_q),
      .radr(yt_rsc_7_26_radr),
      .we(yt_rsc_7_26_we),
      .d(yt_rsc_7_26_d),
      .wadr(yt_rsc_7_26_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_10_i_d_d_iff),
      .q_d(yt_rsc_7_26_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_10_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_258_4_32_16_16_32_1_gen yt_rsc_7_27_i
      (
      .clkr_en(yt_rsc_7_27_clkr_en),
      .clkw_en(yt_rsc_7_27_clkw_en),
      .q(yt_rsc_7_27_q),
      .radr(yt_rsc_7_27_radr),
      .we(yt_rsc_7_27_we),
      .d(yt_rsc_7_27_d),
      .wadr(yt_rsc_7_27_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_11_i_d_d_iff),
      .q_d(yt_rsc_7_27_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_11_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_259_4_32_16_16_32_1_gen yt_rsc_7_28_i
      (
      .clkr_en(yt_rsc_7_28_clkr_en),
      .clkw_en(yt_rsc_7_28_clkw_en),
      .q(yt_rsc_7_28_q),
      .radr(yt_rsc_7_28_radr),
      .we(yt_rsc_7_28_we),
      .d(yt_rsc_7_28_d),
      .wadr(yt_rsc_7_28_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_12_i_d_d_iff),
      .q_d(yt_rsc_7_28_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_3_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_260_4_32_16_16_32_1_gen yt_rsc_7_29_i
      (
      .clkr_en(yt_rsc_7_29_clkr_en),
      .clkw_en(yt_rsc_7_29_clkw_en),
      .q(yt_rsc_7_29_q),
      .radr(yt_rsc_7_29_radr),
      .we(yt_rsc_7_29_we),
      .d(yt_rsc_7_29_d),
      .wadr(yt_rsc_7_29_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_13_i_d_d_iff),
      .q_d(yt_rsc_7_29_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_4_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_261_4_32_16_16_32_1_gen yt_rsc_7_30_i
      (
      .clkr_en(yt_rsc_7_30_clkr_en),
      .clkw_en(yt_rsc_7_30_clkw_en),
      .q(yt_rsc_7_30_q),
      .radr(yt_rsc_7_30_radr),
      .we(yt_rsc_7_30_we),
      .d(yt_rsc_7_30_d),
      .wadr(yt_rsc_7_30_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_14_i_d_d_iff),
      .q_d(yt_rsc_7_30_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_5_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_1R1W_RBW_DUAL_rwport_en_262_4_32_16_16_32_1_gen yt_rsc_7_31_i
      (
      .clkr_en(yt_rsc_7_31_clkr_en),
      .clkw_en(yt_rsc_7_31_clkw_en),
      .q(yt_rsc_7_31_q),
      .radr(yt_rsc_7_31_radr),
      .we(yt_rsc_7_31_we),
      .d(yt_rsc_7_31_d),
      .wadr(yt_rsc_7_31_wadr),
      .clkr(clk),
      .clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .clkw_en_d(yt_rsc_7_16_i_clkr_en_d),
      .d_d(yt_rsc_4_15_i_d_d_iff),
      .q_d(yt_rsc_7_31_i_q_d),
      .radr_d(yt_rsc_0_0_i_radr_d_iff),
      .wadr_d(yt_rsc_4_6_i_wadr_d_iff),
      .we_d(yt_rsc_7_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(yt_rsc_7_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_263_4_32_16_16_32_1_gen xt_rsc_0_0_i
      (
      .qa(xt_rsc_0_0_qa),
      .wea(xt_rsc_0_0_wea),
      .da(xt_rsc_0_0_da),
      .adra(xt_rsc_0_0_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_0_0_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_264_4_32_16_16_32_1_gen xt_rsc_0_1_i
      (
      .qa(xt_rsc_0_1_qa),
      .wea(xt_rsc_0_1_wea),
      .da(xt_rsc_0_1_da),
      .adra(xt_rsc_0_1_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_0_1_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_265_4_32_16_16_32_1_gen xt_rsc_0_2_i
      (
      .qa(xt_rsc_0_2_qa),
      .wea(xt_rsc_0_2_wea),
      .da(xt_rsc_0_2_da),
      .adra(xt_rsc_0_2_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_0_2_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_266_4_32_16_16_32_1_gen xt_rsc_0_3_i
      (
      .qa(xt_rsc_0_3_qa),
      .wea(xt_rsc_0_3_wea),
      .da(xt_rsc_0_3_da),
      .adra(xt_rsc_0_3_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_0_3_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_267_4_32_16_16_32_1_gen xt_rsc_0_4_i
      (
      .qa(xt_rsc_0_4_qa),
      .wea(xt_rsc_0_4_wea),
      .da(xt_rsc_0_4_da),
      .adra(xt_rsc_0_4_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_0_4_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_268_4_32_16_16_32_1_gen xt_rsc_0_5_i
      (
      .qa(xt_rsc_0_5_qa),
      .wea(xt_rsc_0_5_wea),
      .da(xt_rsc_0_5_da),
      .adra(xt_rsc_0_5_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_0_5_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_269_4_32_16_16_32_1_gen xt_rsc_0_6_i
      (
      .qa(xt_rsc_0_6_qa),
      .wea(xt_rsc_0_6_wea),
      .da(xt_rsc_0_6_da),
      .adra(xt_rsc_0_6_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_0_6_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_270_4_32_16_16_32_1_gen xt_rsc_0_7_i
      (
      .qa(xt_rsc_0_7_qa),
      .wea(xt_rsc_0_7_wea),
      .da(xt_rsc_0_7_da),
      .adra(xt_rsc_0_7_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_0_7_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_271_4_32_16_16_32_1_gen xt_rsc_0_8_i
      (
      .qa(xt_rsc_0_8_qa),
      .wea(xt_rsc_0_8_wea),
      .da(xt_rsc_0_8_da),
      .adra(xt_rsc_0_8_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_0_8_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_272_4_32_16_16_32_1_gen xt_rsc_0_9_i
      (
      .qa(xt_rsc_0_9_qa),
      .wea(xt_rsc_0_9_wea),
      .da(xt_rsc_0_9_da),
      .adra(xt_rsc_0_9_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_0_9_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_273_4_32_16_16_32_1_gen xt_rsc_0_10_i
      (
      .qa(xt_rsc_0_10_qa),
      .wea(xt_rsc_0_10_wea),
      .da(xt_rsc_0_10_da),
      .adra(xt_rsc_0_10_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_0_10_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_274_4_32_16_16_32_1_gen xt_rsc_0_11_i
      (
      .qa(xt_rsc_0_11_qa),
      .wea(xt_rsc_0_11_wea),
      .da(xt_rsc_0_11_da),
      .adra(xt_rsc_0_11_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_0_11_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_275_4_32_16_16_32_1_gen xt_rsc_0_12_i
      (
      .qa(xt_rsc_0_12_qa),
      .wea(xt_rsc_0_12_wea),
      .da(xt_rsc_0_12_da),
      .adra(xt_rsc_0_12_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_0_12_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_276_4_32_16_16_32_1_gen xt_rsc_0_13_i
      (
      .qa(xt_rsc_0_13_qa),
      .wea(xt_rsc_0_13_wea),
      .da(xt_rsc_0_13_da),
      .adra(xt_rsc_0_13_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_0_13_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_277_4_32_16_16_32_1_gen xt_rsc_0_14_i
      (
      .qa(xt_rsc_0_14_qa),
      .wea(xt_rsc_0_14_wea),
      .da(xt_rsc_0_14_da),
      .adra(xt_rsc_0_14_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_0_14_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_278_4_32_16_16_32_1_gen xt_rsc_0_15_i
      (
      .qa(xt_rsc_0_15_qa),
      .wea(xt_rsc_0_15_wea),
      .da(xt_rsc_0_15_da),
      .adra(xt_rsc_0_15_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_0_15_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_279_4_32_16_16_32_1_gen xt_rsc_0_16_i
      (
      .qa(xt_rsc_0_16_qa),
      .wea(xt_rsc_0_16_wea),
      .da(xt_rsc_0_16_da),
      .adra(xt_rsc_0_16_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_0_16_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_280_4_32_16_16_32_1_gen xt_rsc_0_17_i
      (
      .qa(xt_rsc_0_17_qa),
      .wea(xt_rsc_0_17_wea),
      .da(xt_rsc_0_17_da),
      .adra(xt_rsc_0_17_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_0_17_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_281_4_32_16_16_32_1_gen xt_rsc_0_18_i
      (
      .qa(xt_rsc_0_18_qa),
      .wea(xt_rsc_0_18_wea),
      .da(xt_rsc_0_18_da),
      .adra(xt_rsc_0_18_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_0_18_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_282_4_32_16_16_32_1_gen xt_rsc_0_19_i
      (
      .qa(xt_rsc_0_19_qa),
      .wea(xt_rsc_0_19_wea),
      .da(xt_rsc_0_19_da),
      .adra(xt_rsc_0_19_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_0_19_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_283_4_32_16_16_32_1_gen xt_rsc_0_20_i
      (
      .qa(xt_rsc_0_20_qa),
      .wea(xt_rsc_0_20_wea),
      .da(xt_rsc_0_20_da),
      .adra(xt_rsc_0_20_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_0_20_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_284_4_32_16_16_32_1_gen xt_rsc_0_21_i
      (
      .qa(xt_rsc_0_21_qa),
      .wea(xt_rsc_0_21_wea),
      .da(xt_rsc_0_21_da),
      .adra(xt_rsc_0_21_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_0_21_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_285_4_32_16_16_32_1_gen xt_rsc_0_22_i
      (
      .qa(xt_rsc_0_22_qa),
      .wea(xt_rsc_0_22_wea),
      .da(xt_rsc_0_22_da),
      .adra(xt_rsc_0_22_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_0_22_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_286_4_32_16_16_32_1_gen xt_rsc_0_23_i
      (
      .qa(xt_rsc_0_23_qa),
      .wea(xt_rsc_0_23_wea),
      .da(xt_rsc_0_23_da),
      .adra(xt_rsc_0_23_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_0_23_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_287_4_32_16_16_32_1_gen xt_rsc_0_24_i
      (
      .qa(xt_rsc_0_24_qa),
      .wea(xt_rsc_0_24_wea),
      .da(xt_rsc_0_24_da),
      .adra(xt_rsc_0_24_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_0_24_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_288_4_32_16_16_32_1_gen xt_rsc_0_25_i
      (
      .qa(xt_rsc_0_25_qa),
      .wea(xt_rsc_0_25_wea),
      .da(xt_rsc_0_25_da),
      .adra(xt_rsc_0_25_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_0_25_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_289_4_32_16_16_32_1_gen xt_rsc_0_26_i
      (
      .qa(xt_rsc_0_26_qa),
      .wea(xt_rsc_0_26_wea),
      .da(xt_rsc_0_26_da),
      .adra(xt_rsc_0_26_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_0_26_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_290_4_32_16_16_32_1_gen xt_rsc_0_27_i
      (
      .qa(xt_rsc_0_27_qa),
      .wea(xt_rsc_0_27_wea),
      .da(xt_rsc_0_27_da),
      .adra(xt_rsc_0_27_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_0_27_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_291_4_32_16_16_32_1_gen xt_rsc_0_28_i
      (
      .qa(xt_rsc_0_28_qa),
      .wea(xt_rsc_0_28_wea),
      .da(xt_rsc_0_28_da),
      .adra(xt_rsc_0_28_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_0_28_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_292_4_32_16_16_32_1_gen xt_rsc_0_29_i
      (
      .qa(xt_rsc_0_29_qa),
      .wea(xt_rsc_0_29_wea),
      .da(xt_rsc_0_29_da),
      .adra(xt_rsc_0_29_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_0_29_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_293_4_32_16_16_32_1_gen xt_rsc_0_30_i
      (
      .qa(xt_rsc_0_30_qa),
      .wea(xt_rsc_0_30_wea),
      .da(xt_rsc_0_30_da),
      .adra(xt_rsc_0_30_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_0_30_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_294_4_32_16_16_32_1_gen xt_rsc_0_31_i
      (
      .qa(xt_rsc_0_31_qa),
      .wea(xt_rsc_0_31_wea),
      .da(xt_rsc_0_31_da),
      .adra(xt_rsc_0_31_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_0_31_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_295_4_32_16_16_32_1_gen xt_rsc_1_0_i
      (
      .qa(xt_rsc_1_0_qa),
      .wea(xt_rsc_1_0_wea),
      .da(xt_rsc_1_0_da),
      .adra(xt_rsc_1_0_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_1_0_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_296_4_32_16_16_32_1_gen xt_rsc_1_1_i
      (
      .qa(xt_rsc_1_1_qa),
      .wea(xt_rsc_1_1_wea),
      .da(xt_rsc_1_1_da),
      .adra(xt_rsc_1_1_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_1_1_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_297_4_32_16_16_32_1_gen xt_rsc_1_2_i
      (
      .qa(xt_rsc_1_2_qa),
      .wea(xt_rsc_1_2_wea),
      .da(xt_rsc_1_2_da),
      .adra(xt_rsc_1_2_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_1_2_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_298_4_32_16_16_32_1_gen xt_rsc_1_3_i
      (
      .qa(xt_rsc_1_3_qa),
      .wea(xt_rsc_1_3_wea),
      .da(xt_rsc_1_3_da),
      .adra(xt_rsc_1_3_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_1_3_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_299_4_32_16_16_32_1_gen xt_rsc_1_4_i
      (
      .qa(xt_rsc_1_4_qa),
      .wea(xt_rsc_1_4_wea),
      .da(xt_rsc_1_4_da),
      .adra(xt_rsc_1_4_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_1_4_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_300_4_32_16_16_32_1_gen xt_rsc_1_5_i
      (
      .qa(xt_rsc_1_5_qa),
      .wea(xt_rsc_1_5_wea),
      .da(xt_rsc_1_5_da),
      .adra(xt_rsc_1_5_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_1_5_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_301_4_32_16_16_32_1_gen xt_rsc_1_6_i
      (
      .qa(xt_rsc_1_6_qa),
      .wea(xt_rsc_1_6_wea),
      .da(xt_rsc_1_6_da),
      .adra(xt_rsc_1_6_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_1_6_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_302_4_32_16_16_32_1_gen xt_rsc_1_7_i
      (
      .qa(xt_rsc_1_7_qa),
      .wea(xt_rsc_1_7_wea),
      .da(xt_rsc_1_7_da),
      .adra(xt_rsc_1_7_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_1_7_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_303_4_32_16_16_32_1_gen xt_rsc_1_8_i
      (
      .qa(xt_rsc_1_8_qa),
      .wea(xt_rsc_1_8_wea),
      .da(xt_rsc_1_8_da),
      .adra(xt_rsc_1_8_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_1_8_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_304_4_32_16_16_32_1_gen xt_rsc_1_9_i
      (
      .qa(xt_rsc_1_9_qa),
      .wea(xt_rsc_1_9_wea),
      .da(xt_rsc_1_9_da),
      .adra(xt_rsc_1_9_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_1_9_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_305_4_32_16_16_32_1_gen xt_rsc_1_10_i
      (
      .qa(xt_rsc_1_10_qa),
      .wea(xt_rsc_1_10_wea),
      .da(xt_rsc_1_10_da),
      .adra(xt_rsc_1_10_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_1_10_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_306_4_32_16_16_32_1_gen xt_rsc_1_11_i
      (
      .qa(xt_rsc_1_11_qa),
      .wea(xt_rsc_1_11_wea),
      .da(xt_rsc_1_11_da),
      .adra(xt_rsc_1_11_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_1_11_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_307_4_32_16_16_32_1_gen xt_rsc_1_12_i
      (
      .qa(xt_rsc_1_12_qa),
      .wea(xt_rsc_1_12_wea),
      .da(xt_rsc_1_12_da),
      .adra(xt_rsc_1_12_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_1_12_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_308_4_32_16_16_32_1_gen xt_rsc_1_13_i
      (
      .qa(xt_rsc_1_13_qa),
      .wea(xt_rsc_1_13_wea),
      .da(xt_rsc_1_13_da),
      .adra(xt_rsc_1_13_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_1_13_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_309_4_32_16_16_32_1_gen xt_rsc_1_14_i
      (
      .qa(xt_rsc_1_14_qa),
      .wea(xt_rsc_1_14_wea),
      .da(xt_rsc_1_14_da),
      .adra(xt_rsc_1_14_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_1_14_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_310_4_32_16_16_32_1_gen xt_rsc_1_15_i
      (
      .qa(xt_rsc_1_15_qa),
      .wea(xt_rsc_1_15_wea),
      .da(xt_rsc_1_15_da),
      .adra(xt_rsc_1_15_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_1_15_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_311_4_32_16_16_32_1_gen xt_rsc_1_16_i
      (
      .qa(xt_rsc_1_16_qa),
      .wea(xt_rsc_1_16_wea),
      .da(xt_rsc_1_16_da),
      .adra(xt_rsc_1_16_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_1_16_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_312_4_32_16_16_32_1_gen xt_rsc_1_17_i
      (
      .qa(xt_rsc_1_17_qa),
      .wea(xt_rsc_1_17_wea),
      .da(xt_rsc_1_17_da),
      .adra(xt_rsc_1_17_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_1_17_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_313_4_32_16_16_32_1_gen xt_rsc_1_18_i
      (
      .qa(xt_rsc_1_18_qa),
      .wea(xt_rsc_1_18_wea),
      .da(xt_rsc_1_18_da),
      .adra(xt_rsc_1_18_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_1_18_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_314_4_32_16_16_32_1_gen xt_rsc_1_19_i
      (
      .qa(xt_rsc_1_19_qa),
      .wea(xt_rsc_1_19_wea),
      .da(xt_rsc_1_19_da),
      .adra(xt_rsc_1_19_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_1_19_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_315_4_32_16_16_32_1_gen xt_rsc_1_20_i
      (
      .qa(xt_rsc_1_20_qa),
      .wea(xt_rsc_1_20_wea),
      .da(xt_rsc_1_20_da),
      .adra(xt_rsc_1_20_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_1_20_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_316_4_32_16_16_32_1_gen xt_rsc_1_21_i
      (
      .qa(xt_rsc_1_21_qa),
      .wea(xt_rsc_1_21_wea),
      .da(xt_rsc_1_21_da),
      .adra(xt_rsc_1_21_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_1_21_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_317_4_32_16_16_32_1_gen xt_rsc_1_22_i
      (
      .qa(xt_rsc_1_22_qa),
      .wea(xt_rsc_1_22_wea),
      .da(xt_rsc_1_22_da),
      .adra(xt_rsc_1_22_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_1_22_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_318_4_32_16_16_32_1_gen xt_rsc_1_23_i
      (
      .qa(xt_rsc_1_23_qa),
      .wea(xt_rsc_1_23_wea),
      .da(xt_rsc_1_23_da),
      .adra(xt_rsc_1_23_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_1_23_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_319_4_32_16_16_32_1_gen xt_rsc_1_24_i
      (
      .qa(xt_rsc_1_24_qa),
      .wea(xt_rsc_1_24_wea),
      .da(xt_rsc_1_24_da),
      .adra(xt_rsc_1_24_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_1_24_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_320_4_32_16_16_32_1_gen xt_rsc_1_25_i
      (
      .qa(xt_rsc_1_25_qa),
      .wea(xt_rsc_1_25_wea),
      .da(xt_rsc_1_25_da),
      .adra(xt_rsc_1_25_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_1_25_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_321_4_32_16_16_32_1_gen xt_rsc_1_26_i
      (
      .qa(xt_rsc_1_26_qa),
      .wea(xt_rsc_1_26_wea),
      .da(xt_rsc_1_26_da),
      .adra(xt_rsc_1_26_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_1_26_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_322_4_32_16_16_32_1_gen xt_rsc_1_27_i
      (
      .qa(xt_rsc_1_27_qa),
      .wea(xt_rsc_1_27_wea),
      .da(xt_rsc_1_27_da),
      .adra(xt_rsc_1_27_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_1_27_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_323_4_32_16_16_32_1_gen xt_rsc_1_28_i
      (
      .qa(xt_rsc_1_28_qa),
      .wea(xt_rsc_1_28_wea),
      .da(xt_rsc_1_28_da),
      .adra(xt_rsc_1_28_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_1_28_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_324_4_32_16_16_32_1_gen xt_rsc_1_29_i
      (
      .qa(xt_rsc_1_29_qa),
      .wea(xt_rsc_1_29_wea),
      .da(xt_rsc_1_29_da),
      .adra(xt_rsc_1_29_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_1_29_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_325_4_32_16_16_32_1_gen xt_rsc_1_30_i
      (
      .qa(xt_rsc_1_30_qa),
      .wea(xt_rsc_1_30_wea),
      .da(xt_rsc_1_30_da),
      .adra(xt_rsc_1_30_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_1_30_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_326_4_32_16_16_32_1_gen xt_rsc_1_31_i
      (
      .qa(xt_rsc_1_31_qa),
      .wea(xt_rsc_1_31_wea),
      .da(xt_rsc_1_31_da),
      .adra(xt_rsc_1_31_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_1_31_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_327_4_32_16_16_32_1_gen xt_rsc_2_0_i
      (
      .qa(xt_rsc_2_0_qa),
      .wea(xt_rsc_2_0_wea),
      .da(xt_rsc_2_0_da),
      .adra(xt_rsc_2_0_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_2_0_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_328_4_32_16_16_32_1_gen xt_rsc_2_1_i
      (
      .qa(xt_rsc_2_1_qa),
      .wea(xt_rsc_2_1_wea),
      .da(xt_rsc_2_1_da),
      .adra(xt_rsc_2_1_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_2_1_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_329_4_32_16_16_32_1_gen xt_rsc_2_2_i
      (
      .qa(xt_rsc_2_2_qa),
      .wea(xt_rsc_2_2_wea),
      .da(xt_rsc_2_2_da),
      .adra(xt_rsc_2_2_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_2_2_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_330_4_32_16_16_32_1_gen xt_rsc_2_3_i
      (
      .qa(xt_rsc_2_3_qa),
      .wea(xt_rsc_2_3_wea),
      .da(xt_rsc_2_3_da),
      .adra(xt_rsc_2_3_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_2_3_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_331_4_32_16_16_32_1_gen xt_rsc_2_4_i
      (
      .qa(xt_rsc_2_4_qa),
      .wea(xt_rsc_2_4_wea),
      .da(xt_rsc_2_4_da),
      .adra(xt_rsc_2_4_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_2_4_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_332_4_32_16_16_32_1_gen xt_rsc_2_5_i
      (
      .qa(xt_rsc_2_5_qa),
      .wea(xt_rsc_2_5_wea),
      .da(xt_rsc_2_5_da),
      .adra(xt_rsc_2_5_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_2_5_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_333_4_32_16_16_32_1_gen xt_rsc_2_6_i
      (
      .qa(xt_rsc_2_6_qa),
      .wea(xt_rsc_2_6_wea),
      .da(xt_rsc_2_6_da),
      .adra(xt_rsc_2_6_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_2_6_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_334_4_32_16_16_32_1_gen xt_rsc_2_7_i
      (
      .qa(xt_rsc_2_7_qa),
      .wea(xt_rsc_2_7_wea),
      .da(xt_rsc_2_7_da),
      .adra(xt_rsc_2_7_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_2_7_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_335_4_32_16_16_32_1_gen xt_rsc_2_8_i
      (
      .qa(xt_rsc_2_8_qa),
      .wea(xt_rsc_2_8_wea),
      .da(xt_rsc_2_8_da),
      .adra(xt_rsc_2_8_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_2_8_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_336_4_32_16_16_32_1_gen xt_rsc_2_9_i
      (
      .qa(xt_rsc_2_9_qa),
      .wea(xt_rsc_2_9_wea),
      .da(xt_rsc_2_9_da),
      .adra(xt_rsc_2_9_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_2_9_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_337_4_32_16_16_32_1_gen xt_rsc_2_10_i
      (
      .qa(xt_rsc_2_10_qa),
      .wea(xt_rsc_2_10_wea),
      .da(xt_rsc_2_10_da),
      .adra(xt_rsc_2_10_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_2_10_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_338_4_32_16_16_32_1_gen xt_rsc_2_11_i
      (
      .qa(xt_rsc_2_11_qa),
      .wea(xt_rsc_2_11_wea),
      .da(xt_rsc_2_11_da),
      .adra(xt_rsc_2_11_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_2_11_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_339_4_32_16_16_32_1_gen xt_rsc_2_12_i
      (
      .qa(xt_rsc_2_12_qa),
      .wea(xt_rsc_2_12_wea),
      .da(xt_rsc_2_12_da),
      .adra(xt_rsc_2_12_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_2_12_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_340_4_32_16_16_32_1_gen xt_rsc_2_13_i
      (
      .qa(xt_rsc_2_13_qa),
      .wea(xt_rsc_2_13_wea),
      .da(xt_rsc_2_13_da),
      .adra(xt_rsc_2_13_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_2_13_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_341_4_32_16_16_32_1_gen xt_rsc_2_14_i
      (
      .qa(xt_rsc_2_14_qa),
      .wea(xt_rsc_2_14_wea),
      .da(xt_rsc_2_14_da),
      .adra(xt_rsc_2_14_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_2_14_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_342_4_32_16_16_32_1_gen xt_rsc_2_15_i
      (
      .qa(xt_rsc_2_15_qa),
      .wea(xt_rsc_2_15_wea),
      .da(xt_rsc_2_15_da),
      .adra(xt_rsc_2_15_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_2_15_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_343_4_32_16_16_32_1_gen xt_rsc_2_16_i
      (
      .qa(xt_rsc_2_16_qa),
      .wea(xt_rsc_2_16_wea),
      .da(xt_rsc_2_16_da),
      .adra(xt_rsc_2_16_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_2_16_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_344_4_32_16_16_32_1_gen xt_rsc_2_17_i
      (
      .qa(xt_rsc_2_17_qa),
      .wea(xt_rsc_2_17_wea),
      .da(xt_rsc_2_17_da),
      .adra(xt_rsc_2_17_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_2_17_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_345_4_32_16_16_32_1_gen xt_rsc_2_18_i
      (
      .qa(xt_rsc_2_18_qa),
      .wea(xt_rsc_2_18_wea),
      .da(xt_rsc_2_18_da),
      .adra(xt_rsc_2_18_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_2_18_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_346_4_32_16_16_32_1_gen xt_rsc_2_19_i
      (
      .qa(xt_rsc_2_19_qa),
      .wea(xt_rsc_2_19_wea),
      .da(xt_rsc_2_19_da),
      .adra(xt_rsc_2_19_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_2_19_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_347_4_32_16_16_32_1_gen xt_rsc_2_20_i
      (
      .qa(xt_rsc_2_20_qa),
      .wea(xt_rsc_2_20_wea),
      .da(xt_rsc_2_20_da),
      .adra(xt_rsc_2_20_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_2_20_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_348_4_32_16_16_32_1_gen xt_rsc_2_21_i
      (
      .qa(xt_rsc_2_21_qa),
      .wea(xt_rsc_2_21_wea),
      .da(xt_rsc_2_21_da),
      .adra(xt_rsc_2_21_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_2_21_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_349_4_32_16_16_32_1_gen xt_rsc_2_22_i
      (
      .qa(xt_rsc_2_22_qa),
      .wea(xt_rsc_2_22_wea),
      .da(xt_rsc_2_22_da),
      .adra(xt_rsc_2_22_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_2_22_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_350_4_32_16_16_32_1_gen xt_rsc_2_23_i
      (
      .qa(xt_rsc_2_23_qa),
      .wea(xt_rsc_2_23_wea),
      .da(xt_rsc_2_23_da),
      .adra(xt_rsc_2_23_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_2_23_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_351_4_32_16_16_32_1_gen xt_rsc_2_24_i
      (
      .qa(xt_rsc_2_24_qa),
      .wea(xt_rsc_2_24_wea),
      .da(xt_rsc_2_24_da),
      .adra(xt_rsc_2_24_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_2_24_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_352_4_32_16_16_32_1_gen xt_rsc_2_25_i
      (
      .qa(xt_rsc_2_25_qa),
      .wea(xt_rsc_2_25_wea),
      .da(xt_rsc_2_25_da),
      .adra(xt_rsc_2_25_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_2_25_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_353_4_32_16_16_32_1_gen xt_rsc_2_26_i
      (
      .qa(xt_rsc_2_26_qa),
      .wea(xt_rsc_2_26_wea),
      .da(xt_rsc_2_26_da),
      .adra(xt_rsc_2_26_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_2_26_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_354_4_32_16_16_32_1_gen xt_rsc_2_27_i
      (
      .qa(xt_rsc_2_27_qa),
      .wea(xt_rsc_2_27_wea),
      .da(xt_rsc_2_27_da),
      .adra(xt_rsc_2_27_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_2_27_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_355_4_32_16_16_32_1_gen xt_rsc_2_28_i
      (
      .qa(xt_rsc_2_28_qa),
      .wea(xt_rsc_2_28_wea),
      .da(xt_rsc_2_28_da),
      .adra(xt_rsc_2_28_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_2_28_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_356_4_32_16_16_32_1_gen xt_rsc_2_29_i
      (
      .qa(xt_rsc_2_29_qa),
      .wea(xt_rsc_2_29_wea),
      .da(xt_rsc_2_29_da),
      .adra(xt_rsc_2_29_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_2_29_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_357_4_32_16_16_32_1_gen xt_rsc_2_30_i
      (
      .qa(xt_rsc_2_30_qa),
      .wea(xt_rsc_2_30_wea),
      .da(xt_rsc_2_30_da),
      .adra(xt_rsc_2_30_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_2_30_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_358_4_32_16_16_32_1_gen xt_rsc_2_31_i
      (
      .qa(xt_rsc_2_31_qa),
      .wea(xt_rsc_2_31_wea),
      .da(xt_rsc_2_31_da),
      .adra(xt_rsc_2_31_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_2_31_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_359_4_32_16_16_32_1_gen xt_rsc_3_0_i
      (
      .qa(xt_rsc_3_0_qa),
      .wea(xt_rsc_3_0_wea),
      .da(xt_rsc_3_0_da),
      .adra(xt_rsc_3_0_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_3_0_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_360_4_32_16_16_32_1_gen xt_rsc_3_1_i
      (
      .qa(xt_rsc_3_1_qa),
      .wea(xt_rsc_3_1_wea),
      .da(xt_rsc_3_1_da),
      .adra(xt_rsc_3_1_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_3_1_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_361_4_32_16_16_32_1_gen xt_rsc_3_2_i
      (
      .qa(xt_rsc_3_2_qa),
      .wea(xt_rsc_3_2_wea),
      .da(xt_rsc_3_2_da),
      .adra(xt_rsc_3_2_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_3_2_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_362_4_32_16_16_32_1_gen xt_rsc_3_3_i
      (
      .qa(xt_rsc_3_3_qa),
      .wea(xt_rsc_3_3_wea),
      .da(xt_rsc_3_3_da),
      .adra(xt_rsc_3_3_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_3_3_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_363_4_32_16_16_32_1_gen xt_rsc_3_4_i
      (
      .qa(xt_rsc_3_4_qa),
      .wea(xt_rsc_3_4_wea),
      .da(xt_rsc_3_4_da),
      .adra(xt_rsc_3_4_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_3_4_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_364_4_32_16_16_32_1_gen xt_rsc_3_5_i
      (
      .qa(xt_rsc_3_5_qa),
      .wea(xt_rsc_3_5_wea),
      .da(xt_rsc_3_5_da),
      .adra(xt_rsc_3_5_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_3_5_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_365_4_32_16_16_32_1_gen xt_rsc_3_6_i
      (
      .qa(xt_rsc_3_6_qa),
      .wea(xt_rsc_3_6_wea),
      .da(xt_rsc_3_6_da),
      .adra(xt_rsc_3_6_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_3_6_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_366_4_32_16_16_32_1_gen xt_rsc_3_7_i
      (
      .qa(xt_rsc_3_7_qa),
      .wea(xt_rsc_3_7_wea),
      .da(xt_rsc_3_7_da),
      .adra(xt_rsc_3_7_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_3_7_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_367_4_32_16_16_32_1_gen xt_rsc_3_8_i
      (
      .qa(xt_rsc_3_8_qa),
      .wea(xt_rsc_3_8_wea),
      .da(xt_rsc_3_8_da),
      .adra(xt_rsc_3_8_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_3_8_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_368_4_32_16_16_32_1_gen xt_rsc_3_9_i
      (
      .qa(xt_rsc_3_9_qa),
      .wea(xt_rsc_3_9_wea),
      .da(xt_rsc_3_9_da),
      .adra(xt_rsc_3_9_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_3_9_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_369_4_32_16_16_32_1_gen xt_rsc_3_10_i
      (
      .qa(xt_rsc_3_10_qa),
      .wea(xt_rsc_3_10_wea),
      .da(xt_rsc_3_10_da),
      .adra(xt_rsc_3_10_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_3_10_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_370_4_32_16_16_32_1_gen xt_rsc_3_11_i
      (
      .qa(xt_rsc_3_11_qa),
      .wea(xt_rsc_3_11_wea),
      .da(xt_rsc_3_11_da),
      .adra(xt_rsc_3_11_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_3_11_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_371_4_32_16_16_32_1_gen xt_rsc_3_12_i
      (
      .qa(xt_rsc_3_12_qa),
      .wea(xt_rsc_3_12_wea),
      .da(xt_rsc_3_12_da),
      .adra(xt_rsc_3_12_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_3_12_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_372_4_32_16_16_32_1_gen xt_rsc_3_13_i
      (
      .qa(xt_rsc_3_13_qa),
      .wea(xt_rsc_3_13_wea),
      .da(xt_rsc_3_13_da),
      .adra(xt_rsc_3_13_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_3_13_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_373_4_32_16_16_32_1_gen xt_rsc_3_14_i
      (
      .qa(xt_rsc_3_14_qa),
      .wea(xt_rsc_3_14_wea),
      .da(xt_rsc_3_14_da),
      .adra(xt_rsc_3_14_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_3_14_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_374_4_32_16_16_32_1_gen xt_rsc_3_15_i
      (
      .qa(xt_rsc_3_15_qa),
      .wea(xt_rsc_3_15_wea),
      .da(xt_rsc_3_15_da),
      .adra(xt_rsc_3_15_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_3_15_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_375_4_32_16_16_32_1_gen xt_rsc_3_16_i
      (
      .qa(xt_rsc_3_16_qa),
      .wea(xt_rsc_3_16_wea),
      .da(xt_rsc_3_16_da),
      .adra(xt_rsc_3_16_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_0_0_i_da_d_iff),
      .qa_d(xt_rsc_3_16_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_376_4_32_16_16_32_1_gen xt_rsc_3_17_i
      (
      .qa(xt_rsc_3_17_qa),
      .wea(xt_rsc_3_17_wea),
      .da(xt_rsc_3_17_da),
      .adra(xt_rsc_3_17_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_0_1_i_da_d_iff),
      .qa_d(xt_rsc_3_17_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_377_4_32_16_16_32_1_gen xt_rsc_3_18_i
      (
      .qa(xt_rsc_3_18_qa),
      .wea(xt_rsc_3_18_wea),
      .da(xt_rsc_3_18_da),
      .adra(xt_rsc_3_18_adra),
      .adra_d(xt_rsc_0_2_i_adra_d_iff),
      .da_d(xt_rsc_0_2_i_da_d_iff),
      .qa_d(xt_rsc_3_18_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_378_4_32_16_16_32_1_gen xt_rsc_3_19_i
      (
      .qa(xt_rsc_3_19_qa),
      .wea(xt_rsc_3_19_wea),
      .da(xt_rsc_3_19_da),
      .adra(xt_rsc_3_19_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_0_3_i_da_d_iff),
      .qa_d(xt_rsc_3_19_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_379_4_32_16_16_32_1_gen xt_rsc_3_20_i
      (
      .qa(xt_rsc_3_20_qa),
      .wea(xt_rsc_3_20_wea),
      .da(xt_rsc_3_20_da),
      .adra(xt_rsc_3_20_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_0_4_i_da_d_iff),
      .qa_d(xt_rsc_3_20_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_380_4_32_16_16_32_1_gen xt_rsc_3_21_i
      (
      .qa(xt_rsc_3_21_qa),
      .wea(xt_rsc_3_21_wea),
      .da(xt_rsc_3_21_da),
      .adra(xt_rsc_3_21_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_0_5_i_da_d_iff),
      .qa_d(xt_rsc_3_21_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_381_4_32_16_16_32_1_gen xt_rsc_3_22_i
      (
      .qa(xt_rsc_3_22_qa),
      .wea(xt_rsc_3_22_wea),
      .da(xt_rsc_3_22_da),
      .adra(xt_rsc_3_22_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_0_6_i_da_d_iff),
      .qa_d(xt_rsc_3_22_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_382_4_32_16_16_32_1_gen xt_rsc_3_23_i
      (
      .qa(xt_rsc_3_23_qa),
      .wea(xt_rsc_3_23_wea),
      .da(xt_rsc_3_23_da),
      .adra(xt_rsc_3_23_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_0_7_i_da_d_iff),
      .qa_d(xt_rsc_3_23_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_383_4_32_16_16_32_1_gen xt_rsc_3_24_i
      (
      .qa(xt_rsc_3_24_qa),
      .wea(xt_rsc_3_24_wea),
      .da(xt_rsc_3_24_da),
      .adra(xt_rsc_3_24_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_0_8_i_da_d_iff),
      .qa_d(xt_rsc_3_24_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_384_4_32_16_16_32_1_gen xt_rsc_3_25_i
      (
      .qa(xt_rsc_3_25_qa),
      .wea(xt_rsc_3_25_wea),
      .da(xt_rsc_3_25_da),
      .adra(xt_rsc_3_25_adra),
      .adra_d(xt_rsc_0_9_i_adra_d_iff),
      .da_d(xt_rsc_0_9_i_da_d_iff),
      .qa_d(xt_rsc_3_25_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_385_4_32_16_16_32_1_gen xt_rsc_3_26_i
      (
      .qa(xt_rsc_3_26_qa),
      .wea(xt_rsc_3_26_wea),
      .da(xt_rsc_3_26_da),
      .adra(xt_rsc_3_26_adra),
      .adra_d(xt_rsc_0_10_i_adra_d_iff),
      .da_d(xt_rsc_0_10_i_da_d_iff),
      .qa_d(xt_rsc_3_26_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_386_4_32_16_16_32_1_gen xt_rsc_3_27_i
      (
      .qa(xt_rsc_3_27_qa),
      .wea(xt_rsc_3_27_wea),
      .da(xt_rsc_3_27_da),
      .adra(xt_rsc_3_27_adra),
      .adra_d(xt_rsc_0_11_i_adra_d_iff),
      .da_d(xt_rsc_0_11_i_da_d_iff),
      .qa_d(xt_rsc_3_27_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_387_4_32_16_16_32_1_gen xt_rsc_3_28_i
      (
      .qa(xt_rsc_3_28_qa),
      .wea(xt_rsc_3_28_wea),
      .da(xt_rsc_3_28_da),
      .adra(xt_rsc_3_28_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_0_12_i_da_d_iff),
      .qa_d(xt_rsc_3_28_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_388_4_32_16_16_32_1_gen xt_rsc_3_29_i
      (
      .qa(xt_rsc_3_29_qa),
      .wea(xt_rsc_3_29_wea),
      .da(xt_rsc_3_29_da),
      .adra(xt_rsc_3_29_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_0_13_i_da_d_iff),
      .qa_d(xt_rsc_3_29_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_389_4_32_16_16_32_1_gen xt_rsc_3_30_i
      (
      .qa(xt_rsc_3_30_qa),
      .wea(xt_rsc_3_30_wea),
      .da(xt_rsc_3_30_da),
      .adra(xt_rsc_3_30_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_0_14_i_da_d_iff),
      .qa_d(xt_rsc_3_30_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_390_4_32_16_16_32_1_gen xt_rsc_3_31_i
      (
      .qa(xt_rsc_3_31_qa),
      .wea(xt_rsc_3_31_wea),
      .da(xt_rsc_3_31_da),
      .adra(xt_rsc_3_31_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_0_15_i_da_d_iff),
      .qa_d(xt_rsc_3_31_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_391_4_32_16_16_32_1_gen xt_rsc_4_0_i
      (
      .qa(xt_rsc_4_0_qa),
      .wea(xt_rsc_4_0_wea),
      .da(xt_rsc_4_0_da),
      .adra(xt_rsc_4_0_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_4_0_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_392_4_32_16_16_32_1_gen xt_rsc_4_1_i
      (
      .qa(xt_rsc_4_1_qa),
      .wea(xt_rsc_4_1_wea),
      .da(xt_rsc_4_1_da),
      .adra(xt_rsc_4_1_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_4_1_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_393_4_32_16_16_32_1_gen xt_rsc_4_2_i
      (
      .qa(xt_rsc_4_2_qa),
      .wea(xt_rsc_4_2_wea),
      .da(xt_rsc_4_2_da),
      .adra(xt_rsc_4_2_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_4_2_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_394_4_32_16_16_32_1_gen xt_rsc_4_3_i
      (
      .qa(xt_rsc_4_3_qa),
      .wea(xt_rsc_4_3_wea),
      .da(xt_rsc_4_3_da),
      .adra(xt_rsc_4_3_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_4_3_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_395_4_32_16_16_32_1_gen xt_rsc_4_4_i
      (
      .qa(xt_rsc_4_4_qa),
      .wea(xt_rsc_4_4_wea),
      .da(xt_rsc_4_4_da),
      .adra(xt_rsc_4_4_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_4_4_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_396_4_32_16_16_32_1_gen xt_rsc_4_5_i
      (
      .qa(xt_rsc_4_5_qa),
      .wea(xt_rsc_4_5_wea),
      .da(xt_rsc_4_5_da),
      .adra(xt_rsc_4_5_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_4_5_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_397_4_32_16_16_32_1_gen xt_rsc_4_6_i
      (
      .qa(xt_rsc_4_6_qa),
      .wea(xt_rsc_4_6_wea),
      .da(xt_rsc_4_6_da),
      .adra(xt_rsc_4_6_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_4_6_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_398_4_32_16_16_32_1_gen xt_rsc_4_7_i
      (
      .qa(xt_rsc_4_7_qa),
      .wea(xt_rsc_4_7_wea),
      .da(xt_rsc_4_7_da),
      .adra(xt_rsc_4_7_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_4_7_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_399_4_32_16_16_32_1_gen xt_rsc_4_8_i
      (
      .qa(xt_rsc_4_8_qa),
      .wea(xt_rsc_4_8_wea),
      .da(xt_rsc_4_8_da),
      .adra(xt_rsc_4_8_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_4_8_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_400_4_32_16_16_32_1_gen xt_rsc_4_9_i
      (
      .qa(xt_rsc_4_9_qa),
      .wea(xt_rsc_4_9_wea),
      .da(xt_rsc_4_9_da),
      .adra(xt_rsc_4_9_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_4_9_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_401_4_32_16_16_32_1_gen xt_rsc_4_10_i
      (
      .qa(xt_rsc_4_10_qa),
      .wea(xt_rsc_4_10_wea),
      .da(xt_rsc_4_10_da),
      .adra(xt_rsc_4_10_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_4_10_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_402_4_32_16_16_32_1_gen xt_rsc_4_11_i
      (
      .qa(xt_rsc_4_11_qa),
      .wea(xt_rsc_4_11_wea),
      .da(xt_rsc_4_11_da),
      .adra(xt_rsc_4_11_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_4_11_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_403_4_32_16_16_32_1_gen xt_rsc_4_12_i
      (
      .qa(xt_rsc_4_12_qa),
      .wea(xt_rsc_4_12_wea),
      .da(xt_rsc_4_12_da),
      .adra(xt_rsc_4_12_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_4_12_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_404_4_32_16_16_32_1_gen xt_rsc_4_13_i
      (
      .qa(xt_rsc_4_13_qa),
      .wea(xt_rsc_4_13_wea),
      .da(xt_rsc_4_13_da),
      .adra(xt_rsc_4_13_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_4_13_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_405_4_32_16_16_32_1_gen xt_rsc_4_14_i
      (
      .qa(xt_rsc_4_14_qa),
      .wea(xt_rsc_4_14_wea),
      .da(xt_rsc_4_14_da),
      .adra(xt_rsc_4_14_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_4_14_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_406_4_32_16_16_32_1_gen xt_rsc_4_15_i
      (
      .qa(xt_rsc_4_15_qa),
      .wea(xt_rsc_4_15_wea),
      .da(xt_rsc_4_15_da),
      .adra(xt_rsc_4_15_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_4_15_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_407_4_32_16_16_32_1_gen xt_rsc_4_16_i
      (
      .qa(xt_rsc_4_16_qa),
      .wea(xt_rsc_4_16_wea),
      .da(xt_rsc_4_16_da),
      .adra(xt_rsc_4_16_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_4_16_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_408_4_32_16_16_32_1_gen xt_rsc_4_17_i
      (
      .qa(xt_rsc_4_17_qa),
      .wea(xt_rsc_4_17_wea),
      .da(xt_rsc_4_17_da),
      .adra(xt_rsc_4_17_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_4_17_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_409_4_32_16_16_32_1_gen xt_rsc_4_18_i
      (
      .qa(xt_rsc_4_18_qa),
      .wea(xt_rsc_4_18_wea),
      .da(xt_rsc_4_18_da),
      .adra(xt_rsc_4_18_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_4_18_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_410_4_32_16_16_32_1_gen xt_rsc_4_19_i
      (
      .qa(xt_rsc_4_19_qa),
      .wea(xt_rsc_4_19_wea),
      .da(xt_rsc_4_19_da),
      .adra(xt_rsc_4_19_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_4_19_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_411_4_32_16_16_32_1_gen xt_rsc_4_20_i
      (
      .qa(xt_rsc_4_20_qa),
      .wea(xt_rsc_4_20_wea),
      .da(xt_rsc_4_20_da),
      .adra(xt_rsc_4_20_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_4_20_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_412_4_32_16_16_32_1_gen xt_rsc_4_21_i
      (
      .qa(xt_rsc_4_21_qa),
      .wea(xt_rsc_4_21_wea),
      .da(xt_rsc_4_21_da),
      .adra(xt_rsc_4_21_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_4_21_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_413_4_32_16_16_32_1_gen xt_rsc_4_22_i
      (
      .qa(xt_rsc_4_22_qa),
      .wea(xt_rsc_4_22_wea),
      .da(xt_rsc_4_22_da),
      .adra(xt_rsc_4_22_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_4_22_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_414_4_32_16_16_32_1_gen xt_rsc_4_23_i
      (
      .qa(xt_rsc_4_23_qa),
      .wea(xt_rsc_4_23_wea),
      .da(xt_rsc_4_23_da),
      .adra(xt_rsc_4_23_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_4_23_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_415_4_32_16_16_32_1_gen xt_rsc_4_24_i
      (
      .qa(xt_rsc_4_24_qa),
      .wea(xt_rsc_4_24_wea),
      .da(xt_rsc_4_24_da),
      .adra(xt_rsc_4_24_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_4_24_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_416_4_32_16_16_32_1_gen xt_rsc_4_25_i
      (
      .qa(xt_rsc_4_25_qa),
      .wea(xt_rsc_4_25_wea),
      .da(xt_rsc_4_25_da),
      .adra(xt_rsc_4_25_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_4_25_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_417_4_32_16_16_32_1_gen xt_rsc_4_26_i
      (
      .qa(xt_rsc_4_26_qa),
      .wea(xt_rsc_4_26_wea),
      .da(xt_rsc_4_26_da),
      .adra(xt_rsc_4_26_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_4_26_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_418_4_32_16_16_32_1_gen xt_rsc_4_27_i
      (
      .qa(xt_rsc_4_27_qa),
      .wea(xt_rsc_4_27_wea),
      .da(xt_rsc_4_27_da),
      .adra(xt_rsc_4_27_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_4_27_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_419_4_32_16_16_32_1_gen xt_rsc_4_28_i
      (
      .qa(xt_rsc_4_28_qa),
      .wea(xt_rsc_4_28_wea),
      .da(xt_rsc_4_28_da),
      .adra(xt_rsc_4_28_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_4_28_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_420_4_32_16_16_32_1_gen xt_rsc_4_29_i
      (
      .qa(xt_rsc_4_29_qa),
      .wea(xt_rsc_4_29_wea),
      .da(xt_rsc_4_29_da),
      .adra(xt_rsc_4_29_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_4_29_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_421_4_32_16_16_32_1_gen xt_rsc_4_30_i
      (
      .qa(xt_rsc_4_30_qa),
      .wea(xt_rsc_4_30_wea),
      .da(xt_rsc_4_30_da),
      .adra(xt_rsc_4_30_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_4_30_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_422_4_32_16_16_32_1_gen xt_rsc_4_31_i
      (
      .qa(xt_rsc_4_31_qa),
      .wea(xt_rsc_4_31_wea),
      .da(xt_rsc_4_31_da),
      .adra(xt_rsc_4_31_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_4_31_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_423_4_32_16_16_32_1_gen xt_rsc_5_0_i
      (
      .qa(xt_rsc_5_0_qa),
      .wea(xt_rsc_5_0_wea),
      .da(xt_rsc_5_0_da),
      .adra(xt_rsc_5_0_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_5_0_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_424_4_32_16_16_32_1_gen xt_rsc_5_1_i
      (
      .qa(xt_rsc_5_1_qa),
      .wea(xt_rsc_5_1_wea),
      .da(xt_rsc_5_1_da),
      .adra(xt_rsc_5_1_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_5_1_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_425_4_32_16_16_32_1_gen xt_rsc_5_2_i
      (
      .qa(xt_rsc_5_2_qa),
      .wea(xt_rsc_5_2_wea),
      .da(xt_rsc_5_2_da),
      .adra(xt_rsc_5_2_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_5_2_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_426_4_32_16_16_32_1_gen xt_rsc_5_3_i
      (
      .qa(xt_rsc_5_3_qa),
      .wea(xt_rsc_5_3_wea),
      .da(xt_rsc_5_3_da),
      .adra(xt_rsc_5_3_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_5_3_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_427_4_32_16_16_32_1_gen xt_rsc_5_4_i
      (
      .qa(xt_rsc_5_4_qa),
      .wea(xt_rsc_5_4_wea),
      .da(xt_rsc_5_4_da),
      .adra(xt_rsc_5_4_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_5_4_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_428_4_32_16_16_32_1_gen xt_rsc_5_5_i
      (
      .qa(xt_rsc_5_5_qa),
      .wea(xt_rsc_5_5_wea),
      .da(xt_rsc_5_5_da),
      .adra(xt_rsc_5_5_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_5_5_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_429_4_32_16_16_32_1_gen xt_rsc_5_6_i
      (
      .qa(xt_rsc_5_6_qa),
      .wea(xt_rsc_5_6_wea),
      .da(xt_rsc_5_6_da),
      .adra(xt_rsc_5_6_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_5_6_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_430_4_32_16_16_32_1_gen xt_rsc_5_7_i
      (
      .qa(xt_rsc_5_7_qa),
      .wea(xt_rsc_5_7_wea),
      .da(xt_rsc_5_7_da),
      .adra(xt_rsc_5_7_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_5_7_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_431_4_32_16_16_32_1_gen xt_rsc_5_8_i
      (
      .qa(xt_rsc_5_8_qa),
      .wea(xt_rsc_5_8_wea),
      .da(xt_rsc_5_8_da),
      .adra(xt_rsc_5_8_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_5_8_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_432_4_32_16_16_32_1_gen xt_rsc_5_9_i
      (
      .qa(xt_rsc_5_9_qa),
      .wea(xt_rsc_5_9_wea),
      .da(xt_rsc_5_9_da),
      .adra(xt_rsc_5_9_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_5_9_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_433_4_32_16_16_32_1_gen xt_rsc_5_10_i
      (
      .qa(xt_rsc_5_10_qa),
      .wea(xt_rsc_5_10_wea),
      .da(xt_rsc_5_10_da),
      .adra(xt_rsc_5_10_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_5_10_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_434_4_32_16_16_32_1_gen xt_rsc_5_11_i
      (
      .qa(xt_rsc_5_11_qa),
      .wea(xt_rsc_5_11_wea),
      .da(xt_rsc_5_11_da),
      .adra(xt_rsc_5_11_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_5_11_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_435_4_32_16_16_32_1_gen xt_rsc_5_12_i
      (
      .qa(xt_rsc_5_12_qa),
      .wea(xt_rsc_5_12_wea),
      .da(xt_rsc_5_12_da),
      .adra(xt_rsc_5_12_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_5_12_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_436_4_32_16_16_32_1_gen xt_rsc_5_13_i
      (
      .qa(xt_rsc_5_13_qa),
      .wea(xt_rsc_5_13_wea),
      .da(xt_rsc_5_13_da),
      .adra(xt_rsc_5_13_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_5_13_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_437_4_32_16_16_32_1_gen xt_rsc_5_14_i
      (
      .qa(xt_rsc_5_14_qa),
      .wea(xt_rsc_5_14_wea),
      .da(xt_rsc_5_14_da),
      .adra(xt_rsc_5_14_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_5_14_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_438_4_32_16_16_32_1_gen xt_rsc_5_15_i
      (
      .qa(xt_rsc_5_15_qa),
      .wea(xt_rsc_5_15_wea),
      .da(xt_rsc_5_15_da),
      .adra(xt_rsc_5_15_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_5_15_i_qa_d),
      .wea_d(xt_rsc_1_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_439_4_32_16_16_32_1_gen xt_rsc_5_16_i
      (
      .qa(xt_rsc_5_16_qa),
      .wea(xt_rsc_5_16_wea),
      .da(xt_rsc_5_16_da),
      .adra(xt_rsc_5_16_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_5_16_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_440_4_32_16_16_32_1_gen xt_rsc_5_17_i
      (
      .qa(xt_rsc_5_17_qa),
      .wea(xt_rsc_5_17_wea),
      .da(xt_rsc_5_17_da),
      .adra(xt_rsc_5_17_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_5_17_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_441_4_32_16_16_32_1_gen xt_rsc_5_18_i
      (
      .qa(xt_rsc_5_18_qa),
      .wea(xt_rsc_5_18_wea),
      .da(xt_rsc_5_18_da),
      .adra(xt_rsc_5_18_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_5_18_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_442_4_32_16_16_32_1_gen xt_rsc_5_19_i
      (
      .qa(xt_rsc_5_19_qa),
      .wea(xt_rsc_5_19_wea),
      .da(xt_rsc_5_19_da),
      .adra(xt_rsc_5_19_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_5_19_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_443_4_32_16_16_32_1_gen xt_rsc_5_20_i
      (
      .qa(xt_rsc_5_20_qa),
      .wea(xt_rsc_5_20_wea),
      .da(xt_rsc_5_20_da),
      .adra(xt_rsc_5_20_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_5_20_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_444_4_32_16_16_32_1_gen xt_rsc_5_21_i
      (
      .qa(xt_rsc_5_21_qa),
      .wea(xt_rsc_5_21_wea),
      .da(xt_rsc_5_21_da),
      .adra(xt_rsc_5_21_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_5_21_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_445_4_32_16_16_32_1_gen xt_rsc_5_22_i
      (
      .qa(xt_rsc_5_22_qa),
      .wea(xt_rsc_5_22_wea),
      .da(xt_rsc_5_22_da),
      .adra(xt_rsc_5_22_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_5_22_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_446_4_32_16_16_32_1_gen xt_rsc_5_23_i
      (
      .qa(xt_rsc_5_23_qa),
      .wea(xt_rsc_5_23_wea),
      .da(xt_rsc_5_23_da),
      .adra(xt_rsc_5_23_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_5_23_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_447_4_32_16_16_32_1_gen xt_rsc_5_24_i
      (
      .qa(xt_rsc_5_24_qa),
      .wea(xt_rsc_5_24_wea),
      .da(xt_rsc_5_24_da),
      .adra(xt_rsc_5_24_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_5_24_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_448_4_32_16_16_32_1_gen xt_rsc_5_25_i
      (
      .qa(xt_rsc_5_25_qa),
      .wea(xt_rsc_5_25_wea),
      .da(xt_rsc_5_25_da),
      .adra(xt_rsc_5_25_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_5_25_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_449_4_32_16_16_32_1_gen xt_rsc_5_26_i
      (
      .qa(xt_rsc_5_26_qa),
      .wea(xt_rsc_5_26_wea),
      .da(xt_rsc_5_26_da),
      .adra(xt_rsc_5_26_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_5_26_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_450_4_32_16_16_32_1_gen xt_rsc_5_27_i
      (
      .qa(xt_rsc_5_27_qa),
      .wea(xt_rsc_5_27_wea),
      .da(xt_rsc_5_27_da),
      .adra(xt_rsc_5_27_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_5_27_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_451_4_32_16_16_32_1_gen xt_rsc_5_28_i
      (
      .qa(xt_rsc_5_28_qa),
      .wea(xt_rsc_5_28_wea),
      .da(xt_rsc_5_28_da),
      .adra(xt_rsc_5_28_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_5_28_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_452_4_32_16_16_32_1_gen xt_rsc_5_29_i
      (
      .qa(xt_rsc_5_29_qa),
      .wea(xt_rsc_5_29_wea),
      .da(xt_rsc_5_29_da),
      .adra(xt_rsc_5_29_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_5_29_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_453_4_32_16_16_32_1_gen xt_rsc_5_30_i
      (
      .qa(xt_rsc_5_30_qa),
      .wea(xt_rsc_5_30_wea),
      .da(xt_rsc_5_30_da),
      .adra(xt_rsc_5_30_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_5_30_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_454_4_32_16_16_32_1_gen xt_rsc_5_31_i
      (
      .qa(xt_rsc_5_31_qa),
      .wea(xt_rsc_5_31_wea),
      .da(xt_rsc_5_31_da),
      .adra(xt_rsc_5_31_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_5_31_i_qa_d),
      .wea_d(xt_rsc_1_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_1_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_455_4_32_16_16_32_1_gen xt_rsc_6_0_i
      (
      .qa(xt_rsc_6_0_qa),
      .wea(xt_rsc_6_0_wea),
      .da(xt_rsc_6_0_da),
      .adra(xt_rsc_6_0_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_6_0_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_456_4_32_16_16_32_1_gen xt_rsc_6_1_i
      (
      .qa(xt_rsc_6_1_qa),
      .wea(xt_rsc_6_1_wea),
      .da(xt_rsc_6_1_da),
      .adra(xt_rsc_6_1_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_6_1_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_457_4_32_16_16_32_1_gen xt_rsc_6_2_i
      (
      .qa(xt_rsc_6_2_qa),
      .wea(xt_rsc_6_2_wea),
      .da(xt_rsc_6_2_da),
      .adra(xt_rsc_6_2_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_6_2_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_458_4_32_16_16_32_1_gen xt_rsc_6_3_i
      (
      .qa(xt_rsc_6_3_qa),
      .wea(xt_rsc_6_3_wea),
      .da(xt_rsc_6_3_da),
      .adra(xt_rsc_6_3_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_6_3_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_459_4_32_16_16_32_1_gen xt_rsc_6_4_i
      (
      .qa(xt_rsc_6_4_qa),
      .wea(xt_rsc_6_4_wea),
      .da(xt_rsc_6_4_da),
      .adra(xt_rsc_6_4_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_6_4_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_460_4_32_16_16_32_1_gen xt_rsc_6_5_i
      (
      .qa(xt_rsc_6_5_qa),
      .wea(xt_rsc_6_5_wea),
      .da(xt_rsc_6_5_da),
      .adra(xt_rsc_6_5_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_6_5_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_461_4_32_16_16_32_1_gen xt_rsc_6_6_i
      (
      .qa(xt_rsc_6_6_qa),
      .wea(xt_rsc_6_6_wea),
      .da(xt_rsc_6_6_da),
      .adra(xt_rsc_6_6_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_6_6_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_462_4_32_16_16_32_1_gen xt_rsc_6_7_i
      (
      .qa(xt_rsc_6_7_qa),
      .wea(xt_rsc_6_7_wea),
      .da(xt_rsc_6_7_da),
      .adra(xt_rsc_6_7_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_6_7_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_463_4_32_16_16_32_1_gen xt_rsc_6_8_i
      (
      .qa(xt_rsc_6_8_qa),
      .wea(xt_rsc_6_8_wea),
      .da(xt_rsc_6_8_da),
      .adra(xt_rsc_6_8_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_6_8_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_464_4_32_16_16_32_1_gen xt_rsc_6_9_i
      (
      .qa(xt_rsc_6_9_qa),
      .wea(xt_rsc_6_9_wea),
      .da(xt_rsc_6_9_da),
      .adra(xt_rsc_6_9_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_6_9_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_465_4_32_16_16_32_1_gen xt_rsc_6_10_i
      (
      .qa(xt_rsc_6_10_qa),
      .wea(xt_rsc_6_10_wea),
      .da(xt_rsc_6_10_da),
      .adra(xt_rsc_6_10_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_6_10_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_466_4_32_16_16_32_1_gen xt_rsc_6_11_i
      (
      .qa(xt_rsc_6_11_qa),
      .wea(xt_rsc_6_11_wea),
      .da(xt_rsc_6_11_da),
      .adra(xt_rsc_6_11_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_6_11_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_467_4_32_16_16_32_1_gen xt_rsc_6_12_i
      (
      .qa(xt_rsc_6_12_qa),
      .wea(xt_rsc_6_12_wea),
      .da(xt_rsc_6_12_da),
      .adra(xt_rsc_6_12_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_6_12_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_468_4_32_16_16_32_1_gen xt_rsc_6_13_i
      (
      .qa(xt_rsc_6_13_qa),
      .wea(xt_rsc_6_13_wea),
      .da(xt_rsc_6_13_da),
      .adra(xt_rsc_6_13_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_6_13_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_469_4_32_16_16_32_1_gen xt_rsc_6_14_i
      (
      .qa(xt_rsc_6_14_qa),
      .wea(xt_rsc_6_14_wea),
      .da(xt_rsc_6_14_da),
      .adra(xt_rsc_6_14_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_6_14_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_470_4_32_16_16_32_1_gen xt_rsc_6_15_i
      (
      .qa(xt_rsc_6_15_qa),
      .wea(xt_rsc_6_15_wea),
      .da(xt_rsc_6_15_da),
      .adra(xt_rsc_6_15_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_6_15_i_qa_d),
      .wea_d(xt_rsc_2_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_471_4_32_16_16_32_1_gen xt_rsc_6_16_i
      (
      .qa(xt_rsc_6_16_qa),
      .wea(xt_rsc_6_16_wea),
      .da(xt_rsc_6_16_da),
      .adra(xt_rsc_6_16_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_6_16_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_472_4_32_16_16_32_1_gen xt_rsc_6_17_i
      (
      .qa(xt_rsc_6_17_qa),
      .wea(xt_rsc_6_17_wea),
      .da(xt_rsc_6_17_da),
      .adra(xt_rsc_6_17_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_6_17_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_473_4_32_16_16_32_1_gen xt_rsc_6_18_i
      (
      .qa(xt_rsc_6_18_qa),
      .wea(xt_rsc_6_18_wea),
      .da(xt_rsc_6_18_da),
      .adra(xt_rsc_6_18_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_6_18_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_474_4_32_16_16_32_1_gen xt_rsc_6_19_i
      (
      .qa(xt_rsc_6_19_qa),
      .wea(xt_rsc_6_19_wea),
      .da(xt_rsc_6_19_da),
      .adra(xt_rsc_6_19_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_6_19_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_475_4_32_16_16_32_1_gen xt_rsc_6_20_i
      (
      .qa(xt_rsc_6_20_qa),
      .wea(xt_rsc_6_20_wea),
      .da(xt_rsc_6_20_da),
      .adra(xt_rsc_6_20_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_6_20_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_476_4_32_16_16_32_1_gen xt_rsc_6_21_i
      (
      .qa(xt_rsc_6_21_qa),
      .wea(xt_rsc_6_21_wea),
      .da(xt_rsc_6_21_da),
      .adra(xt_rsc_6_21_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_6_21_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_477_4_32_16_16_32_1_gen xt_rsc_6_22_i
      (
      .qa(xt_rsc_6_22_qa),
      .wea(xt_rsc_6_22_wea),
      .da(xt_rsc_6_22_da),
      .adra(xt_rsc_6_22_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_6_22_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_478_4_32_16_16_32_1_gen xt_rsc_6_23_i
      (
      .qa(xt_rsc_6_23_qa),
      .wea(xt_rsc_6_23_wea),
      .da(xt_rsc_6_23_da),
      .adra(xt_rsc_6_23_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_6_23_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_479_4_32_16_16_32_1_gen xt_rsc_6_24_i
      (
      .qa(xt_rsc_6_24_qa),
      .wea(xt_rsc_6_24_wea),
      .da(xt_rsc_6_24_da),
      .adra(xt_rsc_6_24_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_6_24_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_480_4_32_16_16_32_1_gen xt_rsc_6_25_i
      (
      .qa(xt_rsc_6_25_qa),
      .wea(xt_rsc_6_25_wea),
      .da(xt_rsc_6_25_da),
      .adra(xt_rsc_6_25_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_6_25_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_481_4_32_16_16_32_1_gen xt_rsc_6_26_i
      (
      .qa(xt_rsc_6_26_qa),
      .wea(xt_rsc_6_26_wea),
      .da(xt_rsc_6_26_da),
      .adra(xt_rsc_6_26_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_6_26_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_482_4_32_16_16_32_1_gen xt_rsc_6_27_i
      (
      .qa(xt_rsc_6_27_qa),
      .wea(xt_rsc_6_27_wea),
      .da(xt_rsc_6_27_da),
      .adra(xt_rsc_6_27_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_6_27_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_483_4_32_16_16_32_1_gen xt_rsc_6_28_i
      (
      .qa(xt_rsc_6_28_qa),
      .wea(xt_rsc_6_28_wea),
      .da(xt_rsc_6_28_da),
      .adra(xt_rsc_6_28_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_6_28_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_484_4_32_16_16_32_1_gen xt_rsc_6_29_i
      (
      .qa(xt_rsc_6_29_qa),
      .wea(xt_rsc_6_29_wea),
      .da(xt_rsc_6_29_da),
      .adra(xt_rsc_6_29_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_6_29_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_485_4_32_16_16_32_1_gen xt_rsc_6_30_i
      (
      .qa(xt_rsc_6_30_qa),
      .wea(xt_rsc_6_30_wea),
      .da(xt_rsc_6_30_da),
      .adra(xt_rsc_6_30_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_6_30_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_486_4_32_16_16_32_1_gen xt_rsc_6_31_i
      (
      .qa(xt_rsc_6_31_qa),
      .wea(xt_rsc_6_31_wea),
      .da(xt_rsc_6_31_da),
      .adra(xt_rsc_6_31_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_6_31_i_qa_d),
      .wea_d(xt_rsc_2_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_2_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_487_4_32_16_16_32_1_gen xt_rsc_7_0_i
      (
      .qa(xt_rsc_7_0_qa),
      .wea(xt_rsc_7_0_wea),
      .da(xt_rsc_7_0_da),
      .adra(xt_rsc_7_0_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_7_0_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_488_4_32_16_16_32_1_gen xt_rsc_7_1_i
      (
      .qa(xt_rsc_7_1_qa),
      .wea(xt_rsc_7_1_wea),
      .da(xt_rsc_7_1_da),
      .adra(xt_rsc_7_1_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_7_1_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_489_4_32_16_16_32_1_gen xt_rsc_7_2_i
      (
      .qa(xt_rsc_7_2_qa),
      .wea(xt_rsc_7_2_wea),
      .da(xt_rsc_7_2_da),
      .adra(xt_rsc_7_2_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_7_2_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_490_4_32_16_16_32_1_gen xt_rsc_7_3_i
      (
      .qa(xt_rsc_7_3_qa),
      .wea(xt_rsc_7_3_wea),
      .da(xt_rsc_7_3_da),
      .adra(xt_rsc_7_3_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_7_3_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_491_4_32_16_16_32_1_gen xt_rsc_7_4_i
      (
      .qa(xt_rsc_7_4_qa),
      .wea(xt_rsc_7_4_wea),
      .da(xt_rsc_7_4_da),
      .adra(xt_rsc_7_4_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_7_4_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_492_4_32_16_16_32_1_gen xt_rsc_7_5_i
      (
      .qa(xt_rsc_7_5_qa),
      .wea(xt_rsc_7_5_wea),
      .da(xt_rsc_7_5_da),
      .adra(xt_rsc_7_5_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_7_5_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_493_4_32_16_16_32_1_gen xt_rsc_7_6_i
      (
      .qa(xt_rsc_7_6_qa),
      .wea(xt_rsc_7_6_wea),
      .da(xt_rsc_7_6_da),
      .adra(xt_rsc_7_6_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_7_6_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_494_4_32_16_16_32_1_gen xt_rsc_7_7_i
      (
      .qa(xt_rsc_7_7_qa),
      .wea(xt_rsc_7_7_wea),
      .da(xt_rsc_7_7_da),
      .adra(xt_rsc_7_7_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_7_7_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_495_4_32_16_16_32_1_gen xt_rsc_7_8_i
      (
      .qa(xt_rsc_7_8_qa),
      .wea(xt_rsc_7_8_wea),
      .da(xt_rsc_7_8_da),
      .adra(xt_rsc_7_8_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_7_8_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_496_4_32_16_16_32_1_gen xt_rsc_7_9_i
      (
      .qa(xt_rsc_7_9_qa),
      .wea(xt_rsc_7_9_wea),
      .da(xt_rsc_7_9_da),
      .adra(xt_rsc_7_9_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_7_9_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_497_4_32_16_16_32_1_gen xt_rsc_7_10_i
      (
      .qa(xt_rsc_7_10_qa),
      .wea(xt_rsc_7_10_wea),
      .da(xt_rsc_7_10_da),
      .adra(xt_rsc_7_10_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_7_10_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_498_4_32_16_16_32_1_gen xt_rsc_7_11_i
      (
      .qa(xt_rsc_7_11_qa),
      .wea(xt_rsc_7_11_wea),
      .da(xt_rsc_7_11_da),
      .adra(xt_rsc_7_11_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_7_11_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_499_4_32_16_16_32_1_gen xt_rsc_7_12_i
      (
      .qa(xt_rsc_7_12_qa),
      .wea(xt_rsc_7_12_wea),
      .da(xt_rsc_7_12_da),
      .adra(xt_rsc_7_12_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_7_12_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_500_4_32_16_16_32_1_gen xt_rsc_7_13_i
      (
      .qa(xt_rsc_7_13_qa),
      .wea(xt_rsc_7_13_wea),
      .da(xt_rsc_7_13_da),
      .adra(xt_rsc_7_13_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_7_13_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_501_4_32_16_16_32_1_gen xt_rsc_7_14_i
      (
      .qa(xt_rsc_7_14_qa),
      .wea(xt_rsc_7_14_wea),
      .da(xt_rsc_7_14_da),
      .adra(xt_rsc_7_14_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_7_14_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_502_4_32_16_16_32_1_gen xt_rsc_7_15_i
      (
      .qa(xt_rsc_7_15_qa),
      .wea(xt_rsc_7_15_wea),
      .da(xt_rsc_7_15_da),
      .adra(xt_rsc_7_15_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_7_15_i_qa_d),
      .wea_d(xt_rsc_3_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_503_4_32_16_16_32_1_gen xt_rsc_7_16_i
      (
      .qa(xt_rsc_7_16_qa),
      .wea(xt_rsc_7_16_wea),
      .da(xt_rsc_7_16_da),
      .adra(xt_rsc_7_16_adra),
      .adra_d(xt_rsc_0_8_i_adra_d_iff),
      .da_d(xt_rsc_4_0_i_da_d_iff),
      .qa_d(xt_rsc_7_16_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_504_4_32_16_16_32_1_gen xt_rsc_7_17_i
      (
      .qa(xt_rsc_7_17_qa),
      .wea(xt_rsc_7_17_wea),
      .da(xt_rsc_7_17_da),
      .adra(xt_rsc_7_17_adra),
      .adra_d(xt_rsc_4_1_i_adra_d_iff),
      .da_d(xt_rsc_4_1_i_da_d_iff),
      .qa_d(xt_rsc_7_17_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_505_4_32_16_16_32_1_gen xt_rsc_7_18_i
      (
      .qa(xt_rsc_7_18_qa),
      .wea(xt_rsc_7_18_wea),
      .da(xt_rsc_7_18_da),
      .adra(xt_rsc_7_18_adra),
      .adra_d(xt_rsc_4_2_i_adra_d_iff),
      .da_d(xt_rsc_4_2_i_da_d_iff),
      .qa_d(xt_rsc_7_18_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_506_4_32_16_16_32_1_gen xt_rsc_7_19_i
      (
      .qa(xt_rsc_7_19_qa),
      .wea(xt_rsc_7_19_wea),
      .da(xt_rsc_7_19_da),
      .adra(xt_rsc_7_19_adra),
      .adra_d(xt_rsc_0_12_i_adra_d_iff),
      .da_d(xt_rsc_4_3_i_da_d_iff),
      .qa_d(xt_rsc_7_19_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_507_4_32_16_16_32_1_gen xt_rsc_7_20_i
      (
      .qa(xt_rsc_7_20_qa),
      .wea(xt_rsc_7_20_wea),
      .da(xt_rsc_7_20_da),
      .adra(xt_rsc_7_20_adra),
      .adra_d(xt_rsc_0_13_i_adra_d_iff),
      .da_d(xt_rsc_4_4_i_da_d_iff),
      .qa_d(xt_rsc_7_20_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_508_4_32_16_16_32_1_gen xt_rsc_7_21_i
      (
      .qa(xt_rsc_7_21_qa),
      .wea(xt_rsc_7_21_wea),
      .da(xt_rsc_7_21_da),
      .adra(xt_rsc_7_21_adra),
      .adra_d(xt_rsc_0_14_i_adra_d_iff),
      .da_d(xt_rsc_4_5_i_da_d_iff),
      .qa_d(xt_rsc_7_21_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_509_4_32_16_16_32_1_gen xt_rsc_7_22_i
      (
      .qa(xt_rsc_7_22_qa),
      .wea(xt_rsc_7_22_wea),
      .da(xt_rsc_7_22_da),
      .adra(xt_rsc_7_22_adra),
      .adra_d(xt_rsc_0_15_i_adra_d_iff),
      .da_d(xt_rsc_4_6_i_da_d_iff),
      .qa_d(xt_rsc_7_22_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_510_4_32_16_16_32_1_gen xt_rsc_7_23_i
      (
      .qa(xt_rsc_7_23_qa),
      .wea(xt_rsc_7_23_wea),
      .da(xt_rsc_7_23_da),
      .adra(xt_rsc_7_23_adra),
      .adra_d(xt_rsc_0_0_i_adra_d_iff),
      .da_d(xt_rsc_4_7_i_da_d_iff),
      .qa_d(xt_rsc_7_23_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_511_4_32_16_16_32_1_gen xt_rsc_7_24_i
      (
      .qa(xt_rsc_7_24_qa),
      .wea(xt_rsc_7_24_wea),
      .da(xt_rsc_7_24_da),
      .adra(xt_rsc_7_24_adra),
      .adra_d(xt_rsc_0_1_i_adra_d_iff),
      .da_d(xt_rsc_4_8_i_da_d_iff),
      .qa_d(xt_rsc_7_24_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_512_4_32_16_16_32_1_gen xt_rsc_7_25_i
      (
      .qa(xt_rsc_7_25_qa),
      .wea(xt_rsc_7_25_wea),
      .da(xt_rsc_7_25_da),
      .adra(xt_rsc_7_25_adra),
      .adra_d(xt_rsc_4_9_i_adra_d_iff),
      .da_d(xt_rsc_4_9_i_da_d_iff),
      .qa_d(xt_rsc_7_25_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_513_4_32_16_16_32_1_gen xt_rsc_7_26_i
      (
      .qa(xt_rsc_7_26_qa),
      .wea(xt_rsc_7_26_wea),
      .da(xt_rsc_7_26_da),
      .adra(xt_rsc_7_26_adra),
      .adra_d(xt_rsc_4_10_i_adra_d_iff),
      .da_d(xt_rsc_4_10_i_da_d_iff),
      .qa_d(xt_rsc_7_26_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_514_4_32_16_16_32_1_gen xt_rsc_7_27_i
      (
      .qa(xt_rsc_7_27_qa),
      .wea(xt_rsc_7_27_wea),
      .da(xt_rsc_7_27_da),
      .adra(xt_rsc_7_27_adra),
      .adra_d(xt_rsc_0_3_i_adra_d_iff),
      .da_d(xt_rsc_4_11_i_da_d_iff),
      .qa_d(xt_rsc_7_27_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_515_4_32_16_16_32_1_gen xt_rsc_7_28_i
      (
      .qa(xt_rsc_7_28_qa),
      .wea(xt_rsc_7_28_wea),
      .da(xt_rsc_7_28_da),
      .adra(xt_rsc_7_28_adra),
      .adra_d(xt_rsc_0_4_i_adra_d_iff),
      .da_d(xt_rsc_4_12_i_da_d_iff),
      .qa_d(xt_rsc_7_28_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_516_4_32_16_16_32_1_gen xt_rsc_7_29_i
      (
      .qa(xt_rsc_7_29_qa),
      .wea(xt_rsc_7_29_wea),
      .da(xt_rsc_7_29_da),
      .adra(xt_rsc_7_29_adra),
      .adra_d(xt_rsc_0_5_i_adra_d_iff),
      .da_d(xt_rsc_4_13_i_da_d_iff),
      .qa_d(xt_rsc_7_29_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_517_4_32_16_16_32_1_gen xt_rsc_7_30_i
      (
      .qa(xt_rsc_7_30_qa),
      .wea(xt_rsc_7_30_wea),
      .da(xt_rsc_7_30_da),
      .adra(xt_rsc_7_30_adra),
      .adra_d(xt_rsc_0_6_i_adra_d_iff),
      .da_d(xt_rsc_4_14_i_da_d_iff),
      .qa_d(xt_rsc_7_30_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_518_4_32_16_16_32_1_gen xt_rsc_7_31_i
      (
      .qa(xt_rsc_7_31_qa),
      .wea(xt_rsc_7_31_wea),
      .da(xt_rsc_7_31_da),
      .adra(xt_rsc_7_31_adra),
      .adra_d(xt_rsc_0_7_i_adra_d_iff),
      .da_d(xt_rsc_4_15_i_da_d_iff),
      .qa_d(xt_rsc_7_31_i_qa_d),
      .wea_d(xt_rsc_3_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_3_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_519_8_32_256_256_32_1_gen twiddle_rsc_0_0_i
      (
      .qb(twiddle_rsc_0_0_qb),
      .web(twiddle_rsc_0_0_web),
      .db(twiddle_rsc_0_0_db),
      .adrb(twiddle_rsc_0_0_adrb),
      .qa(twiddle_rsc_0_0_qa),
      .wea(twiddle_rsc_0_0_wea),
      .da(twiddle_rsc_0_0_da),
      .adra(twiddle_rsc_0_0_adra),
      .adra_d(nl_twiddle_rsc_0_0_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_0_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_520_8_32_256_256_32_1_gen twiddle_rsc_0_1_i
      (
      .qb(twiddle_rsc_0_1_qb),
      .web(twiddle_rsc_0_1_web),
      .db(twiddle_rsc_0_1_db),
      .adrb(twiddle_rsc_0_1_adrb),
      .qa(twiddle_rsc_0_1_qa),
      .wea(twiddle_rsc_0_1_wea),
      .da(twiddle_rsc_0_1_da),
      .adra(twiddle_rsc_0_1_adra),
      .adra_d(nl_twiddle_rsc_0_1_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_1_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_521_8_32_256_256_32_1_gen twiddle_rsc_0_2_i
      (
      .qb(twiddle_rsc_0_2_qb),
      .web(twiddle_rsc_0_2_web),
      .db(twiddle_rsc_0_2_db),
      .adrb(twiddle_rsc_0_2_adrb),
      .qa(twiddle_rsc_0_2_qa),
      .wea(twiddle_rsc_0_2_wea),
      .da(twiddle_rsc_0_2_da),
      .adra(twiddle_rsc_0_2_adra),
      .adra_d(nl_twiddle_rsc_0_2_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_2_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_522_8_32_256_256_32_1_gen twiddle_rsc_0_3_i
      (
      .qb(twiddle_rsc_0_3_qb),
      .web(twiddle_rsc_0_3_web),
      .db(twiddle_rsc_0_3_db),
      .adrb(twiddle_rsc_0_3_adrb),
      .qa(twiddle_rsc_0_3_qa),
      .wea(twiddle_rsc_0_3_wea),
      .da(twiddle_rsc_0_3_da),
      .adra(twiddle_rsc_0_3_adra),
      .adra_d(nl_twiddle_rsc_0_3_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_3_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_523_8_32_256_256_32_1_gen twiddle_rsc_0_4_i
      (
      .qb(twiddle_rsc_0_4_qb),
      .web(twiddle_rsc_0_4_web),
      .db(twiddle_rsc_0_4_db),
      .adrb(twiddle_rsc_0_4_adrb),
      .qa(twiddle_rsc_0_4_qa),
      .wea(twiddle_rsc_0_4_wea),
      .da(twiddle_rsc_0_4_da),
      .adra(twiddle_rsc_0_4_adra),
      .adra_d(nl_twiddle_rsc_0_4_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_4_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_524_8_32_256_256_32_1_gen twiddle_rsc_0_5_i
      (
      .qb(twiddle_rsc_0_5_qb),
      .web(twiddle_rsc_0_5_web),
      .db(twiddle_rsc_0_5_db),
      .adrb(twiddle_rsc_0_5_adrb),
      .qa(twiddle_rsc_0_5_qa),
      .wea(twiddle_rsc_0_5_wea),
      .da(twiddle_rsc_0_5_da),
      .adra(twiddle_rsc_0_5_adra),
      .adra_d(nl_twiddle_rsc_0_5_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_5_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_525_8_32_256_256_32_1_gen twiddle_rsc_0_6_i
      (
      .qb(twiddle_rsc_0_6_qb),
      .web(twiddle_rsc_0_6_web),
      .db(twiddle_rsc_0_6_db),
      .adrb(twiddle_rsc_0_6_adrb),
      .qa(twiddle_rsc_0_6_qa),
      .wea(twiddle_rsc_0_6_wea),
      .da(twiddle_rsc_0_6_da),
      .adra(twiddle_rsc_0_6_adra),
      .adra_d(nl_twiddle_rsc_0_6_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_6_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_526_8_32_256_256_32_1_gen twiddle_rsc_0_7_i
      (
      .qb(twiddle_rsc_0_7_qb),
      .web(twiddle_rsc_0_7_web),
      .db(twiddle_rsc_0_7_db),
      .adrb(twiddle_rsc_0_7_adrb),
      .qa(twiddle_rsc_0_7_qa),
      .wea(twiddle_rsc_0_7_wea),
      .da(twiddle_rsc_0_7_da),
      .adra(twiddle_rsc_0_7_adra),
      .adra_d(nl_twiddle_rsc_0_7_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_7_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_527_8_32_256_256_32_1_gen twiddle_rsc_0_8_i
      (
      .qb(twiddle_rsc_0_8_qb),
      .web(twiddle_rsc_0_8_web),
      .db(twiddle_rsc_0_8_db),
      .adrb(twiddle_rsc_0_8_adrb),
      .qa(twiddle_rsc_0_8_qa),
      .wea(twiddle_rsc_0_8_wea),
      .da(twiddle_rsc_0_8_da),
      .adra(twiddle_rsc_0_8_adra),
      .adra_d(nl_twiddle_rsc_0_8_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_8_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_528_8_32_256_256_32_1_gen twiddle_rsc_0_9_i
      (
      .qb(twiddle_rsc_0_9_qb),
      .web(twiddle_rsc_0_9_web),
      .db(twiddle_rsc_0_9_db),
      .adrb(twiddle_rsc_0_9_adrb),
      .qa(twiddle_rsc_0_9_qa),
      .wea(twiddle_rsc_0_9_wea),
      .da(twiddle_rsc_0_9_da),
      .adra(twiddle_rsc_0_9_adra),
      .adra_d(nl_twiddle_rsc_0_9_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_9_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_529_8_32_256_256_32_1_gen twiddle_rsc_0_10_i
      (
      .qb(twiddle_rsc_0_10_qb),
      .web(twiddle_rsc_0_10_web),
      .db(twiddle_rsc_0_10_db),
      .adrb(twiddle_rsc_0_10_adrb),
      .qa(twiddle_rsc_0_10_qa),
      .wea(twiddle_rsc_0_10_wea),
      .da(twiddle_rsc_0_10_da),
      .adra(twiddle_rsc_0_10_adra),
      .adra_d(nl_twiddle_rsc_0_10_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_10_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_530_8_32_256_256_32_1_gen twiddle_rsc_0_11_i
      (
      .qb(twiddle_rsc_0_11_qb),
      .web(twiddle_rsc_0_11_web),
      .db(twiddle_rsc_0_11_db),
      .adrb(twiddle_rsc_0_11_adrb),
      .qa(twiddle_rsc_0_11_qa),
      .wea(twiddle_rsc_0_11_wea),
      .da(twiddle_rsc_0_11_da),
      .adra(twiddle_rsc_0_11_adra),
      .adra_d(nl_twiddle_rsc_0_11_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_11_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_531_8_32_256_256_32_1_gen twiddle_rsc_0_12_i
      (
      .qb(twiddle_rsc_0_12_qb),
      .web(twiddle_rsc_0_12_web),
      .db(twiddle_rsc_0_12_db),
      .adrb(twiddle_rsc_0_12_adrb),
      .qa(twiddle_rsc_0_12_qa),
      .wea(twiddle_rsc_0_12_wea),
      .da(twiddle_rsc_0_12_da),
      .adra(twiddle_rsc_0_12_adra),
      .adra_d(nl_twiddle_rsc_0_12_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_12_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_532_8_32_256_256_32_1_gen twiddle_rsc_0_13_i
      (
      .qb(twiddle_rsc_0_13_qb),
      .web(twiddle_rsc_0_13_web),
      .db(twiddle_rsc_0_13_db),
      .adrb(twiddle_rsc_0_13_adrb),
      .qa(twiddle_rsc_0_13_qa),
      .wea(twiddle_rsc_0_13_wea),
      .da(twiddle_rsc_0_13_da),
      .adra(twiddle_rsc_0_13_adra),
      .adra_d(nl_twiddle_rsc_0_13_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_13_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_533_8_32_256_256_32_1_gen twiddle_rsc_0_14_i
      (
      .qb(twiddle_rsc_0_14_qb),
      .web(twiddle_rsc_0_14_web),
      .db(twiddle_rsc_0_14_db),
      .adrb(twiddle_rsc_0_14_adrb),
      .qa(twiddle_rsc_0_14_qa),
      .wea(twiddle_rsc_0_14_wea),
      .da(twiddle_rsc_0_14_da),
      .adra(twiddle_rsc_0_14_adra),
      .adra_d(nl_twiddle_rsc_0_14_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_14_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_534_8_32_256_256_32_1_gen twiddle_rsc_0_15_i
      (
      .qb(twiddle_rsc_0_15_qb),
      .web(twiddle_rsc_0_15_web),
      .db(twiddle_rsc_0_15_db),
      .adrb(twiddle_rsc_0_15_adrb),
      .qa(twiddle_rsc_0_15_qa),
      .wea(twiddle_rsc_0_15_wea),
      .da(twiddle_rsc_0_15_da),
      .adra(twiddle_rsc_0_15_adra),
      .adra_d(nl_twiddle_rsc_0_15_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_15_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_535_8_32_256_256_32_1_gen twiddle_h_rsc_0_0_i
      (
      .qb(twiddle_h_rsc_0_0_qb),
      .web(twiddle_h_rsc_0_0_web),
      .db(twiddle_h_rsc_0_0_db),
      .adrb(twiddle_h_rsc_0_0_adrb),
      .qa(twiddle_h_rsc_0_0_qa),
      .wea(twiddle_h_rsc_0_0_wea),
      .da(twiddle_h_rsc_0_0_da),
      .adra(twiddle_h_rsc_0_0_adra),
      .adra_d(nl_twiddle_h_rsc_0_0_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_0_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_536_8_32_256_256_32_1_gen twiddle_h_rsc_0_1_i
      (
      .qb(twiddle_h_rsc_0_1_qb),
      .web(twiddle_h_rsc_0_1_web),
      .db(twiddle_h_rsc_0_1_db),
      .adrb(twiddle_h_rsc_0_1_adrb),
      .qa(twiddle_h_rsc_0_1_qa),
      .wea(twiddle_h_rsc_0_1_wea),
      .da(twiddle_h_rsc_0_1_da),
      .adra(twiddle_h_rsc_0_1_adra),
      .adra_d(nl_twiddle_h_rsc_0_1_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_1_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_537_8_32_256_256_32_1_gen twiddle_h_rsc_0_2_i
      (
      .qb(twiddle_h_rsc_0_2_qb),
      .web(twiddle_h_rsc_0_2_web),
      .db(twiddle_h_rsc_0_2_db),
      .adrb(twiddle_h_rsc_0_2_adrb),
      .qa(twiddle_h_rsc_0_2_qa),
      .wea(twiddle_h_rsc_0_2_wea),
      .da(twiddle_h_rsc_0_2_da),
      .adra(twiddle_h_rsc_0_2_adra),
      .adra_d(nl_twiddle_h_rsc_0_2_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_2_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_538_8_32_256_256_32_1_gen twiddle_h_rsc_0_3_i
      (
      .qb(twiddle_h_rsc_0_3_qb),
      .web(twiddle_h_rsc_0_3_web),
      .db(twiddle_h_rsc_0_3_db),
      .adrb(twiddle_h_rsc_0_3_adrb),
      .qa(twiddle_h_rsc_0_3_qa),
      .wea(twiddle_h_rsc_0_3_wea),
      .da(twiddle_h_rsc_0_3_da),
      .adra(twiddle_h_rsc_0_3_adra),
      .adra_d(nl_twiddle_h_rsc_0_3_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_3_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_539_8_32_256_256_32_1_gen twiddle_h_rsc_0_4_i
      (
      .qb(twiddle_h_rsc_0_4_qb),
      .web(twiddle_h_rsc_0_4_web),
      .db(twiddle_h_rsc_0_4_db),
      .adrb(twiddle_h_rsc_0_4_adrb),
      .qa(twiddle_h_rsc_0_4_qa),
      .wea(twiddle_h_rsc_0_4_wea),
      .da(twiddle_h_rsc_0_4_da),
      .adra(twiddle_h_rsc_0_4_adra),
      .adra_d(nl_twiddle_h_rsc_0_4_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_4_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_540_8_32_256_256_32_1_gen twiddle_h_rsc_0_5_i
      (
      .qb(twiddle_h_rsc_0_5_qb),
      .web(twiddle_h_rsc_0_5_web),
      .db(twiddle_h_rsc_0_5_db),
      .adrb(twiddle_h_rsc_0_5_adrb),
      .qa(twiddle_h_rsc_0_5_qa),
      .wea(twiddle_h_rsc_0_5_wea),
      .da(twiddle_h_rsc_0_5_da),
      .adra(twiddle_h_rsc_0_5_adra),
      .adra_d(nl_twiddle_h_rsc_0_5_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_5_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_541_8_32_256_256_32_1_gen twiddle_h_rsc_0_6_i
      (
      .qb(twiddle_h_rsc_0_6_qb),
      .web(twiddle_h_rsc_0_6_web),
      .db(twiddle_h_rsc_0_6_db),
      .adrb(twiddle_h_rsc_0_6_adrb),
      .qa(twiddle_h_rsc_0_6_qa),
      .wea(twiddle_h_rsc_0_6_wea),
      .da(twiddle_h_rsc_0_6_da),
      .adra(twiddle_h_rsc_0_6_adra),
      .adra_d(nl_twiddle_h_rsc_0_6_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_6_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_542_8_32_256_256_32_1_gen twiddle_h_rsc_0_7_i
      (
      .qb(twiddle_h_rsc_0_7_qb),
      .web(twiddle_h_rsc_0_7_web),
      .db(twiddle_h_rsc_0_7_db),
      .adrb(twiddle_h_rsc_0_7_adrb),
      .qa(twiddle_h_rsc_0_7_qa),
      .wea(twiddle_h_rsc_0_7_wea),
      .da(twiddle_h_rsc_0_7_da),
      .adra(twiddle_h_rsc_0_7_adra),
      .adra_d(nl_twiddle_h_rsc_0_7_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_7_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_543_8_32_256_256_32_1_gen twiddle_h_rsc_0_8_i
      (
      .qb(twiddle_h_rsc_0_8_qb),
      .web(twiddle_h_rsc_0_8_web),
      .db(twiddle_h_rsc_0_8_db),
      .adrb(twiddle_h_rsc_0_8_adrb),
      .qa(twiddle_h_rsc_0_8_qa),
      .wea(twiddle_h_rsc_0_8_wea),
      .da(twiddle_h_rsc_0_8_da),
      .adra(twiddle_h_rsc_0_8_adra),
      .adra_d(nl_twiddle_h_rsc_0_8_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_8_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_544_8_32_256_256_32_1_gen twiddle_h_rsc_0_9_i
      (
      .qb(twiddle_h_rsc_0_9_qb),
      .web(twiddle_h_rsc_0_9_web),
      .db(twiddle_h_rsc_0_9_db),
      .adrb(twiddle_h_rsc_0_9_adrb),
      .qa(twiddle_h_rsc_0_9_qa),
      .wea(twiddle_h_rsc_0_9_wea),
      .da(twiddle_h_rsc_0_9_da),
      .adra(twiddle_h_rsc_0_9_adra),
      .adra_d(nl_twiddle_h_rsc_0_9_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_9_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_545_8_32_256_256_32_1_gen twiddle_h_rsc_0_10_i
      (
      .qb(twiddle_h_rsc_0_10_qb),
      .web(twiddle_h_rsc_0_10_web),
      .db(twiddle_h_rsc_0_10_db),
      .adrb(twiddle_h_rsc_0_10_adrb),
      .qa(twiddle_h_rsc_0_10_qa),
      .wea(twiddle_h_rsc_0_10_wea),
      .da(twiddle_h_rsc_0_10_da),
      .adra(twiddle_h_rsc_0_10_adra),
      .adra_d(nl_twiddle_h_rsc_0_10_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_10_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_546_8_32_256_256_32_1_gen twiddle_h_rsc_0_11_i
      (
      .qb(twiddle_h_rsc_0_11_qb),
      .web(twiddle_h_rsc_0_11_web),
      .db(twiddle_h_rsc_0_11_db),
      .adrb(twiddle_h_rsc_0_11_adrb),
      .qa(twiddle_h_rsc_0_11_qa),
      .wea(twiddle_h_rsc_0_11_wea),
      .da(twiddle_h_rsc_0_11_da),
      .adra(twiddle_h_rsc_0_11_adra),
      .adra_d(nl_twiddle_h_rsc_0_11_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_11_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_547_8_32_256_256_32_1_gen twiddle_h_rsc_0_12_i
      (
      .qb(twiddle_h_rsc_0_12_qb),
      .web(twiddle_h_rsc_0_12_web),
      .db(twiddle_h_rsc_0_12_db),
      .adrb(twiddle_h_rsc_0_12_adrb),
      .qa(twiddle_h_rsc_0_12_qa),
      .wea(twiddle_h_rsc_0_12_wea),
      .da(twiddle_h_rsc_0_12_da),
      .adra(twiddle_h_rsc_0_12_adra),
      .adra_d(nl_twiddle_h_rsc_0_12_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_12_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_548_8_32_256_256_32_1_gen twiddle_h_rsc_0_13_i
      (
      .qb(twiddle_h_rsc_0_13_qb),
      .web(twiddle_h_rsc_0_13_web),
      .db(twiddle_h_rsc_0_13_db),
      .adrb(twiddle_h_rsc_0_13_adrb),
      .qa(twiddle_h_rsc_0_13_qa),
      .wea(twiddle_h_rsc_0_13_wea),
      .da(twiddle_h_rsc_0_13_da),
      .adra(twiddle_h_rsc_0_13_adra),
      .adra_d(nl_twiddle_h_rsc_0_13_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_13_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_549_8_32_256_256_32_1_gen twiddle_h_rsc_0_14_i
      (
      .qb(twiddle_h_rsc_0_14_qb),
      .web(twiddle_h_rsc_0_14_web),
      .db(twiddle_h_rsc_0_14_db),
      .adrb(twiddle_h_rsc_0_14_adrb),
      .qa(twiddle_h_rsc_0_14_qa),
      .wea(twiddle_h_rsc_0_14_wea),
      .da(twiddle_h_rsc_0_14_da),
      .adra(twiddle_h_rsc_0_14_adra),
      .adra_d(nl_twiddle_h_rsc_0_14_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_14_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_550_8_32_256_256_32_1_gen twiddle_h_rsc_0_15_i
      (
      .qb(twiddle_h_rsc_0_15_qb),
      .web(twiddle_h_rsc_0_15_web),
      .db(twiddle_h_rsc_0_15_db),
      .adrb(twiddle_h_rsc_0_15_adrb),
      .qa(twiddle_h_rsc_0_15_qa),
      .wea(twiddle_h_rsc_0_15_wea),
      .da(twiddle_h_rsc_0_15_da),
      .adra(twiddle_h_rsc_0_15_adra),
      .adra_d(nl_twiddle_h_rsc_0_15_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_15_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_core peaseNTT_core_inst (
      .clk(clk),
      .rst(rst),
      .xt_rsc_triosy_0_0_lz(xt_rsc_triosy_0_0_lz),
      .xt_rsc_triosy_0_1_lz(xt_rsc_triosy_0_1_lz),
      .xt_rsc_triosy_0_2_lz(xt_rsc_triosy_0_2_lz),
      .xt_rsc_triosy_0_3_lz(xt_rsc_triosy_0_3_lz),
      .xt_rsc_triosy_0_4_lz(xt_rsc_triosy_0_4_lz),
      .xt_rsc_triosy_0_5_lz(xt_rsc_triosy_0_5_lz),
      .xt_rsc_triosy_0_6_lz(xt_rsc_triosy_0_6_lz),
      .xt_rsc_triosy_0_7_lz(xt_rsc_triosy_0_7_lz),
      .xt_rsc_triosy_0_8_lz(xt_rsc_triosy_0_8_lz),
      .xt_rsc_triosy_0_9_lz(xt_rsc_triosy_0_9_lz),
      .xt_rsc_triosy_0_10_lz(xt_rsc_triosy_0_10_lz),
      .xt_rsc_triosy_0_11_lz(xt_rsc_triosy_0_11_lz),
      .xt_rsc_triosy_0_12_lz(xt_rsc_triosy_0_12_lz),
      .xt_rsc_triosy_0_13_lz(xt_rsc_triosy_0_13_lz),
      .xt_rsc_triosy_0_14_lz(xt_rsc_triosy_0_14_lz),
      .xt_rsc_triosy_0_15_lz(xt_rsc_triosy_0_15_lz),
      .xt_rsc_triosy_0_16_lz(xt_rsc_triosy_0_16_lz),
      .xt_rsc_triosy_0_17_lz(xt_rsc_triosy_0_17_lz),
      .xt_rsc_triosy_0_18_lz(xt_rsc_triosy_0_18_lz),
      .xt_rsc_triosy_0_19_lz(xt_rsc_triosy_0_19_lz),
      .xt_rsc_triosy_0_20_lz(xt_rsc_triosy_0_20_lz),
      .xt_rsc_triosy_0_21_lz(xt_rsc_triosy_0_21_lz),
      .xt_rsc_triosy_0_22_lz(xt_rsc_triosy_0_22_lz),
      .xt_rsc_triosy_0_23_lz(xt_rsc_triosy_0_23_lz),
      .xt_rsc_triosy_0_24_lz(xt_rsc_triosy_0_24_lz),
      .xt_rsc_triosy_0_25_lz(xt_rsc_triosy_0_25_lz),
      .xt_rsc_triosy_0_26_lz(xt_rsc_triosy_0_26_lz),
      .xt_rsc_triosy_0_27_lz(xt_rsc_triosy_0_27_lz),
      .xt_rsc_triosy_0_28_lz(xt_rsc_triosy_0_28_lz),
      .xt_rsc_triosy_0_29_lz(xt_rsc_triosy_0_29_lz),
      .xt_rsc_triosy_0_30_lz(xt_rsc_triosy_0_30_lz),
      .xt_rsc_triosy_0_31_lz(xt_rsc_triosy_0_31_lz),
      .xt_rsc_triosy_1_0_lz(xt_rsc_triosy_1_0_lz),
      .xt_rsc_triosy_1_1_lz(xt_rsc_triosy_1_1_lz),
      .xt_rsc_triosy_1_2_lz(xt_rsc_triosy_1_2_lz),
      .xt_rsc_triosy_1_3_lz(xt_rsc_triosy_1_3_lz),
      .xt_rsc_triosy_1_4_lz(xt_rsc_triosy_1_4_lz),
      .xt_rsc_triosy_1_5_lz(xt_rsc_triosy_1_5_lz),
      .xt_rsc_triosy_1_6_lz(xt_rsc_triosy_1_6_lz),
      .xt_rsc_triosy_1_7_lz(xt_rsc_triosy_1_7_lz),
      .xt_rsc_triosy_1_8_lz(xt_rsc_triosy_1_8_lz),
      .xt_rsc_triosy_1_9_lz(xt_rsc_triosy_1_9_lz),
      .xt_rsc_triosy_1_10_lz(xt_rsc_triosy_1_10_lz),
      .xt_rsc_triosy_1_11_lz(xt_rsc_triosy_1_11_lz),
      .xt_rsc_triosy_1_12_lz(xt_rsc_triosy_1_12_lz),
      .xt_rsc_triosy_1_13_lz(xt_rsc_triosy_1_13_lz),
      .xt_rsc_triosy_1_14_lz(xt_rsc_triosy_1_14_lz),
      .xt_rsc_triosy_1_15_lz(xt_rsc_triosy_1_15_lz),
      .xt_rsc_triosy_1_16_lz(xt_rsc_triosy_1_16_lz),
      .xt_rsc_triosy_1_17_lz(xt_rsc_triosy_1_17_lz),
      .xt_rsc_triosy_1_18_lz(xt_rsc_triosy_1_18_lz),
      .xt_rsc_triosy_1_19_lz(xt_rsc_triosy_1_19_lz),
      .xt_rsc_triosy_1_20_lz(xt_rsc_triosy_1_20_lz),
      .xt_rsc_triosy_1_21_lz(xt_rsc_triosy_1_21_lz),
      .xt_rsc_triosy_1_22_lz(xt_rsc_triosy_1_22_lz),
      .xt_rsc_triosy_1_23_lz(xt_rsc_triosy_1_23_lz),
      .xt_rsc_triosy_1_24_lz(xt_rsc_triosy_1_24_lz),
      .xt_rsc_triosy_1_25_lz(xt_rsc_triosy_1_25_lz),
      .xt_rsc_triosy_1_26_lz(xt_rsc_triosy_1_26_lz),
      .xt_rsc_triosy_1_27_lz(xt_rsc_triosy_1_27_lz),
      .xt_rsc_triosy_1_28_lz(xt_rsc_triosy_1_28_lz),
      .xt_rsc_triosy_1_29_lz(xt_rsc_triosy_1_29_lz),
      .xt_rsc_triosy_1_30_lz(xt_rsc_triosy_1_30_lz),
      .xt_rsc_triosy_1_31_lz(xt_rsc_triosy_1_31_lz),
      .xt_rsc_triosy_2_0_lz(xt_rsc_triosy_2_0_lz),
      .xt_rsc_triosy_2_1_lz(xt_rsc_triosy_2_1_lz),
      .xt_rsc_triosy_2_2_lz(xt_rsc_triosy_2_2_lz),
      .xt_rsc_triosy_2_3_lz(xt_rsc_triosy_2_3_lz),
      .xt_rsc_triosy_2_4_lz(xt_rsc_triosy_2_4_lz),
      .xt_rsc_triosy_2_5_lz(xt_rsc_triosy_2_5_lz),
      .xt_rsc_triosy_2_6_lz(xt_rsc_triosy_2_6_lz),
      .xt_rsc_triosy_2_7_lz(xt_rsc_triosy_2_7_lz),
      .xt_rsc_triosy_2_8_lz(xt_rsc_triosy_2_8_lz),
      .xt_rsc_triosy_2_9_lz(xt_rsc_triosy_2_9_lz),
      .xt_rsc_triosy_2_10_lz(xt_rsc_triosy_2_10_lz),
      .xt_rsc_triosy_2_11_lz(xt_rsc_triosy_2_11_lz),
      .xt_rsc_triosy_2_12_lz(xt_rsc_triosy_2_12_lz),
      .xt_rsc_triosy_2_13_lz(xt_rsc_triosy_2_13_lz),
      .xt_rsc_triosy_2_14_lz(xt_rsc_triosy_2_14_lz),
      .xt_rsc_triosy_2_15_lz(xt_rsc_triosy_2_15_lz),
      .xt_rsc_triosy_2_16_lz(xt_rsc_triosy_2_16_lz),
      .xt_rsc_triosy_2_17_lz(xt_rsc_triosy_2_17_lz),
      .xt_rsc_triosy_2_18_lz(xt_rsc_triosy_2_18_lz),
      .xt_rsc_triosy_2_19_lz(xt_rsc_triosy_2_19_lz),
      .xt_rsc_triosy_2_20_lz(xt_rsc_triosy_2_20_lz),
      .xt_rsc_triosy_2_21_lz(xt_rsc_triosy_2_21_lz),
      .xt_rsc_triosy_2_22_lz(xt_rsc_triosy_2_22_lz),
      .xt_rsc_triosy_2_23_lz(xt_rsc_triosy_2_23_lz),
      .xt_rsc_triosy_2_24_lz(xt_rsc_triosy_2_24_lz),
      .xt_rsc_triosy_2_25_lz(xt_rsc_triosy_2_25_lz),
      .xt_rsc_triosy_2_26_lz(xt_rsc_triosy_2_26_lz),
      .xt_rsc_triosy_2_27_lz(xt_rsc_triosy_2_27_lz),
      .xt_rsc_triosy_2_28_lz(xt_rsc_triosy_2_28_lz),
      .xt_rsc_triosy_2_29_lz(xt_rsc_triosy_2_29_lz),
      .xt_rsc_triosy_2_30_lz(xt_rsc_triosy_2_30_lz),
      .xt_rsc_triosy_2_31_lz(xt_rsc_triosy_2_31_lz),
      .xt_rsc_triosy_3_0_lz(xt_rsc_triosy_3_0_lz),
      .xt_rsc_triosy_3_1_lz(xt_rsc_triosy_3_1_lz),
      .xt_rsc_triosy_3_2_lz(xt_rsc_triosy_3_2_lz),
      .xt_rsc_triosy_3_3_lz(xt_rsc_triosy_3_3_lz),
      .xt_rsc_triosy_3_4_lz(xt_rsc_triosy_3_4_lz),
      .xt_rsc_triosy_3_5_lz(xt_rsc_triosy_3_5_lz),
      .xt_rsc_triosy_3_6_lz(xt_rsc_triosy_3_6_lz),
      .xt_rsc_triosy_3_7_lz(xt_rsc_triosy_3_7_lz),
      .xt_rsc_triosy_3_8_lz(xt_rsc_triosy_3_8_lz),
      .xt_rsc_triosy_3_9_lz(xt_rsc_triosy_3_9_lz),
      .xt_rsc_triosy_3_10_lz(xt_rsc_triosy_3_10_lz),
      .xt_rsc_triosy_3_11_lz(xt_rsc_triosy_3_11_lz),
      .xt_rsc_triosy_3_12_lz(xt_rsc_triosy_3_12_lz),
      .xt_rsc_triosy_3_13_lz(xt_rsc_triosy_3_13_lz),
      .xt_rsc_triosy_3_14_lz(xt_rsc_triosy_3_14_lz),
      .xt_rsc_triosy_3_15_lz(xt_rsc_triosy_3_15_lz),
      .xt_rsc_triosy_3_16_lz(xt_rsc_triosy_3_16_lz),
      .xt_rsc_triosy_3_17_lz(xt_rsc_triosy_3_17_lz),
      .xt_rsc_triosy_3_18_lz(xt_rsc_triosy_3_18_lz),
      .xt_rsc_triosy_3_19_lz(xt_rsc_triosy_3_19_lz),
      .xt_rsc_triosy_3_20_lz(xt_rsc_triosy_3_20_lz),
      .xt_rsc_triosy_3_21_lz(xt_rsc_triosy_3_21_lz),
      .xt_rsc_triosy_3_22_lz(xt_rsc_triosy_3_22_lz),
      .xt_rsc_triosy_3_23_lz(xt_rsc_triosy_3_23_lz),
      .xt_rsc_triosy_3_24_lz(xt_rsc_triosy_3_24_lz),
      .xt_rsc_triosy_3_25_lz(xt_rsc_triosy_3_25_lz),
      .xt_rsc_triosy_3_26_lz(xt_rsc_triosy_3_26_lz),
      .xt_rsc_triosy_3_27_lz(xt_rsc_triosy_3_27_lz),
      .xt_rsc_triosy_3_28_lz(xt_rsc_triosy_3_28_lz),
      .xt_rsc_triosy_3_29_lz(xt_rsc_triosy_3_29_lz),
      .xt_rsc_triosy_3_30_lz(xt_rsc_triosy_3_30_lz),
      .xt_rsc_triosy_3_31_lz(xt_rsc_triosy_3_31_lz),
      .xt_rsc_triosy_4_0_lz(xt_rsc_triosy_4_0_lz),
      .xt_rsc_triosy_4_1_lz(xt_rsc_triosy_4_1_lz),
      .xt_rsc_triosy_4_2_lz(xt_rsc_triosy_4_2_lz),
      .xt_rsc_triosy_4_3_lz(xt_rsc_triosy_4_3_lz),
      .xt_rsc_triosy_4_4_lz(xt_rsc_triosy_4_4_lz),
      .xt_rsc_triosy_4_5_lz(xt_rsc_triosy_4_5_lz),
      .xt_rsc_triosy_4_6_lz(xt_rsc_triosy_4_6_lz),
      .xt_rsc_triosy_4_7_lz(xt_rsc_triosy_4_7_lz),
      .xt_rsc_triosy_4_8_lz(xt_rsc_triosy_4_8_lz),
      .xt_rsc_triosy_4_9_lz(xt_rsc_triosy_4_9_lz),
      .xt_rsc_triosy_4_10_lz(xt_rsc_triosy_4_10_lz),
      .xt_rsc_triosy_4_11_lz(xt_rsc_triosy_4_11_lz),
      .xt_rsc_triosy_4_12_lz(xt_rsc_triosy_4_12_lz),
      .xt_rsc_triosy_4_13_lz(xt_rsc_triosy_4_13_lz),
      .xt_rsc_triosy_4_14_lz(xt_rsc_triosy_4_14_lz),
      .xt_rsc_triosy_4_15_lz(xt_rsc_triosy_4_15_lz),
      .xt_rsc_triosy_4_16_lz(xt_rsc_triosy_4_16_lz),
      .xt_rsc_triosy_4_17_lz(xt_rsc_triosy_4_17_lz),
      .xt_rsc_triosy_4_18_lz(xt_rsc_triosy_4_18_lz),
      .xt_rsc_triosy_4_19_lz(xt_rsc_triosy_4_19_lz),
      .xt_rsc_triosy_4_20_lz(xt_rsc_triosy_4_20_lz),
      .xt_rsc_triosy_4_21_lz(xt_rsc_triosy_4_21_lz),
      .xt_rsc_triosy_4_22_lz(xt_rsc_triosy_4_22_lz),
      .xt_rsc_triosy_4_23_lz(xt_rsc_triosy_4_23_lz),
      .xt_rsc_triosy_4_24_lz(xt_rsc_triosy_4_24_lz),
      .xt_rsc_triosy_4_25_lz(xt_rsc_triosy_4_25_lz),
      .xt_rsc_triosy_4_26_lz(xt_rsc_triosy_4_26_lz),
      .xt_rsc_triosy_4_27_lz(xt_rsc_triosy_4_27_lz),
      .xt_rsc_triosy_4_28_lz(xt_rsc_triosy_4_28_lz),
      .xt_rsc_triosy_4_29_lz(xt_rsc_triosy_4_29_lz),
      .xt_rsc_triosy_4_30_lz(xt_rsc_triosy_4_30_lz),
      .xt_rsc_triosy_4_31_lz(xt_rsc_triosy_4_31_lz),
      .xt_rsc_triosy_5_0_lz(xt_rsc_triosy_5_0_lz),
      .xt_rsc_triosy_5_1_lz(xt_rsc_triosy_5_1_lz),
      .xt_rsc_triosy_5_2_lz(xt_rsc_triosy_5_2_lz),
      .xt_rsc_triosy_5_3_lz(xt_rsc_triosy_5_3_lz),
      .xt_rsc_triosy_5_4_lz(xt_rsc_triosy_5_4_lz),
      .xt_rsc_triosy_5_5_lz(xt_rsc_triosy_5_5_lz),
      .xt_rsc_triosy_5_6_lz(xt_rsc_triosy_5_6_lz),
      .xt_rsc_triosy_5_7_lz(xt_rsc_triosy_5_7_lz),
      .xt_rsc_triosy_5_8_lz(xt_rsc_triosy_5_8_lz),
      .xt_rsc_triosy_5_9_lz(xt_rsc_triosy_5_9_lz),
      .xt_rsc_triosy_5_10_lz(xt_rsc_triosy_5_10_lz),
      .xt_rsc_triosy_5_11_lz(xt_rsc_triosy_5_11_lz),
      .xt_rsc_triosy_5_12_lz(xt_rsc_triosy_5_12_lz),
      .xt_rsc_triosy_5_13_lz(xt_rsc_triosy_5_13_lz),
      .xt_rsc_triosy_5_14_lz(xt_rsc_triosy_5_14_lz),
      .xt_rsc_triosy_5_15_lz(xt_rsc_triosy_5_15_lz),
      .xt_rsc_triosy_5_16_lz(xt_rsc_triosy_5_16_lz),
      .xt_rsc_triosy_5_17_lz(xt_rsc_triosy_5_17_lz),
      .xt_rsc_triosy_5_18_lz(xt_rsc_triosy_5_18_lz),
      .xt_rsc_triosy_5_19_lz(xt_rsc_triosy_5_19_lz),
      .xt_rsc_triosy_5_20_lz(xt_rsc_triosy_5_20_lz),
      .xt_rsc_triosy_5_21_lz(xt_rsc_triosy_5_21_lz),
      .xt_rsc_triosy_5_22_lz(xt_rsc_triosy_5_22_lz),
      .xt_rsc_triosy_5_23_lz(xt_rsc_triosy_5_23_lz),
      .xt_rsc_triosy_5_24_lz(xt_rsc_triosy_5_24_lz),
      .xt_rsc_triosy_5_25_lz(xt_rsc_triosy_5_25_lz),
      .xt_rsc_triosy_5_26_lz(xt_rsc_triosy_5_26_lz),
      .xt_rsc_triosy_5_27_lz(xt_rsc_triosy_5_27_lz),
      .xt_rsc_triosy_5_28_lz(xt_rsc_triosy_5_28_lz),
      .xt_rsc_triosy_5_29_lz(xt_rsc_triosy_5_29_lz),
      .xt_rsc_triosy_5_30_lz(xt_rsc_triosy_5_30_lz),
      .xt_rsc_triosy_5_31_lz(xt_rsc_triosy_5_31_lz),
      .xt_rsc_triosy_6_0_lz(xt_rsc_triosy_6_0_lz),
      .xt_rsc_triosy_6_1_lz(xt_rsc_triosy_6_1_lz),
      .xt_rsc_triosy_6_2_lz(xt_rsc_triosy_6_2_lz),
      .xt_rsc_triosy_6_3_lz(xt_rsc_triosy_6_3_lz),
      .xt_rsc_triosy_6_4_lz(xt_rsc_triosy_6_4_lz),
      .xt_rsc_triosy_6_5_lz(xt_rsc_triosy_6_5_lz),
      .xt_rsc_triosy_6_6_lz(xt_rsc_triosy_6_6_lz),
      .xt_rsc_triosy_6_7_lz(xt_rsc_triosy_6_7_lz),
      .xt_rsc_triosy_6_8_lz(xt_rsc_triosy_6_8_lz),
      .xt_rsc_triosy_6_9_lz(xt_rsc_triosy_6_9_lz),
      .xt_rsc_triosy_6_10_lz(xt_rsc_triosy_6_10_lz),
      .xt_rsc_triosy_6_11_lz(xt_rsc_triosy_6_11_lz),
      .xt_rsc_triosy_6_12_lz(xt_rsc_triosy_6_12_lz),
      .xt_rsc_triosy_6_13_lz(xt_rsc_triosy_6_13_lz),
      .xt_rsc_triosy_6_14_lz(xt_rsc_triosy_6_14_lz),
      .xt_rsc_triosy_6_15_lz(xt_rsc_triosy_6_15_lz),
      .xt_rsc_triosy_6_16_lz(xt_rsc_triosy_6_16_lz),
      .xt_rsc_triosy_6_17_lz(xt_rsc_triosy_6_17_lz),
      .xt_rsc_triosy_6_18_lz(xt_rsc_triosy_6_18_lz),
      .xt_rsc_triosy_6_19_lz(xt_rsc_triosy_6_19_lz),
      .xt_rsc_triosy_6_20_lz(xt_rsc_triosy_6_20_lz),
      .xt_rsc_triosy_6_21_lz(xt_rsc_triosy_6_21_lz),
      .xt_rsc_triosy_6_22_lz(xt_rsc_triosy_6_22_lz),
      .xt_rsc_triosy_6_23_lz(xt_rsc_triosy_6_23_lz),
      .xt_rsc_triosy_6_24_lz(xt_rsc_triosy_6_24_lz),
      .xt_rsc_triosy_6_25_lz(xt_rsc_triosy_6_25_lz),
      .xt_rsc_triosy_6_26_lz(xt_rsc_triosy_6_26_lz),
      .xt_rsc_triosy_6_27_lz(xt_rsc_triosy_6_27_lz),
      .xt_rsc_triosy_6_28_lz(xt_rsc_triosy_6_28_lz),
      .xt_rsc_triosy_6_29_lz(xt_rsc_triosy_6_29_lz),
      .xt_rsc_triosy_6_30_lz(xt_rsc_triosy_6_30_lz),
      .xt_rsc_triosy_6_31_lz(xt_rsc_triosy_6_31_lz),
      .xt_rsc_triosy_7_0_lz(xt_rsc_triosy_7_0_lz),
      .xt_rsc_triosy_7_1_lz(xt_rsc_triosy_7_1_lz),
      .xt_rsc_triosy_7_2_lz(xt_rsc_triosy_7_2_lz),
      .xt_rsc_triosy_7_3_lz(xt_rsc_triosy_7_3_lz),
      .xt_rsc_triosy_7_4_lz(xt_rsc_triosy_7_4_lz),
      .xt_rsc_triosy_7_5_lz(xt_rsc_triosy_7_5_lz),
      .xt_rsc_triosy_7_6_lz(xt_rsc_triosy_7_6_lz),
      .xt_rsc_triosy_7_7_lz(xt_rsc_triosy_7_7_lz),
      .xt_rsc_triosy_7_8_lz(xt_rsc_triosy_7_8_lz),
      .xt_rsc_triosy_7_9_lz(xt_rsc_triosy_7_9_lz),
      .xt_rsc_triosy_7_10_lz(xt_rsc_triosy_7_10_lz),
      .xt_rsc_triosy_7_11_lz(xt_rsc_triosy_7_11_lz),
      .xt_rsc_triosy_7_12_lz(xt_rsc_triosy_7_12_lz),
      .xt_rsc_triosy_7_13_lz(xt_rsc_triosy_7_13_lz),
      .xt_rsc_triosy_7_14_lz(xt_rsc_triosy_7_14_lz),
      .xt_rsc_triosy_7_15_lz(xt_rsc_triosy_7_15_lz),
      .xt_rsc_triosy_7_16_lz(xt_rsc_triosy_7_16_lz),
      .xt_rsc_triosy_7_17_lz(xt_rsc_triosy_7_17_lz),
      .xt_rsc_triosy_7_18_lz(xt_rsc_triosy_7_18_lz),
      .xt_rsc_triosy_7_19_lz(xt_rsc_triosy_7_19_lz),
      .xt_rsc_triosy_7_20_lz(xt_rsc_triosy_7_20_lz),
      .xt_rsc_triosy_7_21_lz(xt_rsc_triosy_7_21_lz),
      .xt_rsc_triosy_7_22_lz(xt_rsc_triosy_7_22_lz),
      .xt_rsc_triosy_7_23_lz(xt_rsc_triosy_7_23_lz),
      .xt_rsc_triosy_7_24_lz(xt_rsc_triosy_7_24_lz),
      .xt_rsc_triosy_7_25_lz(xt_rsc_triosy_7_25_lz),
      .xt_rsc_triosy_7_26_lz(xt_rsc_triosy_7_26_lz),
      .xt_rsc_triosy_7_27_lz(xt_rsc_triosy_7_27_lz),
      .xt_rsc_triosy_7_28_lz(xt_rsc_triosy_7_28_lz),
      .xt_rsc_triosy_7_29_lz(xt_rsc_triosy_7_29_lz),
      .xt_rsc_triosy_7_30_lz(xt_rsc_triosy_7_30_lz),
      .xt_rsc_triosy_7_31_lz(xt_rsc_triosy_7_31_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_0_0_lz(twiddle_rsc_triosy_0_0_lz),
      .twiddle_rsc_triosy_0_1_lz(twiddle_rsc_triosy_0_1_lz),
      .twiddle_rsc_triosy_0_2_lz(twiddle_rsc_triosy_0_2_lz),
      .twiddle_rsc_triosy_0_3_lz(twiddle_rsc_triosy_0_3_lz),
      .twiddle_rsc_triosy_0_4_lz(twiddle_rsc_triosy_0_4_lz),
      .twiddle_rsc_triosy_0_5_lz(twiddle_rsc_triosy_0_5_lz),
      .twiddle_rsc_triosy_0_6_lz(twiddle_rsc_triosy_0_6_lz),
      .twiddle_rsc_triosy_0_7_lz(twiddle_rsc_triosy_0_7_lz),
      .twiddle_rsc_triosy_0_8_lz(twiddle_rsc_triosy_0_8_lz),
      .twiddle_rsc_triosy_0_9_lz(twiddle_rsc_triosy_0_9_lz),
      .twiddle_rsc_triosy_0_10_lz(twiddle_rsc_triosy_0_10_lz),
      .twiddle_rsc_triosy_0_11_lz(twiddle_rsc_triosy_0_11_lz),
      .twiddle_rsc_triosy_0_12_lz(twiddle_rsc_triosy_0_12_lz),
      .twiddle_rsc_triosy_0_13_lz(twiddle_rsc_triosy_0_13_lz),
      .twiddle_rsc_triosy_0_14_lz(twiddle_rsc_triosy_0_14_lz),
      .twiddle_rsc_triosy_0_15_lz(twiddle_rsc_triosy_0_15_lz),
      .twiddle_h_rsc_triosy_0_0_lz(twiddle_h_rsc_triosy_0_0_lz),
      .twiddle_h_rsc_triosy_0_1_lz(twiddle_h_rsc_triosy_0_1_lz),
      .twiddle_h_rsc_triosy_0_2_lz(twiddle_h_rsc_triosy_0_2_lz),
      .twiddle_h_rsc_triosy_0_3_lz(twiddle_h_rsc_triosy_0_3_lz),
      .twiddle_h_rsc_triosy_0_4_lz(twiddle_h_rsc_triosy_0_4_lz),
      .twiddle_h_rsc_triosy_0_5_lz(twiddle_h_rsc_triosy_0_5_lz),
      .twiddle_h_rsc_triosy_0_6_lz(twiddle_h_rsc_triosy_0_6_lz),
      .twiddle_h_rsc_triosy_0_7_lz(twiddle_h_rsc_triosy_0_7_lz),
      .twiddle_h_rsc_triosy_0_8_lz(twiddle_h_rsc_triosy_0_8_lz),
      .twiddle_h_rsc_triosy_0_9_lz(twiddle_h_rsc_triosy_0_9_lz),
      .twiddle_h_rsc_triosy_0_10_lz(twiddle_h_rsc_triosy_0_10_lz),
      .twiddle_h_rsc_triosy_0_11_lz(twiddle_h_rsc_triosy_0_11_lz),
      .twiddle_h_rsc_triosy_0_12_lz(twiddle_h_rsc_triosy_0_12_lz),
      .twiddle_h_rsc_triosy_0_13_lz(twiddle_h_rsc_triosy_0_13_lz),
      .twiddle_h_rsc_triosy_0_14_lz(twiddle_h_rsc_triosy_0_14_lz),
      .twiddle_h_rsc_triosy_0_15_lz(twiddle_h_rsc_triosy_0_15_lz),
      .yt_rsc_0_0_i_clkr_en_d(yt_rsc_0_0_i_clkr_en_d),
      .yt_rsc_0_0_i_q_d(yt_rsc_0_0_i_q_d),
      .yt_rsc_0_1_i_q_d(yt_rsc_0_1_i_q_d),
      .yt_rsc_0_2_i_q_d(yt_rsc_0_2_i_q_d),
      .yt_rsc_0_3_i_q_d(yt_rsc_0_3_i_q_d),
      .yt_rsc_0_4_i_q_d(yt_rsc_0_4_i_q_d),
      .yt_rsc_0_5_i_q_d(yt_rsc_0_5_i_q_d),
      .yt_rsc_0_6_i_q_d(yt_rsc_0_6_i_q_d),
      .yt_rsc_0_7_i_q_d(yt_rsc_0_7_i_q_d),
      .yt_rsc_0_8_i_q_d(yt_rsc_0_8_i_q_d),
      .yt_rsc_0_9_i_q_d(yt_rsc_0_9_i_q_d),
      .yt_rsc_0_10_i_q_d(yt_rsc_0_10_i_q_d),
      .yt_rsc_0_11_i_q_d(yt_rsc_0_11_i_q_d),
      .yt_rsc_0_12_i_q_d(yt_rsc_0_12_i_q_d),
      .yt_rsc_0_13_i_q_d(yt_rsc_0_13_i_q_d),
      .yt_rsc_0_14_i_q_d(yt_rsc_0_14_i_q_d),
      .yt_rsc_0_15_i_q_d(yt_rsc_0_15_i_q_d),
      .yt_rsc_0_16_i_clkr_en_d(yt_rsc_0_16_i_clkr_en_d),
      .yt_rsc_0_16_i_q_d(yt_rsc_0_16_i_q_d),
      .yt_rsc_0_17_i_q_d(yt_rsc_0_17_i_q_d),
      .yt_rsc_0_18_i_q_d(yt_rsc_0_18_i_q_d),
      .yt_rsc_0_19_i_q_d(yt_rsc_0_19_i_q_d),
      .yt_rsc_0_20_i_q_d(yt_rsc_0_20_i_q_d),
      .yt_rsc_0_21_i_q_d(yt_rsc_0_21_i_q_d),
      .yt_rsc_0_22_i_q_d(yt_rsc_0_22_i_q_d),
      .yt_rsc_0_23_i_q_d(yt_rsc_0_23_i_q_d),
      .yt_rsc_0_24_i_q_d(yt_rsc_0_24_i_q_d),
      .yt_rsc_0_25_i_q_d(yt_rsc_0_25_i_q_d),
      .yt_rsc_0_26_i_q_d(yt_rsc_0_26_i_q_d),
      .yt_rsc_0_27_i_q_d(yt_rsc_0_27_i_q_d),
      .yt_rsc_0_28_i_q_d(yt_rsc_0_28_i_q_d),
      .yt_rsc_0_29_i_q_d(yt_rsc_0_29_i_q_d),
      .yt_rsc_0_30_i_q_d(yt_rsc_0_30_i_q_d),
      .yt_rsc_0_31_i_q_d(yt_rsc_0_31_i_q_d),
      .yt_rsc_1_0_i_clkr_en_d(yt_rsc_1_0_i_clkr_en_d),
      .yt_rsc_1_0_i_q_d(yt_rsc_1_0_i_q_d),
      .yt_rsc_1_1_i_q_d(yt_rsc_1_1_i_q_d),
      .yt_rsc_1_2_i_q_d(yt_rsc_1_2_i_q_d),
      .yt_rsc_1_3_i_q_d(yt_rsc_1_3_i_q_d),
      .yt_rsc_1_4_i_q_d(yt_rsc_1_4_i_q_d),
      .yt_rsc_1_5_i_q_d(yt_rsc_1_5_i_q_d),
      .yt_rsc_1_6_i_q_d(yt_rsc_1_6_i_q_d),
      .yt_rsc_1_7_i_q_d(yt_rsc_1_7_i_q_d),
      .yt_rsc_1_8_i_q_d(yt_rsc_1_8_i_q_d),
      .yt_rsc_1_9_i_q_d(yt_rsc_1_9_i_q_d),
      .yt_rsc_1_10_i_q_d(yt_rsc_1_10_i_q_d),
      .yt_rsc_1_11_i_q_d(yt_rsc_1_11_i_q_d),
      .yt_rsc_1_12_i_q_d(yt_rsc_1_12_i_q_d),
      .yt_rsc_1_13_i_q_d(yt_rsc_1_13_i_q_d),
      .yt_rsc_1_14_i_q_d(yt_rsc_1_14_i_q_d),
      .yt_rsc_1_15_i_q_d(yt_rsc_1_15_i_q_d),
      .yt_rsc_1_16_i_clkr_en_d(yt_rsc_1_16_i_clkr_en_d),
      .yt_rsc_1_16_i_q_d(yt_rsc_1_16_i_q_d),
      .yt_rsc_1_17_i_q_d(yt_rsc_1_17_i_q_d),
      .yt_rsc_1_18_i_q_d(yt_rsc_1_18_i_q_d),
      .yt_rsc_1_19_i_q_d(yt_rsc_1_19_i_q_d),
      .yt_rsc_1_20_i_q_d(yt_rsc_1_20_i_q_d),
      .yt_rsc_1_21_i_q_d(yt_rsc_1_21_i_q_d),
      .yt_rsc_1_22_i_q_d(yt_rsc_1_22_i_q_d),
      .yt_rsc_1_23_i_q_d(yt_rsc_1_23_i_q_d),
      .yt_rsc_1_24_i_q_d(yt_rsc_1_24_i_q_d),
      .yt_rsc_1_25_i_q_d(yt_rsc_1_25_i_q_d),
      .yt_rsc_1_26_i_q_d(yt_rsc_1_26_i_q_d),
      .yt_rsc_1_27_i_q_d(yt_rsc_1_27_i_q_d),
      .yt_rsc_1_28_i_q_d(yt_rsc_1_28_i_q_d),
      .yt_rsc_1_29_i_q_d(yt_rsc_1_29_i_q_d),
      .yt_rsc_1_30_i_q_d(yt_rsc_1_30_i_q_d),
      .yt_rsc_1_31_i_q_d(yt_rsc_1_31_i_q_d),
      .yt_rsc_2_0_i_clkr_en_d(yt_rsc_2_0_i_clkr_en_d),
      .yt_rsc_2_0_i_q_d(yt_rsc_2_0_i_q_d),
      .yt_rsc_2_1_i_q_d(yt_rsc_2_1_i_q_d),
      .yt_rsc_2_2_i_q_d(yt_rsc_2_2_i_q_d),
      .yt_rsc_2_3_i_q_d(yt_rsc_2_3_i_q_d),
      .yt_rsc_2_4_i_q_d(yt_rsc_2_4_i_q_d),
      .yt_rsc_2_5_i_q_d(yt_rsc_2_5_i_q_d),
      .yt_rsc_2_6_i_q_d(yt_rsc_2_6_i_q_d),
      .yt_rsc_2_7_i_q_d(yt_rsc_2_7_i_q_d),
      .yt_rsc_2_8_i_q_d(yt_rsc_2_8_i_q_d),
      .yt_rsc_2_9_i_q_d(yt_rsc_2_9_i_q_d),
      .yt_rsc_2_10_i_q_d(yt_rsc_2_10_i_q_d),
      .yt_rsc_2_11_i_q_d(yt_rsc_2_11_i_q_d),
      .yt_rsc_2_12_i_q_d(yt_rsc_2_12_i_q_d),
      .yt_rsc_2_13_i_q_d(yt_rsc_2_13_i_q_d),
      .yt_rsc_2_14_i_q_d(yt_rsc_2_14_i_q_d),
      .yt_rsc_2_15_i_q_d(yt_rsc_2_15_i_q_d),
      .yt_rsc_2_16_i_clkr_en_d(yt_rsc_2_16_i_clkr_en_d),
      .yt_rsc_2_16_i_q_d(yt_rsc_2_16_i_q_d),
      .yt_rsc_2_17_i_q_d(yt_rsc_2_17_i_q_d),
      .yt_rsc_2_18_i_q_d(yt_rsc_2_18_i_q_d),
      .yt_rsc_2_19_i_q_d(yt_rsc_2_19_i_q_d),
      .yt_rsc_2_20_i_q_d(yt_rsc_2_20_i_q_d),
      .yt_rsc_2_21_i_q_d(yt_rsc_2_21_i_q_d),
      .yt_rsc_2_22_i_q_d(yt_rsc_2_22_i_q_d),
      .yt_rsc_2_23_i_q_d(yt_rsc_2_23_i_q_d),
      .yt_rsc_2_24_i_q_d(yt_rsc_2_24_i_q_d),
      .yt_rsc_2_25_i_q_d(yt_rsc_2_25_i_q_d),
      .yt_rsc_2_26_i_q_d(yt_rsc_2_26_i_q_d),
      .yt_rsc_2_27_i_q_d(yt_rsc_2_27_i_q_d),
      .yt_rsc_2_28_i_q_d(yt_rsc_2_28_i_q_d),
      .yt_rsc_2_29_i_q_d(yt_rsc_2_29_i_q_d),
      .yt_rsc_2_30_i_q_d(yt_rsc_2_30_i_q_d),
      .yt_rsc_2_31_i_q_d(yt_rsc_2_31_i_q_d),
      .yt_rsc_3_0_i_clkr_en_d(yt_rsc_3_0_i_clkr_en_d),
      .yt_rsc_3_0_i_q_d(yt_rsc_3_0_i_q_d),
      .yt_rsc_3_1_i_q_d(yt_rsc_3_1_i_q_d),
      .yt_rsc_3_2_i_q_d(yt_rsc_3_2_i_q_d),
      .yt_rsc_3_3_i_q_d(yt_rsc_3_3_i_q_d),
      .yt_rsc_3_4_i_q_d(yt_rsc_3_4_i_q_d),
      .yt_rsc_3_5_i_q_d(yt_rsc_3_5_i_q_d),
      .yt_rsc_3_6_i_q_d(yt_rsc_3_6_i_q_d),
      .yt_rsc_3_7_i_q_d(yt_rsc_3_7_i_q_d),
      .yt_rsc_3_8_i_q_d(yt_rsc_3_8_i_q_d),
      .yt_rsc_3_9_i_q_d(yt_rsc_3_9_i_q_d),
      .yt_rsc_3_10_i_q_d(yt_rsc_3_10_i_q_d),
      .yt_rsc_3_11_i_q_d(yt_rsc_3_11_i_q_d),
      .yt_rsc_3_12_i_q_d(yt_rsc_3_12_i_q_d),
      .yt_rsc_3_13_i_q_d(yt_rsc_3_13_i_q_d),
      .yt_rsc_3_14_i_q_d(yt_rsc_3_14_i_q_d),
      .yt_rsc_3_15_i_q_d(yt_rsc_3_15_i_q_d),
      .yt_rsc_3_16_i_clkr_en_d(yt_rsc_3_16_i_clkr_en_d),
      .yt_rsc_3_16_i_q_d(yt_rsc_3_16_i_q_d),
      .yt_rsc_3_17_i_q_d(yt_rsc_3_17_i_q_d),
      .yt_rsc_3_18_i_q_d(yt_rsc_3_18_i_q_d),
      .yt_rsc_3_19_i_q_d(yt_rsc_3_19_i_q_d),
      .yt_rsc_3_20_i_q_d(yt_rsc_3_20_i_q_d),
      .yt_rsc_3_21_i_q_d(yt_rsc_3_21_i_q_d),
      .yt_rsc_3_22_i_q_d(yt_rsc_3_22_i_q_d),
      .yt_rsc_3_23_i_q_d(yt_rsc_3_23_i_q_d),
      .yt_rsc_3_24_i_q_d(yt_rsc_3_24_i_q_d),
      .yt_rsc_3_25_i_q_d(yt_rsc_3_25_i_q_d),
      .yt_rsc_3_26_i_q_d(yt_rsc_3_26_i_q_d),
      .yt_rsc_3_27_i_q_d(yt_rsc_3_27_i_q_d),
      .yt_rsc_3_28_i_q_d(yt_rsc_3_28_i_q_d),
      .yt_rsc_3_29_i_q_d(yt_rsc_3_29_i_q_d),
      .yt_rsc_3_30_i_q_d(yt_rsc_3_30_i_q_d),
      .yt_rsc_3_31_i_q_d(yt_rsc_3_31_i_q_d),
      .yt_rsc_4_0_i_clkr_en_d(yt_rsc_4_0_i_clkr_en_d),
      .yt_rsc_4_0_i_q_d(yt_rsc_4_0_i_q_d),
      .yt_rsc_4_1_i_q_d(yt_rsc_4_1_i_q_d),
      .yt_rsc_4_2_i_q_d(yt_rsc_4_2_i_q_d),
      .yt_rsc_4_3_i_q_d(yt_rsc_4_3_i_q_d),
      .yt_rsc_4_4_i_q_d(yt_rsc_4_4_i_q_d),
      .yt_rsc_4_5_i_q_d(yt_rsc_4_5_i_q_d),
      .yt_rsc_4_6_i_q_d(yt_rsc_4_6_i_q_d),
      .yt_rsc_4_7_i_q_d(yt_rsc_4_7_i_q_d),
      .yt_rsc_4_8_i_q_d(yt_rsc_4_8_i_q_d),
      .yt_rsc_4_9_i_q_d(yt_rsc_4_9_i_q_d),
      .yt_rsc_4_10_i_q_d(yt_rsc_4_10_i_q_d),
      .yt_rsc_4_11_i_q_d(yt_rsc_4_11_i_q_d),
      .yt_rsc_4_12_i_q_d(yt_rsc_4_12_i_q_d),
      .yt_rsc_4_13_i_q_d(yt_rsc_4_13_i_q_d),
      .yt_rsc_4_14_i_q_d(yt_rsc_4_14_i_q_d),
      .yt_rsc_4_15_i_q_d(yt_rsc_4_15_i_q_d),
      .yt_rsc_4_16_i_clkr_en_d(yt_rsc_4_16_i_clkr_en_d),
      .yt_rsc_4_16_i_q_d(yt_rsc_4_16_i_q_d),
      .yt_rsc_4_17_i_q_d(yt_rsc_4_17_i_q_d),
      .yt_rsc_4_18_i_q_d(yt_rsc_4_18_i_q_d),
      .yt_rsc_4_19_i_q_d(yt_rsc_4_19_i_q_d),
      .yt_rsc_4_20_i_q_d(yt_rsc_4_20_i_q_d),
      .yt_rsc_4_21_i_q_d(yt_rsc_4_21_i_q_d),
      .yt_rsc_4_22_i_q_d(yt_rsc_4_22_i_q_d),
      .yt_rsc_4_23_i_q_d(yt_rsc_4_23_i_q_d),
      .yt_rsc_4_24_i_q_d(yt_rsc_4_24_i_q_d),
      .yt_rsc_4_25_i_q_d(yt_rsc_4_25_i_q_d),
      .yt_rsc_4_26_i_q_d(yt_rsc_4_26_i_q_d),
      .yt_rsc_4_27_i_q_d(yt_rsc_4_27_i_q_d),
      .yt_rsc_4_28_i_q_d(yt_rsc_4_28_i_q_d),
      .yt_rsc_4_29_i_q_d(yt_rsc_4_29_i_q_d),
      .yt_rsc_4_30_i_q_d(yt_rsc_4_30_i_q_d),
      .yt_rsc_4_31_i_q_d(yt_rsc_4_31_i_q_d),
      .yt_rsc_5_0_i_clkr_en_d(yt_rsc_5_0_i_clkr_en_d),
      .yt_rsc_5_0_i_q_d(yt_rsc_5_0_i_q_d),
      .yt_rsc_5_1_i_q_d(yt_rsc_5_1_i_q_d),
      .yt_rsc_5_2_i_q_d(yt_rsc_5_2_i_q_d),
      .yt_rsc_5_3_i_q_d(yt_rsc_5_3_i_q_d),
      .yt_rsc_5_4_i_q_d(yt_rsc_5_4_i_q_d),
      .yt_rsc_5_5_i_q_d(yt_rsc_5_5_i_q_d),
      .yt_rsc_5_6_i_q_d(yt_rsc_5_6_i_q_d),
      .yt_rsc_5_7_i_q_d(yt_rsc_5_7_i_q_d),
      .yt_rsc_5_8_i_q_d(yt_rsc_5_8_i_q_d),
      .yt_rsc_5_9_i_q_d(yt_rsc_5_9_i_q_d),
      .yt_rsc_5_10_i_q_d(yt_rsc_5_10_i_q_d),
      .yt_rsc_5_11_i_q_d(yt_rsc_5_11_i_q_d),
      .yt_rsc_5_12_i_q_d(yt_rsc_5_12_i_q_d),
      .yt_rsc_5_13_i_q_d(yt_rsc_5_13_i_q_d),
      .yt_rsc_5_14_i_q_d(yt_rsc_5_14_i_q_d),
      .yt_rsc_5_15_i_q_d(yt_rsc_5_15_i_q_d),
      .yt_rsc_5_16_i_clkr_en_d(yt_rsc_5_16_i_clkr_en_d),
      .yt_rsc_5_16_i_q_d(yt_rsc_5_16_i_q_d),
      .yt_rsc_5_17_i_q_d(yt_rsc_5_17_i_q_d),
      .yt_rsc_5_18_i_q_d(yt_rsc_5_18_i_q_d),
      .yt_rsc_5_19_i_q_d(yt_rsc_5_19_i_q_d),
      .yt_rsc_5_20_i_q_d(yt_rsc_5_20_i_q_d),
      .yt_rsc_5_21_i_q_d(yt_rsc_5_21_i_q_d),
      .yt_rsc_5_22_i_q_d(yt_rsc_5_22_i_q_d),
      .yt_rsc_5_23_i_q_d(yt_rsc_5_23_i_q_d),
      .yt_rsc_5_24_i_q_d(yt_rsc_5_24_i_q_d),
      .yt_rsc_5_25_i_q_d(yt_rsc_5_25_i_q_d),
      .yt_rsc_5_26_i_q_d(yt_rsc_5_26_i_q_d),
      .yt_rsc_5_27_i_q_d(yt_rsc_5_27_i_q_d),
      .yt_rsc_5_28_i_q_d(yt_rsc_5_28_i_q_d),
      .yt_rsc_5_29_i_q_d(yt_rsc_5_29_i_q_d),
      .yt_rsc_5_30_i_q_d(yt_rsc_5_30_i_q_d),
      .yt_rsc_5_31_i_q_d(yt_rsc_5_31_i_q_d),
      .yt_rsc_6_0_i_clkr_en_d(yt_rsc_6_0_i_clkr_en_d),
      .yt_rsc_6_0_i_q_d(yt_rsc_6_0_i_q_d),
      .yt_rsc_6_1_i_q_d(yt_rsc_6_1_i_q_d),
      .yt_rsc_6_2_i_q_d(yt_rsc_6_2_i_q_d),
      .yt_rsc_6_3_i_q_d(yt_rsc_6_3_i_q_d),
      .yt_rsc_6_4_i_q_d(yt_rsc_6_4_i_q_d),
      .yt_rsc_6_5_i_q_d(yt_rsc_6_5_i_q_d),
      .yt_rsc_6_6_i_q_d(yt_rsc_6_6_i_q_d),
      .yt_rsc_6_7_i_q_d(yt_rsc_6_7_i_q_d),
      .yt_rsc_6_8_i_q_d(yt_rsc_6_8_i_q_d),
      .yt_rsc_6_9_i_q_d(yt_rsc_6_9_i_q_d),
      .yt_rsc_6_10_i_q_d(yt_rsc_6_10_i_q_d),
      .yt_rsc_6_11_i_q_d(yt_rsc_6_11_i_q_d),
      .yt_rsc_6_12_i_q_d(yt_rsc_6_12_i_q_d),
      .yt_rsc_6_13_i_q_d(yt_rsc_6_13_i_q_d),
      .yt_rsc_6_14_i_q_d(yt_rsc_6_14_i_q_d),
      .yt_rsc_6_15_i_q_d(yt_rsc_6_15_i_q_d),
      .yt_rsc_6_16_i_clkr_en_d(yt_rsc_6_16_i_clkr_en_d),
      .yt_rsc_6_16_i_q_d(yt_rsc_6_16_i_q_d),
      .yt_rsc_6_17_i_q_d(yt_rsc_6_17_i_q_d),
      .yt_rsc_6_18_i_q_d(yt_rsc_6_18_i_q_d),
      .yt_rsc_6_19_i_q_d(yt_rsc_6_19_i_q_d),
      .yt_rsc_6_20_i_q_d(yt_rsc_6_20_i_q_d),
      .yt_rsc_6_21_i_q_d(yt_rsc_6_21_i_q_d),
      .yt_rsc_6_22_i_q_d(yt_rsc_6_22_i_q_d),
      .yt_rsc_6_23_i_q_d(yt_rsc_6_23_i_q_d),
      .yt_rsc_6_24_i_q_d(yt_rsc_6_24_i_q_d),
      .yt_rsc_6_25_i_q_d(yt_rsc_6_25_i_q_d),
      .yt_rsc_6_26_i_q_d(yt_rsc_6_26_i_q_d),
      .yt_rsc_6_27_i_q_d(yt_rsc_6_27_i_q_d),
      .yt_rsc_6_28_i_q_d(yt_rsc_6_28_i_q_d),
      .yt_rsc_6_29_i_q_d(yt_rsc_6_29_i_q_d),
      .yt_rsc_6_30_i_q_d(yt_rsc_6_30_i_q_d),
      .yt_rsc_6_31_i_q_d(yt_rsc_6_31_i_q_d),
      .yt_rsc_7_0_i_clkr_en_d(yt_rsc_7_0_i_clkr_en_d),
      .yt_rsc_7_0_i_q_d(yt_rsc_7_0_i_q_d),
      .yt_rsc_7_1_i_q_d(yt_rsc_7_1_i_q_d),
      .yt_rsc_7_2_i_q_d(yt_rsc_7_2_i_q_d),
      .yt_rsc_7_3_i_q_d(yt_rsc_7_3_i_q_d),
      .yt_rsc_7_4_i_q_d(yt_rsc_7_4_i_q_d),
      .yt_rsc_7_5_i_q_d(yt_rsc_7_5_i_q_d),
      .yt_rsc_7_6_i_q_d(yt_rsc_7_6_i_q_d),
      .yt_rsc_7_7_i_q_d(yt_rsc_7_7_i_q_d),
      .yt_rsc_7_8_i_q_d(yt_rsc_7_8_i_q_d),
      .yt_rsc_7_9_i_q_d(yt_rsc_7_9_i_q_d),
      .yt_rsc_7_10_i_q_d(yt_rsc_7_10_i_q_d),
      .yt_rsc_7_11_i_q_d(yt_rsc_7_11_i_q_d),
      .yt_rsc_7_12_i_q_d(yt_rsc_7_12_i_q_d),
      .yt_rsc_7_13_i_q_d(yt_rsc_7_13_i_q_d),
      .yt_rsc_7_14_i_q_d(yt_rsc_7_14_i_q_d),
      .yt_rsc_7_15_i_q_d(yt_rsc_7_15_i_q_d),
      .yt_rsc_7_16_i_clkr_en_d(yt_rsc_7_16_i_clkr_en_d),
      .yt_rsc_7_16_i_q_d(yt_rsc_7_16_i_q_d),
      .yt_rsc_7_17_i_q_d(yt_rsc_7_17_i_q_d),
      .yt_rsc_7_18_i_q_d(yt_rsc_7_18_i_q_d),
      .yt_rsc_7_19_i_q_d(yt_rsc_7_19_i_q_d),
      .yt_rsc_7_20_i_q_d(yt_rsc_7_20_i_q_d),
      .yt_rsc_7_21_i_q_d(yt_rsc_7_21_i_q_d),
      .yt_rsc_7_22_i_q_d(yt_rsc_7_22_i_q_d),
      .yt_rsc_7_23_i_q_d(yt_rsc_7_23_i_q_d),
      .yt_rsc_7_24_i_q_d(yt_rsc_7_24_i_q_d),
      .yt_rsc_7_25_i_q_d(yt_rsc_7_25_i_q_d),
      .yt_rsc_7_26_i_q_d(yt_rsc_7_26_i_q_d),
      .yt_rsc_7_27_i_q_d(yt_rsc_7_27_i_q_d),
      .yt_rsc_7_28_i_q_d(yt_rsc_7_28_i_q_d),
      .yt_rsc_7_29_i_q_d(yt_rsc_7_29_i_q_d),
      .yt_rsc_7_30_i_q_d(yt_rsc_7_30_i_q_d),
      .yt_rsc_7_31_i_q_d(yt_rsc_7_31_i_q_d),
      .xt_rsc_0_0_i_qa_d(xt_rsc_0_0_i_qa_d),
      .xt_rsc_0_1_i_qa_d(xt_rsc_0_1_i_qa_d),
      .xt_rsc_0_2_i_qa_d(xt_rsc_0_2_i_qa_d),
      .xt_rsc_0_3_i_qa_d(xt_rsc_0_3_i_qa_d),
      .xt_rsc_0_4_i_qa_d(xt_rsc_0_4_i_qa_d),
      .xt_rsc_0_5_i_qa_d(xt_rsc_0_5_i_qa_d),
      .xt_rsc_0_6_i_qa_d(xt_rsc_0_6_i_qa_d),
      .xt_rsc_0_7_i_qa_d(xt_rsc_0_7_i_qa_d),
      .xt_rsc_0_8_i_qa_d(xt_rsc_0_8_i_qa_d),
      .xt_rsc_0_9_i_qa_d(xt_rsc_0_9_i_qa_d),
      .xt_rsc_0_10_i_qa_d(xt_rsc_0_10_i_qa_d),
      .xt_rsc_0_11_i_qa_d(xt_rsc_0_11_i_qa_d),
      .xt_rsc_0_12_i_qa_d(xt_rsc_0_12_i_qa_d),
      .xt_rsc_0_13_i_qa_d(xt_rsc_0_13_i_qa_d),
      .xt_rsc_0_14_i_qa_d(xt_rsc_0_14_i_qa_d),
      .xt_rsc_0_15_i_qa_d(xt_rsc_0_15_i_qa_d),
      .xt_rsc_0_16_i_qa_d(xt_rsc_0_16_i_qa_d),
      .xt_rsc_0_17_i_qa_d(xt_rsc_0_17_i_qa_d),
      .xt_rsc_0_18_i_qa_d(xt_rsc_0_18_i_qa_d),
      .xt_rsc_0_19_i_qa_d(xt_rsc_0_19_i_qa_d),
      .xt_rsc_0_20_i_qa_d(xt_rsc_0_20_i_qa_d),
      .xt_rsc_0_21_i_qa_d(xt_rsc_0_21_i_qa_d),
      .xt_rsc_0_22_i_qa_d(xt_rsc_0_22_i_qa_d),
      .xt_rsc_0_23_i_qa_d(xt_rsc_0_23_i_qa_d),
      .xt_rsc_0_24_i_qa_d(xt_rsc_0_24_i_qa_d),
      .xt_rsc_0_25_i_qa_d(xt_rsc_0_25_i_qa_d),
      .xt_rsc_0_26_i_qa_d(xt_rsc_0_26_i_qa_d),
      .xt_rsc_0_27_i_qa_d(xt_rsc_0_27_i_qa_d),
      .xt_rsc_0_28_i_qa_d(xt_rsc_0_28_i_qa_d),
      .xt_rsc_0_29_i_qa_d(xt_rsc_0_29_i_qa_d),
      .xt_rsc_0_30_i_qa_d(xt_rsc_0_30_i_qa_d),
      .xt_rsc_0_31_i_qa_d(xt_rsc_0_31_i_qa_d),
      .xt_rsc_1_0_i_qa_d(xt_rsc_1_0_i_qa_d),
      .xt_rsc_1_1_i_qa_d(xt_rsc_1_1_i_qa_d),
      .xt_rsc_1_2_i_qa_d(xt_rsc_1_2_i_qa_d),
      .xt_rsc_1_3_i_qa_d(xt_rsc_1_3_i_qa_d),
      .xt_rsc_1_4_i_qa_d(xt_rsc_1_4_i_qa_d),
      .xt_rsc_1_5_i_qa_d(xt_rsc_1_5_i_qa_d),
      .xt_rsc_1_6_i_qa_d(xt_rsc_1_6_i_qa_d),
      .xt_rsc_1_7_i_qa_d(xt_rsc_1_7_i_qa_d),
      .xt_rsc_1_8_i_qa_d(xt_rsc_1_8_i_qa_d),
      .xt_rsc_1_9_i_qa_d(xt_rsc_1_9_i_qa_d),
      .xt_rsc_1_10_i_qa_d(xt_rsc_1_10_i_qa_d),
      .xt_rsc_1_11_i_qa_d(xt_rsc_1_11_i_qa_d),
      .xt_rsc_1_12_i_qa_d(xt_rsc_1_12_i_qa_d),
      .xt_rsc_1_13_i_qa_d(xt_rsc_1_13_i_qa_d),
      .xt_rsc_1_14_i_qa_d(xt_rsc_1_14_i_qa_d),
      .xt_rsc_1_15_i_qa_d(xt_rsc_1_15_i_qa_d),
      .xt_rsc_1_16_i_qa_d(xt_rsc_1_16_i_qa_d),
      .xt_rsc_1_17_i_qa_d(xt_rsc_1_17_i_qa_d),
      .xt_rsc_1_18_i_qa_d(xt_rsc_1_18_i_qa_d),
      .xt_rsc_1_19_i_qa_d(xt_rsc_1_19_i_qa_d),
      .xt_rsc_1_20_i_qa_d(xt_rsc_1_20_i_qa_d),
      .xt_rsc_1_21_i_qa_d(xt_rsc_1_21_i_qa_d),
      .xt_rsc_1_22_i_qa_d(xt_rsc_1_22_i_qa_d),
      .xt_rsc_1_23_i_qa_d(xt_rsc_1_23_i_qa_d),
      .xt_rsc_1_24_i_qa_d(xt_rsc_1_24_i_qa_d),
      .xt_rsc_1_25_i_qa_d(xt_rsc_1_25_i_qa_d),
      .xt_rsc_1_26_i_qa_d(xt_rsc_1_26_i_qa_d),
      .xt_rsc_1_27_i_qa_d(xt_rsc_1_27_i_qa_d),
      .xt_rsc_1_28_i_qa_d(xt_rsc_1_28_i_qa_d),
      .xt_rsc_1_29_i_qa_d(xt_rsc_1_29_i_qa_d),
      .xt_rsc_1_30_i_qa_d(xt_rsc_1_30_i_qa_d),
      .xt_rsc_1_31_i_qa_d(xt_rsc_1_31_i_qa_d),
      .xt_rsc_2_0_i_qa_d(xt_rsc_2_0_i_qa_d),
      .xt_rsc_2_1_i_qa_d(xt_rsc_2_1_i_qa_d),
      .xt_rsc_2_2_i_qa_d(xt_rsc_2_2_i_qa_d),
      .xt_rsc_2_3_i_qa_d(xt_rsc_2_3_i_qa_d),
      .xt_rsc_2_4_i_qa_d(xt_rsc_2_4_i_qa_d),
      .xt_rsc_2_5_i_qa_d(xt_rsc_2_5_i_qa_d),
      .xt_rsc_2_6_i_qa_d(xt_rsc_2_6_i_qa_d),
      .xt_rsc_2_7_i_qa_d(xt_rsc_2_7_i_qa_d),
      .xt_rsc_2_8_i_qa_d(xt_rsc_2_8_i_qa_d),
      .xt_rsc_2_9_i_qa_d(xt_rsc_2_9_i_qa_d),
      .xt_rsc_2_10_i_qa_d(xt_rsc_2_10_i_qa_d),
      .xt_rsc_2_11_i_qa_d(xt_rsc_2_11_i_qa_d),
      .xt_rsc_2_12_i_qa_d(xt_rsc_2_12_i_qa_d),
      .xt_rsc_2_13_i_qa_d(xt_rsc_2_13_i_qa_d),
      .xt_rsc_2_14_i_qa_d(xt_rsc_2_14_i_qa_d),
      .xt_rsc_2_15_i_qa_d(xt_rsc_2_15_i_qa_d),
      .xt_rsc_2_16_i_qa_d(xt_rsc_2_16_i_qa_d),
      .xt_rsc_2_17_i_qa_d(xt_rsc_2_17_i_qa_d),
      .xt_rsc_2_18_i_qa_d(xt_rsc_2_18_i_qa_d),
      .xt_rsc_2_19_i_qa_d(xt_rsc_2_19_i_qa_d),
      .xt_rsc_2_20_i_qa_d(xt_rsc_2_20_i_qa_d),
      .xt_rsc_2_21_i_qa_d(xt_rsc_2_21_i_qa_d),
      .xt_rsc_2_22_i_qa_d(xt_rsc_2_22_i_qa_d),
      .xt_rsc_2_23_i_qa_d(xt_rsc_2_23_i_qa_d),
      .xt_rsc_2_24_i_qa_d(xt_rsc_2_24_i_qa_d),
      .xt_rsc_2_25_i_qa_d(xt_rsc_2_25_i_qa_d),
      .xt_rsc_2_26_i_qa_d(xt_rsc_2_26_i_qa_d),
      .xt_rsc_2_27_i_qa_d(xt_rsc_2_27_i_qa_d),
      .xt_rsc_2_28_i_qa_d(xt_rsc_2_28_i_qa_d),
      .xt_rsc_2_29_i_qa_d(xt_rsc_2_29_i_qa_d),
      .xt_rsc_2_30_i_qa_d(xt_rsc_2_30_i_qa_d),
      .xt_rsc_2_31_i_qa_d(xt_rsc_2_31_i_qa_d),
      .xt_rsc_3_0_i_qa_d(xt_rsc_3_0_i_qa_d),
      .xt_rsc_3_1_i_qa_d(xt_rsc_3_1_i_qa_d),
      .xt_rsc_3_2_i_qa_d(xt_rsc_3_2_i_qa_d),
      .xt_rsc_3_3_i_qa_d(xt_rsc_3_3_i_qa_d),
      .xt_rsc_3_4_i_qa_d(xt_rsc_3_4_i_qa_d),
      .xt_rsc_3_5_i_qa_d(xt_rsc_3_5_i_qa_d),
      .xt_rsc_3_6_i_qa_d(xt_rsc_3_6_i_qa_d),
      .xt_rsc_3_7_i_qa_d(xt_rsc_3_7_i_qa_d),
      .xt_rsc_3_8_i_qa_d(xt_rsc_3_8_i_qa_d),
      .xt_rsc_3_9_i_qa_d(xt_rsc_3_9_i_qa_d),
      .xt_rsc_3_10_i_qa_d(xt_rsc_3_10_i_qa_d),
      .xt_rsc_3_11_i_qa_d(xt_rsc_3_11_i_qa_d),
      .xt_rsc_3_12_i_qa_d(xt_rsc_3_12_i_qa_d),
      .xt_rsc_3_13_i_qa_d(xt_rsc_3_13_i_qa_d),
      .xt_rsc_3_14_i_qa_d(xt_rsc_3_14_i_qa_d),
      .xt_rsc_3_15_i_qa_d(xt_rsc_3_15_i_qa_d),
      .xt_rsc_3_16_i_qa_d(xt_rsc_3_16_i_qa_d),
      .xt_rsc_3_17_i_qa_d(xt_rsc_3_17_i_qa_d),
      .xt_rsc_3_18_i_qa_d(xt_rsc_3_18_i_qa_d),
      .xt_rsc_3_19_i_qa_d(xt_rsc_3_19_i_qa_d),
      .xt_rsc_3_20_i_qa_d(xt_rsc_3_20_i_qa_d),
      .xt_rsc_3_21_i_qa_d(xt_rsc_3_21_i_qa_d),
      .xt_rsc_3_22_i_qa_d(xt_rsc_3_22_i_qa_d),
      .xt_rsc_3_23_i_qa_d(xt_rsc_3_23_i_qa_d),
      .xt_rsc_3_24_i_qa_d(xt_rsc_3_24_i_qa_d),
      .xt_rsc_3_25_i_qa_d(xt_rsc_3_25_i_qa_d),
      .xt_rsc_3_26_i_qa_d(xt_rsc_3_26_i_qa_d),
      .xt_rsc_3_27_i_qa_d(xt_rsc_3_27_i_qa_d),
      .xt_rsc_3_28_i_qa_d(xt_rsc_3_28_i_qa_d),
      .xt_rsc_3_29_i_qa_d(xt_rsc_3_29_i_qa_d),
      .xt_rsc_3_30_i_qa_d(xt_rsc_3_30_i_qa_d),
      .xt_rsc_3_31_i_qa_d(xt_rsc_3_31_i_qa_d),
      .xt_rsc_4_0_i_qa_d(xt_rsc_4_0_i_qa_d),
      .xt_rsc_4_1_i_qa_d(xt_rsc_4_1_i_qa_d),
      .xt_rsc_4_2_i_qa_d(xt_rsc_4_2_i_qa_d),
      .xt_rsc_4_3_i_qa_d(xt_rsc_4_3_i_qa_d),
      .xt_rsc_4_4_i_qa_d(xt_rsc_4_4_i_qa_d),
      .xt_rsc_4_5_i_qa_d(xt_rsc_4_5_i_qa_d),
      .xt_rsc_4_6_i_qa_d(xt_rsc_4_6_i_qa_d),
      .xt_rsc_4_7_i_qa_d(xt_rsc_4_7_i_qa_d),
      .xt_rsc_4_8_i_qa_d(xt_rsc_4_8_i_qa_d),
      .xt_rsc_4_9_i_qa_d(xt_rsc_4_9_i_qa_d),
      .xt_rsc_4_10_i_qa_d(xt_rsc_4_10_i_qa_d),
      .xt_rsc_4_11_i_qa_d(xt_rsc_4_11_i_qa_d),
      .xt_rsc_4_12_i_qa_d(xt_rsc_4_12_i_qa_d),
      .xt_rsc_4_13_i_qa_d(xt_rsc_4_13_i_qa_d),
      .xt_rsc_4_14_i_qa_d(xt_rsc_4_14_i_qa_d),
      .xt_rsc_4_15_i_qa_d(xt_rsc_4_15_i_qa_d),
      .xt_rsc_4_16_i_qa_d(xt_rsc_4_16_i_qa_d),
      .xt_rsc_4_17_i_qa_d(xt_rsc_4_17_i_qa_d),
      .xt_rsc_4_18_i_qa_d(xt_rsc_4_18_i_qa_d),
      .xt_rsc_4_19_i_qa_d(xt_rsc_4_19_i_qa_d),
      .xt_rsc_4_20_i_qa_d(xt_rsc_4_20_i_qa_d),
      .xt_rsc_4_21_i_qa_d(xt_rsc_4_21_i_qa_d),
      .xt_rsc_4_22_i_qa_d(xt_rsc_4_22_i_qa_d),
      .xt_rsc_4_23_i_qa_d(xt_rsc_4_23_i_qa_d),
      .xt_rsc_4_24_i_qa_d(xt_rsc_4_24_i_qa_d),
      .xt_rsc_4_25_i_qa_d(xt_rsc_4_25_i_qa_d),
      .xt_rsc_4_26_i_qa_d(xt_rsc_4_26_i_qa_d),
      .xt_rsc_4_27_i_qa_d(xt_rsc_4_27_i_qa_d),
      .xt_rsc_4_28_i_qa_d(xt_rsc_4_28_i_qa_d),
      .xt_rsc_4_29_i_qa_d(xt_rsc_4_29_i_qa_d),
      .xt_rsc_4_30_i_qa_d(xt_rsc_4_30_i_qa_d),
      .xt_rsc_4_31_i_qa_d(xt_rsc_4_31_i_qa_d),
      .xt_rsc_5_0_i_qa_d(xt_rsc_5_0_i_qa_d),
      .xt_rsc_5_1_i_qa_d(xt_rsc_5_1_i_qa_d),
      .xt_rsc_5_2_i_qa_d(xt_rsc_5_2_i_qa_d),
      .xt_rsc_5_3_i_qa_d(xt_rsc_5_3_i_qa_d),
      .xt_rsc_5_4_i_qa_d(xt_rsc_5_4_i_qa_d),
      .xt_rsc_5_5_i_qa_d(xt_rsc_5_5_i_qa_d),
      .xt_rsc_5_6_i_qa_d(xt_rsc_5_6_i_qa_d),
      .xt_rsc_5_7_i_qa_d(xt_rsc_5_7_i_qa_d),
      .xt_rsc_5_8_i_qa_d(xt_rsc_5_8_i_qa_d),
      .xt_rsc_5_9_i_qa_d(xt_rsc_5_9_i_qa_d),
      .xt_rsc_5_10_i_qa_d(xt_rsc_5_10_i_qa_d),
      .xt_rsc_5_11_i_qa_d(xt_rsc_5_11_i_qa_d),
      .xt_rsc_5_12_i_qa_d(xt_rsc_5_12_i_qa_d),
      .xt_rsc_5_13_i_qa_d(xt_rsc_5_13_i_qa_d),
      .xt_rsc_5_14_i_qa_d(xt_rsc_5_14_i_qa_d),
      .xt_rsc_5_15_i_qa_d(xt_rsc_5_15_i_qa_d),
      .xt_rsc_5_16_i_qa_d(xt_rsc_5_16_i_qa_d),
      .xt_rsc_5_17_i_qa_d(xt_rsc_5_17_i_qa_d),
      .xt_rsc_5_18_i_qa_d(xt_rsc_5_18_i_qa_d),
      .xt_rsc_5_19_i_qa_d(xt_rsc_5_19_i_qa_d),
      .xt_rsc_5_20_i_qa_d(xt_rsc_5_20_i_qa_d),
      .xt_rsc_5_21_i_qa_d(xt_rsc_5_21_i_qa_d),
      .xt_rsc_5_22_i_qa_d(xt_rsc_5_22_i_qa_d),
      .xt_rsc_5_23_i_qa_d(xt_rsc_5_23_i_qa_d),
      .xt_rsc_5_24_i_qa_d(xt_rsc_5_24_i_qa_d),
      .xt_rsc_5_25_i_qa_d(xt_rsc_5_25_i_qa_d),
      .xt_rsc_5_26_i_qa_d(xt_rsc_5_26_i_qa_d),
      .xt_rsc_5_27_i_qa_d(xt_rsc_5_27_i_qa_d),
      .xt_rsc_5_28_i_qa_d(xt_rsc_5_28_i_qa_d),
      .xt_rsc_5_29_i_qa_d(xt_rsc_5_29_i_qa_d),
      .xt_rsc_5_30_i_qa_d(xt_rsc_5_30_i_qa_d),
      .xt_rsc_5_31_i_qa_d(xt_rsc_5_31_i_qa_d),
      .xt_rsc_6_0_i_qa_d(xt_rsc_6_0_i_qa_d),
      .xt_rsc_6_1_i_qa_d(xt_rsc_6_1_i_qa_d),
      .xt_rsc_6_2_i_qa_d(xt_rsc_6_2_i_qa_d),
      .xt_rsc_6_3_i_qa_d(xt_rsc_6_3_i_qa_d),
      .xt_rsc_6_4_i_qa_d(xt_rsc_6_4_i_qa_d),
      .xt_rsc_6_5_i_qa_d(xt_rsc_6_5_i_qa_d),
      .xt_rsc_6_6_i_qa_d(xt_rsc_6_6_i_qa_d),
      .xt_rsc_6_7_i_qa_d(xt_rsc_6_7_i_qa_d),
      .xt_rsc_6_8_i_qa_d(xt_rsc_6_8_i_qa_d),
      .xt_rsc_6_9_i_qa_d(xt_rsc_6_9_i_qa_d),
      .xt_rsc_6_10_i_qa_d(xt_rsc_6_10_i_qa_d),
      .xt_rsc_6_11_i_qa_d(xt_rsc_6_11_i_qa_d),
      .xt_rsc_6_12_i_qa_d(xt_rsc_6_12_i_qa_d),
      .xt_rsc_6_13_i_qa_d(xt_rsc_6_13_i_qa_d),
      .xt_rsc_6_14_i_qa_d(xt_rsc_6_14_i_qa_d),
      .xt_rsc_6_15_i_qa_d(xt_rsc_6_15_i_qa_d),
      .xt_rsc_6_16_i_qa_d(xt_rsc_6_16_i_qa_d),
      .xt_rsc_6_17_i_qa_d(xt_rsc_6_17_i_qa_d),
      .xt_rsc_6_18_i_qa_d(xt_rsc_6_18_i_qa_d),
      .xt_rsc_6_19_i_qa_d(xt_rsc_6_19_i_qa_d),
      .xt_rsc_6_20_i_qa_d(xt_rsc_6_20_i_qa_d),
      .xt_rsc_6_21_i_qa_d(xt_rsc_6_21_i_qa_d),
      .xt_rsc_6_22_i_qa_d(xt_rsc_6_22_i_qa_d),
      .xt_rsc_6_23_i_qa_d(xt_rsc_6_23_i_qa_d),
      .xt_rsc_6_24_i_qa_d(xt_rsc_6_24_i_qa_d),
      .xt_rsc_6_25_i_qa_d(xt_rsc_6_25_i_qa_d),
      .xt_rsc_6_26_i_qa_d(xt_rsc_6_26_i_qa_d),
      .xt_rsc_6_27_i_qa_d(xt_rsc_6_27_i_qa_d),
      .xt_rsc_6_28_i_qa_d(xt_rsc_6_28_i_qa_d),
      .xt_rsc_6_29_i_qa_d(xt_rsc_6_29_i_qa_d),
      .xt_rsc_6_30_i_qa_d(xt_rsc_6_30_i_qa_d),
      .xt_rsc_6_31_i_qa_d(xt_rsc_6_31_i_qa_d),
      .xt_rsc_7_0_i_qa_d(xt_rsc_7_0_i_qa_d),
      .xt_rsc_7_1_i_qa_d(xt_rsc_7_1_i_qa_d),
      .xt_rsc_7_2_i_qa_d(xt_rsc_7_2_i_qa_d),
      .xt_rsc_7_3_i_qa_d(xt_rsc_7_3_i_qa_d),
      .xt_rsc_7_4_i_qa_d(xt_rsc_7_4_i_qa_d),
      .xt_rsc_7_5_i_qa_d(xt_rsc_7_5_i_qa_d),
      .xt_rsc_7_6_i_qa_d(xt_rsc_7_6_i_qa_d),
      .xt_rsc_7_7_i_qa_d(xt_rsc_7_7_i_qa_d),
      .xt_rsc_7_8_i_qa_d(xt_rsc_7_8_i_qa_d),
      .xt_rsc_7_9_i_qa_d(xt_rsc_7_9_i_qa_d),
      .xt_rsc_7_10_i_qa_d(xt_rsc_7_10_i_qa_d),
      .xt_rsc_7_11_i_qa_d(xt_rsc_7_11_i_qa_d),
      .xt_rsc_7_12_i_qa_d(xt_rsc_7_12_i_qa_d),
      .xt_rsc_7_13_i_qa_d(xt_rsc_7_13_i_qa_d),
      .xt_rsc_7_14_i_qa_d(xt_rsc_7_14_i_qa_d),
      .xt_rsc_7_15_i_qa_d(xt_rsc_7_15_i_qa_d),
      .xt_rsc_7_16_i_qa_d(xt_rsc_7_16_i_qa_d),
      .xt_rsc_7_17_i_qa_d(xt_rsc_7_17_i_qa_d),
      .xt_rsc_7_18_i_qa_d(xt_rsc_7_18_i_qa_d),
      .xt_rsc_7_19_i_qa_d(xt_rsc_7_19_i_qa_d),
      .xt_rsc_7_20_i_qa_d(xt_rsc_7_20_i_qa_d),
      .xt_rsc_7_21_i_qa_d(xt_rsc_7_21_i_qa_d),
      .xt_rsc_7_22_i_qa_d(xt_rsc_7_22_i_qa_d),
      .xt_rsc_7_23_i_qa_d(xt_rsc_7_23_i_qa_d),
      .xt_rsc_7_24_i_qa_d(xt_rsc_7_24_i_qa_d),
      .xt_rsc_7_25_i_qa_d(xt_rsc_7_25_i_qa_d),
      .xt_rsc_7_26_i_qa_d(xt_rsc_7_26_i_qa_d),
      .xt_rsc_7_27_i_qa_d(xt_rsc_7_27_i_qa_d),
      .xt_rsc_7_28_i_qa_d(xt_rsc_7_28_i_qa_d),
      .xt_rsc_7_29_i_qa_d(xt_rsc_7_29_i_qa_d),
      .xt_rsc_7_30_i_qa_d(xt_rsc_7_30_i_qa_d),
      .xt_rsc_7_31_i_qa_d(xt_rsc_7_31_i_qa_d),
      .twiddle_rsc_0_0_i_adra_d(twiddle_rsc_0_0_i_adra_d),
      .twiddle_rsc_0_0_i_qa_d(twiddle_rsc_0_0_i_qa_d),
      .twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_1_i_adra_d(twiddle_rsc_0_1_i_adra_d),
      .twiddle_rsc_0_1_i_qa_d(twiddle_rsc_0_1_i_qa_d),
      .twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_2_i_adra_d(twiddle_rsc_0_2_i_adra_d),
      .twiddle_rsc_0_2_i_qa_d(twiddle_rsc_0_2_i_qa_d),
      .twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_3_i_adra_d(twiddle_rsc_0_3_i_adra_d),
      .twiddle_rsc_0_3_i_qa_d(twiddle_rsc_0_3_i_qa_d),
      .twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_4_i_adra_d(twiddle_rsc_0_4_i_adra_d),
      .twiddle_rsc_0_4_i_qa_d(twiddle_rsc_0_4_i_qa_d),
      .twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_5_i_adra_d(twiddle_rsc_0_5_i_adra_d),
      .twiddle_rsc_0_5_i_qa_d(twiddle_rsc_0_5_i_qa_d),
      .twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_6_i_adra_d(twiddle_rsc_0_6_i_adra_d),
      .twiddle_rsc_0_6_i_qa_d(twiddle_rsc_0_6_i_qa_d),
      .twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_7_i_adra_d(twiddle_rsc_0_7_i_adra_d),
      .twiddle_rsc_0_7_i_qa_d(twiddle_rsc_0_7_i_qa_d),
      .twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_8_i_adra_d(twiddle_rsc_0_8_i_adra_d),
      .twiddle_rsc_0_8_i_qa_d(twiddle_rsc_0_8_i_qa_d),
      .twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_9_i_adra_d(twiddle_rsc_0_9_i_adra_d),
      .twiddle_rsc_0_9_i_qa_d(twiddle_rsc_0_9_i_qa_d),
      .twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_10_i_adra_d(twiddle_rsc_0_10_i_adra_d),
      .twiddle_rsc_0_10_i_qa_d(twiddle_rsc_0_10_i_qa_d),
      .twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_11_i_adra_d(twiddle_rsc_0_11_i_adra_d),
      .twiddle_rsc_0_11_i_qa_d(twiddle_rsc_0_11_i_qa_d),
      .twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_12_i_adra_d(twiddle_rsc_0_12_i_adra_d),
      .twiddle_rsc_0_12_i_qa_d(twiddle_rsc_0_12_i_qa_d),
      .twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_13_i_adra_d(twiddle_rsc_0_13_i_adra_d),
      .twiddle_rsc_0_13_i_qa_d(twiddle_rsc_0_13_i_qa_d),
      .twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_14_i_adra_d(twiddle_rsc_0_14_i_adra_d),
      .twiddle_rsc_0_14_i_qa_d(twiddle_rsc_0_14_i_qa_d),
      .twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_15_i_adra_d(twiddle_rsc_0_15_i_adra_d),
      .twiddle_rsc_0_15_i_qa_d(twiddle_rsc_0_15_i_qa_d),
      .twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_0_i_adra_d(twiddle_h_rsc_0_0_i_adra_d),
      .twiddle_h_rsc_0_0_i_qa_d(twiddle_h_rsc_0_0_i_qa_d),
      .twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_1_i_adra_d(twiddle_h_rsc_0_1_i_adra_d),
      .twiddle_h_rsc_0_1_i_qa_d(twiddle_h_rsc_0_1_i_qa_d),
      .twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_2_i_adra_d(twiddle_h_rsc_0_2_i_adra_d),
      .twiddle_h_rsc_0_2_i_qa_d(twiddle_h_rsc_0_2_i_qa_d),
      .twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_3_i_adra_d(twiddle_h_rsc_0_3_i_adra_d),
      .twiddle_h_rsc_0_3_i_qa_d(twiddle_h_rsc_0_3_i_qa_d),
      .twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_4_i_adra_d(twiddle_h_rsc_0_4_i_adra_d),
      .twiddle_h_rsc_0_4_i_qa_d(twiddle_h_rsc_0_4_i_qa_d),
      .twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_5_i_adra_d(twiddle_h_rsc_0_5_i_adra_d),
      .twiddle_h_rsc_0_5_i_qa_d(twiddle_h_rsc_0_5_i_qa_d),
      .twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_6_i_adra_d(twiddle_h_rsc_0_6_i_adra_d),
      .twiddle_h_rsc_0_6_i_qa_d(twiddle_h_rsc_0_6_i_qa_d),
      .twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_7_i_adra_d(twiddle_h_rsc_0_7_i_adra_d),
      .twiddle_h_rsc_0_7_i_qa_d(twiddle_h_rsc_0_7_i_qa_d),
      .twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_8_i_adra_d(twiddle_h_rsc_0_8_i_adra_d),
      .twiddle_h_rsc_0_8_i_qa_d(twiddle_h_rsc_0_8_i_qa_d),
      .twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_9_i_adra_d(twiddle_h_rsc_0_9_i_adra_d),
      .twiddle_h_rsc_0_9_i_qa_d(twiddle_h_rsc_0_9_i_qa_d),
      .twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_10_i_adra_d(twiddle_h_rsc_0_10_i_adra_d),
      .twiddle_h_rsc_0_10_i_qa_d(twiddle_h_rsc_0_10_i_qa_d),
      .twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_11_i_adra_d(twiddle_h_rsc_0_11_i_adra_d),
      .twiddle_h_rsc_0_11_i_qa_d(twiddle_h_rsc_0_11_i_qa_d),
      .twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_12_i_adra_d(twiddle_h_rsc_0_12_i_adra_d),
      .twiddle_h_rsc_0_12_i_qa_d(twiddle_h_rsc_0_12_i_qa_d),
      .twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_13_i_adra_d(twiddle_h_rsc_0_13_i_adra_d),
      .twiddle_h_rsc_0_13_i_qa_d(twiddle_h_rsc_0_13_i_qa_d),
      .twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_14_i_adra_d(twiddle_h_rsc_0_14_i_adra_d),
      .twiddle_h_rsc_0_14_i_qa_d(twiddle_h_rsc_0_14_i_qa_d),
      .twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_15_i_adra_d(twiddle_h_rsc_0_15_i_adra_d),
      .twiddle_h_rsc_0_15_i_qa_d(twiddle_h_rsc_0_15_i_qa_d),
      .twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_0_i_d_d_pff(yt_rsc_0_0_i_d_d_iff),
      .yt_rsc_0_0_i_radr_d_pff(yt_rsc_0_0_i_radr_d_iff),
      .yt_rsc_0_0_i_wadr_d_pff(yt_rsc_0_0_i_wadr_d_iff),
      .yt_rsc_0_0_i_we_d_pff(yt_rsc_0_0_i_we_d_iff),
      .yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_0_1_i_d_d_pff(yt_rsc_0_1_i_d_d_iff),
      .yt_rsc_0_1_i_wadr_d_pff(yt_rsc_0_1_i_wadr_d_iff),
      .yt_rsc_0_2_i_d_d_pff(yt_rsc_0_2_i_d_d_iff),
      .yt_rsc_0_2_i_wadr_d_pff(yt_rsc_0_2_i_wadr_d_iff),
      .yt_rsc_0_3_i_d_d_pff(yt_rsc_0_3_i_d_d_iff),
      .yt_rsc_0_3_i_wadr_d_pff(yt_rsc_0_3_i_wadr_d_iff),
      .yt_rsc_0_4_i_d_d_pff(yt_rsc_0_4_i_d_d_iff),
      .yt_rsc_0_4_i_wadr_d_pff(yt_rsc_0_4_i_wadr_d_iff),
      .yt_rsc_0_5_i_d_d_pff(yt_rsc_0_5_i_d_d_iff),
      .yt_rsc_0_5_i_wadr_d_pff(yt_rsc_0_5_i_wadr_d_iff),
      .yt_rsc_0_6_i_d_d_pff(yt_rsc_0_6_i_d_d_iff),
      .yt_rsc_0_6_i_wadr_d_pff(yt_rsc_0_6_i_wadr_d_iff),
      .yt_rsc_0_7_i_d_d_pff(yt_rsc_0_7_i_d_d_iff),
      .yt_rsc_0_8_i_d_d_pff(yt_rsc_0_8_i_d_d_iff),
      .yt_rsc_0_9_i_d_d_pff(yt_rsc_0_9_i_d_d_iff),
      .yt_rsc_0_10_i_d_d_pff(yt_rsc_0_10_i_d_d_iff),
      .yt_rsc_0_10_i_wadr_d_pff(yt_rsc_0_10_i_wadr_d_iff),
      .yt_rsc_0_11_i_d_d_pff(yt_rsc_0_11_i_d_d_iff),
      .yt_rsc_0_11_i_wadr_d_pff(yt_rsc_0_11_i_wadr_d_iff),
      .yt_rsc_0_12_i_d_d_pff(yt_rsc_0_12_i_d_d_iff),
      .yt_rsc_0_13_i_d_d_pff(yt_rsc_0_13_i_d_d_iff),
      .yt_rsc_0_14_i_d_d_pff(yt_rsc_0_14_i_d_d_iff),
      .yt_rsc_0_15_i_d_d_pff(yt_rsc_0_15_i_d_d_iff),
      .yt_rsc_0_16_i_we_d_pff(yt_rsc_0_16_i_we_d_iff),
      .yt_rsc_1_0_i_we_d_pff(yt_rsc_1_0_i_we_d_iff),
      .yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_1_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_1_16_i_we_d_pff(yt_rsc_1_16_i_we_d_iff),
      .yt_rsc_2_0_i_we_d_pff(yt_rsc_2_0_i_we_d_iff),
      .yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_2_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_2_16_i_we_d_pff(yt_rsc_2_16_i_we_d_iff),
      .yt_rsc_3_0_i_we_d_pff(yt_rsc_3_0_i_we_d_iff),
      .yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_3_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_3_16_i_we_d_pff(yt_rsc_3_16_i_we_d_iff),
      .yt_rsc_4_0_i_d_d_pff(yt_rsc_4_0_i_d_d_iff),
      .yt_rsc_4_0_i_wadr_d_pff(yt_rsc_4_0_i_wadr_d_iff),
      .yt_rsc_4_0_i_we_d_pff(yt_rsc_4_0_i_we_d_iff),
      .yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_4_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_4_1_i_d_d_pff(yt_rsc_4_1_i_d_d_iff),
      .yt_rsc_4_1_i_wadr_d_pff(yt_rsc_4_1_i_wadr_d_iff),
      .yt_rsc_4_2_i_d_d_pff(yt_rsc_4_2_i_d_d_iff),
      .yt_rsc_4_2_i_wadr_d_pff(yt_rsc_4_2_i_wadr_d_iff),
      .yt_rsc_4_3_i_d_d_pff(yt_rsc_4_3_i_d_d_iff),
      .yt_rsc_4_3_i_wadr_d_pff(yt_rsc_4_3_i_wadr_d_iff),
      .yt_rsc_4_4_i_d_d_pff(yt_rsc_4_4_i_d_d_iff),
      .yt_rsc_4_4_i_wadr_d_pff(yt_rsc_4_4_i_wadr_d_iff),
      .yt_rsc_4_5_i_d_d_pff(yt_rsc_4_5_i_d_d_iff),
      .yt_rsc_4_5_i_wadr_d_pff(yt_rsc_4_5_i_wadr_d_iff),
      .yt_rsc_4_6_i_d_d_pff(yt_rsc_4_6_i_d_d_iff),
      .yt_rsc_4_6_i_wadr_d_pff(yt_rsc_4_6_i_wadr_d_iff),
      .yt_rsc_4_7_i_d_d_pff(yt_rsc_4_7_i_d_d_iff),
      .yt_rsc_4_8_i_d_d_pff(yt_rsc_4_8_i_d_d_iff),
      .yt_rsc_4_9_i_d_d_pff(yt_rsc_4_9_i_d_d_iff),
      .yt_rsc_4_9_i_wadr_d_pff(yt_rsc_4_9_i_wadr_d_iff),
      .yt_rsc_4_10_i_d_d_pff(yt_rsc_4_10_i_d_d_iff),
      .yt_rsc_4_10_i_wadr_d_pff(yt_rsc_4_10_i_wadr_d_iff),
      .yt_rsc_4_11_i_d_d_pff(yt_rsc_4_11_i_d_d_iff),
      .yt_rsc_4_11_i_wadr_d_pff(yt_rsc_4_11_i_wadr_d_iff),
      .yt_rsc_4_12_i_d_d_pff(yt_rsc_4_12_i_d_d_iff),
      .yt_rsc_4_13_i_d_d_pff(yt_rsc_4_13_i_d_d_iff),
      .yt_rsc_4_14_i_d_d_pff(yt_rsc_4_14_i_d_d_iff),
      .yt_rsc_4_15_i_d_d_pff(yt_rsc_4_15_i_d_d_iff),
      .yt_rsc_4_16_i_we_d_pff(yt_rsc_4_16_i_we_d_iff),
      .yt_rsc_5_0_i_we_d_pff(yt_rsc_5_0_i_we_d_iff),
      .yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_5_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_5_16_i_we_d_pff(yt_rsc_5_16_i_we_d_iff),
      .yt_rsc_6_0_i_we_d_pff(yt_rsc_6_0_i_we_d_iff),
      .yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_6_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_6_16_i_we_d_pff(yt_rsc_6_16_i_we_d_iff),
      .yt_rsc_7_0_i_we_d_pff(yt_rsc_7_0_i_we_d_iff),
      .yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_pff(yt_rsc_7_0_i_readA_r_ram_ir_internal_RMASK_B_d_iff),
      .yt_rsc_7_16_i_we_d_pff(yt_rsc_7_16_i_we_d_iff),
      .xt_rsc_0_0_i_adra_d_pff(xt_rsc_0_0_i_adra_d_iff),
      .xt_rsc_0_0_i_da_d_pff(xt_rsc_0_0_i_da_d_iff),
      .xt_rsc_0_0_i_wea_d_pff(xt_rsc_0_0_i_wea_d_iff),
      .xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_0_1_i_adra_d_pff(xt_rsc_0_1_i_adra_d_iff),
      .xt_rsc_0_1_i_da_d_pff(xt_rsc_0_1_i_da_d_iff),
      .xt_rsc_0_2_i_adra_d_pff(xt_rsc_0_2_i_adra_d_iff),
      .xt_rsc_0_2_i_da_d_pff(xt_rsc_0_2_i_da_d_iff),
      .xt_rsc_0_3_i_adra_d_pff(xt_rsc_0_3_i_adra_d_iff),
      .xt_rsc_0_3_i_da_d_pff(xt_rsc_0_3_i_da_d_iff),
      .xt_rsc_0_4_i_adra_d_pff(xt_rsc_0_4_i_adra_d_iff),
      .xt_rsc_0_4_i_da_d_pff(xt_rsc_0_4_i_da_d_iff),
      .xt_rsc_0_5_i_adra_d_pff(xt_rsc_0_5_i_adra_d_iff),
      .xt_rsc_0_5_i_da_d_pff(xt_rsc_0_5_i_da_d_iff),
      .xt_rsc_0_6_i_adra_d_pff(xt_rsc_0_6_i_adra_d_iff),
      .xt_rsc_0_6_i_da_d_pff(xt_rsc_0_6_i_da_d_iff),
      .xt_rsc_0_7_i_adra_d_pff(xt_rsc_0_7_i_adra_d_iff),
      .xt_rsc_0_7_i_da_d_pff(xt_rsc_0_7_i_da_d_iff),
      .xt_rsc_0_8_i_adra_d_pff(xt_rsc_0_8_i_adra_d_iff),
      .xt_rsc_0_8_i_da_d_pff(xt_rsc_0_8_i_da_d_iff),
      .xt_rsc_0_9_i_adra_d_pff(xt_rsc_0_9_i_adra_d_iff),
      .xt_rsc_0_9_i_da_d_pff(xt_rsc_0_9_i_da_d_iff),
      .xt_rsc_0_10_i_adra_d_pff(xt_rsc_0_10_i_adra_d_iff),
      .xt_rsc_0_10_i_da_d_pff(xt_rsc_0_10_i_da_d_iff),
      .xt_rsc_0_11_i_adra_d_pff(xt_rsc_0_11_i_adra_d_iff),
      .xt_rsc_0_11_i_da_d_pff(xt_rsc_0_11_i_da_d_iff),
      .xt_rsc_0_12_i_adra_d_pff(xt_rsc_0_12_i_adra_d_iff),
      .xt_rsc_0_12_i_da_d_pff(xt_rsc_0_12_i_da_d_iff),
      .xt_rsc_0_13_i_adra_d_pff(xt_rsc_0_13_i_adra_d_iff),
      .xt_rsc_0_13_i_da_d_pff(xt_rsc_0_13_i_da_d_iff),
      .xt_rsc_0_14_i_adra_d_pff(xt_rsc_0_14_i_adra_d_iff),
      .xt_rsc_0_14_i_da_d_pff(xt_rsc_0_14_i_da_d_iff),
      .xt_rsc_0_15_i_adra_d_pff(xt_rsc_0_15_i_adra_d_iff),
      .xt_rsc_0_15_i_da_d_pff(xt_rsc_0_15_i_da_d_iff),
      .xt_rsc_0_16_i_wea_d_pff(xt_rsc_0_16_i_wea_d_iff),
      .xt_rsc_1_0_i_wea_d_pff(xt_rsc_1_0_i_wea_d_iff),
      .xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_1_16_i_wea_d_pff(xt_rsc_1_16_i_wea_d_iff),
      .xt_rsc_2_0_i_wea_d_pff(xt_rsc_2_0_i_wea_d_iff),
      .xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_2_16_i_wea_d_pff(xt_rsc_2_16_i_wea_d_iff),
      .xt_rsc_3_0_i_wea_d_pff(xt_rsc_3_0_i_wea_d_iff),
      .xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_3_16_i_wea_d_pff(xt_rsc_3_16_i_wea_d_iff),
      .xt_rsc_4_0_i_da_d_pff(xt_rsc_4_0_i_da_d_iff),
      .xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_4_1_i_adra_d_pff(xt_rsc_4_1_i_adra_d_iff),
      .xt_rsc_4_1_i_da_d_pff(xt_rsc_4_1_i_da_d_iff),
      .xt_rsc_4_2_i_adra_d_pff(xt_rsc_4_2_i_adra_d_iff),
      .xt_rsc_4_2_i_da_d_pff(xt_rsc_4_2_i_da_d_iff),
      .xt_rsc_4_3_i_da_d_pff(xt_rsc_4_3_i_da_d_iff),
      .xt_rsc_4_4_i_da_d_pff(xt_rsc_4_4_i_da_d_iff),
      .xt_rsc_4_5_i_da_d_pff(xt_rsc_4_5_i_da_d_iff),
      .xt_rsc_4_6_i_da_d_pff(xt_rsc_4_6_i_da_d_iff),
      .xt_rsc_4_7_i_da_d_pff(xt_rsc_4_7_i_da_d_iff),
      .xt_rsc_4_8_i_da_d_pff(xt_rsc_4_8_i_da_d_iff),
      .xt_rsc_4_9_i_adra_d_pff(xt_rsc_4_9_i_adra_d_iff),
      .xt_rsc_4_9_i_da_d_pff(xt_rsc_4_9_i_da_d_iff),
      .xt_rsc_4_10_i_adra_d_pff(xt_rsc_4_10_i_adra_d_iff),
      .xt_rsc_4_10_i_da_d_pff(xt_rsc_4_10_i_da_d_iff),
      .xt_rsc_4_11_i_da_d_pff(xt_rsc_4_11_i_da_d_iff),
      .xt_rsc_4_12_i_da_d_pff(xt_rsc_4_12_i_da_d_iff),
      .xt_rsc_4_13_i_da_d_pff(xt_rsc_4_13_i_da_d_iff),
      .xt_rsc_4_14_i_da_d_pff(xt_rsc_4_14_i_da_d_iff),
      .xt_rsc_4_15_i_da_d_pff(xt_rsc_4_15_i_da_d_iff),
      .xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff),
      .xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff(xt_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff)
    );
endmodule



