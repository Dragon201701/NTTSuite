
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_libs/interfaces/amba/amba_comps.vhd 
--//////////////////////////////////////////////////////////////////////////////
-- Catapult Synthesis - Custom Interfaces
--
-- Copyright (c) 2016 Mentor Graphics Corp.
--       All Rights Reserved
-- 
-- This document contains information that is proprietary to Mentor Graphics
-- Corp. The original recipient of this document may duplicate this  
-- document in whole or in part for internal business purposes only, provided  
-- that this entire notice appears in all copies. In duplicating any part of  
-- this document, the recipient agrees to make every reasonable effort to  
-- prevent the unauthorized use and distribution of the proprietary information.
-- 
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in prepartion for creating
-- their own custom interfaces. This design does not present a complete
-- implementation of the named protocol or standard.
--
-- NO WARRANTY.
-- MENTOR GRAPHICS CORP. EXPRESSLY DISCLAIMS ALL WARRANTY
-- FOR THE SOFTWARE. TO THE MAXIMUM EXTENT PERMITTED BY APPLICABLE
-- LAW, THE SOFTWARE AND ANY RELATED DOCUMENTATION IS PROVIDED "AS IS"
-- AND WITH ALL FAULTS AND WITHOUT WARRANTIES OR CONDITIONS OF ANY
-- KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, WITHOUT LIMITATION, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR
-- PURPOSE, OR NONINFRINGEMENT. THE ENTIRE RISK ARISING OUT OF USE OR
-- DISTRIBUTION OF THE SOFTWARE REMAINS WITH YOU.
-- 
--//////////////////////////////////////////////////////////////////////////////

-- --------------------------------------------------------------------------
-- LIBRARY: amba
--
-- CONTENTS:
--    axi4stream_w_wire, axi4stream_r_wire, axi4svideo_w_wire, axi4svideo_r_wire
--      Catapult AXI-4 Stream bus definitions
--    ccs_axi4stream_in
--      AXI4-Streaming input interface
--    ccs_axi4stream_out
--      AXI4-Streaming output interface
--    ccs_axi4stream_pipe
--      AXI4-Streaming FIFO interconnect component
--    ccs_axi4svideo_in
--      AXI4-Streaming video input interface
--    ccs_axi4svideo_out
--      AXI4-Streaming video output interface
--    ccs_axi4svideo_pipe
--      AXI4-Streaming video FIFO interconnect component
--
--    axi4_busdef
--      Catapult AXI-4 bus definition
--
--    ccs_axi4_slave_mem
--      Catapult AXI-4 slave memory
---
--    ccs_axi4_master
--      Catapult AXI4 master interface for read/write data
--
--    apb_busdef
--      Catapult APB bus definition
--    apb_slave_mem
--      APB Slave Memory interface
--
-- CHANGE LOG:
--
--  10/01/16 - dgb - Initial implementation
--
-- --------------------------------------------------------------------------

-- --------------------------------------------------------------------------
-- PACKAGE:     amba_comps
--
-- DESCRIPTION:
--   Contains component declarations for all design units in this file.
--
-- CHANGE LOG:
--
--  10/01/16 - dgb - Initial implementation
--
-- --------------------------------------------------------------------------

LIBRARY ieee;

   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_arith.all;
   USE ieee.std_logic_unsigned.all;

PACKAGE amba_comps IS

  -- ==============================================================
  -- AXI-4 Stream Components
  -- ------------------------------ TSTRB/TKEEP controls --------------------
  --    TKEEP   TSTRB   Data Type         Description
  --    high    high    Data byte         Valid data byte (supported in these models)
  --    high    low     Position byte     Byte is position not data/null (not supported)
  --    low     low     Null byte         Byte is null (not supported)
  --    low     high    Reserved          Do not use (not supported)

  COMPONENT axi4stream_w_wire -- slave interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 16;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : IN   std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : IN   std_logic_vector(AXI4_USER_WIDTH-1 downto 0)      -- M->S      Optional user-defined sideband data
    );
  END COMPONENT;

  COMPONENT axi4stream_r_wire -- master interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 16;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : OUT  std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : OUT  std_logic_vector(AXI4_USER_WIDTH-1 downto 0)      -- M->S      Optional user-defined sideband data
    );
  END COMPONENT;

  COMPONENT axi4svideo_w_wire -- slave interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1024 := 33;           -- Catapult read/write operator width
      AXI4_DATA_WIDTH  : INTEGER                 := 16            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TUSER     : IN   std_logic;                                        -- M->S      Start of Frame
      TLAST     : IN   std_logic                                         -- M->S      End of Line
    );
  END COMPONENT;

  COMPONENT axi4svideo_r_wire -- master interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1024 := 33;           -- Catapult read/write operator width
      AXI4_DATA_WIDTH  : INTEGER                 := 16            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TUSER     : OUT  std_logic;                                        -- M->S      Start of Frame
      TLAST     : OUT  std_logic                                         -- M->S      End of Line
    );
  END COMPONENT;

  COMPONENT ccs_axi4stream_in
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW synchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : IN   std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : IN   std_logic_vector(AXI4_USER_WIDTH-1 downto 0);     -- M->S      Optional user-defined sideband data
      -- Catapult interface (equiv to mgc_in_wire_wait)
      d         : OUT  std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER(...) TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TVALID
      ld        : IN   std_logic                                         -- ld - TREADY
    );
  END COMPONENT;

  COMPONENT ccs_axi4stream_out
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW synchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : OUT  std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : OUT  std_logic_vector(AXI4_USER_WIDTH-1 downto 0);     -- M->S      Optional user-defined sideband data
      -- Catapult interface (equiv to mgc_out_stdreg_wait)
      d         : IN   std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER(...) TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TREADY
      ld        : IN   std_logic                                         -- ld - TVALID
    );
  END COMPONENT;

  -- This implementation currently does not work - the 'width' parameter is not configured properly
  COMPONENT ccs_axi4stream_pipe
    GENERIC(
      rscid            : INTEGER := 1;                            -- Resource ID from Catapult
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      fifo_sz          : INTEGER RANGE 0 TO 128 := 0;            -- Fifo size
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                          -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                          -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface input                                      -- Src->Dst  Description
      sTVALID   : IN   std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      sTREADY   : OUT  std_logic;                                          -- S->M      Indicates slave can accept a transfer
      sTDATA    : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      sTSTRB    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      sTKEEP    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      sTLAST    : IN   std_logic;                                          -- M->S      Indicates boundary of a packet
      sTUSER    : IN   std_logic_vector(AXI4_USER_WIDTH-1 downto 0);       -- M->S      Optional user-defined sideband data
      -- AXI-4 Stream interface output                                     -- Src->Dst  Description
      mTVALID   : OUT  std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      mTREADY   : IN   std_logic;                                          -- S->M      Indicates slave can accept a transfer
      mTDATA    : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      mTSTRB    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      mTKEEP    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      mTLAST    : OUT  std_logic;                                          -- M->S      Indicates boundary of a packet
      mTUSER    : OUT  std_logic_vector(AXI4_USER_WIDTH-1 downto 0)        -- M->S      Optional user-defined sideband data
    );
  END COMPONENT;

  COMPONENT ccs_axi4svideo_in
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : IN   std_logic;                                        -- M->S      End-of-line
      TUSER     : IN   std_logic;                                        -- M->S      Start-of-frame
      -- Catapult interface (equiv to mgc_in_wire_wait)
      d         : OUT  std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TVALID
      ld        : IN   std_logic                                         -- ld - TREADY
    );
  END COMPONENT;

  COMPONENT ccs_axi4svideo_out
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : OUT  std_logic;                                        -- M->S      End-of-line
      TUSER     : OUT  std_logic;                                        -- M->S      Start-of-frame
      -- Catapult interface (equiv to mgc_out_stdreg_wait)
      d         : IN   std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TREADY
      ld        : IN   std_logic                                         -- ld - TVALID
    );
  END COMPONENT;

  COMPONENT ccs_axi4svideo_pipe
    GENERIC(
      rscid            : INTEGER := 1;                                 -- Resource ID from Catapult
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      fifo_sz          : INTEGER RANGE 0 TO 128 := 0;            -- Fifo size
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                          -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                          -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface input                                      -- Src->Dst  Description
      sTVALID   : IN   std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      sTREADY   : OUT  std_logic;                                          -- S->M      Indicates slave can accept a transfer
      sTDATA    : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      sTSTRB    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      sTKEEP    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      sTLAST    : IN   std_logic;                                          -- M->S      End-of-line
      sTUSER    : IN   std_logic;                                          -- M->S      Start-of-frame
      -- AXI-4 Stream interface output                                     -- Src->Dst  Description
      mTVALID   : OUT  std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      mTREADY   : IN   std_logic;                                          -- S->M      Indicates slave can accept a transfer
      mTDATA    : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      mTSTRB    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      mTKEEP    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      mTLAST    : OUT  std_logic;                                          -- M->S      End-of-line
      mTUSER    : OUT  std_logic                                           -- M->S      Start-of-frame
    );
  END COMPONENT;

  -- ==============================================================
  -- AXI-4 Bus Components

  -- Used to define the AXI-4 bus definition (direction of signals is from the slave's perspective)
    -- Pin directions are based on the usage of this busdef as a "master" driving an input slave.
    -- To use the bus in the reverse direction set the interface to "slave".
  COMPONENT axi4_busdef -- 
    GENERIC(   
      host_tidw      : INTEGER RANGE 1 TO 11 := 4;            -- Width of transaction ID fields
      host_userw     : INTEGER RANGE 1 TO 16 := 4;            -- Width of user-defined signals
      ADDR_WIDTH     : INTEGER RANGE 1 TO 64 := 32;           -- Host address width
      DATA_WIDTH     : INTEGER RANGE 8 TO 64 := 8             -- Host data width
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                 -- Rising edge clock
      ARESETn    : IN   std_logic;                                 -- Active LOW synchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(host_tidw-1 downto 0);    -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);      -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);              -- Write burst length    - must always be 0 in AXI4-Lite
      AWSIZE     : OUT  std_logic_vector(1 downto 0);              -- Write burst size      - must equal host_dw_bytes-2
      AWBURST    : OUT  std_logic_vector(1 downto 0);              -- Write burst mode      - must always be 0 (fixed mode) in AXI4-Lite
      AWLOCK     : OUT  std_logic;                                 -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      AWCACHE    : OUT  std_logic_vector(3 downto 0);              -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      AWPROT     : OUT  std_logic_vector(2 downto 0);              -- Protection Type       - ignored in this model
      AWQOS      : OUT  std_logic_vector(3 downto 0);              -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);              -- Region identifier
      AWUSER     : OUT  std_logic_vector(host_userw-1 downto 0);   -- User signal
      AWVALID    : OUT  std_logic;                                 -- Write address valid
      AWREADY    : IN   std_logic;                                 -- Write address ready (slave is ready to accept AWADDR)
      
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0); -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise) - ignored in AXI-4 Lite
      WLAST      : OUT  std_logic;                                        -- Write last
      WUSER      : OUT  std_logic_vector(host_userw-1 downto 0);          -- User signal
      WVALID     : OUT  std_logic;                                        -- Write data is valid
      WREADY     : IN   std_logic;                                        -- Write ready (slave is ready to accept WDATA)
      
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(host_tidw-1 downto 0);    -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);              -- Write response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      BUSER      : IN   std_logic_vector(host_userw-1 downto 0);   -- User signal
      BVALID     : IN   std_logic;                                 -- Write response valid (slave accepted WDATA)
      BREADY     : OUT  std_logic;                                 -- Response ready (master can accept slave's write response)
      
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(host_tidw-1 downto 0);    -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);      -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);              -- Read burst length     - must always be 0 in AXI4-Lite
      ARSIZE     : OUT  std_logic_vector(1 downto 0);              -- Read burst size       - must equal host_dw_bytes-2
      ARBURST    : OUT  std_logic_vector(1 downto 0);              -- Read burst mode       - must always be 0 (fixed mode) in AXI4-Lite
      ARLOCK     : OUT  std_logic;                                 -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      ARCACHE    : OUT  std_logic_vector(3 downto 0);              -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      ARPROT     : OUT  std_logic_vector(2 downto 0);              -- Protection Type       - ignored in this model
      ARQOS      : OUT  std_logic_vector(3 downto 0);              -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);              -- Region identifier
      ARUSER     : OUT  std_logic_vector(host_userw-1 downto 0);   -- User signal
      ARVALID    : OUT  std_logic;                                 -- Read address valid
      ARREADY    : IN   std_logic;                                 -- Read address ready (slave is ready to accept ARADDR)
      
      -- ============== AXI4 Read Data Channel Signals
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0); -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                      -- Read response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      RVALID     : IN   std_logic;                                         -- Read valid (slave providing RDATA)
      RREADY     : OUT  std_logic;                                         -- Read ready (master ready to receive RDATA)
      RID        : OUT  std_logic_vector(host_tidw-1 downto 0);            -- Read ID tag
      RLAST      : IN   std_logic;                                         -- Read last
      RUSER      : IN   std_logic_vector(host_userw-1 downto 0)            -- User signal
    );
  END COMPONENT;

  -- AXI4 Lite GPIO with CDC
  COMPONENT ccs_axi4_lite_slave_cdc
    GENERIC(
      rscid          : INTEGER               := 1;            -- Required resource ID parameter
      op_width       : INTEGER RANGE 1 TO 64 := 1;            -- Operator width (dummy parameter)
      cwidth         : INTEGER RANGE 1 TO 256 := 32;          -- Internal register width
      nopreload      : INTEGER RANGE 0 TO 1 := 0;             -- 1=disable required preload before Catapult can read
      ADDR_WIDTH     : INTEGER RANGE 12 TO 32 := 32;          -- AXI4-Lite host address width
      DATA_WIDTH     : INTEGER RANGE 32 TO 64 := 32           -- AXI4-Lite host data width (must be 32 or 64)
    );
    PORT(
      -- AXI-4 Lite Interface
      ACLK       : IN   std_logic;                                 -- AXI-4 Bus Clock - Rising edge
      ARESETn    : IN   std_logic;                                 -- Active LOW synchronous reset
      -- ============== AXI4-Lite Write Address Channel Signals
      AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);               -- Write address
      AWVALID    : IN   std_logic;                                          -- Write address valid
      AWREADY    : OUT  std_logic;                                          -- Write address ready (slave is ready to accept AWADDR)
      -- ============== AXI4-Lite Write Data Channel
      WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0); -- Write data
      WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise) - ignored in AXI-4 Lite
      WVALID     : IN   std_logic;                                          -- Write data is valid
      WREADY     : OUT  std_logic;                                          -- Write ready (slave is ready to accept WDATA)
      -- ============== AXI4-Lite Write Response Channel Signals
      BRESP      : OUT  std_logic_vector(1 downto 0);                       -- Write response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      BVALID     : OUT  std_logic;                                          -- Write response valid (slave accepted WDATA)
      BREADY     : IN   std_logic;                                          -- Response ready (master can accept slave's write response)
      -- ============== AXI4-Lite Read Address Channel Signals
      ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);               -- Read address
      ARVALID    : IN   std_logic;                                          -- Read address valid
      ARREADY    : OUT  std_logic;                                          -- Read address ready (slave is ready to accept ARADDR)
      -- ============== AXI4-Lite Read Data Channel Signals
      RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0); -- Read data
      RRESP      : OUT  std_logic_vector(1 downto 0);                       -- Read response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      RVALID     : OUT  std_logic;                                          -- Read valid (slave providing RDATA)
      RREADY     : IN   std_logic;                                          -- Read ready (master ready to receive RDATA)

      -- Catapult interface assuming sidebyside packing 
      clk        : IN   std_logic;                                     -- Catapult Clock
      arst_n     : IN   std_logic;                                     -- Reset
--    d_from_ccs : IN   std_logic_vector(cwidth-1 downto 0);           -- Data out of Catapult block
--    d_from_vld : IN   std_logic;                                     -- Data out is valid
      d_to_ccs   : OUT  std_logic_vector(cwidth-1 downto 0)            -- Data into Catapult bloc
    );
  END COMPONENT;

  
  -- AXI4 Lite Slave Output
  COMPONENT ccs_axi4_lite_slave_out
    GENERIC(
      rscid          : INTEGER               := 1;            -- Required resource ID parameter
      op_width       : INTEGER RANGE 1 TO 64 := 1;            -- Operator width (dummy parameter)
      cwidth         : INTEGER RANGE 1 TO 256 := 32;          -- Internal register width
      nopreload      : INTEGER RANGE 0 TO 1 := 0;             -- 1=disable required preload before Catapult can read
      ADDR_WIDTH     : INTEGER RANGE 12 TO 32 := 32;          -- AXI4-Lite host address width
      DATA_WIDTH     : INTEGER RANGE 32 TO 64 := 32           -- AXI4-Lite host data width (must be 32 or 64)
    );
    PORT(
      -- AXI-4 Lite Interface
      ACLK       : IN   std_logic;                                     -- AXI-4 Bus Clock - Rising edge
      ARESETn    : IN   std_logic;                                     -- Active LOW synchronous reset
      -- ============== AXI4-Lite Write Address Channel Signals
      AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
      AWVALID    : IN   std_logic;                                     -- Write address valid
      AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
      --AWLEN      : IN   std_logic_vector(7 downto 0);                -- Write burst length    - must always be 0 in AXI4-Lite
      --AWSIZE     : IN   std_logic_vector(1 downto 0);                -- Write burst size      - must equal host_dw_bytes-2
      --AWBURST    : IN   std_logic_vector(1 downto 0);                -- Write burst mode      - must always be 0 (fixed mode) in AXI4-Lite
      --AWLOCK     : IN   std_logic;                                   -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      --AWCACHE    : IN   std_logic_vector(3 downto 0);                -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      --AWPROT     : IN   std_logic_vector(2 downto 0);                -- Protection Type       - ignored in this model
      -- ============== AXI4-Lite Write Data Channel
      WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
      WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise) - ignored in AXI-4 Lite
      WVALID     : IN   std_logic;                                     -- Write data is valid
      WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
      -- ============== AXI4-Lite Write Response Channel Signals
      BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
      BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
      -- ============== AXI4-Lite Read Address Channel Signals
      ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
      ARVALID    : IN   std_logic;                                     -- Read address valid
      ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
      --ARLEN      : IN   std_logic_vector(7 downto 0);                -- Read burst length     - must always be 0 in AXI4-Lite
      --ARSIZE     : IN   std_logic_vector(1 downto 0);                -- Read burst size       - must equal host_dw_bytes-2
      --ARBURST    : IN   std_logic_vector(1 downto 0);                -- Read burst mode       - must always be 0 (fixed mode) in AXI4-Lite
      --ARLOCK     : IN   std_logic;                                   -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      --ARCACHE    : IN   std_logic_vector(3 downto 0);                -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      --ARPROT     : IN   std_logic_vector(2 downto 0);                -- Protection Type       - ignored in this model
      -- ============== AXI4-Lite Read Data Channel Signals
      RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
      RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
      RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)

      -- Catapult interface assuming sidebyside packing 
      d_from_ccs : IN   std_logic_vector(cwidth-1 downto 0);           -- Data out of Catapult block
      d_from_vld : IN   std_logic                                      -- Data out is valid
--    d_to_ccs   : OUT  std_logic_vector(cwidth-1 downto 0)            -- Data into Catapult bloc
    );
  END COMPONENT;

  COMPONENT ccs_axi4_slave_mem
    GENERIC(
      rscid           : integer                 := 1;    -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;   -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
      cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
      addr_w          : integer range 1 to 64   := 4;    -- Catapult address bus widths
      nopreload       : integer range 0 to 1    := 0;    -- 1= no preload before Catapult can read
      rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;    -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;    -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;    -- AXI4 Region Map (ignored in this model)
      wBASE_ADDRESS   : integer                 := 0;    -- AXI4 write channel base address alignment based on data bus width
      rBASE_ADDRESS   : integer                 := 0     -- AXI4 read channel base address alignment based on data bus width
     );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                     -- Rising edge clock
      ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Write address ID
      AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
      AWLEN      : IN   std_logic_vector(7 downto 0);                  -- Write burst length
      AWSIZE     : IN   std_logic_vector(2 downto 0);                  -- Write burst size
      AWBURST    : IN   std_logic_vector(1 downto 0);                  -- Write burst mode
      AWLOCK     : IN   std_logic;                                     -- Lock type
      AWCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
      AWPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
      AWQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
      AWREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
      AWUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      AWVALID    : IN   std_logic;                                     -- Write address valid
      AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)

      -- ============== AXI4 Write Data Channel
      WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
      WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
      WLAST      : IN   std_logic;                                     -- Write last
      WUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      WVALID     : IN   std_logic;                                     -- Write data is valid
      WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
      
      -- ============== AXI4 Write Response Channel Signals
      BID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Response ID tag
      BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
      BUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
      BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
      
      -- ============== AXI4 Read Address Channel Signals
      ARID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Read address ID
      ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
      ARLEN      : IN   std_logic_vector(7 downto 0);                  -- Read burst length
      ARSIZE     : IN   std_logic_vector(2 downto 0);                  -- Read burst size
      ARBURST    : IN   std_logic_vector(1 downto 0);                  -- Read burst mode
      ARLOCK     : IN   std_logic;                                     -- Lock type
      ARCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
      ARPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
      ARQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
      ARREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
      ARUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      ARVALID    : IN   std_logic;                                     -- Read address valid
      ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
      
      -- ============== AXI4 Read Data Channel Signals
      RID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Read ID tag
      RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
      RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
      RLAST      : OUT  std_logic;                                     -- Read last
      RUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
      RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
      
      -- Catapult interface
      s_re      : IN   std_logic;                                      -- Catapult attempting read of slave memory
      s_we      : IN   std_logic;                                      -- Catapult attempting write to slave memory
      s_raddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_raddr)
      s_waddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_waddr)
      s_din     : OUT  std_logic_vector(cwidth-1 downto 0);            -- Data into catapult block through this interface
      s_dout    : IN   std_logic_vector(cwidth-1 downto 0);            -- Data out to slave from catapult
      s_rrdy    : OUT  std_logic;                                      -- Read data is valid
      s_wrdy    : OUT  std_logic;                                      -- Slave memory ready for write by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                      -- component is idle - clock can be suppressed
      tr_write_done : IN std_logic;                                    -- transactor resource preload write done
      s_tdone   : IN   std_logic                                       -- Transaction_done in scverify
    );  
  END COMPONENT;

  COMPONENT ccs_axi4_master_read_core
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic                                        -- The component is idle. The next clk can be suppressed
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_read
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                 := 0;      -- Base address 
      BASE_ADDRESSU   : integer                 := 0       -- Upper word for 64-bit Base address 
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic                                        -- The component is idle. The next clk can be suppressed
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_write_core
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_write
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for write burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                 := 0;      -- Base address
      BASE_ADDRESSU   : integer                 := 0       -- Upper word for 64-bit Base address
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Catapult interface
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_core
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xwburstsize     : integer                 := 0;      -- wBurst size for scverify transactor
      xrburstsize     : integer                 := 0;      -- rBurst size for scverify transactor
      xwBASE_ADDRESS  : integer                 := 0;      -- wBase address for scverify transactor
      xrBASE_ADDRESS  : integer                 := 0;      -- rBase address for scverify transactor
      xwBASE_ADDRESSU : integer                 := 0;      -- Upper word for 64-bit wBase address for scverify transactor
      xrBASE_ADDRESSU : integer                 := 0       -- Upper word for 64-bit rBase address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgwBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgrBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgwBurstSize  : IN  std_logic_vector(31 downto 0);            
      cfgrBurstSize  : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;

  COMPONENT ccs_axi4_master_cfg
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      cburst_mode     : integer range 0 to 2    := 0;      -- Burst mode (0==use w/rburstsize, 1==configuration port)
      wburstsize      : integer                 := 0;      -- Catapult configuration option for Write burst size
      rburstsize      : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      use_go          : integer range 0 to 1    := 0;      -- Use the cfgBus stop/go mechanism.  Default not.

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      base_addr_mode  : integer range 0 to 2    := 0;      -- Where base address is specified (0=param, 1=cfg, 2=port)
      wBASE_ADDRESS   : integer                 := 0;      -- AXI4 write channel base address
      rBASE_ADDRESS   : integer                 := 0;      -- AXI4 read channel base address
      wBASE_ADDRESSU  : integer                 := 0;      -- Upper word of 64-bit AXI4 write channel base address
      rBASE_ADDRESSU  : integer                 := 0       -- Upper word of 64-bit AXI4 read channel base address
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- AXI-lite slave interface to program base_addr - address 0, 1, 2
      cfgAWADDR  : IN  std_logic_vector(31 downto 0);
      cfgAWVALID : IN  std_logic;
      cfgAWREADY : OUT std_logic;
      cfgWDATA   : IN  std_logic_vector(31 downto 0);
      cfgWSTRB   : IN  std_logic_vector(3 downto 0);
      cfgWVALID  : IN  std_logic;
      cfgWREADY  : OUT std_logic;
      cfgBRESP   : OUT std_logic_vector(1 downto 0);
      cfgBVALID  : OUT std_logic;
      cfgBREADY  : IN  std_logic;
      cfgARADDR  : IN  std_logic_vector(31 downto 0);
      cfgARVALID : IN  std_logic;
      cfgARREADY : OUT std_logic;
      cfgRDATA   : OUT std_logic_vector(31 downto 0);
      cfgRRESP   : OUT std_logic_vector(1 downto 0);
      cfgRVALID  : OUT std_logic;
      cfgRREADY  : IN  std_logic;

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;

  COMPONENT ccs_axi4_master
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      wburstsize      : integer                 := 0;      -- Catapult configuration option for Write burst size
      rburstsize      : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      wBASE_ADDRESS    : integer                := 0;      -- AXI4 write channel base address
      rBASE_ADDRESS    : integer                := 0;      -- AXI4 read channel base address
      wBASE_ADDRESSU   : integer                := 0;      -- Upper word for 64-bit AXI4 write channel base address
      rBASE_ADDRESSU   : integer                := 0       -- Upper word for 64-bit AXI4 read channel base addressable
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;

COMPONENT ccs_axi4_master_instream_core
    GENERIC(
      rscid           : integer                 := 1;     -- Resource ID
      -- Catapult Bus Configuration generics
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      fpga            : integer range 0 to 1    := 0;      -- Choose the fpga better-route version
      
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xframe_size      : integer                := 16;     -- Number of elements in the frame to be streamed
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready

      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            
      cfgFrameSize   : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      rdy       : OUT  std_logic                                        -- For transactor
    );

END COMPONENT;

COMPONENT ccs_axi4_master_outstream_core
    GENERIC(
      rscid           : integer;                           -- Resource ID
      -- Catapult Bus Configuration generics
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16   := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize       : integer                := 0;      -- Burst size for scverify transactor
      xframe_size      : integer                := 16;     -- Number of elements in the frame to be streamed
      xBASE_ADDRESS    : integer                := 0;      -- Base addess  for scverify transactor
      xBASE_ADDRESSU   : integer                := 0       -- Upper word for 64-bit Base addess  for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Catapult interface
      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            
      cfgFrameSize   : IN  std_logic_vector(31 downto 0);            

      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      vld       : OUT  std_logic                                        -- Core produced data.  Written into transactor "row"
    );

END COMPONENT;

COMPONENT ccs_axi4_master_instream
    GENERIC(
      rscid           : integer                 := 1;     -- Resource ID
      -- Catapult Bus Configuration generics
      frame_size      : integer                 := 16;     -- Number of elements in the frame to be streamed
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      fpga            : integer range 0 to 1    := 0;      -- Choose the fpga better-route version
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall
      
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                 := 0;      -- Base address 
      BASE_ADDRESSU   : integer                 := 0       -- Upper word for 64-bit Base address 
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready

      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      rdy       : OUT  std_logic                                        -- For transactor
    );

END COMPONENT;

COMPONENT ccs_axi4_master_outstream
    GENERIC(
      rscid           : integer;                           -- Resource ID
      -- Catapult Bus Configuration generics
      frame_size      : integer                 := 16;     -- Number of elements in the frame to be streamed
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for Write burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16   := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;     -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                := 0;      -- AXI4 write channel base address
      BASE_ADDRESSU   : integer                := 0       -- Upper word for 64-bit AXI4 write channel base address
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Catapult interface
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      vld       : OUT  std_logic                                        -- Core produced data.  Written into transactor "row"
    );

END COMPONENT;

COMPONENT ccs_axi4_lite_slave_outreg
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS   : integer                  := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    ivld      : IN   std_logic;                                      -- Catapult data ready
    idat      : in   std_logic_vector(cwidth-1 downto 0);            -- Data from catapult

    -- External valid flag
    vld       : OUT  std_logic                                       -- Data valid for AXI read
    );

END COMPONENT;

COMPONENT ccs_axi4_lite_slave_inreg 
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    disable_vld     : integer range 0 to 1    := 0;    -- Disable use of vld signal to stall I/O
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS    : integer                 := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- Catapult interface
    ivld      : OUT   std_logic;                                      -- Data valid.  Duration 1 cycle
    idat      : OUT   std_logic_vector(cwidth-1 downto 0)             -- Data into catapult block through this interface
    );
END COMPONENT;

COMPONENT ccs_axi4_lite_slave_indirect
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS    : integer                 := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    idat      : OUT   std_logic_vector(cwidth-1 downto 0)             -- Data into catapult block through this interface
    );
END COMPONENT;

COMPONENT ccs_axi4_lite_slave_outsync
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 32  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 32 to 64  := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS   : integer                  := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)

    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe - not used in LITE
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    irdy      : OUT  std_logic;                                      -- Catapult data ready
    ivld      : IN   std_logic;                                      -- Catapult data ready
    triosy    : OUT  std_logic                                       -- Data from catapult
    );

END COMPONENT;

COMPONENT ccs_axi4_lite_slave_insync
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 32  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 32 to 64  := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS    : integer                 := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)

    -- Catapult interface
    irdy      : IN    std_logic;
    ivld      : OUT   std_logic;
    triosy    : OUT   std_logic                                       -- // transactor uses 
    );
END COMPONENT;


  -- ==============================================================
  -- APB Components

  -- Used to define the APB bus definition (direction of signals is from the slave's perspective)
  COMPONENT apb_busdef
    GENERIC(
      width        : INTEGER RANGE 1 TO 32 := 32;           -- Number of bits in an element
      addr_width   : INTEGER RANGE 1 TO 32 := 1             -- Number of address bits to address 'words' elements
    );
    PORT(
      -- APB interface
      PCLK      : IN   std_logic;                           -- Rising edge clock
      PRESETn   : IN   std_logic;                           -- Active LOW synchronous reset
      PADDR     : IN   std_logic_vector(addr_width-1 downto 0);  -- APB Bridge driven address bus (32 bit max)
      PSELx     : IN   std_logic;                           -- APB Bridge driven select for this slave
      PWRITE    : IN   std_logic;                           -- APB Bridge driven read/write signal (0=read)
      PENABLE   : IN   std_logic;                           -- APB Bridge driven enable signal
      PWDATA    : IN   std_logic_vector(width-1 downto 0);  -- APB Bridge driven data to write to slave (32 bit max)
      PRDATA    : OUT  std_logic_vector(width-1 downto 0);  -- Slave driven data back to APB Bridge (32 bit max)
      PREADY    : OUT  std_logic;                           -- Slave driven signal to extend transfer cycles (1=ready)
      PSLVERR   : OUT  std_logic                            -- Slave driven signal indicating transfer failed (1=fail)
    );
  END COMPONENT;

  COMPONENT apb_master
    GENERIC(
      words        : INTEGER RANGE 1 TO 256 := 1;           -- Number of addressable elements
      width        : INTEGER RANGE 1 TO 32 := 32;           -- Number of bits in an element
      addr_width   : INTEGER RANGE 1 TO 32 := 1             -- Number of address bits to address 'words' elements
    );
    PORT(
      -- APB interface
      PCLK      : IN   std_logic;                           -- Rising edge clock
      PRESETn   : IN   std_logic;                           -- Active LOW synchronous reset
      PADDR     : OUT  std_logic_vector(30 downto 0);       -- APB Bridge driven address bus (32 bit max)
      PSELx     : OUT  std_logic;                           -- APB Bridge driven select for this slave
      PWRITE    : OUT  std_logic;                           -- APB Bridge driven read/write signal (0=read)
      PENABLE   : OUT  std_logic;                           -- APB Bridge driven enable signal
      PWDATA    : OUT  std_logic_vector(width-1 downto 0);  -- APB Bridge driven data to write to slave (32 bit max)
      PRDATA    : IN   std_logic_vector(width-1 downto 0);  -- Slave driven data back to APB Bridge (32 bit max)
      PREADY    : IN   std_logic;                           -- Slave driven signal to extend transfer cycles (1=ready)
      PSLVERR   : IN   std_logic;                           -- Slave driven signal indicating transfer failed (1=fail)
      -- Catapult interface
      m_rw      : IN   std_logic;                           -- read/write
      m_strobe  : IN   std_logic;                           -- initiate a bus transfer
      m_adr     : IN   std_logic_vector(addr_width-1 downto 0); -- target address
      m_din     : OUT  std_logic_vector(width-1 downto 0);  -- data in from slave
      m_dout    : IN   std_logic_vector(width-1 downto 0);  -- data out to slave
      m_rdy     : OUT  std_logic                            -- ready for transfer (1=ready)
    );
  END COMPONENT;

  -- APB slave memory
  COMPONENT apb_slave_mem
    GENERIC(
      words          : INTEGER RANGE 1 TO 256 := 1;            -- Number of addressable elements
      width          : INTEGER RANGE 1 TO 32 := 32;           -- Number of bits in an element
      addr_width     : INTEGER RANGE 1 TO 32 := 1;            -- Number of address bits to address 'words' elements
      num_rwports    : INTEGER RANGE 1 TO 100 := 1;           -- Number of register file "ports"
      nopreload      : INTEGER RANGE 0 TO 1 := 0              -- 1=disable required preload before Catapult can read
    );
    PORT(
      -- APB interface
      PCLK      : IN   std_logic;                           -- Rising edge clock
      PRESETn   : IN   std_logic;                           -- Active LOW synchronous reset
      PADDR     : IN   std_logic_vector(30 downto 0);       -- APB Bridge driven address bus (32 bit max)
      PSELx     : IN   std_logic;                           -- APB Bridge driven select for this slave
      PWRITE    : IN   std_logic;                           -- APB Bridge driven read/write signal (0=read)
      PENABLE   : IN   std_logic;                           -- APB Bridge driven enable signal
      PWDATA    : IN   std_logic_vector(width-1 downto 0);  -- APB Bridge driven data to write to slave (32 bit max)
      PRDATA    : OUT  std_logic_vector(width-1 downto 0);  -- Slave driven data back to APB Bridge (32 bit max)
      PREADY    : OUT  std_logic;                           -- Slave driven signal to extend transfer cycles (1=ready)
      PSLVERR   : OUT  std_logic;                           -- Slave driven signal indicating transfer failed (1=fail)
      -- Catapult interface
      s_rw      : IN   std_logic_vector(num_rwports-1 downto 0);            -- read/write
      s_strobe  : IN   std_logic_vector(num_rwports-1 downto 0);            -- Catapult attempting read of slave
      s_adr     : IN   std_logic_vector(num_rwports*addr_width-1 downto 0); -- Catapult addressing into memory
      s_din     : OUT  std_logic_vector(num_rwports*width-1 downto 0);      -- Data into catapult block through this interface
      s_dout    : IN   std_logic_vector(num_rwports*width-1 downto 0);      -- Data out to slave from catapult
      s_rdy     : OUT  std_logic_vector(num_rwports-1 downto 0)             -- Slave memory ready for read (1=ready)
    );
  END COMPONENT;

  -- ==============================================================
  -- Internally referenced components

  COMPONENT amba_generic_reg
    GENERIC (
      width    : INTEGER := 1;
      ph_en    : INTEGER RANGE 0 TO 1 := 1;
      has_en   : INTEGER RANGE 0 TO 1 := 1
    );
    PORT (
      clk     : IN  std_logic;
      en      : IN  std_logic;
      arst    : IN  std_logic;
      srst    : IN  std_logic;
      d       : IN  std_logic_vector(width-1 DOWNTO 0);
      z       : OUT std_logic_vector(width-1 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT amba_pipe_ctrl
    GENERIC (
      rscid    : INTEGER := 0;
      width    : INTEGER := 8;
      sz_width : INTEGER := 8;
      fifo_sz  : INTEGER RANGE 0 TO 128 := 8;
      ph_en    : INTEGER RANGE 0 TO 1 := 1
    );
    PORT (
      clk      : IN  std_logic;
      en       : IN  std_logic;
      arst     : IN  std_logic;
      srst     : IN  std_logic;
      din_vld  : IN  std_logic;
      din_rdy  : OUT std_logic;
      din      : IN  std_logic_vector(width-1 DOWNTO 0);
      dout_vld : OUT std_logic;
      dout_rdy : IN  std_logic;
      dout     : OUT std_logic_vector(width-1 DOWNTO 0);
      sd       : OUT std_logic_vector(sz_width-1 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT amba_pipe
    GENERIC (
      rscid    : INTEGER := 0;
      width    : INTEGER := 8;
      sz_width : INTEGER := 8;
      fifo_sz  : INTEGER RANGE 0 TO 128 := 8;
      ph_en    : INTEGER RANGE 0 TO 1 := 1
    );
    PORT (
      -- clock
      clk      : IN  std_logic;
      en       : IN  std_logic;
      arst     : IN  std_logic;
      srst     : IN  std_logic;
      -- writer
      din_rdy  : OUT std_logic;
      din_vld  : IN  std_logic;
      din      : IN  std_logic_vector(width-1 DOWNTO 0);
      -- reader
      dout_rdy : IN  std_logic;
      dout_vld : OUT std_logic;
      dout     : OUT std_logic_vector(width-1 DOWNTO 0);
      -- size
      sz       : OUT std_logic_vector(sz_width-1 DOWNTO 0);
      sz_req   : in  std_logic
    );
  END COMPONENT;

  COMPONENT amba_ctrl_in_buf_wait
    GENERIC (
      width    : INTEGER := 8
    );
    PORT (
      clk      : IN  std_logic;
      arst     : IN  std_logic;
      irdy   : IN  std_logic;
      ivld   : OUT std_logic;
      idat   : OUT std_logic_vector(width-1 DOWNTO 0);
      rdy    : OUT std_logic;
      vld    : IN  std_logic;
      dat    : IN  std_logic_vector(width-1 DOWNTO 0);
      is_idle : out std_logic
    );
  END COMPONENT;

  COMPONENT ML_amba_ctrl_in_buf_wait
    GENERIC (
      width    : INTEGER := 8
    );
    PORT (
      clk      : IN  std_logic;
      arst     : IN  std_logic;
      irdy   : IN  std_logic;
      ivld   : OUT std_logic;
      idat   : OUT std_logic_vector(width-1 DOWNTO 0);
      rdy    : OUT std_logic;
      vld    : IN  std_logic;
      dat    : IN  std_logic_vector(width-1 DOWNTO 0);
      is_idle : out std_logic
    );
  END COMPONENT;

COMPONENT ML_ccs_axi4_master_fpga_instream_core
    GENERIC(
      rscid           : integer                 := 1;     -- Resource ID
      -- Catapult Bus Configuration generics
      frame_size      : integer                 := 16;     -- Number of elements in the frame to be streamed
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready

      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      rdy       : OUT  std_logic                                        -- For transactor
    );
END COMPONENT;

  
  -- ==============================================================
  -- AMBA Protocol Constants

  -- AxBURST modes
  CONSTANT AXI4_AxBURST_FIXED    : std_logic_vector(1 downto 0) := "00";
  CONSTANT AXI4_AxBURST_INCR     : std_logic_vector(1 downto 0) := "01";
  CONSTANT AXI4_AxBURST_WRAP     : std_logic_vector(1 downto 0) := "10";
  CONSTANT AXI4_AxBURST_RESERVED : std_logic_vector(1 downto 0) := "11";
  -- AxLOCK modes
  CONSTANT AXI4_AxLOCK_NORMAL    : std_logic                    := '0';
  CONSTANT AXI4_AxLOCK_EXCLUSIVE : std_logic                    := '1';
  -- Memory types W and R mostly the xame
  CONSTANT AXI4_AWCACHE_NB        : std_logic_vector(3 downto 0) := "0000";
  CONSTANT AXI4_AWCACHE_B         : std_logic_vector(3 downto 0) := "0001";
  CONSTANT AXI4_AWCACHE_NORM_NCNB : std_logic_vector(3 downto 0) := "0010"; --
  CONSTANT AXI4_AWCACHE_NORM_NCB  : std_logic_vector(3 downto 0) := "0011" ;
  CONSTANT AXI4_AWCACHE_WTNA      : std_logic_vector(3 downto 0) := "0110";
  CONSTANT AXI4_AWCACHE_WTRA      : std_logic_vector(3 downto 0) := "0110";
  CONSTANT AXI4_AWCACHE_WTWA      : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_AWCACHE_WTRWA     : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_AWCACHE_WBNA      : std_logic_vector(3 downto 0) := "0111";
  CONSTANT AXI4_AWCACHE_WBRA      : std_logic_vector(3 downto 0) := "0111";
  CONSTANT AXI4_WACACHE_WBWA      : std_logic_vector(3 downto 0) := "1111";
  CONSTANT AXI4_AWCACHE_WBRWA     : std_logic_vector(3 downto 0) := "1111";
  CONSTANT AXI4_ARCACHE_NB        : std_logic_vector(3 downto 0) := "0000";
  CONSTANT AXI4_ARCACHE_B         : std_logic_vector(3 downto 0) := "0001";
  CONSTANT AXI4_ARCACHE_NORM_NCNB : std_logic_vector(3 downto 0) := "0010"; --
  CONSTANT AXI4_ARCACHE_NORM_NCB  : std_logic_vector(3 downto 0) := "0011" ;
  CONSTANT AXI4_ARCACHE_WTNA      : std_logic_vector(3 downto 0) := "1010";
  CONSTANT AXI4_ARCACHE_WTRA      : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_ARCACHE_WTWA      : std_logic_vector(3 downto 0) := "1010";
  CONSTANT AXI4_ARCACHE_WTRWA     : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_ARCACHE_WBNA      : std_logic_vector(3 downto 0) := "1011";
  CONSTANT AXI4_ARCACHE_WBRA      : std_logic_vector(3 downto 0) := "1111";
  CONSTANT AXI4_ARCACHE_WBWA      : std_logic_vector(3 downto 0) := "1011";
  CONSTANT AXI4_ARCACHE_WBRWA     : std_logic_vector(3 downto 0) := "1111";
  -- QOS pre-defines
  CONSTANT AXI4_AxQOS_NONE        : std_logic_vector(3 downto 0) := "0000";
  -- AxSIZE byte sizes
  CONSTANT AXI4_AxSIZE_001_BYTE  : std_logic_vector(2 downto 0) := "000";
  CONSTANT AXI4_AxSIZE_002_BYTE  : std_logic_vector(2 downto 0) := "001";
  CONSTANT AXI4_AxSIZE_004_BYTE  : std_logic_vector(2 downto 0) := "010";
  CONSTANT AXI4_AxSIZE_008_BYTE  : std_logic_vector(2 downto 0) := "011";
  CONSTANT AXI4_AxSIZE_016_BYTE  : std_logic_vector(2 downto 0) := "100";
  CONSTANT AXI4_AxSIZE_032_BYTE  : std_logic_vector(2 downto 0) := "101";
  CONSTANT AXI4_AxSIZE_064_BYTE  : std_logic_vector(2 downto 0) := "110";
  CONSTANT AXI4_AxSIZE_128_BYTE  : std_logic_vector(2 downto 0) := "111";
  -- AxPROT bit fields
  CONSTANT AXI4_AxPROT_b0_UNPRIV   : std_logic := '0';
  CONSTANT AXI4_AxPROT_b0_PRIV     : std_logic := '1';
  CONSTANT AXI4_AxPROT_b1_SECURE   : std_logic := '0';
  CONSTANT AXI4_AxPROT_b1_UNSECURE : std_logic := '1';
  CONSTANT AXI4_AxPROT_b2_DATA     : std_logic := '0';
  CONSTANT AXI4_AxPROT_b2_INSTR    : std_logic := '1';
  -- xRESP response codes
  CONSTANT AXI4_xRESP_OKAY         : std_logic_vector(1 downto 0) := "00";
  CONSTANT AXI4_xRESP_EXOKAY       : std_logic_vector(1 downto 0) := "01";
  CONSTANT AXI4_xRESP_SLVERR       : std_logic_vector(1 downto 0) := "10";
  CONSTANT AXI4_xRESP_DECERR       : std_logic_vector(1 downto 0) := "11";

  -- Utility function(s) to support debug needs
  FUNCTION bits ( size : INTEGER) RETURN INTEGER;
  FUNCTION slv2bin(vec: std_logic_vector) RETURN string;
  FUNCTION slv2hex(vec: std_logic_vector) RETURN string;

END PACKAGE amba_comps;

PACKAGE BODY amba_comps IS

   -- Find the number of bits required to represent an unsigned
   -- number less than size
  FUNCTION bits (size : integer) RETURN INTEGER IS
  BEGIN
    IF (size < 0) THEN RETURN 0;
    ELSIF (size = 0) THEN RETURN 1;
    ELSE
      FOR i IN 1 TO size LOOP
        IF (2**i >= size) THEN
          RETURN i;
        END IF;
      END LOOP;
      RETURN 0;
    END IF;
  END;

   -- Convert an std_logic_vector to a (hex)string for printing
   -- vec needs to be a multiple of 4 in size
  FUNCTION slv2hex(vec: std_logic_vector) RETURN string IS
      variable quad : std_logic_vector(3 downto 0);
      constant ne: integer := vec'length/4;
      variable s: string(1 to ne);
   BEGIN
      if vec'length mod 4 /= 0 then
         assert false
         report "slv2hex called with slv lenght that is not a multiple of 4";
         return s;
      end if;
      for i in 0 to ne-1 loop
         quad := vec(4*i+3 downto 4*i);
         case quad is
            when x"0" => s(ne-i) := '0';
            when x"1" => s(ne-i) := '1';
            when x"2" => s(ne-i) := '2';
            when x"3" => s(ne-i) := '3';
            when x"4" => s(ne-i) := '4';
            when x"5" => s(ne-i) := '5';
            when x"6" => s(ne-i) := '6';
            when x"7" => s(ne-i) := '7';
            when x"8" => s(ne-i) := '8';
            when x"9" => s(ne-i) := '9';
            when x"A" => s(ne-i) := 'A';
            when x"B" => s(ne-i) := 'B';
            when x"C" => s(ne-i) := 'C';
            when x"D" => s(ne-i) := 'D';
            when x"E" => s(ne-i) := 'E';
            when x"F" => s(ne-i) := 'F';
            when others => s(ne-i) := '-';
         end case;
      end loop;
      return s;
   END;

   -- Convert an std_logic_vector to a (binary)string for printing
   FUNCTION slv2bin(vec: std_logic_vector) RETURN string IS
      VARIABLE stmp: string(vec'left+1 downto 1);
   BEGIN
      FOR i in vec'reverse_range LOOP
         IF (vec(i) = 'U') THEN
            stmp(i+1) := 'U';
         ELSIF (vec(i) = 'X') THEN
            stmp(i+1) := 'X';
         ELSIF (vec(i) = '0') THEN
            stmp(i+1) := '0';
         ELSIF (vec(i) = '1') THEN
            stmp(i+1) := '1';
         ELSIF (vec(i) = 'Z') THEN
            stmp(i+1) := 'Z';
         ELSIF (vec(i) = 'W') THEN
            stmp(i+1) := 'W';
         ELSIF (vec(i) = 'L') THEN
            stmp(i+1) := 'L';
         ELSIF (vec(i) = 'H') THEN
            stmp(i+1) := 'H';
         ELSE
            stmp(i+1) := '-';
         END IF;
      END LOOP;
      RETURN stmp;
   END;

END amba_comps;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_libs/interfaces/amba/ccs_axi4_slave_mem.vhd 

-- --------------------------------------------------------------------------
-- DESIGN UNIT:        ccs_axi4_slave_mem
--
-- DESCRIPTION:
--   This model implements an AXI-4 Slave memory interface for use in 
--   Interface Synthesis in Catapult. The component details are described in the datasheet.
--
--   AXI/Catapult read/write to the same address in the same cycle is non-determinant
--
-- Notes:
--  1. This model implements a local memory of size {cwidth x depth}.
--     If the Catapult operation requires a memory width cwidth <= AXI bus width
--     this model will zero-pad the high end bits as necessary.
-- CHANGE LOG:
--  01/29/19 - Add reset phase and separate base address for read/write channels
--  11/26/18 - Add burst and other tweaks
--  02/28/18 - Initial implementation
--
-- -------------------------------------------------------------------------------
--  Memory Organization
--   This model is designed to provide storage for only the bits/elements that
--   the Catapult core actually interacts with.
--   The user supplies a base address for the AXI memory store via BASE_ADDRESS
--   parameter.  
-- Example:
--   C++ array declared as "ac_int<7,false>  coeffs[4];"
--   results in a Catapult operator width (op_width) of 7,
--   and cwidth=7 and addr_w=2 (addressing 4 element locations).
--   The library forces DATA_WIDTH to be big enough to hold
--   cwidth bits, rounded up to power-of-2 as needed.
--
--   The AXI address scheme addresses bytes and so increments
--   by number-of-bytes per data transaction, plus the BASE_ADDRESS. 
--   The top and left describe the AXI view of the memory. 
--   The bottom and right describe the Catapult view of the memory.
--
--      AXI-4 SIGNALS
--      ADDR_WIDTH=4        DATA_WIDTH=32
--        AxADDR               xDATA
--                    31                       0
--                    +------------+-----------+
--      BA+0000       |            |           |
--                    +------------+-----------+
--      BA+0000       |            |           |
--                    +------------+===========+
--      BA+1100       |            |  elem3    |    11
--                    +------------+===========+
--      BA+1000       |            |  elem2    |    10
--                    +------------+===========+
--      BA+0100       |            |  elem1    |    01
--                    +------------+===========+
--      BA+0000       |            |  elem0    |    00
--                    +------------+===========+
--                                 6           0
--                                   s_din/out     s_addr
--                                   cwidth=7      addr_w=2
--                                         CATAPULT SIGNALS
--
-- -------------------------------------------------------------------------------

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;       
  USE std.textio.all;
  USE ieee.std_logic_textio.all;
  USE ieee.math_real.all;


USE work.amba_comps.all;

ENTITY ccs_axi4_slave_mem IS
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    depth           : integer                 := 16;   -- Number of addressable elements (up to 20bit address)
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    addr_w          : integer range 1 to 64   := 4;    -- Catapult address bus widths
    nopreload       : integer range 0 to 1    := 0;    -- 1= no preload before Catapult can read
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    ID_WIDTH        : integer range 1 to 16   := 1;    -- AXI4 ID field width (ignored in this model)
    USER_WIDTH      : integer range 1 to 32   := 1;    -- AXI4 User field width (ignored in this model)
    REGION_MAP_SIZE : integer range 1 to 15   := 1;    -- AXI4 Region Map (ignored in this model)
    wBASE_ADDRESS   : integer                 := 0;    -- AXI4 write channel base address alignment based on data bus width
    rBASE_ADDRESS   : integer                 := 0     -- AXI4 read channel base address alignment based on data bus width
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Write address ID
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWLEN      : IN   std_logic_vector(7 downto 0);                  -- Write burst length
    AWSIZE     : IN   std_logic_vector(2 downto 0);                  -- Write burst size
    AWBURST    : IN   std_logic_vector(1 downto 0);                  -- Write burst mode
    AWLOCK     : IN   std_logic;                                     -- Lock type
    AWCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
    AWPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
    AWQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
    AWREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
    AWUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WLAST      : IN   std_logic;                                     -- Write last
    WUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Response ID tag
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Read address ID
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARLEN      : IN   std_logic_vector(7 downto 0);                  -- Read burst length
    ARSIZE     : IN   std_logic_vector(2 downto 0);                  -- Read burst size
    ARBURST    : IN   std_logic_vector(1 downto 0);                  -- Read burst mode
    ARLOCK     : IN   std_logic;                                     -- Lock type
    ARCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
    ARPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
    ARQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
    ARREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
    ARUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Read ID tag
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RLAST      : OUT  std_logic;                                     -- Read last
    RUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    s_re      : IN   std_logic;                                      -- Catapult attempting read of slave memory
    s_we      : IN   std_logic;                                      -- Catapult attempting write to slave memory
    s_raddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_raddr)
    s_waddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_waddr)
    s_din     : OUT  std_logic_vector(cwidth-1 downto 0);            -- Data into catapult block through this interface
    s_dout    : IN   std_logic_vector(cwidth-1 downto 0);            -- Data out to slave from catapult
    s_rrdy    : OUT  std_logic;                                      -- Read data is valid
    s_wrdy    : OUT  std_logic;                                      -- Slave memory ready for write by Catapult (1=ready)
    is_idle   : OUT  std_logic;                                      -- component is idle - clock can be suppressed
    -- Transactor/scverify support
    tr_write_done : IN std_logic;                                    -- transactor resource preload write done
    s_tdone       : IN std_logic                                     -- Transaction_done in scverify
    );
  

    -- Always rule for checking component parameter values
    --  addr_w == bits(depth)
    --    used to ensure that the width of the address bus on the Catapult side
    --    is capable of addressing 'depth' number of elements. 'depth' will be
    --    determined by the array size operator parameter 'size'
    --    (see the PROP_MAP_size attribute)
    --  ADDR_WIDTH >= addr_w
    --    used to ensure that the address width of the Catapult side is
    --    large enough to accommodate the address width of the AXI-4 bus.
    --    (may need some work to align byte addresses)
    --  ADDR_WIDTH >= 32
    --    ensure that the minimum address space is 4k (AXI requirement)
    --  cwidth == 8 + (op_width>8)*8 + (op_width>16)*16 + (op_width>32)*32 + 
    --                (op_width>64)*64 + (op_width>128)*128 + (op_width>256)*256 +
    --                (op_width>512)*512
    --    used to "round up" the operator width 'op_width' to the next power
    --    of two value (8, 16, 32, 64, 128, 256, 512, 1024)
    --    (see the PROP_MAP_width attribute)
    --  DATA_WIDTH >= cwidth
    --    used to ensure that the Catapult data width is large enough to
    --    accommodate the data width of the AXI-4 bus.
    --    - must be power-of-2 bytes.
    --    - #bits must be some positive integer number of bytes.
    --     Note: user can override DATA_WIDTH from the MAP_TO_MODULE
    --     directive during interface synthesis. No checking is done
    --     to ensure that the override value is a power-of-2 bytes.

END ccs_axi4_slave_mem;

ARCHITECTURE rtl of ccs_axi4_slave_mem IS

  -- Signals for current and next state values
  TYPE   read_state_t IS (axi4r_idle, axi4r_read);
  TYPE   write_state_t IS (axi4w_idle, axi4w_write, axi4w_write_done,  axi4w_catwrite, axi4w_catwrite_done);
  SIGNAL read_state       : read_state_t;
  SIGNAL write_state      : write_state_t;

  -- Memory embedded in this slave
  TYPE   mem_type IS ARRAY (depth-1 downto 0) of std_logic_vector(cwidth-1 downto 0);
  SIGNAL mem                : mem_type;


  -- In/out connections and constant outputs  
  SIGNAL AWREADY_reg : std_logic;
  SIGNAL AWID_reg    : std_logic_vector(ID_WIDTH-1 downto 0);
  SIGNAL WREADY_reg  : std_logic;
  SIGNAL BRESP_reg   : std_logic_vector(1 downto 0);
  SIGNAL BVALID_reg  : std_logic;
  SIGNAL ARREADY_reg : std_logic;
  SIGNAL ARID_reg    : std_logic_vector(ID_WIDTH-1 downto 0);
  SIGNAL RDATA_reg   : std_logic_vector(DATA_WIDTH-1 downto 0);
  SIGNAL RRESP_reg   : std_logic_vector(1 downto 0);
  SIGNAL RLAST_reg   : std_logic;
  SIGNAL RVALID_reg  : std_logic;
  SIGNAL s_din_reg   : std_logic_vector(cwidth-1 downto 0);
  SIGNAL s_rrdy_reg  : std_logic;
  SIGNAL s_wrdy_reg  : std_logic;

  SIGNAL rCatOutOfOrder : std_logic;
  SIGNAL catIsReading   : std_logic;
  SIGNAL next_raddr     : integer;
  
  SIGNAL readBurstCnt: std_logic_vector(7 downto 0);   -- how many are left
  SIGNAL wbase_addr   : std_logic_vector(ADDR_WIDTH-1 downto 0);
  SIGNAL rbase_addr   : std_logic_vector(ADDR_WIDTH-1 downto 0);
  SIGNAL address     : std_logic_vector(ADDR_WIDTH-1 downto 0);
  SIGNAL addrShift : integer;
  SIGNAL readAddr : integer;
  SIGNAL writeAddr : integer;
  SIGNAL int_ARESETn : std_logic;
  
-- catapult address sizes are smaller and cause problems used with axi address sizes
  function extCatAddr(catAddr : std_logic_vector(addr_w -1 downto 0))
    return std_logic_vector is
  
    variable axiAddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
  
  begin
    axiAddr := (others => '0');
    axiAddr(addr_w -1 downto 0) := catAddr;
    return axiAddr;
  end function extCatAddr;

BEGIN
  
  int_ARESETn <= ARESETn when (rst_ph = 0) else (not ARESETn);

  addrShift <= 0 when (DATA_WIDTH/8 <= 1)   else 
               1 when (DATA_WIDTH/8 <= 2)   else
               2 when (DATA_WIDTH/8 <= 4)   else
               3 when (DATA_WIDTH/8 <= 8)   else
               4 when (DATA_WIDTH/8 <= 16)  else
               5 when (DATA_WIDTH/8 <= 32)  else
               6 when (DATA_WIDTH/8 <= 64)  else
               7 when (DATA_WIDTH/8 <= 128) else
               0;

  -- unused outputs
  BUSER   <= (others => '0');
  RUSER   <= (others => '0');
  is_idle <= '0';
  
  AWREADY <= AWREADY_reg;
  WREADY  <= WREADY_reg ;
  BID     <= AWID_reg;
  BRESP   <= BRESP_reg  ;
  BVALID  <= BVALID_reg ;
  ARREADY <= ARREADY_reg;
  RID     <= ARID_reg;
  RDATA   <= RDATA_reg  ;
  RRESP   <= RRESP_reg  ;
  RLAST   <= RLAST_reg  ;
  RVALID  <= RVALID_reg ;
  s_din   <= s_din_reg  ;
  s_wrdy  <= s_wrdy_reg and (not s_tdone);
  s_rrdy  <= s_rrdy_reg and (not rCatOutOfOrder);

  wbase_addr <= std_logic_vector(to_unsigned(wBASE_ADDRESS, wbase_addr'length));
  rbase_addr <= std_logic_vector(to_unsigned(rBASE_ADDRESS, rbase_addr'length));
  
  -- pragma translate_off
  -- error checks.  Keep consistent with axi4_master.v/vhd
  -- all data widths the same
  errChk: process
    variable nBytes : std_logic_vector(31 downto 0);
    variable nBytes2 : std_logic_vector(31 downto 0);
  begin  -- process errChk
    nBytes := std_logic_vector(to_unsigned(DATA_WIDTH/8, 32));
    if (cwidth > DATA_WIDTH) then
      report  "Catapult(cwidth=" & integer'image(cwidth) & ") cannot be greater than AXI(DATA_BUS="
        & integer'image(DATA_WIDTH) & ")."
        severity error;
    end if;
    if ( (DATA_WIDTH mod 8) /= 0) then
      report  "Data bus width(DATA_WIDTH=" & integer'image(DATA_WIDTH) & ") not a discrete number of bytes."
        severity error;
    end if;
    if (to_integer(unsigned(nBytes)) = 0) then 
      report  "Data bus width(DATA_WIDTH=" & integer'image(DATA_WIDTH) & ") must be at least 1 byte."
        severity error;
    end if;
    nBytes2 := std_logic_vector(to_unsigned((DATA_WIDTH/8) - 1, 32));
    nBytes2 := nBytes  and nBytes2;
    if ( to_integer(unsigned(nBytes2)) /= 0) then
      report  "Data bus width must be power-of-2 number of bytes(DATA_WIDTH/8=" & integer'image(DATA_WIDTH/8) & ")"
        severity error;
    end if;
    if (ADDR_WIDTH < 12) then
      report  "AXI bus address width(ADDR_WIDTH=" & integer'image(ADDR_WIDTH) & ") must be at least 12 to address 4K memory space."
        severity error;
    end if;
    wait;
  end process errChk;
  -- pragma translate_on
  
  -- AXI4 Bus Read processing
  axiRead: process(ACLK, int_ARESETn)
    -- pragma translate_off
    variable buf : line;
    -- pragma translate_on
    variable useAddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
    variable useAddr2 : std_logic_vector(ADDR_WIDTH-1 downto 0);
  begin
    if (int_ARESETn = '0') then
      read_state <= axi4r_idle;
      ARREADY_reg <= '1';
      ARID_reg <= (others => '0');
      RDATA_reg <= (others => '0');
      RRESP_reg <= AXI4_xRESP_OKAY;
      RLAST_reg <= '0';
      RVALID_reg <= '0';
      readAddr <= 0;
      readBurstCnt <= (others => '0');
    elsif rising_edge(ACLK) then
      if ((read_state = axi4r_idle) and (ARVALID = '1')) then
        useAddr := std_logic_vector(shift_right(unsigned(ARADDR) - unsigned(rbase_addr), addrShift));
        -- Protect from out of range addressing
        if (unsigned(useAddr) < depth) then
          if (cwidth < DATA_WIDTH) then
            RDATA_reg(DATA_WIDTH-1 downto cwidth) <= (others => '0');
            RDATA_reg(cwidth-1 downto 0) <= mem(to_integer(unsigned(useAddr)));
          else
            RDATA_reg <= mem(to_integer(unsigned(useAddr)));
          end if;
          --write(buf, string'("Slave AXI1 read:mem[0x"));
          --write(buf,  slv2hex(useAddr));
          --write(buf, string'("]=0x"));
          --write(buf,  slv2hex(mem(to_integer(unsigned(useAddr)))));
          --write(buf, string'(" at T="));
          --write(buf, now);
          --writeline(output, buf);
        else
          -- pragma translate_off
          write(buf, string'("Error:  Out-of-range AXI memory read access:0x"));
          write(buf,  slv2hex(ARADDR));
          write(buf, string'(" at T="));
          write(buf, now);
          writeline(output, buf);
          -- pragma translate_on
        end if;
        RRESP_reg <= AXI4_xRESP_OKAY;
        readAddr <= to_integer(unsigned(useAddr));
        readBurstCnt <= ARLEN;
        if (unsigned(ARLEN) = 0) then
          ARREADY_reg <= '0';
          RLAST_reg <= '1';
        end if;
        RVALID_reg <= '1';
        ARID_reg <= ARID;
        read_state <= axi4r_read;
      elsif (read_state = axi4r_read) then
        if (RREADY = '1') then
          if (unsigned(readBurstCnt) = 0) then
            -- we already sent the last data
            ARREADY_reg <= '1';
            RRESP_reg <= AXI4_xRESP_OKAY;
            RLAST_reg <= '0';
            RVALID_reg <= '0';
            read_state <= axi4r_idle;               
          else
            useAddr2 := std_logic_vector(to_unsigned(readAddr + 1, useAddr2'length));
            readAddr <= readAddr + 1;
            -- Protect from out of range addressing
            if (unsigned(useAddr2) < depth) then
              if (cwidth < DATA_WIDTH) then
                RDATA_reg(DATA_WIDTH-1 downto cwidth) <= (others => '0');
                RDATA_reg(cwidth-1 downto 0) <=  mem(to_integer(unsigned(useAddr2)));
              else
                RDATA_reg <=  mem(to_integer(unsigned(useAddr2)));
              end if;
              --write(buf, string'("Slave AXI2 read:mem[0x"));
              --write(buf,  slv2hex(useAddr2));
              --write(buf, string'("]=0x"));
              --write(buf,  slv2hex(mem(to_integer(unsigned(useAddr2)))));
              --write(buf, string'(" at T="));
              --write(buf, now);
              --writeline(output, buf);
            else
              -- We bursted right off the end of the array
              -- pragma translate_off
              write(buf, string'("Error:  Out-of-range AXI memory read access:0x"));
              write(buf,  slv2hex(ARADDR));
              write(buf, string'(" at T="));
              write(buf, now);
              writeline(output, buf);
              -- pragma translate_on
            end if;
            readBurstCnt <= std_logic_vector(unsigned(readBurstCnt) - 1);
            if ((unsigned(readBurstCnt) - 1) = 0) then
              ARREADY_reg <= '0';        
              RRESP_reg <= AXI4_xRESP_OKAY;
              RLAST_reg <= '1';
            end if;
            RVALID_reg <= '1';
          end if;
        end if;
      end if;
    end if;
  end process;  -- axiRead process

   -- AXI and catapult write processing.
   -- Catapult write is one-cycle long so basically a write can happen
   -- in any axi state.  AXI has precedence in that catapult write is processed
   -- first at each cycle
  axiWrite: process(ACLK, int_ARESETn)
    -- pragma translate_off
    variable buf : line;
    -- pragma translate_on
    variable i : integer;
    variable useAddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
    variable useAddr2 : std_logic_vector(ADDR_WIDTH-1 downto 0);
  begin
    if (int_ARESETn = '0') then
      AWREADY_reg <= '1';
      AWID_reg <= (others => '0');
      WREADY_reg <= '1';
      BRESP_reg <= AXI4_xRESP_OKAY;
      BVALID_reg <= '0';
      write_state <= axi4w_idle;
      writeAddr <= 0;
      s_wrdy_reg <= '0';
      -- pragma translate_off
      for i in 0 to depth-1 loop 
        mem(i) <= (others => '0');
      end loop;
      -- pragma translate_on
    elsif rising_edge(ACLK) then
      -- When in idle state, catapult and AXI can both initiate writes.
      -- If to the same address, then AXI wins... in this implementation
      if ((s_we = '1') and (write_state = axi4w_idle) and (s_tdone = '0')) then
        mem(to_integer(unsigned(s_waddr))) <= s_dout;
        --write(buf, string'("Slave CAT1 write:mem[0x"));
        --write(buf,  slv2hex(s_waddr));
        --write(buf, string'("]=0x"));
        --write(buf,  slv2hex(s_dout));
        --write(buf, string'(" at T="));
        --write(buf, now);
        --writeline(output, buf);
      end if;
      if ((write_state = axi4w_idle) and (AWVALID = '1')) then
        s_wrdy_reg <= '0';
        AWREADY_reg <= '0';
        AWID_reg <= AWID;
        useAddr := std_logic_vector(shift_right(unsigned(AWADDR) - unsigned(wbase_addr), addrShift));
        -- $display("AWADDR=%d base_address=%d addrShift=%d useAddr=%d at T=%t",
        -- AWADDR, base_address, addrShift, useAddr, $time);
        if (WVALID = '1') then
          -- allow for address and data to be presented in one cycle
          -- Check for the write to be masked
          if (unsigned(WSTRB) /= 0) then -- a byte at a time.  Watch for cwidth much less than DATA_WIDTH
            if (unsigned(useAddr) < depth) then
              for i in 0 to (DATA_WIDTH/8)-1 loop 
                if (WSTRB(i) = '1') then
                  if ((8*i) < cwidth) then
                    if (8*(i+1) <= cwidth) then
                      mem(to_integer(unsigned(useAddr))) (8*(i+1)-1 downto (8*i)) <= WDATA(8*(i+1)-1 downto (8*i));
                    else
                      mem(to_integer(unsigned(useAddr))) (cwidth-1 downto (8*i)) <= WDATA(cwidth-1 downto (8*i));
                    end if;
                  end if;
                end if;
              end loop;
              
              --write(buf, string'("Slave AXI1 write:mem[0x"));
              --write(buf,  slv2hex(useAddr));
              --write(buf, string'("]=0x"));
              --write(buf,  slv2hex(WDATA));
              --write(buf, string'(" at T="));
              --write(buf, now);
              --writeline(output, buf);
            else
              -- pragma translate_off
              write(buf, string'("Error:  Out-of-range AXI memory write access:0x"));
              write(buf,  slv2hex(AWADDR));
              write(buf, string'(" at T="));
              write(buf, now);
              writeline(output, buf);
              -- pragma translate_on
            end if;
          end if;
        end if;
        writeAddr <= to_integer(unsigned(useAddr));
        if ((WLAST = '1') and (WVALID = '1')) then
          write_state <= axi4w_write_done;
          WREADY_reg <= '0';
          BRESP_reg <= AXI4_xRESP_OKAY;
          BVALID_reg <= '1';
        else
          write_state <= axi4w_write;
        end if;
      elsif (write_state = axi4w_write) then
        if (WVALID = '1') then
          useAddr2 := std_logic_vector(to_unsigned(writeAddr+1, useAddr2'length));
          if (unsigned(WSTRB) /= 0) then
            if (unsigned(useAddr2) < depth) then
              for i in 0 to (DATA_WIDTH/8)-1 loop 
                if (WSTRB(i) = '1') then
                  if ((8*i) < cwidth) then
                    if (8*(i+1) <= cwidth) then
                      mem(to_integer(unsigned(useAddr2))) (8*(i+1)-1 downto (8*i)) <= WDATA(8*(i+1)-1 downto (8*i));
                    else
                      mem(to_integer(unsigned(useAddr2))) (cwidth-1 downto (8*i)) <= WDATA(cwidth-1 downto (8*i));
                    end if;
                  end if;
                end if;
              end loop;
              --write(buf, string'("Slave AXI2 write:mem[0x"));
              --write(buf,  slv2hex(useAddr2));
              --write(buf, string'("]=0x"));
              --write(buf,  slv2hex(WDATA));
              --write(buf, string'(" at T="));
              --write(buf, now);
              --writeline(output, buf);
            else 
              -- pragma translate_off
              write(buf, string'("Error:  Out-of-range AXI memory write access:0x"));
              write(buf,  slv2hex(AWADDR));
              write(buf, string'(" at T="));
              write(buf, now);
              writeline(output, buf);
              -- pragma translate_on
            end if;
          end if;
          writeAddr <= to_integer(unsigned(useAddr2));
          if (WLAST = '1') then
            write_state <= axi4w_write_done;
            WREADY_reg <= '0';
            BRESP_reg <= AXI4_xRESP_OKAY;
            BVALID_reg <= '1';
          end if;
        end if;
      elsif (write_state = axi4w_write_done) then
        if (BREADY = '1') then
          AWREADY_reg <= '1';
          WREADY_reg <= '1';
          BRESP_reg <= AXI4_xRESP_OKAY;
          BVALID_reg <= '0';
          write_state <= axi4w_idle;
          s_wrdy_reg <= '1';
        end if;
      else
        s_wrdy_reg <= '1';
      end if;
    end if;
  end process; -- axiWrite

  rCatOutOfOrder <= '1' when (s_re = '1') and
                             (s_rrdy_reg = '1') and
                             (catIsReading = '1') and
                             (next_raddr /= to_integer(unsigned(extCatAddr(s_raddr)))+1)
                  else '0';
  
  -- Catapult read processing
  catRead : process(ACLK, int_ARESETn)
    -- pragma translate_off
    variable buf : line;
    -- pragma translate_on
  begin
    if (int_ARESETn = '0') then
      s_din_reg <= (others => '0');
      s_rrdy_reg <= '0';
      catIsReading <= '0';
      next_raddr <= 0;
    elsif rising_edge(ACLK) then
      -- Catapult has read access to memory
      if (tr_write_done = '1') then
        if ( s_re = '1') then
          --$display("Slave CAT read.  Addr=%x Data=%d T=%t", s_raddr, mem[s_raddr], $time);
          --write(buf, string'("Slave CAT read.  Addr=0x"));
          --write(buf,  slv2hex(s_raddr));
          --write(buf, string'(" Data=0x"));
          --write(buf,  slv2hex(mem(to_integer(unsigned(s_raddr)))));
          --write(buf, string'(" T="));
          --write(buf, now);
          --writeline(output, buf);
          if ((catIsReading = '1') and (rCatOutOfOrder /= '1')) then
            -- Make sure next_addr hasnt incremented off the end
            if (next_raddr < depth) then 
              s_din_reg <= mem(next_raddr);
              next_raddr <= next_raddr+1;
            else
              s_rrdy_reg <= '0';
              catIsReading <= '0';
              next_raddr <= 0;                  
            end if;
          else
            s_din_reg <= mem(to_integer(unsigned(s_raddr)));
            s_rrdy_reg <= '1';
            next_raddr <= to_integer(unsigned(extCatAddr(s_raddr)))+1;
            if ((catIsReading = '1') and (rCatOutOfOrder = '1')) then
              catIsReading <= '0';
            else
              catIsReading <= '1';
            end if;
          end if;
        else
          s_rrdy_reg <= '0';
          catIsReading <= '0';
          next_raddr <= 0;
        end if;
      else
        s_rrdy_reg <= '0';
        catIsReading <= '0';
        next_raddr <= 0;
      end if;
    end if;
  end process;    -- catRead 
  
END rtl;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_mul_pipe IS
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_mul_pipe;

LIBRARY IEEE;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_mul_pipe IS
  TYPE reg_array_type is array(natural range<>) of std_logic_vector(width_z-1 DOWNTO 0); 
  SIGNAL xz : std_logic_vector(width_a+width_b DOWNTO 0);

--MF Added pipelined input
    signal a_f     : STD_LOGIC_VECTOR(width_a-1 downto 0); 
    signal b_f     : STD_LOGIC_VECTOR(width_b-1 downto 0);
   type a_array is array (natural range <>) of STD_LOGIC_VECTOR(width_a-1 downto 0);
   type b_array is array (natural range <>) of STD_LOGIC_VECTOR(width_b-1 downto 0);
BEGIN
  n_inreg_gt_0: if n_inreg > 0 generate
    GENPOS_INREG: IF clock_edge = 1 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '1' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;

            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);    
                                                   
          end if;
        end if;
      end process;
    END GENERATE;
  
   GENNEG_INREG: IF clock_edge = 0 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '0' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;            
                                 
            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);
                                                        
          end if;
        end if;
      end process;
    END GENERATE;
  END GENERATE;

  n_inreg_eq_0: if n_inreg = 0 generate
    a_f <= a;
    b_f <= b;
  end generate n_inreg_eq_0;

  xz <= '0'&(unsigned(a_f) * unsigned(b_f)) WHEN signd_a = 0 AND signd_b = 0 ELSE
            (  signed(a_f) * unsigned(b_f)) WHEN signd_a = 1 AND signd_b = 0 ELSE
            (unsigned(a_f) *   signed(b_f)) WHEN signd_a = 0 AND signd_b = 1 ELSE
        '0'&(  signed(a_f) *   signed(b_f));

  GENPOS: IF clock_edge = 1 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '1') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;

  GENNEG: IF clock_edge = 0 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '0') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_bl_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_bl_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_bl_v5 IS

  FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
    CONSTANT len: INTEGER := input1'LENGTH;
    ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
    ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
    VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
  BEGIN
    result := (others => '0');
    --synopsys translate_off
    FOR i IN len-1 DOWNTO 0 LOOP
      result(i) := resolved(input1a(i) & input2a(i));
    END LOOP;
    --synopsys translate_on
    RETURN result;
  END;

  FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED)
  RETURN UNSIGNED IS
  BEGIN
    RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                             STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED)
  RETURN SIGNED IS
  BEGIN
    RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                           STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
    BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

 FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
    --synopsys translate_off
           | 'L'
    --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
    --synopsys translate_off
           | 'H'
    --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_unsigned(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: SIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
      --synopsys translate_off
           | 'L'
      --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
      --synopsys translate_off
           | 'H'
      --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_signed(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), signed(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), signed(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_DPRAM_RBW_DUAL.vhd 
-- Memory Type:            BLOCK
-- Operating Mode:         True Dual Port (2-Port)
-- Clock Mode:             Dual Clock
-- 
-- RTL Code RW Resolution: RBW
-- Catapult RW Resolution: RBW
-- 
-- HDL Work Library:       Xilinx_RAMS_lib
-- Component Name:         BLOCK_DPRAM_RBW_DUAL
-- Latency = 1:            RAM with no registers on inputs or outputs
--         = 2:            adds embedded register on RAM output
--         = 3:            adds fabric registers to non-clock input RAM pins
--         = 4:            adds fabric register to output (driven by embedded register from latency=2)

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
PACKAGE BLOCK_DPRAM_RBW_DUAL_pkg IS
  COMPONENT BLOCK_DPRAM_RBW_DUAL IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    adra : in std_logic_vector(addr_width-1 downto 0) ;
    adrb : in std_logic_vector(addr_width-1 downto 0) ;
    clka : in std_logic ;
    clka_en : in std_logic ;
    clkb : in std_logic ;
    clkb_en : in std_logic ;
    da : in std_logic_vector(data_width-1 downto 0) ;
    db : in std_logic_vector(data_width-1 downto 0) ;
    qa : out std_logic_vector(data_width-1 downto 0) ;
    qb : out std_logic_vector(data_width-1 downto 0) ;
    wea : in std_logic ;
    web : in std_logic 
    
  );
  END COMPONENT;
END BLOCK_DPRAM_RBW_DUAL_pkg;
LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
ENTITY BLOCK_DPRAM_RBW_DUAL IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    adra : in std_logic_vector(addr_width-1 downto 0) ;
    adrb : in std_logic_vector(addr_width-1 downto 0) ;
    clka : in std_logic ;
    clka_en : in std_logic ;
    clkb : in std_logic ;
    clkb_en : in std_logic ;
    da : in std_logic_vector(data_width-1 downto 0) ;
    db : in std_logic_vector(data_width-1 downto 0) ;
    qa : out std_logic_vector(data_width-1 downto 0) ;
    qb : out std_logic_vector(data_width-1 downto 0) ;
    wea : in std_logic ;
    web : in std_logic 
    
  );
 END BLOCK_DPRAM_RBW_DUAL;
ARCHITECTURE rtl OF BLOCK_DPRAM_RBW_DUAL IS
  TYPE ram_t IS ARRAY (depth-1 DOWNTO 0) OF std_logic_vector(data_width-1 DOWNTO 0);
  SHARED VARIABLE mem : ram_t := (OTHERS => (OTHERS => '0'));
  ATTRIBUTE ram_style: STRING;
  ATTRIBUTE ram_style OF mem : VARIABLE IS "block";
  ATTRIBUTE syn_ramstyle: STRING;
  ATTRIBUTE syn_ramstyle OF mem : VARIABLE IS "block";
  
  SIGNAL ramqa : std_logic_vector(data_width-1 downto 0);
  SIGNAL ramqb : std_logic_vector(data_width-1 downto 0);
  
BEGIN
-- Port Map
-- rwA :: ADDRESS adra CLOCK clka ENABLE clka_en DATA_IN da DATA_OUT qa WRITE_ENABLE wea
-- rwB :: ADDRESS adrb CLOCK clkb ENABLE clkb_en DATA_IN db DATA_OUT qb WRITE_ENABLE web

-- Access memory with non-registered inputs (latency = 1||2)
  IN_PIN :  IF latency < 3 GENERATE
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adra)) < depth) THEN
          --pragma translate_on
          ramqa <= mem(to_integer(unsigned(adra)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (wea = '1') THEN
            mem(to_integer(unsigned(adra))) := da;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adrb)) < depth) THEN
          --pragma translate_on
          ramqb <= mem(to_integer(unsigned(adrb)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (web = '1') THEN
            mem(to_integer(unsigned(adrb))) := db;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_PIN; 

-- Register all non-clock inputs (latency = 3||4)
  IN_REG :  IF latency > 2 GENERATE
    SIGNAL adra_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL da_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL wea_reg : std_logic;
    SIGNAL adrb_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL db_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL web_reg : std_logic;
    
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          adra_reg <= adra;
          da_reg <= da;
          wea_reg <= wea;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          adrb_reg <= adrb;
          db_reg <= db;
          web_reg <= web;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adra_reg)) < depth) THEN
          --pragma translate_on
          ramqa <= mem(to_integer(unsigned(adra_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (wea_reg = '1') THEN
            mem(to_integer(unsigned(adra_reg))) := da_reg;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
         IF (clka_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
         IF (clkb_en = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adrb_reg)) < depth) THEN
          --pragma translate_on
          ramqb <= mem(to_integer(unsigned(adrb_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (web_reg = '1') THEN
            mem(to_integer(unsigned(adrb_reg))) := db_reg;
          END IF;
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_REG;

  out_ram : IF latency = 1 GENERATE
  BEGIN
    qa <= ramqa;
    qb <= ramqb;
    
  END GENERATE out_ram;

  out_reg1 : IF ((latency = 2) OR (latency = 3)) GENERATE
    SIGNAL tmpqa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmpqb : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          tmpqa <= ramqa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          tmpqb <= ramqb;
        END IF;
      END IF;
    END PROCESS;
    
    qa <= tmpqa;
    qb <= tmpqb;
    
  END GENERATE out_reg1;

  out_reg2 : IF latency = 4 GENERATE
    SIGNAL tmp1qa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmp1qb : std_logic_vector(data_width-1 downto 0);
    
    SIGNAL tmp2qa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmp2qb : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          tmp1qa <= ramqa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          tmp1qb <= ramqb;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clka)
    BEGIN
      IF (rising_edge(clka)) THEN
        IF (clka_en = '1') THEN
          tmp2qa <= tmp1qa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clkb)
    BEGIN
      IF (rising_edge(clkb)) THEN
        IF (clkb_en = '1') THEN
          tmp2qb <= tmp1qb;
        END IF;
      END IF;
    END PROCESS;
    
    qa <= tmp2qa;
    qb <= tmp2qb;
    
  END GENERATE out_reg2;


END rtl;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   jd4691@newnano.poly.edu
--  Generated date: Tue Sep 14 10:11:16 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_73_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_73_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_73_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_73_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_72_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_72_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_72_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_72_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_71_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_71_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_71_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_71_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_70_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_70_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_70_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_70_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_69_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_69_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_69_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_69_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_68_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_68_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_68_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_68_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_67_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_67_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_67_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_67_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_66_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_66_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_66_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_66_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_65_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_65_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_65_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_65_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_64_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_64_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_64_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_64_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_63_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_63_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_63_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_63_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_62_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_62_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_62_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_62_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_61_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_61_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_61_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_61_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_60_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_60_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_60_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_60_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_59_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_59_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_59_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_59_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_58_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_58_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_58_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_58_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_57_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_57_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_57_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_57_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_56_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_56_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_56_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_56_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_55_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_55_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_55_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_55_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_54_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_54_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_54_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_54_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_53_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_53_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_53_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_53_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_52_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_52_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_52_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_52_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_47_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_47_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_47_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_47_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_46_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_46_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_46_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_46_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_45_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_45_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_45_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_45_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_44_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_44_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_44_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_44_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_43_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_43_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_43_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_43_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_42_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_42_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_42_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_42_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_41_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_41_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_41_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_41_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_40_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_40_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_40_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_40_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_39_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_39_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_39_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_39_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_5_32_32_32_32_1_gen IS
  PORT(
    clkb_en : OUT STD_LOGIC;
    clka_en : OUT STD_LOGIC;
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    web : OUT STD_LOGIC;
    db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    clka : IN STD_LOGIC;
    clka_en_d : IN STD_LOGIC;
    clkb_en_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
  );
END hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  clkb_en <= clkb_en_d;
  clka_en <= clka_en_d;
  qa_d(63 DOWNTO 32) <= qb;
  web <= (rwA_rw_ram_ir_internal_WMASK_B_d(1));
  db <= (da_d(63 DOWNTO 32));
  adrb <= (adra_d(9 DOWNTO 5));
  qa_d(31 DOWNTO 0) <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d(0));
  da <= (da_d(31 DOWNTO 0));
  adra <= (adra_d(4 DOWNTO 0));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_4_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_4_5_32_32_32_32_1_gen IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_4_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_4_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_3_5_32_32_32_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_3_5_32_32_32_32_1_gen IS
  PORT(
    qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    adrb_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_3_5_32_32_32_32_1_gen;

ARCHITECTURE v14 OF hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_3_5_32_32_32_32_1_gen
    IS
  -- Default Constants

BEGIN
  qb_d <= qb;
  adrb <= (adrb_d);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
    S1_OUTER_LOOP_for_C_5_tr0 : IN STD_LOGIC;
    S1_OUTER_LOOP_C_0_tr0 : IN STD_LOGIC;
    S2_COPY_LOOP_for_C_4_tr0 : IN STD_LOGIC;
    S2_COPY_LOOP_C_0_tr0 : IN STD_LOGIC;
    S2_INNER_LOOP1_for_C_20_tr0 : IN STD_LOGIC;
    S2_INNER_LOOP1_C_2_tr0 : IN STD_LOGIC;
    S2_INNER_LOOP2_for_C_20_tr0 : IN STD_LOGIC;
    S2_INNER_LOOP2_C_2_tr0 : IN STD_LOGIC;
    S2_INNER_LOOP2_C_2_tr1 : IN STD_LOGIC;
    S2_INNER_LOOP3_for_C_20_tr0 : IN STD_LOGIC;
    S2_INNER_LOOP3_C_2_tr0 : IN STD_LOGIC;
    S34_OUTER_LOOP_for_C_12_tr0 : IN STD_LOGIC;
    S34_OUTER_LOOP_C_0_tr0 : IN STD_LOGIC;
    S5_COPY_LOOP_for_C_4_tr0 : IN STD_LOGIC;
    S5_COPY_LOOP_C_0_tr0 : IN STD_LOGIC;
    S5_INNER_LOOP1_for_C_20_tr0 : IN STD_LOGIC;
    S5_INNER_LOOP1_C_2_tr0 : IN STD_LOGIC;
    S5_INNER_LOOP2_for_C_20_tr0 : IN STD_LOGIC;
    S5_INNER_LOOP2_C_2_tr0 : IN STD_LOGIC;
    S5_INNER_LOOP2_C_2_tr1 : IN STD_LOGIC;
    S5_INNER_LOOP3_for_C_20_tr0 : IN STD_LOGIC;
    S5_INNER_LOOP3_C_2_tr0 : IN STD_LOGIC;
    S6_OUTER_LOOP_for_C_4_tr0 : IN STD_LOGIC;
    S6_OUTER_LOOP_C_0_tr0 : IN STD_LOGIC
  );
END hybrid_core_core_fsm;

ARCHITECTURE v14 OF hybrid_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for hybrid_core_core_fsm_1
  TYPE hybrid_core_core_fsm_1_ST IS (main_C_0, S1_OUTER_LOOP_for_C_0, S1_OUTER_LOOP_for_C_1,
      S1_OUTER_LOOP_for_C_2, S1_OUTER_LOOP_for_C_3, S1_OUTER_LOOP_for_C_4, S1_OUTER_LOOP_for_C_5,
      S1_OUTER_LOOP_C_0, S2_COPY_LOOP_for_C_0, S2_COPY_LOOP_for_C_1, S2_COPY_LOOP_for_C_2,
      S2_COPY_LOOP_for_C_3, S2_COPY_LOOP_for_C_4, S2_COPY_LOOP_C_0, S2_OUTER_LOOP_C_0,
      S2_INNER_LOOP1_C_0, S2_INNER_LOOP1_C_1, S2_INNER_LOOP1_for_C_0, S2_INNER_LOOP1_for_C_1,
      S2_INNER_LOOP1_for_C_2, S2_INNER_LOOP1_for_C_3, S2_INNER_LOOP1_for_C_4, S2_INNER_LOOP1_for_C_5,
      S2_INNER_LOOP1_for_C_6, S2_INNER_LOOP1_for_C_7, S2_INNER_LOOP1_for_C_8, S2_INNER_LOOP1_for_C_9,
      S2_INNER_LOOP1_for_C_10, S2_INNER_LOOP1_for_C_11, S2_INNER_LOOP1_for_C_12,
      S2_INNER_LOOP1_for_C_13, S2_INNER_LOOP1_for_C_14, S2_INNER_LOOP1_for_C_15,
      S2_INNER_LOOP1_for_C_16, S2_INNER_LOOP1_for_C_17, S2_INNER_LOOP1_for_C_18,
      S2_INNER_LOOP1_for_C_19, S2_INNER_LOOP1_for_C_20, S2_INNER_LOOP1_C_2, S2_OUTER_LOOP_C_1,
      S2_INNER_LOOP2_C_0, S2_INNER_LOOP2_C_1, S2_INNER_LOOP2_for_C_0, S2_INNER_LOOP2_for_C_1,
      S2_INNER_LOOP2_for_C_2, S2_INNER_LOOP2_for_C_3, S2_INNER_LOOP2_for_C_4, S2_INNER_LOOP2_for_C_5,
      S2_INNER_LOOP2_for_C_6, S2_INNER_LOOP2_for_C_7, S2_INNER_LOOP2_for_C_8, S2_INNER_LOOP2_for_C_9,
      S2_INNER_LOOP2_for_C_10, S2_INNER_LOOP2_for_C_11, S2_INNER_LOOP2_for_C_12,
      S2_INNER_LOOP2_for_C_13, S2_INNER_LOOP2_for_C_14, S2_INNER_LOOP2_for_C_15,
      S2_INNER_LOOP2_for_C_16, S2_INNER_LOOP2_for_C_17, S2_INNER_LOOP2_for_C_18,
      S2_INNER_LOOP2_for_C_19, S2_INNER_LOOP2_for_C_20, S2_INNER_LOOP2_C_2, S2_INNER_LOOP3_C_0,
      S2_INNER_LOOP3_C_1, S2_INNER_LOOP3_for_C_0, S2_INNER_LOOP3_for_C_1, S2_INNER_LOOP3_for_C_2,
      S2_INNER_LOOP3_for_C_3, S2_INNER_LOOP3_for_C_4, S2_INNER_LOOP3_for_C_5, S2_INNER_LOOP3_for_C_6,
      S2_INNER_LOOP3_for_C_7, S2_INNER_LOOP3_for_C_8, S2_INNER_LOOP3_for_C_9, S2_INNER_LOOP3_for_C_10,
      S2_INNER_LOOP3_for_C_11, S2_INNER_LOOP3_for_C_12, S2_INNER_LOOP3_for_C_13,
      S2_INNER_LOOP3_for_C_14, S2_INNER_LOOP3_for_C_15, S2_INNER_LOOP3_for_C_16,
      S2_INNER_LOOP3_for_C_17, S2_INNER_LOOP3_for_C_18, S2_INNER_LOOP3_for_C_19,
      S2_INNER_LOOP3_for_C_20, S2_INNER_LOOP3_C_2, S34_OUTER_LOOP_for_C_0, S34_OUTER_LOOP_for_C_1,
      S34_OUTER_LOOP_for_C_2, S34_OUTER_LOOP_for_C_3, S34_OUTER_LOOP_for_C_4, S34_OUTER_LOOP_for_C_5,
      S34_OUTER_LOOP_for_C_6, S34_OUTER_LOOP_for_C_7, S34_OUTER_LOOP_for_C_8, S34_OUTER_LOOP_for_C_9,
      S34_OUTER_LOOP_for_C_10, S34_OUTER_LOOP_for_C_11, S34_OUTER_LOOP_for_C_12,
      S34_OUTER_LOOP_C_0, S5_COPY_LOOP_for_C_0, S5_COPY_LOOP_for_C_1, S5_COPY_LOOP_for_C_2,
      S5_COPY_LOOP_for_C_3, S5_COPY_LOOP_for_C_4, S5_COPY_LOOP_C_0, S5_OUTER_LOOP_C_0,
      S5_INNER_LOOP1_C_0, S5_INNER_LOOP1_C_1, S5_INNER_LOOP1_for_C_0, S5_INNER_LOOP1_for_C_1,
      S5_INNER_LOOP1_for_C_2, S5_INNER_LOOP1_for_C_3, S5_INNER_LOOP1_for_C_4, S5_INNER_LOOP1_for_C_5,
      S5_INNER_LOOP1_for_C_6, S5_INNER_LOOP1_for_C_7, S5_INNER_LOOP1_for_C_8, S5_INNER_LOOP1_for_C_9,
      S5_INNER_LOOP1_for_C_10, S5_INNER_LOOP1_for_C_11, S5_INNER_LOOP1_for_C_12,
      S5_INNER_LOOP1_for_C_13, S5_INNER_LOOP1_for_C_14, S5_INNER_LOOP1_for_C_15,
      S5_INNER_LOOP1_for_C_16, S5_INNER_LOOP1_for_C_17, S5_INNER_LOOP1_for_C_18,
      S5_INNER_LOOP1_for_C_19, S5_INNER_LOOP1_for_C_20, S5_INNER_LOOP1_C_2, S5_OUTER_LOOP_C_1,
      S5_INNER_LOOP2_C_0, S5_INNER_LOOP2_C_1, S5_INNER_LOOP2_for_C_0, S5_INNER_LOOP2_for_C_1,
      S5_INNER_LOOP2_for_C_2, S5_INNER_LOOP2_for_C_3, S5_INNER_LOOP2_for_C_4, S5_INNER_LOOP2_for_C_5,
      S5_INNER_LOOP2_for_C_6, S5_INNER_LOOP2_for_C_7, S5_INNER_LOOP2_for_C_8, S5_INNER_LOOP2_for_C_9,
      S5_INNER_LOOP2_for_C_10, S5_INNER_LOOP2_for_C_11, S5_INNER_LOOP2_for_C_12,
      S5_INNER_LOOP2_for_C_13, S5_INNER_LOOP2_for_C_14, S5_INNER_LOOP2_for_C_15,
      S5_INNER_LOOP2_for_C_16, S5_INNER_LOOP2_for_C_17, S5_INNER_LOOP2_for_C_18,
      S5_INNER_LOOP2_for_C_19, S5_INNER_LOOP2_for_C_20, S5_INNER_LOOP2_C_2, S5_INNER_LOOP3_C_0,
      S5_INNER_LOOP3_C_1, S5_INNER_LOOP3_for_C_0, S5_INNER_LOOP3_for_C_1, S5_INNER_LOOP3_for_C_2,
      S5_INNER_LOOP3_for_C_3, S5_INNER_LOOP3_for_C_4, S5_INNER_LOOP3_for_C_5, S5_INNER_LOOP3_for_C_6,
      S5_INNER_LOOP3_for_C_7, S5_INNER_LOOP3_for_C_8, S5_INNER_LOOP3_for_C_9, S5_INNER_LOOP3_for_C_10,
      S5_INNER_LOOP3_for_C_11, S5_INNER_LOOP3_for_C_12, S5_INNER_LOOP3_for_C_13,
      S5_INNER_LOOP3_for_C_14, S5_INNER_LOOP3_for_C_15, S5_INNER_LOOP3_for_C_16,
      S5_INNER_LOOP3_for_C_17, S5_INNER_LOOP3_for_C_18, S5_INNER_LOOP3_for_C_19,
      S5_INNER_LOOP3_for_C_20, S5_INNER_LOOP3_C_2, S6_OUTER_LOOP_for_C_0, S6_OUTER_LOOP_for_C_1,
      S6_OUTER_LOOP_for_C_2, S6_OUTER_LOOP_for_C_3, S6_OUTER_LOOP_for_C_4, S6_OUTER_LOOP_C_0,
      main_C_1);

  SIGNAL state_var : hybrid_core_core_fsm_1_ST;
  SIGNAL state_var_NS : hybrid_core_core_fsm_1_ST;

BEGIN
  hybrid_core_core_fsm_1 : PROCESS (S1_OUTER_LOOP_for_C_5_tr0, S1_OUTER_LOOP_C_0_tr0,
      S2_COPY_LOOP_for_C_4_tr0, S2_COPY_LOOP_C_0_tr0, S2_INNER_LOOP1_for_C_20_tr0,
      S2_INNER_LOOP1_C_2_tr0, S2_INNER_LOOP2_for_C_20_tr0, S2_INNER_LOOP2_C_2_tr0,
      S2_INNER_LOOP2_C_2_tr1, S2_INNER_LOOP3_for_C_20_tr0, S2_INNER_LOOP3_C_2_tr0,
      S34_OUTER_LOOP_for_C_12_tr0, S34_OUTER_LOOP_C_0_tr0, S5_COPY_LOOP_for_C_4_tr0,
      S5_COPY_LOOP_C_0_tr0, S5_INNER_LOOP1_for_C_20_tr0, S5_INNER_LOOP1_C_2_tr0,
      S5_INNER_LOOP2_for_C_20_tr0, S5_INNER_LOOP2_C_2_tr0, S5_INNER_LOOP2_C_2_tr1,
      S5_INNER_LOOP3_for_C_20_tr0, S5_INNER_LOOP3_C_2_tr0, S6_OUTER_LOOP_for_C_4_tr0,
      S6_OUTER_LOOP_C_0_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN S1_OUTER_LOOP_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000001");
        state_var_NS <= S1_OUTER_LOOP_for_C_1;
      WHEN S1_OUTER_LOOP_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000010");
        state_var_NS <= S1_OUTER_LOOP_for_C_2;
      WHEN S1_OUTER_LOOP_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000011");
        state_var_NS <= S1_OUTER_LOOP_for_C_3;
      WHEN S1_OUTER_LOOP_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000100");
        state_var_NS <= S1_OUTER_LOOP_for_C_4;
      WHEN S1_OUTER_LOOP_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000101");
        state_var_NS <= S1_OUTER_LOOP_for_C_5;
      WHEN S1_OUTER_LOOP_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000110");
        IF ( S1_OUTER_LOOP_for_C_5_tr0 = '1' ) THEN
          state_var_NS <= S1_OUTER_LOOP_C_0;
        ELSE
          state_var_NS <= S1_OUTER_LOOP_for_C_0;
        END IF;
      WHEN S1_OUTER_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000111");
        IF ( S1_OUTER_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= S2_COPY_LOOP_for_C_0;
        ELSE
          state_var_NS <= S1_OUTER_LOOP_for_C_0;
        END IF;
      WHEN S2_COPY_LOOP_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001000");
        state_var_NS <= S2_COPY_LOOP_for_C_1;
      WHEN S2_COPY_LOOP_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001001");
        state_var_NS <= S2_COPY_LOOP_for_C_2;
      WHEN S2_COPY_LOOP_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001010");
        state_var_NS <= S2_COPY_LOOP_for_C_3;
      WHEN S2_COPY_LOOP_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001011");
        state_var_NS <= S2_COPY_LOOP_for_C_4;
      WHEN S2_COPY_LOOP_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001100");
        IF ( S2_COPY_LOOP_for_C_4_tr0 = '1' ) THEN
          state_var_NS <= S2_COPY_LOOP_C_0;
        ELSE
          state_var_NS <= S2_COPY_LOOP_for_C_0;
        END IF;
      WHEN S2_COPY_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001101");
        IF ( S2_COPY_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= S2_OUTER_LOOP_C_0;
        ELSE
          state_var_NS <= S2_COPY_LOOP_for_C_0;
        END IF;
      WHEN S2_OUTER_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001110");
        state_var_NS <= S2_INNER_LOOP1_C_0;
      WHEN S2_INNER_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00001111");
        state_var_NS <= S2_INNER_LOOP1_C_1;
      WHEN S2_INNER_LOOP1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010000");
        state_var_NS <= S2_INNER_LOOP1_for_C_0;
      WHEN S2_INNER_LOOP1_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010001");
        state_var_NS <= S2_INNER_LOOP1_for_C_1;
      WHEN S2_INNER_LOOP1_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010010");
        state_var_NS <= S2_INNER_LOOP1_for_C_2;
      WHEN S2_INNER_LOOP1_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010011");
        state_var_NS <= S2_INNER_LOOP1_for_C_3;
      WHEN S2_INNER_LOOP1_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010100");
        state_var_NS <= S2_INNER_LOOP1_for_C_4;
      WHEN S2_INNER_LOOP1_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010101");
        state_var_NS <= S2_INNER_LOOP1_for_C_5;
      WHEN S2_INNER_LOOP1_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010110");
        state_var_NS <= S2_INNER_LOOP1_for_C_6;
      WHEN S2_INNER_LOOP1_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00010111");
        state_var_NS <= S2_INNER_LOOP1_for_C_7;
      WHEN S2_INNER_LOOP1_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011000");
        state_var_NS <= S2_INNER_LOOP1_for_C_8;
      WHEN S2_INNER_LOOP1_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011001");
        state_var_NS <= S2_INNER_LOOP1_for_C_9;
      WHEN S2_INNER_LOOP1_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011010");
        state_var_NS <= S2_INNER_LOOP1_for_C_10;
      WHEN S2_INNER_LOOP1_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011011");
        state_var_NS <= S2_INNER_LOOP1_for_C_11;
      WHEN S2_INNER_LOOP1_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011100");
        state_var_NS <= S2_INNER_LOOP1_for_C_12;
      WHEN S2_INNER_LOOP1_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011101");
        state_var_NS <= S2_INNER_LOOP1_for_C_13;
      WHEN S2_INNER_LOOP1_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011110");
        state_var_NS <= S2_INNER_LOOP1_for_C_14;
      WHEN S2_INNER_LOOP1_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00011111");
        state_var_NS <= S2_INNER_LOOP1_for_C_15;
      WHEN S2_INNER_LOOP1_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100000");
        state_var_NS <= S2_INNER_LOOP1_for_C_16;
      WHEN S2_INNER_LOOP1_for_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100001");
        state_var_NS <= S2_INNER_LOOP1_for_C_17;
      WHEN S2_INNER_LOOP1_for_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100010");
        state_var_NS <= S2_INNER_LOOP1_for_C_18;
      WHEN S2_INNER_LOOP1_for_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100011");
        state_var_NS <= S2_INNER_LOOP1_for_C_19;
      WHEN S2_INNER_LOOP1_for_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100100");
        state_var_NS <= S2_INNER_LOOP1_for_C_20;
      WHEN S2_INNER_LOOP1_for_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100101");
        IF ( S2_INNER_LOOP1_for_C_20_tr0 = '1' ) THEN
          state_var_NS <= S2_INNER_LOOP1_C_2;
        ELSE
          state_var_NS <= S2_INNER_LOOP1_for_C_0;
        END IF;
      WHEN S2_INNER_LOOP1_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100110");
        IF ( S2_INNER_LOOP1_C_2_tr0 = '1' ) THEN
          state_var_NS <= S2_OUTER_LOOP_C_1;
        ELSE
          state_var_NS <= S2_INNER_LOOP1_C_0;
        END IF;
      WHEN S2_OUTER_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00100111");
        state_var_NS <= S2_INNER_LOOP2_C_0;
      WHEN S2_INNER_LOOP2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101000");
        state_var_NS <= S2_INNER_LOOP2_C_1;
      WHEN S2_INNER_LOOP2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101001");
        state_var_NS <= S2_INNER_LOOP2_for_C_0;
      WHEN S2_INNER_LOOP2_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101010");
        state_var_NS <= S2_INNER_LOOP2_for_C_1;
      WHEN S2_INNER_LOOP2_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101011");
        state_var_NS <= S2_INNER_LOOP2_for_C_2;
      WHEN S2_INNER_LOOP2_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101100");
        state_var_NS <= S2_INNER_LOOP2_for_C_3;
      WHEN S2_INNER_LOOP2_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101101");
        state_var_NS <= S2_INNER_LOOP2_for_C_4;
      WHEN S2_INNER_LOOP2_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101110");
        state_var_NS <= S2_INNER_LOOP2_for_C_5;
      WHEN S2_INNER_LOOP2_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00101111");
        state_var_NS <= S2_INNER_LOOP2_for_C_6;
      WHEN S2_INNER_LOOP2_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110000");
        state_var_NS <= S2_INNER_LOOP2_for_C_7;
      WHEN S2_INNER_LOOP2_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110001");
        state_var_NS <= S2_INNER_LOOP2_for_C_8;
      WHEN S2_INNER_LOOP2_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110010");
        state_var_NS <= S2_INNER_LOOP2_for_C_9;
      WHEN S2_INNER_LOOP2_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110011");
        state_var_NS <= S2_INNER_LOOP2_for_C_10;
      WHEN S2_INNER_LOOP2_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110100");
        state_var_NS <= S2_INNER_LOOP2_for_C_11;
      WHEN S2_INNER_LOOP2_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110101");
        state_var_NS <= S2_INNER_LOOP2_for_C_12;
      WHEN S2_INNER_LOOP2_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110110");
        state_var_NS <= S2_INNER_LOOP2_for_C_13;
      WHEN S2_INNER_LOOP2_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00110111");
        state_var_NS <= S2_INNER_LOOP2_for_C_14;
      WHEN S2_INNER_LOOP2_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111000");
        state_var_NS <= S2_INNER_LOOP2_for_C_15;
      WHEN S2_INNER_LOOP2_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111001");
        state_var_NS <= S2_INNER_LOOP2_for_C_16;
      WHEN S2_INNER_LOOP2_for_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111010");
        state_var_NS <= S2_INNER_LOOP2_for_C_17;
      WHEN S2_INNER_LOOP2_for_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111011");
        state_var_NS <= S2_INNER_LOOP2_for_C_18;
      WHEN S2_INNER_LOOP2_for_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111100");
        state_var_NS <= S2_INNER_LOOP2_for_C_19;
      WHEN S2_INNER_LOOP2_for_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111101");
        state_var_NS <= S2_INNER_LOOP2_for_C_20;
      WHEN S2_INNER_LOOP2_for_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111110");
        IF ( S2_INNER_LOOP2_for_C_20_tr0 = '1' ) THEN
          state_var_NS <= S2_INNER_LOOP2_C_2;
        ELSE
          state_var_NS <= S2_INNER_LOOP2_for_C_0;
        END IF;
      WHEN S2_INNER_LOOP2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "00111111");
        IF ( S2_INNER_LOOP2_C_2_tr0 = '1' ) THEN
          state_var_NS <= S2_INNER_LOOP3_C_0;
        ELSIF ( S2_INNER_LOOP2_C_2_tr1 = '1' ) THEN
          state_var_NS <= S2_INNER_LOOP2_C_0;
        ELSE
          state_var_NS <= S2_OUTER_LOOP_C_0;
        END IF;
      WHEN S2_INNER_LOOP3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000000");
        state_var_NS <= S2_INNER_LOOP3_C_1;
      WHEN S2_INNER_LOOP3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000001");
        state_var_NS <= S2_INNER_LOOP3_for_C_0;
      WHEN S2_INNER_LOOP3_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000010");
        state_var_NS <= S2_INNER_LOOP3_for_C_1;
      WHEN S2_INNER_LOOP3_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000011");
        state_var_NS <= S2_INNER_LOOP3_for_C_2;
      WHEN S2_INNER_LOOP3_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000100");
        state_var_NS <= S2_INNER_LOOP3_for_C_3;
      WHEN S2_INNER_LOOP3_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000101");
        state_var_NS <= S2_INNER_LOOP3_for_C_4;
      WHEN S2_INNER_LOOP3_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000110");
        state_var_NS <= S2_INNER_LOOP3_for_C_5;
      WHEN S2_INNER_LOOP3_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01000111");
        state_var_NS <= S2_INNER_LOOP3_for_C_6;
      WHEN S2_INNER_LOOP3_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001000");
        state_var_NS <= S2_INNER_LOOP3_for_C_7;
      WHEN S2_INNER_LOOP3_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001001");
        state_var_NS <= S2_INNER_LOOP3_for_C_8;
      WHEN S2_INNER_LOOP3_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001010");
        state_var_NS <= S2_INNER_LOOP3_for_C_9;
      WHEN S2_INNER_LOOP3_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001011");
        state_var_NS <= S2_INNER_LOOP3_for_C_10;
      WHEN S2_INNER_LOOP3_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001100");
        state_var_NS <= S2_INNER_LOOP3_for_C_11;
      WHEN S2_INNER_LOOP3_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001101");
        state_var_NS <= S2_INNER_LOOP3_for_C_12;
      WHEN S2_INNER_LOOP3_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001110");
        state_var_NS <= S2_INNER_LOOP3_for_C_13;
      WHEN S2_INNER_LOOP3_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01001111");
        state_var_NS <= S2_INNER_LOOP3_for_C_14;
      WHEN S2_INNER_LOOP3_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010000");
        state_var_NS <= S2_INNER_LOOP3_for_C_15;
      WHEN S2_INNER_LOOP3_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010001");
        state_var_NS <= S2_INNER_LOOP3_for_C_16;
      WHEN S2_INNER_LOOP3_for_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010010");
        state_var_NS <= S2_INNER_LOOP3_for_C_17;
      WHEN S2_INNER_LOOP3_for_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010011");
        state_var_NS <= S2_INNER_LOOP3_for_C_18;
      WHEN S2_INNER_LOOP3_for_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010100");
        state_var_NS <= S2_INNER_LOOP3_for_C_19;
      WHEN S2_INNER_LOOP3_for_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010101");
        state_var_NS <= S2_INNER_LOOP3_for_C_20;
      WHEN S2_INNER_LOOP3_for_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010110");
        IF ( S2_INNER_LOOP3_for_C_20_tr0 = '1' ) THEN
          state_var_NS <= S2_INNER_LOOP3_C_2;
        ELSE
          state_var_NS <= S2_INNER_LOOP3_for_C_0;
        END IF;
      WHEN S2_INNER_LOOP3_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01010111");
        IF ( S2_INNER_LOOP3_C_2_tr0 = '1' ) THEN
          state_var_NS <= S34_OUTER_LOOP_for_C_0;
        ELSE
          state_var_NS <= S2_INNER_LOOP3_C_0;
        END IF;
      WHEN S34_OUTER_LOOP_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011000");
        state_var_NS <= S34_OUTER_LOOP_for_C_1;
      WHEN S34_OUTER_LOOP_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011001");
        state_var_NS <= S34_OUTER_LOOP_for_C_2;
      WHEN S34_OUTER_LOOP_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011010");
        state_var_NS <= S34_OUTER_LOOP_for_C_3;
      WHEN S34_OUTER_LOOP_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011011");
        state_var_NS <= S34_OUTER_LOOP_for_C_4;
      WHEN S34_OUTER_LOOP_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011100");
        state_var_NS <= S34_OUTER_LOOP_for_C_5;
      WHEN S34_OUTER_LOOP_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011101");
        state_var_NS <= S34_OUTER_LOOP_for_C_6;
      WHEN S34_OUTER_LOOP_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011110");
        state_var_NS <= S34_OUTER_LOOP_for_C_7;
      WHEN S34_OUTER_LOOP_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01011111");
        state_var_NS <= S34_OUTER_LOOP_for_C_8;
      WHEN S34_OUTER_LOOP_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100000");
        state_var_NS <= S34_OUTER_LOOP_for_C_9;
      WHEN S34_OUTER_LOOP_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100001");
        state_var_NS <= S34_OUTER_LOOP_for_C_10;
      WHEN S34_OUTER_LOOP_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100010");
        state_var_NS <= S34_OUTER_LOOP_for_C_11;
      WHEN S34_OUTER_LOOP_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100011");
        state_var_NS <= S34_OUTER_LOOP_for_C_12;
      WHEN S34_OUTER_LOOP_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100100");
        IF ( S34_OUTER_LOOP_for_C_12_tr0 = '1' ) THEN
          state_var_NS <= S34_OUTER_LOOP_C_0;
        ELSE
          state_var_NS <= S34_OUTER_LOOP_for_C_0;
        END IF;
      WHEN S34_OUTER_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100101");
        IF ( S34_OUTER_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= S5_COPY_LOOP_for_C_0;
        ELSE
          state_var_NS <= S34_OUTER_LOOP_for_C_0;
        END IF;
      WHEN S5_COPY_LOOP_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100110");
        state_var_NS <= S5_COPY_LOOP_for_C_1;
      WHEN S5_COPY_LOOP_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01100111");
        state_var_NS <= S5_COPY_LOOP_for_C_2;
      WHEN S5_COPY_LOOP_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101000");
        state_var_NS <= S5_COPY_LOOP_for_C_3;
      WHEN S5_COPY_LOOP_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101001");
        state_var_NS <= S5_COPY_LOOP_for_C_4;
      WHEN S5_COPY_LOOP_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101010");
        IF ( S5_COPY_LOOP_for_C_4_tr0 = '1' ) THEN
          state_var_NS <= S5_COPY_LOOP_C_0;
        ELSE
          state_var_NS <= S5_COPY_LOOP_for_C_0;
        END IF;
      WHEN S5_COPY_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101011");
        IF ( S5_COPY_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= S5_OUTER_LOOP_C_0;
        ELSE
          state_var_NS <= S5_COPY_LOOP_for_C_0;
        END IF;
      WHEN S5_OUTER_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101100");
        state_var_NS <= S5_INNER_LOOP1_C_0;
      WHEN S5_INNER_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101101");
        state_var_NS <= S5_INNER_LOOP1_C_1;
      WHEN S5_INNER_LOOP1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101110");
        state_var_NS <= S5_INNER_LOOP1_for_C_0;
      WHEN S5_INNER_LOOP1_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01101111");
        state_var_NS <= S5_INNER_LOOP1_for_C_1;
      WHEN S5_INNER_LOOP1_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110000");
        state_var_NS <= S5_INNER_LOOP1_for_C_2;
      WHEN S5_INNER_LOOP1_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110001");
        state_var_NS <= S5_INNER_LOOP1_for_C_3;
      WHEN S5_INNER_LOOP1_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110010");
        state_var_NS <= S5_INNER_LOOP1_for_C_4;
      WHEN S5_INNER_LOOP1_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110011");
        state_var_NS <= S5_INNER_LOOP1_for_C_5;
      WHEN S5_INNER_LOOP1_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110100");
        state_var_NS <= S5_INNER_LOOP1_for_C_6;
      WHEN S5_INNER_LOOP1_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110101");
        state_var_NS <= S5_INNER_LOOP1_for_C_7;
      WHEN S5_INNER_LOOP1_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110110");
        state_var_NS <= S5_INNER_LOOP1_for_C_8;
      WHEN S5_INNER_LOOP1_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01110111");
        state_var_NS <= S5_INNER_LOOP1_for_C_9;
      WHEN S5_INNER_LOOP1_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111000");
        state_var_NS <= S5_INNER_LOOP1_for_C_10;
      WHEN S5_INNER_LOOP1_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111001");
        state_var_NS <= S5_INNER_LOOP1_for_C_11;
      WHEN S5_INNER_LOOP1_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111010");
        state_var_NS <= S5_INNER_LOOP1_for_C_12;
      WHEN S5_INNER_LOOP1_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111011");
        state_var_NS <= S5_INNER_LOOP1_for_C_13;
      WHEN S5_INNER_LOOP1_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111100");
        state_var_NS <= S5_INNER_LOOP1_for_C_14;
      WHEN S5_INNER_LOOP1_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111101");
        state_var_NS <= S5_INNER_LOOP1_for_C_15;
      WHEN S5_INNER_LOOP1_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111110");
        state_var_NS <= S5_INNER_LOOP1_for_C_16;
      WHEN S5_INNER_LOOP1_for_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "01111111");
        state_var_NS <= S5_INNER_LOOP1_for_C_17;
      WHEN S5_INNER_LOOP1_for_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000000");
        state_var_NS <= S5_INNER_LOOP1_for_C_18;
      WHEN S5_INNER_LOOP1_for_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000001");
        state_var_NS <= S5_INNER_LOOP1_for_C_19;
      WHEN S5_INNER_LOOP1_for_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000010");
        state_var_NS <= S5_INNER_LOOP1_for_C_20;
      WHEN S5_INNER_LOOP1_for_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000011");
        IF ( S5_INNER_LOOP1_for_C_20_tr0 = '1' ) THEN
          state_var_NS <= S5_INNER_LOOP1_C_2;
        ELSE
          state_var_NS <= S5_INNER_LOOP1_for_C_0;
        END IF;
      WHEN S5_INNER_LOOP1_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000100");
        IF ( S5_INNER_LOOP1_C_2_tr0 = '1' ) THEN
          state_var_NS <= S5_OUTER_LOOP_C_1;
        ELSE
          state_var_NS <= S5_INNER_LOOP1_C_0;
        END IF;
      WHEN S5_OUTER_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000101");
        state_var_NS <= S5_INNER_LOOP2_C_0;
      WHEN S5_INNER_LOOP2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000110");
        state_var_NS <= S5_INNER_LOOP2_C_1;
      WHEN S5_INNER_LOOP2_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10000111");
        state_var_NS <= S5_INNER_LOOP2_for_C_0;
      WHEN S5_INNER_LOOP2_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001000");
        state_var_NS <= S5_INNER_LOOP2_for_C_1;
      WHEN S5_INNER_LOOP2_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001001");
        state_var_NS <= S5_INNER_LOOP2_for_C_2;
      WHEN S5_INNER_LOOP2_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001010");
        state_var_NS <= S5_INNER_LOOP2_for_C_3;
      WHEN S5_INNER_LOOP2_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001011");
        state_var_NS <= S5_INNER_LOOP2_for_C_4;
      WHEN S5_INNER_LOOP2_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001100");
        state_var_NS <= S5_INNER_LOOP2_for_C_5;
      WHEN S5_INNER_LOOP2_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001101");
        state_var_NS <= S5_INNER_LOOP2_for_C_6;
      WHEN S5_INNER_LOOP2_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001110");
        state_var_NS <= S5_INNER_LOOP2_for_C_7;
      WHEN S5_INNER_LOOP2_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10001111");
        state_var_NS <= S5_INNER_LOOP2_for_C_8;
      WHEN S5_INNER_LOOP2_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010000");
        state_var_NS <= S5_INNER_LOOP2_for_C_9;
      WHEN S5_INNER_LOOP2_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010001");
        state_var_NS <= S5_INNER_LOOP2_for_C_10;
      WHEN S5_INNER_LOOP2_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010010");
        state_var_NS <= S5_INNER_LOOP2_for_C_11;
      WHEN S5_INNER_LOOP2_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010011");
        state_var_NS <= S5_INNER_LOOP2_for_C_12;
      WHEN S5_INNER_LOOP2_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010100");
        state_var_NS <= S5_INNER_LOOP2_for_C_13;
      WHEN S5_INNER_LOOP2_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010101");
        state_var_NS <= S5_INNER_LOOP2_for_C_14;
      WHEN S5_INNER_LOOP2_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010110");
        state_var_NS <= S5_INNER_LOOP2_for_C_15;
      WHEN S5_INNER_LOOP2_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10010111");
        state_var_NS <= S5_INNER_LOOP2_for_C_16;
      WHEN S5_INNER_LOOP2_for_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011000");
        state_var_NS <= S5_INNER_LOOP2_for_C_17;
      WHEN S5_INNER_LOOP2_for_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011001");
        state_var_NS <= S5_INNER_LOOP2_for_C_18;
      WHEN S5_INNER_LOOP2_for_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011010");
        state_var_NS <= S5_INNER_LOOP2_for_C_19;
      WHEN S5_INNER_LOOP2_for_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011011");
        state_var_NS <= S5_INNER_LOOP2_for_C_20;
      WHEN S5_INNER_LOOP2_for_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011100");
        IF ( S5_INNER_LOOP2_for_C_20_tr0 = '1' ) THEN
          state_var_NS <= S5_INNER_LOOP2_C_2;
        ELSE
          state_var_NS <= S5_INNER_LOOP2_for_C_0;
        END IF;
      WHEN S5_INNER_LOOP2_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011101");
        IF ( S5_INNER_LOOP2_C_2_tr0 = '1' ) THEN
          state_var_NS <= S5_INNER_LOOP3_C_0;
        ELSIF ( S5_INNER_LOOP2_C_2_tr1 = '1' ) THEN
          state_var_NS <= S5_INNER_LOOP2_C_0;
        ELSE
          state_var_NS <= S5_OUTER_LOOP_C_0;
        END IF;
      WHEN S5_INNER_LOOP3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011110");
        state_var_NS <= S5_INNER_LOOP3_C_1;
      WHEN S5_INNER_LOOP3_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10011111");
        state_var_NS <= S5_INNER_LOOP3_for_C_0;
      WHEN S5_INNER_LOOP3_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100000");
        state_var_NS <= S5_INNER_LOOP3_for_C_1;
      WHEN S5_INNER_LOOP3_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100001");
        state_var_NS <= S5_INNER_LOOP3_for_C_2;
      WHEN S5_INNER_LOOP3_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100010");
        state_var_NS <= S5_INNER_LOOP3_for_C_3;
      WHEN S5_INNER_LOOP3_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100011");
        state_var_NS <= S5_INNER_LOOP3_for_C_4;
      WHEN S5_INNER_LOOP3_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100100");
        state_var_NS <= S5_INNER_LOOP3_for_C_5;
      WHEN S5_INNER_LOOP3_for_C_5 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100101");
        state_var_NS <= S5_INNER_LOOP3_for_C_6;
      WHEN S5_INNER_LOOP3_for_C_6 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100110");
        state_var_NS <= S5_INNER_LOOP3_for_C_7;
      WHEN S5_INNER_LOOP3_for_C_7 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10100111");
        state_var_NS <= S5_INNER_LOOP3_for_C_8;
      WHEN S5_INNER_LOOP3_for_C_8 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101000");
        state_var_NS <= S5_INNER_LOOP3_for_C_9;
      WHEN S5_INNER_LOOP3_for_C_9 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101001");
        state_var_NS <= S5_INNER_LOOP3_for_C_10;
      WHEN S5_INNER_LOOP3_for_C_10 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101010");
        state_var_NS <= S5_INNER_LOOP3_for_C_11;
      WHEN S5_INNER_LOOP3_for_C_11 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101011");
        state_var_NS <= S5_INNER_LOOP3_for_C_12;
      WHEN S5_INNER_LOOP3_for_C_12 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101100");
        state_var_NS <= S5_INNER_LOOP3_for_C_13;
      WHEN S5_INNER_LOOP3_for_C_13 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101101");
        state_var_NS <= S5_INNER_LOOP3_for_C_14;
      WHEN S5_INNER_LOOP3_for_C_14 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101110");
        state_var_NS <= S5_INNER_LOOP3_for_C_15;
      WHEN S5_INNER_LOOP3_for_C_15 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10101111");
        state_var_NS <= S5_INNER_LOOP3_for_C_16;
      WHEN S5_INNER_LOOP3_for_C_16 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110000");
        state_var_NS <= S5_INNER_LOOP3_for_C_17;
      WHEN S5_INNER_LOOP3_for_C_17 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110001");
        state_var_NS <= S5_INNER_LOOP3_for_C_18;
      WHEN S5_INNER_LOOP3_for_C_18 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110010");
        state_var_NS <= S5_INNER_LOOP3_for_C_19;
      WHEN S5_INNER_LOOP3_for_C_19 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110011");
        state_var_NS <= S5_INNER_LOOP3_for_C_20;
      WHEN S5_INNER_LOOP3_for_C_20 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110100");
        IF ( S5_INNER_LOOP3_for_C_20_tr0 = '1' ) THEN
          state_var_NS <= S5_INNER_LOOP3_C_2;
        ELSE
          state_var_NS <= S5_INNER_LOOP3_for_C_0;
        END IF;
      WHEN S5_INNER_LOOP3_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110101");
        IF ( S5_INNER_LOOP3_C_2_tr0 = '1' ) THEN
          state_var_NS <= S6_OUTER_LOOP_for_C_0;
        ELSE
          state_var_NS <= S5_INNER_LOOP3_C_0;
        END IF;
      WHEN S6_OUTER_LOOP_for_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110110");
        state_var_NS <= S6_OUTER_LOOP_for_C_1;
      WHEN S6_OUTER_LOOP_for_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10110111");
        state_var_NS <= S6_OUTER_LOOP_for_C_2;
      WHEN S6_OUTER_LOOP_for_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111000");
        state_var_NS <= S6_OUTER_LOOP_for_C_3;
      WHEN S6_OUTER_LOOP_for_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111001");
        state_var_NS <= S6_OUTER_LOOP_for_C_4;
      WHEN S6_OUTER_LOOP_for_C_4 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111010");
        IF ( S6_OUTER_LOOP_for_C_4_tr0 = '1' ) THEN
          state_var_NS <= S6_OUTER_LOOP_C_0;
        ELSE
          state_var_NS <= S6_OUTER_LOOP_for_C_0;
        END IF;
      WHEN S6_OUTER_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111011");
        IF ( S6_OUTER_LOOP_C_0_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSE
          state_var_NS <= S6_OUTER_LOOP_for_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "10111100");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "00000000");
        state_var_NS <= S1_OUTER_LOOP_for_C_0;
    END CASE;
  END PROCESS hybrid_core_core_fsm_1;

  hybrid_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        IF ( core_wen = '1' ) THEN
          state_var <= state_var_NS;
        END IF;
      END IF;
    END IF;
  END PROCESS hybrid_core_core_fsm_1_REG;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_staller
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_staller IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    core_wen : OUT STD_LOGIC;
    core_wten : OUT STD_LOGIC;
    revArr_rsci_wen_comp : IN STD_LOGIC;
    tw_rsci_wen_comp : IN STD_LOGIC;
    tw_h_rsci_wen_comp : IN STD_LOGIC;
    x_rsc_0_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_0_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_1_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_1_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_2_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_2_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_3_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_3_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_4_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_4_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_5_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_5_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_6_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_6_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_7_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_7_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_8_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_8_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_9_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_9_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_10_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_10_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_11_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_11_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_12_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_12_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_13_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_13_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_14_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_14_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_15_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_15_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_16_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_16_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_17_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_17_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_18_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_18_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_19_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_19_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_20_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_20_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_21_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_21_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_22_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_22_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_23_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_23_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_24_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_24_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_25_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_25_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_26_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_26_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_27_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_27_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_28_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_28_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_29_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_29_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_30_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_30_0_i_wen_comp_1 : IN STD_LOGIC;
    x_rsc_31_0_i_wen_comp : IN STD_LOGIC;
    x_rsc_31_0_i_wen_comp_1 : IN STD_LOGIC
  );
END hybrid_core_staller;

ARCHITECTURE v14 OF hybrid_core_staller IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL core_wen_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL core_wten_reg : STD_LOGIC;

BEGIN
  -- Output Reader Assignments
  core_wen <= core_wen_drv;

  core_wen_drv <= revArr_rsci_wen_comp AND tw_rsci_wen_comp AND tw_h_rsci_wen_comp
      AND x_rsc_0_0_i_wen_comp AND x_rsc_0_0_i_wen_comp_1 AND x_rsc_1_0_i_wen_comp
      AND x_rsc_1_0_i_wen_comp_1 AND x_rsc_2_0_i_wen_comp AND x_rsc_2_0_i_wen_comp_1
      AND x_rsc_3_0_i_wen_comp AND x_rsc_3_0_i_wen_comp_1 AND x_rsc_4_0_i_wen_comp
      AND x_rsc_4_0_i_wen_comp_1 AND x_rsc_5_0_i_wen_comp AND x_rsc_5_0_i_wen_comp_1
      AND x_rsc_6_0_i_wen_comp AND x_rsc_6_0_i_wen_comp_1 AND x_rsc_7_0_i_wen_comp
      AND x_rsc_7_0_i_wen_comp_1 AND x_rsc_8_0_i_wen_comp AND x_rsc_8_0_i_wen_comp_1
      AND x_rsc_9_0_i_wen_comp AND x_rsc_9_0_i_wen_comp_1 AND x_rsc_10_0_i_wen_comp
      AND x_rsc_10_0_i_wen_comp_1 AND x_rsc_11_0_i_wen_comp AND x_rsc_11_0_i_wen_comp_1
      AND x_rsc_12_0_i_wen_comp AND x_rsc_12_0_i_wen_comp_1 AND x_rsc_13_0_i_wen_comp
      AND x_rsc_13_0_i_wen_comp_1 AND x_rsc_14_0_i_wen_comp AND x_rsc_14_0_i_wen_comp_1
      AND x_rsc_15_0_i_wen_comp AND x_rsc_15_0_i_wen_comp_1 AND x_rsc_16_0_i_wen_comp
      AND x_rsc_16_0_i_wen_comp_1 AND x_rsc_17_0_i_wen_comp AND x_rsc_17_0_i_wen_comp_1
      AND x_rsc_18_0_i_wen_comp AND x_rsc_18_0_i_wen_comp_1 AND x_rsc_19_0_i_wen_comp
      AND x_rsc_19_0_i_wen_comp_1 AND x_rsc_20_0_i_wen_comp AND x_rsc_20_0_i_wen_comp_1
      AND x_rsc_21_0_i_wen_comp AND x_rsc_21_0_i_wen_comp_1 AND x_rsc_22_0_i_wen_comp
      AND x_rsc_22_0_i_wen_comp_1 AND x_rsc_23_0_i_wen_comp AND x_rsc_23_0_i_wen_comp_1
      AND x_rsc_24_0_i_wen_comp AND x_rsc_24_0_i_wen_comp_1 AND x_rsc_25_0_i_wen_comp
      AND x_rsc_25_0_i_wen_comp_1 AND x_rsc_26_0_i_wen_comp AND x_rsc_26_0_i_wen_comp_1
      AND x_rsc_27_0_i_wen_comp AND x_rsc_27_0_i_wen_comp_1 AND x_rsc_28_0_i_wen_comp
      AND x_rsc_28_0_i_wen_comp_1 AND x_rsc_29_0_i_wen_comp AND x_rsc_29_0_i_wen_comp_1
      AND x_rsc_30_0_i_wen_comp AND x_rsc_30_0_i_wen_comp_1 AND x_rsc_31_0_i_wen_comp
      AND x_rsc_31_0_i_wen_comp_1;
  core_wten <= core_wten_reg;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        core_wten_reg <= '0';
      ELSE
        core_wten_reg <= NOT core_wen_drv;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    tw_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    tw_h_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl IS
  -- Default Constants

BEGIN
  tw_h_rsc_triosy_obj_ld_core_sct <= tw_h_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    tw_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    tw_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl IS
  -- Default Constants

BEGIN
  tw_rsc_triosy_obj_ld_core_sct <= tw_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    revArr_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    revArr_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl
    IS
  -- Default Constants

BEGIN
  revArr_rsc_triosy_obj_ld_core_sct <= revArr_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_obj_ld_core_sct <= twiddle_h_rsc_triosy_obj_iswt0 AND (NOT
      core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_obj_ld_core_sct <= twiddle_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    m_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    m_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl IS
  -- Default Constants

BEGIN
  m_rsc_triosy_obj_ld_core_sct <= m_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_0_0_obj_ld_core_sct <= x_rsc_triosy_0_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_1_0_obj_ld_core_sct <= x_rsc_triosy_1_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_2_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_2_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_2_0_obj_ld_core_sct <= x_rsc_triosy_2_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_3_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_3_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_3_0_obj_ld_core_sct <= x_rsc_triosy_3_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_4_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_4_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_4_0_obj_ld_core_sct <= x_rsc_triosy_4_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_5_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_5_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_5_0_obj_ld_core_sct <= x_rsc_triosy_5_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_6_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_6_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_6_0_obj_ld_core_sct <= x_rsc_triosy_6_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_7_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_7_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_7_0_obj_ld_core_sct <= x_rsc_triosy_7_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_8_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_8_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_8_0_obj_ld_core_sct <= x_rsc_triosy_8_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_9_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_9_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl IS
  -- Default Constants

BEGIN
  x_rsc_triosy_9_0_obj_ld_core_sct <= x_rsc_triosy_9_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_10_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_10_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_10_0_obj_ld_core_sct <= x_rsc_triosy_10_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_11_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_11_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_11_0_obj_ld_core_sct <= x_rsc_triosy_11_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_12_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_12_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_12_0_obj_ld_core_sct <= x_rsc_triosy_12_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_13_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_13_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_13_0_obj_ld_core_sct <= x_rsc_triosy_13_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_14_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_14_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_14_0_obj_ld_core_sct <= x_rsc_triosy_14_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_15_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_15_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_15_0_obj_ld_core_sct <= x_rsc_triosy_15_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_16_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_16_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_16_0_obj_ld_core_sct <= x_rsc_triosy_16_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_17_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_17_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_17_0_obj_ld_core_sct <= x_rsc_triosy_17_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_18_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_18_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_18_0_obj_ld_core_sct <= x_rsc_triosy_18_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_19_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_19_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_19_0_obj_ld_core_sct <= x_rsc_triosy_19_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_20_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_20_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_20_0_obj_ld_core_sct <= x_rsc_triosy_20_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_21_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_21_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_21_0_obj_ld_core_sct <= x_rsc_triosy_21_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_22_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_22_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_22_0_obj_ld_core_sct <= x_rsc_triosy_22_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_23_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_23_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_23_0_obj_ld_core_sct <= x_rsc_triosy_23_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_24_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_24_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_24_0_obj_ld_core_sct <= x_rsc_triosy_24_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_25_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_25_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_25_0_obj_ld_core_sct <= x_rsc_triosy_25_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_26_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_26_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_26_0_obj_ld_core_sct <= x_rsc_triosy_26_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_27_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_27_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_27_0_obj_ld_core_sct <= x_rsc_triosy_27_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_28_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_28_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_28_0_obj_ld_core_sct <= x_rsc_triosy_28_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_29_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_29_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_29_0_obj_ld_core_sct <= x_rsc_triosy_29_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_30_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_30_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_30_0_obj_ld_core_sct <= x_rsc_triosy_30_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_31_0_obj_iswt0 : IN STD_LOGIC;
    x_rsc_triosy_31_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  x_rsc_triosy_31_0_obj_ld_core_sct <= x_rsc_triosy_31_0_obj_iswt0 AND (NOT core_wten);
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_31_0_i_oswt : IN STD_LOGIC;
    x_rsc_31_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_31_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_31_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_31_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_31_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_31_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_i_biwt : IN STD_LOGIC;
    x_rsc_31_0_i_bdwt : IN STD_LOGIC;
    x_rsc_31_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_31_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_31_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_31_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_31_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_31_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_31_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_31_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_31_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_31_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_31_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_31_0_i_bcwt <= x_rsc_31_0_i_bcwt_drv;
  x_rsc_31_0_i_bcwt_1 <= x_rsc_31_0_i_bcwt_1_drv;

  x_rsc_31_0_i_wen_comp <= (NOT x_rsc_31_0_i_oswt) OR x_rsc_31_0_i_biwt OR x_rsc_31_0_i_bcwt_drv;
  x_rsc_31_0_i_wen_comp_1 <= (NOT x_rsc_31_0_i_oswt_1) OR x_rsc_31_0_i_biwt_1 OR
      x_rsc_31_0_i_bcwt_1_drv;
  x_rsc_31_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_31_0_i_s_raddr_core,
      x_rsc_31_0_i_s_raddr_core_sct);
  x_rsc_31_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_31_0_i_s_waddr_core,
      x_rsc_31_0_i_s_waddr_core_sct);
  x_rsc_31_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_31_0_i_s_din, x_rsc_31_0_i_s_din_bfwt,
      x_rsc_31_0_i_bcwt_drv);
  x_rsc_31_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_31_0_i_s_dout_core, x_rsc_31_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_31_0_i_bcwt_drv <= '0';
        x_rsc_31_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_31_0_i_bcwt_drv <= NOT((NOT(x_rsc_31_0_i_bcwt_drv OR x_rsc_31_0_i_biwt))
            OR x_rsc_31_0_i_bdwt);
        x_rsc_31_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_31_0_i_bcwt_1_drv OR x_rsc_31_0_i_biwt_1))
            OR x_rsc_31_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_31_0_i_biwt = '1' ) THEN
        x_rsc_31_0_i_s_din_bfwt <= x_rsc_31_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_31_0_i_oswt : IN STD_LOGIC;
    x_rsc_31_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_31_0_i_biwt : OUT STD_LOGIC;
    x_rsc_31_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_31_0_i_bcwt : IN STD_LOGIC;
    x_rsc_31_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_31_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_31_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_31_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_31_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_31_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_31_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_31_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_31_0_i_bdwt <= x_rsc_31_0_i_oswt AND core_wen;
  x_rsc_31_0_i_biwt <= x_rsc_31_0_i_ogwt AND x_rsc_31_0_i_s_rrdy;
  x_rsc_31_0_i_ogwt <= x_rsc_31_0_i_oswt AND (NOT x_rsc_31_0_i_bcwt);
  x_rsc_31_0_i_s_re_core_sct <= x_rsc_31_0_i_ogwt;
  x_rsc_31_0_i_bdwt_2 <= x_rsc_31_0_i_oswt_1 AND core_wen;
  x_rsc_31_0_i_biwt_1 <= x_rsc_31_0_i_ogwt_1 AND x_rsc_31_0_i_s_wrdy;
  x_rsc_31_0_i_ogwt_1 <= x_rsc_31_0_i_oswt_1 AND (NOT x_rsc_31_0_i_bcwt_1);
  x_rsc_31_0_i_s_we_core_sct <= x_rsc_31_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_30_0_i_oswt : IN STD_LOGIC;
    x_rsc_30_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_30_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_30_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_30_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_30_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_30_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_i_biwt : IN STD_LOGIC;
    x_rsc_30_0_i_bdwt : IN STD_LOGIC;
    x_rsc_30_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_30_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_30_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_30_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_30_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_30_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_30_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_30_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_30_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_30_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_30_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_30_0_i_bcwt <= x_rsc_30_0_i_bcwt_drv;
  x_rsc_30_0_i_bcwt_1 <= x_rsc_30_0_i_bcwt_1_drv;

  x_rsc_30_0_i_wen_comp <= (NOT x_rsc_30_0_i_oswt) OR x_rsc_30_0_i_biwt OR x_rsc_30_0_i_bcwt_drv;
  x_rsc_30_0_i_wen_comp_1 <= (NOT x_rsc_30_0_i_oswt_1) OR x_rsc_30_0_i_biwt_1 OR
      x_rsc_30_0_i_bcwt_1_drv;
  x_rsc_30_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_30_0_i_s_raddr_core,
      x_rsc_30_0_i_s_raddr_core_sct);
  x_rsc_30_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_30_0_i_s_waddr_core,
      x_rsc_30_0_i_s_waddr_core_sct);
  x_rsc_30_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_30_0_i_s_din, x_rsc_30_0_i_s_din_bfwt,
      x_rsc_30_0_i_bcwt_drv);
  x_rsc_30_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_30_0_i_s_dout_core, x_rsc_30_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_30_0_i_bcwt_drv <= '0';
        x_rsc_30_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_30_0_i_bcwt_drv <= NOT((NOT(x_rsc_30_0_i_bcwt_drv OR x_rsc_30_0_i_biwt))
            OR x_rsc_30_0_i_bdwt);
        x_rsc_30_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_30_0_i_bcwt_1_drv OR x_rsc_30_0_i_biwt_1))
            OR x_rsc_30_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_30_0_i_biwt = '1' ) THEN
        x_rsc_30_0_i_s_din_bfwt <= x_rsc_30_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_30_0_i_oswt : IN STD_LOGIC;
    x_rsc_30_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_30_0_i_biwt : OUT STD_LOGIC;
    x_rsc_30_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_30_0_i_bcwt : IN STD_LOGIC;
    x_rsc_30_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_30_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_30_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_30_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_30_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_30_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_30_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_30_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_30_0_i_bdwt <= x_rsc_30_0_i_oswt AND core_wen;
  x_rsc_30_0_i_biwt <= x_rsc_30_0_i_ogwt AND x_rsc_30_0_i_s_rrdy;
  x_rsc_30_0_i_ogwt <= x_rsc_30_0_i_oswt AND (NOT x_rsc_30_0_i_bcwt);
  x_rsc_30_0_i_s_re_core_sct <= x_rsc_30_0_i_ogwt;
  x_rsc_30_0_i_bdwt_2 <= x_rsc_30_0_i_oswt_1 AND core_wen;
  x_rsc_30_0_i_biwt_1 <= x_rsc_30_0_i_ogwt_1 AND x_rsc_30_0_i_s_wrdy;
  x_rsc_30_0_i_ogwt_1 <= x_rsc_30_0_i_oswt_1 AND (NOT x_rsc_30_0_i_bcwt_1);
  x_rsc_30_0_i_s_we_core_sct <= x_rsc_30_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_29_0_i_oswt : IN STD_LOGIC;
    x_rsc_29_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_29_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_29_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_29_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_29_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_29_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_i_biwt : IN STD_LOGIC;
    x_rsc_29_0_i_bdwt : IN STD_LOGIC;
    x_rsc_29_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_29_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_29_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_29_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_29_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_29_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_29_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_29_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_29_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_29_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_29_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_29_0_i_bcwt <= x_rsc_29_0_i_bcwt_drv;
  x_rsc_29_0_i_bcwt_1 <= x_rsc_29_0_i_bcwt_1_drv;

  x_rsc_29_0_i_wen_comp <= (NOT x_rsc_29_0_i_oswt) OR x_rsc_29_0_i_biwt OR x_rsc_29_0_i_bcwt_drv;
  x_rsc_29_0_i_wen_comp_1 <= (NOT x_rsc_29_0_i_oswt_1) OR x_rsc_29_0_i_biwt_1 OR
      x_rsc_29_0_i_bcwt_1_drv;
  x_rsc_29_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_29_0_i_s_raddr_core,
      x_rsc_29_0_i_s_raddr_core_sct);
  x_rsc_29_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_29_0_i_s_waddr_core,
      x_rsc_29_0_i_s_waddr_core_sct);
  x_rsc_29_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_29_0_i_s_din, x_rsc_29_0_i_s_din_bfwt,
      x_rsc_29_0_i_bcwt_drv);
  x_rsc_29_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_29_0_i_s_dout_core, x_rsc_29_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_29_0_i_bcwt_drv <= '0';
        x_rsc_29_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_29_0_i_bcwt_drv <= NOT((NOT(x_rsc_29_0_i_bcwt_drv OR x_rsc_29_0_i_biwt))
            OR x_rsc_29_0_i_bdwt);
        x_rsc_29_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_29_0_i_bcwt_1_drv OR x_rsc_29_0_i_biwt_1))
            OR x_rsc_29_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_29_0_i_biwt = '1' ) THEN
        x_rsc_29_0_i_s_din_bfwt <= x_rsc_29_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_29_0_i_oswt : IN STD_LOGIC;
    x_rsc_29_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_29_0_i_biwt : OUT STD_LOGIC;
    x_rsc_29_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_29_0_i_bcwt : IN STD_LOGIC;
    x_rsc_29_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_29_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_29_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_29_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_29_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_29_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_29_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_29_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_29_0_i_bdwt <= x_rsc_29_0_i_oswt AND core_wen;
  x_rsc_29_0_i_biwt <= x_rsc_29_0_i_ogwt AND x_rsc_29_0_i_s_rrdy;
  x_rsc_29_0_i_ogwt <= x_rsc_29_0_i_oswt AND (NOT x_rsc_29_0_i_bcwt);
  x_rsc_29_0_i_s_re_core_sct <= x_rsc_29_0_i_ogwt;
  x_rsc_29_0_i_bdwt_2 <= x_rsc_29_0_i_oswt_1 AND core_wen;
  x_rsc_29_0_i_biwt_1 <= x_rsc_29_0_i_ogwt_1 AND x_rsc_29_0_i_s_wrdy;
  x_rsc_29_0_i_ogwt_1 <= x_rsc_29_0_i_oswt_1 AND (NOT x_rsc_29_0_i_bcwt_1);
  x_rsc_29_0_i_s_we_core_sct <= x_rsc_29_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_28_0_i_oswt : IN STD_LOGIC;
    x_rsc_28_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_28_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_28_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_28_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_28_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_28_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_i_biwt : IN STD_LOGIC;
    x_rsc_28_0_i_bdwt : IN STD_LOGIC;
    x_rsc_28_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_28_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_28_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_28_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_28_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_28_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_28_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_28_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_28_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_28_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_28_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_28_0_i_bcwt <= x_rsc_28_0_i_bcwt_drv;
  x_rsc_28_0_i_bcwt_1 <= x_rsc_28_0_i_bcwt_1_drv;

  x_rsc_28_0_i_wen_comp <= (NOT x_rsc_28_0_i_oswt) OR x_rsc_28_0_i_biwt OR x_rsc_28_0_i_bcwt_drv;
  x_rsc_28_0_i_wen_comp_1 <= (NOT x_rsc_28_0_i_oswt_1) OR x_rsc_28_0_i_biwt_1 OR
      x_rsc_28_0_i_bcwt_1_drv;
  x_rsc_28_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_28_0_i_s_raddr_core,
      x_rsc_28_0_i_s_raddr_core_sct);
  x_rsc_28_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_28_0_i_s_waddr_core,
      x_rsc_28_0_i_s_waddr_core_sct);
  x_rsc_28_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_28_0_i_s_din, x_rsc_28_0_i_s_din_bfwt,
      x_rsc_28_0_i_bcwt_drv);
  x_rsc_28_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_28_0_i_s_dout_core, x_rsc_28_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_28_0_i_bcwt_drv <= '0';
        x_rsc_28_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_28_0_i_bcwt_drv <= NOT((NOT(x_rsc_28_0_i_bcwt_drv OR x_rsc_28_0_i_biwt))
            OR x_rsc_28_0_i_bdwt);
        x_rsc_28_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_28_0_i_bcwt_1_drv OR x_rsc_28_0_i_biwt_1))
            OR x_rsc_28_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_28_0_i_biwt = '1' ) THEN
        x_rsc_28_0_i_s_din_bfwt <= x_rsc_28_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_28_0_i_oswt : IN STD_LOGIC;
    x_rsc_28_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_28_0_i_biwt : OUT STD_LOGIC;
    x_rsc_28_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_28_0_i_bcwt : IN STD_LOGIC;
    x_rsc_28_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_28_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_28_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_28_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_28_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_28_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_28_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_28_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_28_0_i_bdwt <= x_rsc_28_0_i_oswt AND core_wen;
  x_rsc_28_0_i_biwt <= x_rsc_28_0_i_ogwt AND x_rsc_28_0_i_s_rrdy;
  x_rsc_28_0_i_ogwt <= x_rsc_28_0_i_oswt AND (NOT x_rsc_28_0_i_bcwt);
  x_rsc_28_0_i_s_re_core_sct <= x_rsc_28_0_i_ogwt;
  x_rsc_28_0_i_bdwt_2 <= x_rsc_28_0_i_oswt_1 AND core_wen;
  x_rsc_28_0_i_biwt_1 <= x_rsc_28_0_i_ogwt_1 AND x_rsc_28_0_i_s_wrdy;
  x_rsc_28_0_i_ogwt_1 <= x_rsc_28_0_i_oswt_1 AND (NOT x_rsc_28_0_i_bcwt_1);
  x_rsc_28_0_i_s_we_core_sct <= x_rsc_28_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_27_0_i_oswt : IN STD_LOGIC;
    x_rsc_27_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_27_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_27_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_27_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_27_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_27_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_i_biwt : IN STD_LOGIC;
    x_rsc_27_0_i_bdwt : IN STD_LOGIC;
    x_rsc_27_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_27_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_27_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_27_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_27_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_27_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_27_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_27_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_27_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_27_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_27_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_27_0_i_bcwt <= x_rsc_27_0_i_bcwt_drv;
  x_rsc_27_0_i_bcwt_1 <= x_rsc_27_0_i_bcwt_1_drv;

  x_rsc_27_0_i_wen_comp <= (NOT x_rsc_27_0_i_oswt) OR x_rsc_27_0_i_biwt OR x_rsc_27_0_i_bcwt_drv;
  x_rsc_27_0_i_wen_comp_1 <= (NOT x_rsc_27_0_i_oswt_1) OR x_rsc_27_0_i_biwt_1 OR
      x_rsc_27_0_i_bcwt_1_drv;
  x_rsc_27_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_27_0_i_s_raddr_core,
      x_rsc_27_0_i_s_raddr_core_sct);
  x_rsc_27_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_27_0_i_s_waddr_core,
      x_rsc_27_0_i_s_waddr_core_sct);
  x_rsc_27_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_27_0_i_s_din, x_rsc_27_0_i_s_din_bfwt,
      x_rsc_27_0_i_bcwt_drv);
  x_rsc_27_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_27_0_i_s_dout_core, x_rsc_27_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_27_0_i_bcwt_drv <= '0';
        x_rsc_27_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_27_0_i_bcwt_drv <= NOT((NOT(x_rsc_27_0_i_bcwt_drv OR x_rsc_27_0_i_biwt))
            OR x_rsc_27_0_i_bdwt);
        x_rsc_27_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_27_0_i_bcwt_1_drv OR x_rsc_27_0_i_biwt_1))
            OR x_rsc_27_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_27_0_i_biwt = '1' ) THEN
        x_rsc_27_0_i_s_din_bfwt <= x_rsc_27_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_27_0_i_oswt : IN STD_LOGIC;
    x_rsc_27_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_27_0_i_biwt : OUT STD_LOGIC;
    x_rsc_27_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_27_0_i_bcwt : IN STD_LOGIC;
    x_rsc_27_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_27_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_27_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_27_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_27_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_27_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_27_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_27_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_27_0_i_bdwt <= x_rsc_27_0_i_oswt AND core_wen;
  x_rsc_27_0_i_biwt <= x_rsc_27_0_i_ogwt AND x_rsc_27_0_i_s_rrdy;
  x_rsc_27_0_i_ogwt <= x_rsc_27_0_i_oswt AND (NOT x_rsc_27_0_i_bcwt);
  x_rsc_27_0_i_s_re_core_sct <= x_rsc_27_0_i_ogwt;
  x_rsc_27_0_i_bdwt_2 <= x_rsc_27_0_i_oswt_1 AND core_wen;
  x_rsc_27_0_i_biwt_1 <= x_rsc_27_0_i_ogwt_1 AND x_rsc_27_0_i_s_wrdy;
  x_rsc_27_0_i_ogwt_1 <= x_rsc_27_0_i_oswt_1 AND (NOT x_rsc_27_0_i_bcwt_1);
  x_rsc_27_0_i_s_we_core_sct <= x_rsc_27_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_26_0_i_oswt : IN STD_LOGIC;
    x_rsc_26_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_26_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_26_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_26_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_26_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_26_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_i_biwt : IN STD_LOGIC;
    x_rsc_26_0_i_bdwt : IN STD_LOGIC;
    x_rsc_26_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_26_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_26_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_26_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_26_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_26_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_26_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_26_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_26_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_26_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_26_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_26_0_i_bcwt <= x_rsc_26_0_i_bcwt_drv;
  x_rsc_26_0_i_bcwt_1 <= x_rsc_26_0_i_bcwt_1_drv;

  x_rsc_26_0_i_wen_comp <= (NOT x_rsc_26_0_i_oswt) OR x_rsc_26_0_i_biwt OR x_rsc_26_0_i_bcwt_drv;
  x_rsc_26_0_i_wen_comp_1 <= (NOT x_rsc_26_0_i_oswt_1) OR x_rsc_26_0_i_biwt_1 OR
      x_rsc_26_0_i_bcwt_1_drv;
  x_rsc_26_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_26_0_i_s_raddr_core,
      x_rsc_26_0_i_s_raddr_core_sct);
  x_rsc_26_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_26_0_i_s_waddr_core,
      x_rsc_26_0_i_s_waddr_core_sct);
  x_rsc_26_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_26_0_i_s_din, x_rsc_26_0_i_s_din_bfwt,
      x_rsc_26_0_i_bcwt_drv);
  x_rsc_26_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_26_0_i_s_dout_core, x_rsc_26_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_26_0_i_bcwt_drv <= '0';
        x_rsc_26_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_26_0_i_bcwt_drv <= NOT((NOT(x_rsc_26_0_i_bcwt_drv OR x_rsc_26_0_i_biwt))
            OR x_rsc_26_0_i_bdwt);
        x_rsc_26_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_26_0_i_bcwt_1_drv OR x_rsc_26_0_i_biwt_1))
            OR x_rsc_26_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_26_0_i_biwt = '1' ) THEN
        x_rsc_26_0_i_s_din_bfwt <= x_rsc_26_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_26_0_i_oswt : IN STD_LOGIC;
    x_rsc_26_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_26_0_i_biwt : OUT STD_LOGIC;
    x_rsc_26_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_26_0_i_bcwt : IN STD_LOGIC;
    x_rsc_26_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_26_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_26_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_26_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_26_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_26_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_26_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_26_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_26_0_i_bdwt <= x_rsc_26_0_i_oswt AND core_wen;
  x_rsc_26_0_i_biwt <= x_rsc_26_0_i_ogwt AND x_rsc_26_0_i_s_rrdy;
  x_rsc_26_0_i_ogwt <= x_rsc_26_0_i_oswt AND (NOT x_rsc_26_0_i_bcwt);
  x_rsc_26_0_i_s_re_core_sct <= x_rsc_26_0_i_ogwt;
  x_rsc_26_0_i_bdwt_2 <= x_rsc_26_0_i_oswt_1 AND core_wen;
  x_rsc_26_0_i_biwt_1 <= x_rsc_26_0_i_ogwt_1 AND x_rsc_26_0_i_s_wrdy;
  x_rsc_26_0_i_ogwt_1 <= x_rsc_26_0_i_oswt_1 AND (NOT x_rsc_26_0_i_bcwt_1);
  x_rsc_26_0_i_s_we_core_sct <= x_rsc_26_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_25_0_i_oswt : IN STD_LOGIC;
    x_rsc_25_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_25_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_25_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_25_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_25_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_25_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_i_biwt : IN STD_LOGIC;
    x_rsc_25_0_i_bdwt : IN STD_LOGIC;
    x_rsc_25_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_25_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_25_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_25_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_25_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_25_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_25_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_25_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_25_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_25_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_25_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_25_0_i_bcwt <= x_rsc_25_0_i_bcwt_drv;
  x_rsc_25_0_i_bcwt_1 <= x_rsc_25_0_i_bcwt_1_drv;

  x_rsc_25_0_i_wen_comp <= (NOT x_rsc_25_0_i_oswt) OR x_rsc_25_0_i_biwt OR x_rsc_25_0_i_bcwt_drv;
  x_rsc_25_0_i_wen_comp_1 <= (NOT x_rsc_25_0_i_oswt_1) OR x_rsc_25_0_i_biwt_1 OR
      x_rsc_25_0_i_bcwt_1_drv;
  x_rsc_25_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_25_0_i_s_raddr_core,
      x_rsc_25_0_i_s_raddr_core_sct);
  x_rsc_25_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_25_0_i_s_waddr_core,
      x_rsc_25_0_i_s_waddr_core_sct);
  x_rsc_25_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_25_0_i_s_din, x_rsc_25_0_i_s_din_bfwt,
      x_rsc_25_0_i_bcwt_drv);
  x_rsc_25_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_25_0_i_s_dout_core, x_rsc_25_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_25_0_i_bcwt_drv <= '0';
        x_rsc_25_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_25_0_i_bcwt_drv <= NOT((NOT(x_rsc_25_0_i_bcwt_drv OR x_rsc_25_0_i_biwt))
            OR x_rsc_25_0_i_bdwt);
        x_rsc_25_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_25_0_i_bcwt_1_drv OR x_rsc_25_0_i_biwt_1))
            OR x_rsc_25_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_25_0_i_biwt = '1' ) THEN
        x_rsc_25_0_i_s_din_bfwt <= x_rsc_25_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_25_0_i_oswt : IN STD_LOGIC;
    x_rsc_25_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_25_0_i_biwt : OUT STD_LOGIC;
    x_rsc_25_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_25_0_i_bcwt : IN STD_LOGIC;
    x_rsc_25_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_25_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_25_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_25_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_25_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_25_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_25_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_25_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_25_0_i_bdwt <= x_rsc_25_0_i_oswt AND core_wen;
  x_rsc_25_0_i_biwt <= x_rsc_25_0_i_ogwt AND x_rsc_25_0_i_s_rrdy;
  x_rsc_25_0_i_ogwt <= x_rsc_25_0_i_oswt AND (NOT x_rsc_25_0_i_bcwt);
  x_rsc_25_0_i_s_re_core_sct <= x_rsc_25_0_i_ogwt;
  x_rsc_25_0_i_bdwt_2 <= x_rsc_25_0_i_oswt_1 AND core_wen;
  x_rsc_25_0_i_biwt_1 <= x_rsc_25_0_i_ogwt_1 AND x_rsc_25_0_i_s_wrdy;
  x_rsc_25_0_i_ogwt_1 <= x_rsc_25_0_i_oswt_1 AND (NOT x_rsc_25_0_i_bcwt_1);
  x_rsc_25_0_i_s_we_core_sct <= x_rsc_25_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_24_0_i_oswt : IN STD_LOGIC;
    x_rsc_24_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_24_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_24_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_24_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_24_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_24_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_i_biwt : IN STD_LOGIC;
    x_rsc_24_0_i_bdwt : IN STD_LOGIC;
    x_rsc_24_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_24_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_24_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_24_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_24_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_24_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_24_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_24_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_24_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_24_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_24_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_24_0_i_bcwt <= x_rsc_24_0_i_bcwt_drv;
  x_rsc_24_0_i_bcwt_1 <= x_rsc_24_0_i_bcwt_1_drv;

  x_rsc_24_0_i_wen_comp <= (NOT x_rsc_24_0_i_oswt) OR x_rsc_24_0_i_biwt OR x_rsc_24_0_i_bcwt_drv;
  x_rsc_24_0_i_wen_comp_1 <= (NOT x_rsc_24_0_i_oswt_1) OR x_rsc_24_0_i_biwt_1 OR
      x_rsc_24_0_i_bcwt_1_drv;
  x_rsc_24_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_24_0_i_s_raddr_core,
      x_rsc_24_0_i_s_raddr_core_sct);
  x_rsc_24_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_24_0_i_s_waddr_core,
      x_rsc_24_0_i_s_waddr_core_sct);
  x_rsc_24_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_24_0_i_s_din, x_rsc_24_0_i_s_din_bfwt,
      x_rsc_24_0_i_bcwt_drv);
  x_rsc_24_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_24_0_i_s_dout_core, x_rsc_24_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_24_0_i_bcwt_drv <= '0';
        x_rsc_24_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_24_0_i_bcwt_drv <= NOT((NOT(x_rsc_24_0_i_bcwt_drv OR x_rsc_24_0_i_biwt))
            OR x_rsc_24_0_i_bdwt);
        x_rsc_24_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_24_0_i_bcwt_1_drv OR x_rsc_24_0_i_biwt_1))
            OR x_rsc_24_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_24_0_i_biwt = '1' ) THEN
        x_rsc_24_0_i_s_din_bfwt <= x_rsc_24_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_24_0_i_oswt : IN STD_LOGIC;
    x_rsc_24_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_24_0_i_biwt : OUT STD_LOGIC;
    x_rsc_24_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_24_0_i_bcwt : IN STD_LOGIC;
    x_rsc_24_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_24_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_24_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_24_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_24_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_24_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_24_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_24_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_24_0_i_bdwt <= x_rsc_24_0_i_oswt AND core_wen;
  x_rsc_24_0_i_biwt <= x_rsc_24_0_i_ogwt AND x_rsc_24_0_i_s_rrdy;
  x_rsc_24_0_i_ogwt <= x_rsc_24_0_i_oswt AND (NOT x_rsc_24_0_i_bcwt);
  x_rsc_24_0_i_s_re_core_sct <= x_rsc_24_0_i_ogwt;
  x_rsc_24_0_i_bdwt_2 <= x_rsc_24_0_i_oswt_1 AND core_wen;
  x_rsc_24_0_i_biwt_1 <= x_rsc_24_0_i_ogwt_1 AND x_rsc_24_0_i_s_wrdy;
  x_rsc_24_0_i_ogwt_1 <= x_rsc_24_0_i_oswt_1 AND (NOT x_rsc_24_0_i_bcwt_1);
  x_rsc_24_0_i_s_we_core_sct <= x_rsc_24_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_23_0_i_oswt : IN STD_LOGIC;
    x_rsc_23_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_23_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_23_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_23_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_23_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_23_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_i_biwt : IN STD_LOGIC;
    x_rsc_23_0_i_bdwt : IN STD_LOGIC;
    x_rsc_23_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_23_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_23_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_23_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_23_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_23_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_23_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_23_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_23_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_23_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_23_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_23_0_i_bcwt <= x_rsc_23_0_i_bcwt_drv;
  x_rsc_23_0_i_bcwt_1 <= x_rsc_23_0_i_bcwt_1_drv;

  x_rsc_23_0_i_wen_comp <= (NOT x_rsc_23_0_i_oswt) OR x_rsc_23_0_i_biwt OR x_rsc_23_0_i_bcwt_drv;
  x_rsc_23_0_i_wen_comp_1 <= (NOT x_rsc_23_0_i_oswt_1) OR x_rsc_23_0_i_biwt_1 OR
      x_rsc_23_0_i_bcwt_1_drv;
  x_rsc_23_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_23_0_i_s_raddr_core,
      x_rsc_23_0_i_s_raddr_core_sct);
  x_rsc_23_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_23_0_i_s_waddr_core,
      x_rsc_23_0_i_s_waddr_core_sct);
  x_rsc_23_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_23_0_i_s_din, x_rsc_23_0_i_s_din_bfwt,
      x_rsc_23_0_i_bcwt_drv);
  x_rsc_23_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_23_0_i_s_dout_core, x_rsc_23_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_23_0_i_bcwt_drv <= '0';
        x_rsc_23_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_23_0_i_bcwt_drv <= NOT((NOT(x_rsc_23_0_i_bcwt_drv OR x_rsc_23_0_i_biwt))
            OR x_rsc_23_0_i_bdwt);
        x_rsc_23_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_23_0_i_bcwt_1_drv OR x_rsc_23_0_i_biwt_1))
            OR x_rsc_23_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_23_0_i_biwt = '1' ) THEN
        x_rsc_23_0_i_s_din_bfwt <= x_rsc_23_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_23_0_i_oswt : IN STD_LOGIC;
    x_rsc_23_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_23_0_i_biwt : OUT STD_LOGIC;
    x_rsc_23_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_23_0_i_bcwt : IN STD_LOGIC;
    x_rsc_23_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_23_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_23_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_23_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_23_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_23_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_23_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_23_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_23_0_i_bdwt <= x_rsc_23_0_i_oswt AND core_wen;
  x_rsc_23_0_i_biwt <= x_rsc_23_0_i_ogwt AND x_rsc_23_0_i_s_rrdy;
  x_rsc_23_0_i_ogwt <= x_rsc_23_0_i_oswt AND (NOT x_rsc_23_0_i_bcwt);
  x_rsc_23_0_i_s_re_core_sct <= x_rsc_23_0_i_ogwt;
  x_rsc_23_0_i_bdwt_2 <= x_rsc_23_0_i_oswt_1 AND core_wen;
  x_rsc_23_0_i_biwt_1 <= x_rsc_23_0_i_ogwt_1 AND x_rsc_23_0_i_s_wrdy;
  x_rsc_23_0_i_ogwt_1 <= x_rsc_23_0_i_oswt_1 AND (NOT x_rsc_23_0_i_bcwt_1);
  x_rsc_23_0_i_s_we_core_sct <= x_rsc_23_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_22_0_i_oswt : IN STD_LOGIC;
    x_rsc_22_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_22_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_22_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_22_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_22_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_22_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_i_biwt : IN STD_LOGIC;
    x_rsc_22_0_i_bdwt : IN STD_LOGIC;
    x_rsc_22_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_22_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_22_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_22_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_22_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_22_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_22_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_22_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_22_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_22_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_22_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_22_0_i_bcwt <= x_rsc_22_0_i_bcwt_drv;
  x_rsc_22_0_i_bcwt_1 <= x_rsc_22_0_i_bcwt_1_drv;

  x_rsc_22_0_i_wen_comp <= (NOT x_rsc_22_0_i_oswt) OR x_rsc_22_0_i_biwt OR x_rsc_22_0_i_bcwt_drv;
  x_rsc_22_0_i_wen_comp_1 <= (NOT x_rsc_22_0_i_oswt_1) OR x_rsc_22_0_i_biwt_1 OR
      x_rsc_22_0_i_bcwt_1_drv;
  x_rsc_22_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_22_0_i_s_raddr_core,
      x_rsc_22_0_i_s_raddr_core_sct);
  x_rsc_22_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_22_0_i_s_waddr_core,
      x_rsc_22_0_i_s_waddr_core_sct);
  x_rsc_22_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_22_0_i_s_din, x_rsc_22_0_i_s_din_bfwt,
      x_rsc_22_0_i_bcwt_drv);
  x_rsc_22_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_22_0_i_s_dout_core, x_rsc_22_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_22_0_i_bcwt_drv <= '0';
        x_rsc_22_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_22_0_i_bcwt_drv <= NOT((NOT(x_rsc_22_0_i_bcwt_drv OR x_rsc_22_0_i_biwt))
            OR x_rsc_22_0_i_bdwt);
        x_rsc_22_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_22_0_i_bcwt_1_drv OR x_rsc_22_0_i_biwt_1))
            OR x_rsc_22_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_22_0_i_biwt = '1' ) THEN
        x_rsc_22_0_i_s_din_bfwt <= x_rsc_22_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_22_0_i_oswt : IN STD_LOGIC;
    x_rsc_22_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_22_0_i_biwt : OUT STD_LOGIC;
    x_rsc_22_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_22_0_i_bcwt : IN STD_LOGIC;
    x_rsc_22_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_22_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_22_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_22_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_22_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_22_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_22_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_22_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_22_0_i_bdwt <= x_rsc_22_0_i_oswt AND core_wen;
  x_rsc_22_0_i_biwt <= x_rsc_22_0_i_ogwt AND x_rsc_22_0_i_s_rrdy;
  x_rsc_22_0_i_ogwt <= x_rsc_22_0_i_oswt AND (NOT x_rsc_22_0_i_bcwt);
  x_rsc_22_0_i_s_re_core_sct <= x_rsc_22_0_i_ogwt;
  x_rsc_22_0_i_bdwt_2 <= x_rsc_22_0_i_oswt_1 AND core_wen;
  x_rsc_22_0_i_biwt_1 <= x_rsc_22_0_i_ogwt_1 AND x_rsc_22_0_i_s_wrdy;
  x_rsc_22_0_i_ogwt_1 <= x_rsc_22_0_i_oswt_1 AND (NOT x_rsc_22_0_i_bcwt_1);
  x_rsc_22_0_i_s_we_core_sct <= x_rsc_22_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_21_0_i_oswt : IN STD_LOGIC;
    x_rsc_21_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_21_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_21_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_21_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_21_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_21_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_i_biwt : IN STD_LOGIC;
    x_rsc_21_0_i_bdwt : IN STD_LOGIC;
    x_rsc_21_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_21_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_21_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_21_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_21_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_21_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_21_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_21_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_21_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_21_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_21_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_21_0_i_bcwt <= x_rsc_21_0_i_bcwt_drv;
  x_rsc_21_0_i_bcwt_1 <= x_rsc_21_0_i_bcwt_1_drv;

  x_rsc_21_0_i_wen_comp <= (NOT x_rsc_21_0_i_oswt) OR x_rsc_21_0_i_biwt OR x_rsc_21_0_i_bcwt_drv;
  x_rsc_21_0_i_wen_comp_1 <= (NOT x_rsc_21_0_i_oswt_1) OR x_rsc_21_0_i_biwt_1 OR
      x_rsc_21_0_i_bcwt_1_drv;
  x_rsc_21_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_21_0_i_s_raddr_core,
      x_rsc_21_0_i_s_raddr_core_sct);
  x_rsc_21_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_21_0_i_s_waddr_core,
      x_rsc_21_0_i_s_waddr_core_sct);
  x_rsc_21_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_21_0_i_s_din, x_rsc_21_0_i_s_din_bfwt,
      x_rsc_21_0_i_bcwt_drv);
  x_rsc_21_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_21_0_i_s_dout_core, x_rsc_21_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_21_0_i_bcwt_drv <= '0';
        x_rsc_21_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_21_0_i_bcwt_drv <= NOT((NOT(x_rsc_21_0_i_bcwt_drv OR x_rsc_21_0_i_biwt))
            OR x_rsc_21_0_i_bdwt);
        x_rsc_21_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_21_0_i_bcwt_1_drv OR x_rsc_21_0_i_biwt_1))
            OR x_rsc_21_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_21_0_i_biwt = '1' ) THEN
        x_rsc_21_0_i_s_din_bfwt <= x_rsc_21_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_21_0_i_oswt : IN STD_LOGIC;
    x_rsc_21_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_21_0_i_biwt : OUT STD_LOGIC;
    x_rsc_21_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_21_0_i_bcwt : IN STD_LOGIC;
    x_rsc_21_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_21_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_21_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_21_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_21_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_21_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_21_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_21_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_21_0_i_bdwt <= x_rsc_21_0_i_oswt AND core_wen;
  x_rsc_21_0_i_biwt <= x_rsc_21_0_i_ogwt AND x_rsc_21_0_i_s_rrdy;
  x_rsc_21_0_i_ogwt <= x_rsc_21_0_i_oswt AND (NOT x_rsc_21_0_i_bcwt);
  x_rsc_21_0_i_s_re_core_sct <= x_rsc_21_0_i_ogwt;
  x_rsc_21_0_i_bdwt_2 <= x_rsc_21_0_i_oswt_1 AND core_wen;
  x_rsc_21_0_i_biwt_1 <= x_rsc_21_0_i_ogwt_1 AND x_rsc_21_0_i_s_wrdy;
  x_rsc_21_0_i_ogwt_1 <= x_rsc_21_0_i_oswt_1 AND (NOT x_rsc_21_0_i_bcwt_1);
  x_rsc_21_0_i_s_we_core_sct <= x_rsc_21_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_20_0_i_oswt : IN STD_LOGIC;
    x_rsc_20_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_20_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_20_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_20_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_20_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_20_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_i_biwt : IN STD_LOGIC;
    x_rsc_20_0_i_bdwt : IN STD_LOGIC;
    x_rsc_20_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_20_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_20_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_20_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_20_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_20_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_20_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_20_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_20_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_20_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_20_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_20_0_i_bcwt <= x_rsc_20_0_i_bcwt_drv;
  x_rsc_20_0_i_bcwt_1 <= x_rsc_20_0_i_bcwt_1_drv;

  x_rsc_20_0_i_wen_comp <= (NOT x_rsc_20_0_i_oswt) OR x_rsc_20_0_i_biwt OR x_rsc_20_0_i_bcwt_drv;
  x_rsc_20_0_i_wen_comp_1 <= (NOT x_rsc_20_0_i_oswt_1) OR x_rsc_20_0_i_biwt_1 OR
      x_rsc_20_0_i_bcwt_1_drv;
  x_rsc_20_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_20_0_i_s_raddr_core,
      x_rsc_20_0_i_s_raddr_core_sct);
  x_rsc_20_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_20_0_i_s_waddr_core,
      x_rsc_20_0_i_s_waddr_core_sct);
  x_rsc_20_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_20_0_i_s_din, x_rsc_20_0_i_s_din_bfwt,
      x_rsc_20_0_i_bcwt_drv);
  x_rsc_20_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_20_0_i_s_dout_core, x_rsc_20_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_20_0_i_bcwt_drv <= '0';
        x_rsc_20_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_20_0_i_bcwt_drv <= NOT((NOT(x_rsc_20_0_i_bcwt_drv OR x_rsc_20_0_i_biwt))
            OR x_rsc_20_0_i_bdwt);
        x_rsc_20_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_20_0_i_bcwt_1_drv OR x_rsc_20_0_i_biwt_1))
            OR x_rsc_20_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_20_0_i_biwt = '1' ) THEN
        x_rsc_20_0_i_s_din_bfwt <= x_rsc_20_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_20_0_i_oswt : IN STD_LOGIC;
    x_rsc_20_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_20_0_i_biwt : OUT STD_LOGIC;
    x_rsc_20_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_20_0_i_bcwt : IN STD_LOGIC;
    x_rsc_20_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_20_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_20_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_20_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_20_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_20_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_20_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_20_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_20_0_i_bdwt <= x_rsc_20_0_i_oswt AND core_wen;
  x_rsc_20_0_i_biwt <= x_rsc_20_0_i_ogwt AND x_rsc_20_0_i_s_rrdy;
  x_rsc_20_0_i_ogwt <= x_rsc_20_0_i_oswt AND (NOT x_rsc_20_0_i_bcwt);
  x_rsc_20_0_i_s_re_core_sct <= x_rsc_20_0_i_ogwt;
  x_rsc_20_0_i_bdwt_2 <= x_rsc_20_0_i_oswt_1 AND core_wen;
  x_rsc_20_0_i_biwt_1 <= x_rsc_20_0_i_ogwt_1 AND x_rsc_20_0_i_s_wrdy;
  x_rsc_20_0_i_ogwt_1 <= x_rsc_20_0_i_oswt_1 AND (NOT x_rsc_20_0_i_bcwt_1);
  x_rsc_20_0_i_s_we_core_sct <= x_rsc_20_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_19_0_i_oswt : IN STD_LOGIC;
    x_rsc_19_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_19_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_19_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_19_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_19_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_19_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_i_biwt : IN STD_LOGIC;
    x_rsc_19_0_i_bdwt : IN STD_LOGIC;
    x_rsc_19_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_19_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_19_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_19_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_19_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_19_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_19_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_19_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_19_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_19_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_19_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_19_0_i_bcwt <= x_rsc_19_0_i_bcwt_drv;
  x_rsc_19_0_i_bcwt_1 <= x_rsc_19_0_i_bcwt_1_drv;

  x_rsc_19_0_i_wen_comp <= (NOT x_rsc_19_0_i_oswt) OR x_rsc_19_0_i_biwt OR x_rsc_19_0_i_bcwt_drv;
  x_rsc_19_0_i_wen_comp_1 <= (NOT x_rsc_19_0_i_oswt_1) OR x_rsc_19_0_i_biwt_1 OR
      x_rsc_19_0_i_bcwt_1_drv;
  x_rsc_19_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_19_0_i_s_raddr_core,
      x_rsc_19_0_i_s_raddr_core_sct);
  x_rsc_19_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_19_0_i_s_waddr_core,
      x_rsc_19_0_i_s_waddr_core_sct);
  x_rsc_19_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_19_0_i_s_din, x_rsc_19_0_i_s_din_bfwt,
      x_rsc_19_0_i_bcwt_drv);
  x_rsc_19_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_19_0_i_s_dout_core, x_rsc_19_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_19_0_i_bcwt_drv <= '0';
        x_rsc_19_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_19_0_i_bcwt_drv <= NOT((NOT(x_rsc_19_0_i_bcwt_drv OR x_rsc_19_0_i_biwt))
            OR x_rsc_19_0_i_bdwt);
        x_rsc_19_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_19_0_i_bcwt_1_drv OR x_rsc_19_0_i_biwt_1))
            OR x_rsc_19_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_19_0_i_biwt = '1' ) THEN
        x_rsc_19_0_i_s_din_bfwt <= x_rsc_19_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_19_0_i_oswt : IN STD_LOGIC;
    x_rsc_19_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_19_0_i_biwt : OUT STD_LOGIC;
    x_rsc_19_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_19_0_i_bcwt : IN STD_LOGIC;
    x_rsc_19_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_19_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_19_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_19_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_19_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_19_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_19_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_19_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_19_0_i_bdwt <= x_rsc_19_0_i_oswt AND core_wen;
  x_rsc_19_0_i_biwt <= x_rsc_19_0_i_ogwt AND x_rsc_19_0_i_s_rrdy;
  x_rsc_19_0_i_ogwt <= x_rsc_19_0_i_oswt AND (NOT x_rsc_19_0_i_bcwt);
  x_rsc_19_0_i_s_re_core_sct <= x_rsc_19_0_i_ogwt;
  x_rsc_19_0_i_bdwt_2 <= x_rsc_19_0_i_oswt_1 AND core_wen;
  x_rsc_19_0_i_biwt_1 <= x_rsc_19_0_i_ogwt_1 AND x_rsc_19_0_i_s_wrdy;
  x_rsc_19_0_i_ogwt_1 <= x_rsc_19_0_i_oswt_1 AND (NOT x_rsc_19_0_i_bcwt_1);
  x_rsc_19_0_i_s_we_core_sct <= x_rsc_19_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_18_0_i_oswt : IN STD_LOGIC;
    x_rsc_18_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_18_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_18_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_18_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_18_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_18_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_i_biwt : IN STD_LOGIC;
    x_rsc_18_0_i_bdwt : IN STD_LOGIC;
    x_rsc_18_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_18_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_18_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_18_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_18_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_18_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_18_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_18_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_18_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_18_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_18_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_18_0_i_bcwt <= x_rsc_18_0_i_bcwt_drv;
  x_rsc_18_0_i_bcwt_1 <= x_rsc_18_0_i_bcwt_1_drv;

  x_rsc_18_0_i_wen_comp <= (NOT x_rsc_18_0_i_oswt) OR x_rsc_18_0_i_biwt OR x_rsc_18_0_i_bcwt_drv;
  x_rsc_18_0_i_wen_comp_1 <= (NOT x_rsc_18_0_i_oswt_1) OR x_rsc_18_0_i_biwt_1 OR
      x_rsc_18_0_i_bcwt_1_drv;
  x_rsc_18_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_18_0_i_s_raddr_core,
      x_rsc_18_0_i_s_raddr_core_sct);
  x_rsc_18_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_18_0_i_s_waddr_core,
      x_rsc_18_0_i_s_waddr_core_sct);
  x_rsc_18_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_18_0_i_s_din, x_rsc_18_0_i_s_din_bfwt,
      x_rsc_18_0_i_bcwt_drv);
  x_rsc_18_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_18_0_i_s_dout_core, x_rsc_18_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_18_0_i_bcwt_drv <= '0';
        x_rsc_18_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_18_0_i_bcwt_drv <= NOT((NOT(x_rsc_18_0_i_bcwt_drv OR x_rsc_18_0_i_biwt))
            OR x_rsc_18_0_i_bdwt);
        x_rsc_18_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_18_0_i_bcwt_1_drv OR x_rsc_18_0_i_biwt_1))
            OR x_rsc_18_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_18_0_i_biwt = '1' ) THEN
        x_rsc_18_0_i_s_din_bfwt <= x_rsc_18_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_18_0_i_oswt : IN STD_LOGIC;
    x_rsc_18_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_18_0_i_biwt : OUT STD_LOGIC;
    x_rsc_18_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_18_0_i_bcwt : IN STD_LOGIC;
    x_rsc_18_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_18_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_18_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_18_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_18_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_18_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_18_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_18_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_18_0_i_bdwt <= x_rsc_18_0_i_oswt AND core_wen;
  x_rsc_18_0_i_biwt <= x_rsc_18_0_i_ogwt AND x_rsc_18_0_i_s_rrdy;
  x_rsc_18_0_i_ogwt <= x_rsc_18_0_i_oswt AND (NOT x_rsc_18_0_i_bcwt);
  x_rsc_18_0_i_s_re_core_sct <= x_rsc_18_0_i_ogwt;
  x_rsc_18_0_i_bdwt_2 <= x_rsc_18_0_i_oswt_1 AND core_wen;
  x_rsc_18_0_i_biwt_1 <= x_rsc_18_0_i_ogwt_1 AND x_rsc_18_0_i_s_wrdy;
  x_rsc_18_0_i_ogwt_1 <= x_rsc_18_0_i_oswt_1 AND (NOT x_rsc_18_0_i_bcwt_1);
  x_rsc_18_0_i_s_we_core_sct <= x_rsc_18_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_17_0_i_oswt : IN STD_LOGIC;
    x_rsc_17_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_17_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_17_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_17_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_17_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_17_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_i_biwt : IN STD_LOGIC;
    x_rsc_17_0_i_bdwt : IN STD_LOGIC;
    x_rsc_17_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_17_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_17_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_17_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_17_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_17_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_17_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_17_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_17_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_17_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_17_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_17_0_i_bcwt <= x_rsc_17_0_i_bcwt_drv;
  x_rsc_17_0_i_bcwt_1 <= x_rsc_17_0_i_bcwt_1_drv;

  x_rsc_17_0_i_wen_comp <= (NOT x_rsc_17_0_i_oswt) OR x_rsc_17_0_i_biwt OR x_rsc_17_0_i_bcwt_drv;
  x_rsc_17_0_i_wen_comp_1 <= (NOT x_rsc_17_0_i_oswt_1) OR x_rsc_17_0_i_biwt_1 OR
      x_rsc_17_0_i_bcwt_1_drv;
  x_rsc_17_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_17_0_i_s_raddr_core,
      x_rsc_17_0_i_s_raddr_core_sct);
  x_rsc_17_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_17_0_i_s_waddr_core,
      x_rsc_17_0_i_s_waddr_core_sct);
  x_rsc_17_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_17_0_i_s_din, x_rsc_17_0_i_s_din_bfwt,
      x_rsc_17_0_i_bcwt_drv);
  x_rsc_17_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_17_0_i_s_dout_core, x_rsc_17_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_17_0_i_bcwt_drv <= '0';
        x_rsc_17_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_17_0_i_bcwt_drv <= NOT((NOT(x_rsc_17_0_i_bcwt_drv OR x_rsc_17_0_i_biwt))
            OR x_rsc_17_0_i_bdwt);
        x_rsc_17_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_17_0_i_bcwt_1_drv OR x_rsc_17_0_i_biwt_1))
            OR x_rsc_17_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_17_0_i_biwt = '1' ) THEN
        x_rsc_17_0_i_s_din_bfwt <= x_rsc_17_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_17_0_i_oswt : IN STD_LOGIC;
    x_rsc_17_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_17_0_i_biwt : OUT STD_LOGIC;
    x_rsc_17_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_17_0_i_bcwt : IN STD_LOGIC;
    x_rsc_17_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_17_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_17_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_17_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_17_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_17_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_17_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_17_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_17_0_i_bdwt <= x_rsc_17_0_i_oswt AND core_wen;
  x_rsc_17_0_i_biwt <= x_rsc_17_0_i_ogwt AND x_rsc_17_0_i_s_rrdy;
  x_rsc_17_0_i_ogwt <= x_rsc_17_0_i_oswt AND (NOT x_rsc_17_0_i_bcwt);
  x_rsc_17_0_i_s_re_core_sct <= x_rsc_17_0_i_ogwt;
  x_rsc_17_0_i_bdwt_2 <= x_rsc_17_0_i_oswt_1 AND core_wen;
  x_rsc_17_0_i_biwt_1 <= x_rsc_17_0_i_ogwt_1 AND x_rsc_17_0_i_s_wrdy;
  x_rsc_17_0_i_ogwt_1 <= x_rsc_17_0_i_oswt_1 AND (NOT x_rsc_17_0_i_bcwt_1);
  x_rsc_17_0_i_s_we_core_sct <= x_rsc_17_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_16_0_i_oswt : IN STD_LOGIC;
    x_rsc_16_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_16_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_16_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_16_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_16_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_16_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_i_biwt : IN STD_LOGIC;
    x_rsc_16_0_i_bdwt : IN STD_LOGIC;
    x_rsc_16_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_16_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_16_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_16_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_16_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_16_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_16_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_16_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_16_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_16_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_16_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_16_0_i_bcwt <= x_rsc_16_0_i_bcwt_drv;
  x_rsc_16_0_i_bcwt_1 <= x_rsc_16_0_i_bcwt_1_drv;

  x_rsc_16_0_i_wen_comp <= (NOT x_rsc_16_0_i_oswt) OR x_rsc_16_0_i_biwt OR x_rsc_16_0_i_bcwt_drv;
  x_rsc_16_0_i_wen_comp_1 <= (NOT x_rsc_16_0_i_oswt_1) OR x_rsc_16_0_i_biwt_1 OR
      x_rsc_16_0_i_bcwt_1_drv;
  x_rsc_16_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_16_0_i_s_raddr_core,
      x_rsc_16_0_i_s_raddr_core_sct);
  x_rsc_16_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_16_0_i_s_waddr_core,
      x_rsc_16_0_i_s_waddr_core_sct);
  x_rsc_16_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_16_0_i_s_din, x_rsc_16_0_i_s_din_bfwt,
      x_rsc_16_0_i_bcwt_drv);
  x_rsc_16_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_16_0_i_s_dout_core, x_rsc_16_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_16_0_i_bcwt_drv <= '0';
        x_rsc_16_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_16_0_i_bcwt_drv <= NOT((NOT(x_rsc_16_0_i_bcwt_drv OR x_rsc_16_0_i_biwt))
            OR x_rsc_16_0_i_bdwt);
        x_rsc_16_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_16_0_i_bcwt_1_drv OR x_rsc_16_0_i_biwt_1))
            OR x_rsc_16_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_16_0_i_biwt = '1' ) THEN
        x_rsc_16_0_i_s_din_bfwt <= x_rsc_16_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_16_0_i_oswt : IN STD_LOGIC;
    x_rsc_16_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_16_0_i_biwt : OUT STD_LOGIC;
    x_rsc_16_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_16_0_i_bcwt : IN STD_LOGIC;
    x_rsc_16_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_16_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_16_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_16_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_16_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_16_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_16_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_16_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_16_0_i_bdwt <= x_rsc_16_0_i_oswt AND core_wen;
  x_rsc_16_0_i_biwt <= x_rsc_16_0_i_ogwt AND x_rsc_16_0_i_s_rrdy;
  x_rsc_16_0_i_ogwt <= x_rsc_16_0_i_oswt AND (NOT x_rsc_16_0_i_bcwt);
  x_rsc_16_0_i_s_re_core_sct <= x_rsc_16_0_i_ogwt;
  x_rsc_16_0_i_bdwt_2 <= x_rsc_16_0_i_oswt_1 AND core_wen;
  x_rsc_16_0_i_biwt_1 <= x_rsc_16_0_i_ogwt_1 AND x_rsc_16_0_i_s_wrdy;
  x_rsc_16_0_i_ogwt_1 <= x_rsc_16_0_i_oswt_1 AND (NOT x_rsc_16_0_i_bcwt_1);
  x_rsc_16_0_i_s_we_core_sct <= x_rsc_16_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_15_0_i_oswt : IN STD_LOGIC;
    x_rsc_15_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_15_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_15_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_15_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_15_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_15_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_i_biwt : IN STD_LOGIC;
    x_rsc_15_0_i_bdwt : IN STD_LOGIC;
    x_rsc_15_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_15_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_15_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_15_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_15_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_15_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_15_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_15_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_15_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_15_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_15_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_15_0_i_bcwt <= x_rsc_15_0_i_bcwt_drv;
  x_rsc_15_0_i_bcwt_1 <= x_rsc_15_0_i_bcwt_1_drv;

  x_rsc_15_0_i_wen_comp <= (NOT x_rsc_15_0_i_oswt) OR x_rsc_15_0_i_biwt OR x_rsc_15_0_i_bcwt_drv;
  x_rsc_15_0_i_wen_comp_1 <= (NOT x_rsc_15_0_i_oswt_1) OR x_rsc_15_0_i_biwt_1 OR
      x_rsc_15_0_i_bcwt_1_drv;
  x_rsc_15_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_15_0_i_s_raddr_core,
      x_rsc_15_0_i_s_raddr_core_sct);
  x_rsc_15_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_15_0_i_s_waddr_core,
      x_rsc_15_0_i_s_waddr_core_sct);
  x_rsc_15_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_15_0_i_s_din, x_rsc_15_0_i_s_din_bfwt,
      x_rsc_15_0_i_bcwt_drv);
  x_rsc_15_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_15_0_i_s_dout_core, x_rsc_15_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_15_0_i_bcwt_drv <= '0';
        x_rsc_15_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_15_0_i_bcwt_drv <= NOT((NOT(x_rsc_15_0_i_bcwt_drv OR x_rsc_15_0_i_biwt))
            OR x_rsc_15_0_i_bdwt);
        x_rsc_15_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_15_0_i_bcwt_1_drv OR x_rsc_15_0_i_biwt_1))
            OR x_rsc_15_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_15_0_i_biwt = '1' ) THEN
        x_rsc_15_0_i_s_din_bfwt <= x_rsc_15_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_15_0_i_oswt : IN STD_LOGIC;
    x_rsc_15_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_15_0_i_biwt : OUT STD_LOGIC;
    x_rsc_15_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_15_0_i_bcwt : IN STD_LOGIC;
    x_rsc_15_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_15_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_15_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_15_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_15_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_15_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_15_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_15_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_15_0_i_bdwt <= x_rsc_15_0_i_oswt AND core_wen;
  x_rsc_15_0_i_biwt <= x_rsc_15_0_i_ogwt AND x_rsc_15_0_i_s_rrdy;
  x_rsc_15_0_i_ogwt <= x_rsc_15_0_i_oswt AND (NOT x_rsc_15_0_i_bcwt);
  x_rsc_15_0_i_s_re_core_sct <= x_rsc_15_0_i_ogwt;
  x_rsc_15_0_i_bdwt_2 <= x_rsc_15_0_i_oswt_1 AND core_wen;
  x_rsc_15_0_i_biwt_1 <= x_rsc_15_0_i_ogwt_1 AND x_rsc_15_0_i_s_wrdy;
  x_rsc_15_0_i_ogwt_1 <= x_rsc_15_0_i_oswt_1 AND (NOT x_rsc_15_0_i_bcwt_1);
  x_rsc_15_0_i_s_we_core_sct <= x_rsc_15_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_14_0_i_oswt : IN STD_LOGIC;
    x_rsc_14_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_14_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_14_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_14_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_14_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_14_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_i_biwt : IN STD_LOGIC;
    x_rsc_14_0_i_bdwt : IN STD_LOGIC;
    x_rsc_14_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_14_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_14_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_14_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_14_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_14_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_14_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_14_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_14_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_14_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_14_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_14_0_i_bcwt <= x_rsc_14_0_i_bcwt_drv;
  x_rsc_14_0_i_bcwt_1 <= x_rsc_14_0_i_bcwt_1_drv;

  x_rsc_14_0_i_wen_comp <= (NOT x_rsc_14_0_i_oswt) OR x_rsc_14_0_i_biwt OR x_rsc_14_0_i_bcwt_drv;
  x_rsc_14_0_i_wen_comp_1 <= (NOT x_rsc_14_0_i_oswt_1) OR x_rsc_14_0_i_biwt_1 OR
      x_rsc_14_0_i_bcwt_1_drv;
  x_rsc_14_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_14_0_i_s_raddr_core,
      x_rsc_14_0_i_s_raddr_core_sct);
  x_rsc_14_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_14_0_i_s_waddr_core,
      x_rsc_14_0_i_s_waddr_core_sct);
  x_rsc_14_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_14_0_i_s_din, x_rsc_14_0_i_s_din_bfwt,
      x_rsc_14_0_i_bcwt_drv);
  x_rsc_14_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_14_0_i_s_dout_core, x_rsc_14_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_14_0_i_bcwt_drv <= '0';
        x_rsc_14_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_14_0_i_bcwt_drv <= NOT((NOT(x_rsc_14_0_i_bcwt_drv OR x_rsc_14_0_i_biwt))
            OR x_rsc_14_0_i_bdwt);
        x_rsc_14_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_14_0_i_bcwt_1_drv OR x_rsc_14_0_i_biwt_1))
            OR x_rsc_14_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_14_0_i_biwt = '1' ) THEN
        x_rsc_14_0_i_s_din_bfwt <= x_rsc_14_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_14_0_i_oswt : IN STD_LOGIC;
    x_rsc_14_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_14_0_i_biwt : OUT STD_LOGIC;
    x_rsc_14_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_14_0_i_bcwt : IN STD_LOGIC;
    x_rsc_14_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_14_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_14_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_14_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_14_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_14_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_14_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_14_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_14_0_i_bdwt <= x_rsc_14_0_i_oswt AND core_wen;
  x_rsc_14_0_i_biwt <= x_rsc_14_0_i_ogwt AND x_rsc_14_0_i_s_rrdy;
  x_rsc_14_0_i_ogwt <= x_rsc_14_0_i_oswt AND (NOT x_rsc_14_0_i_bcwt);
  x_rsc_14_0_i_s_re_core_sct <= x_rsc_14_0_i_ogwt;
  x_rsc_14_0_i_bdwt_2 <= x_rsc_14_0_i_oswt_1 AND core_wen;
  x_rsc_14_0_i_biwt_1 <= x_rsc_14_0_i_ogwt_1 AND x_rsc_14_0_i_s_wrdy;
  x_rsc_14_0_i_ogwt_1 <= x_rsc_14_0_i_oswt_1 AND (NOT x_rsc_14_0_i_bcwt_1);
  x_rsc_14_0_i_s_we_core_sct <= x_rsc_14_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_13_0_i_oswt : IN STD_LOGIC;
    x_rsc_13_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_13_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_13_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_13_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_13_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_13_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_i_biwt : IN STD_LOGIC;
    x_rsc_13_0_i_bdwt : IN STD_LOGIC;
    x_rsc_13_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_13_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_13_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_13_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_13_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_13_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_13_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_13_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_13_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_13_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_13_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_13_0_i_bcwt <= x_rsc_13_0_i_bcwt_drv;
  x_rsc_13_0_i_bcwt_1 <= x_rsc_13_0_i_bcwt_1_drv;

  x_rsc_13_0_i_wen_comp <= (NOT x_rsc_13_0_i_oswt) OR x_rsc_13_0_i_biwt OR x_rsc_13_0_i_bcwt_drv;
  x_rsc_13_0_i_wen_comp_1 <= (NOT x_rsc_13_0_i_oswt_1) OR x_rsc_13_0_i_biwt_1 OR
      x_rsc_13_0_i_bcwt_1_drv;
  x_rsc_13_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_13_0_i_s_raddr_core,
      x_rsc_13_0_i_s_raddr_core_sct);
  x_rsc_13_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_13_0_i_s_waddr_core,
      x_rsc_13_0_i_s_waddr_core_sct);
  x_rsc_13_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_13_0_i_s_din, x_rsc_13_0_i_s_din_bfwt,
      x_rsc_13_0_i_bcwt_drv);
  x_rsc_13_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_13_0_i_s_dout_core, x_rsc_13_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_13_0_i_bcwt_drv <= '0';
        x_rsc_13_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_13_0_i_bcwt_drv <= NOT((NOT(x_rsc_13_0_i_bcwt_drv OR x_rsc_13_0_i_biwt))
            OR x_rsc_13_0_i_bdwt);
        x_rsc_13_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_13_0_i_bcwt_1_drv OR x_rsc_13_0_i_biwt_1))
            OR x_rsc_13_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_13_0_i_biwt = '1' ) THEN
        x_rsc_13_0_i_s_din_bfwt <= x_rsc_13_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_13_0_i_oswt : IN STD_LOGIC;
    x_rsc_13_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_13_0_i_biwt : OUT STD_LOGIC;
    x_rsc_13_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_13_0_i_bcwt : IN STD_LOGIC;
    x_rsc_13_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_13_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_13_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_13_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_13_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_13_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_13_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_13_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_13_0_i_bdwt <= x_rsc_13_0_i_oswt AND core_wen;
  x_rsc_13_0_i_biwt <= x_rsc_13_0_i_ogwt AND x_rsc_13_0_i_s_rrdy;
  x_rsc_13_0_i_ogwt <= x_rsc_13_0_i_oswt AND (NOT x_rsc_13_0_i_bcwt);
  x_rsc_13_0_i_s_re_core_sct <= x_rsc_13_0_i_ogwt;
  x_rsc_13_0_i_bdwt_2 <= x_rsc_13_0_i_oswt_1 AND core_wen;
  x_rsc_13_0_i_biwt_1 <= x_rsc_13_0_i_ogwt_1 AND x_rsc_13_0_i_s_wrdy;
  x_rsc_13_0_i_ogwt_1 <= x_rsc_13_0_i_oswt_1 AND (NOT x_rsc_13_0_i_bcwt_1);
  x_rsc_13_0_i_s_we_core_sct <= x_rsc_13_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_12_0_i_oswt : IN STD_LOGIC;
    x_rsc_12_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_12_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_12_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_12_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_12_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_12_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_i_biwt : IN STD_LOGIC;
    x_rsc_12_0_i_bdwt : IN STD_LOGIC;
    x_rsc_12_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_12_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_12_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_12_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_12_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_12_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_12_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_12_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_12_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_12_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_12_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_12_0_i_bcwt <= x_rsc_12_0_i_bcwt_drv;
  x_rsc_12_0_i_bcwt_1 <= x_rsc_12_0_i_bcwt_1_drv;

  x_rsc_12_0_i_wen_comp <= (NOT x_rsc_12_0_i_oswt) OR x_rsc_12_0_i_biwt OR x_rsc_12_0_i_bcwt_drv;
  x_rsc_12_0_i_wen_comp_1 <= (NOT x_rsc_12_0_i_oswt_1) OR x_rsc_12_0_i_biwt_1 OR
      x_rsc_12_0_i_bcwt_1_drv;
  x_rsc_12_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_12_0_i_s_raddr_core,
      x_rsc_12_0_i_s_raddr_core_sct);
  x_rsc_12_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_12_0_i_s_waddr_core,
      x_rsc_12_0_i_s_waddr_core_sct);
  x_rsc_12_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_12_0_i_s_din, x_rsc_12_0_i_s_din_bfwt,
      x_rsc_12_0_i_bcwt_drv);
  x_rsc_12_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_12_0_i_s_dout_core, x_rsc_12_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_12_0_i_bcwt_drv <= '0';
        x_rsc_12_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_12_0_i_bcwt_drv <= NOT((NOT(x_rsc_12_0_i_bcwt_drv OR x_rsc_12_0_i_biwt))
            OR x_rsc_12_0_i_bdwt);
        x_rsc_12_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_12_0_i_bcwt_1_drv OR x_rsc_12_0_i_biwt_1))
            OR x_rsc_12_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_12_0_i_biwt = '1' ) THEN
        x_rsc_12_0_i_s_din_bfwt <= x_rsc_12_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_12_0_i_oswt : IN STD_LOGIC;
    x_rsc_12_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_12_0_i_biwt : OUT STD_LOGIC;
    x_rsc_12_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_12_0_i_bcwt : IN STD_LOGIC;
    x_rsc_12_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_12_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_12_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_12_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_12_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_12_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_12_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_12_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_12_0_i_bdwt <= x_rsc_12_0_i_oswt AND core_wen;
  x_rsc_12_0_i_biwt <= x_rsc_12_0_i_ogwt AND x_rsc_12_0_i_s_rrdy;
  x_rsc_12_0_i_ogwt <= x_rsc_12_0_i_oswt AND (NOT x_rsc_12_0_i_bcwt);
  x_rsc_12_0_i_s_re_core_sct <= x_rsc_12_0_i_ogwt;
  x_rsc_12_0_i_bdwt_2 <= x_rsc_12_0_i_oswt_1 AND core_wen;
  x_rsc_12_0_i_biwt_1 <= x_rsc_12_0_i_ogwt_1 AND x_rsc_12_0_i_s_wrdy;
  x_rsc_12_0_i_ogwt_1 <= x_rsc_12_0_i_oswt_1 AND (NOT x_rsc_12_0_i_bcwt_1);
  x_rsc_12_0_i_s_we_core_sct <= x_rsc_12_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_11_0_i_oswt : IN STD_LOGIC;
    x_rsc_11_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_11_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_11_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_11_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_11_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_11_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_i_biwt : IN STD_LOGIC;
    x_rsc_11_0_i_bdwt : IN STD_LOGIC;
    x_rsc_11_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_11_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_11_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_11_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_11_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_11_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_11_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_11_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_11_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_11_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_11_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_11_0_i_bcwt <= x_rsc_11_0_i_bcwt_drv;
  x_rsc_11_0_i_bcwt_1 <= x_rsc_11_0_i_bcwt_1_drv;

  x_rsc_11_0_i_wen_comp <= (NOT x_rsc_11_0_i_oswt) OR x_rsc_11_0_i_biwt OR x_rsc_11_0_i_bcwt_drv;
  x_rsc_11_0_i_wen_comp_1 <= (NOT x_rsc_11_0_i_oswt_1) OR x_rsc_11_0_i_biwt_1 OR
      x_rsc_11_0_i_bcwt_1_drv;
  x_rsc_11_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_11_0_i_s_raddr_core,
      x_rsc_11_0_i_s_raddr_core_sct);
  x_rsc_11_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_11_0_i_s_waddr_core,
      x_rsc_11_0_i_s_waddr_core_sct);
  x_rsc_11_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_11_0_i_s_din, x_rsc_11_0_i_s_din_bfwt,
      x_rsc_11_0_i_bcwt_drv);
  x_rsc_11_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_11_0_i_s_dout_core, x_rsc_11_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_11_0_i_bcwt_drv <= '0';
        x_rsc_11_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_11_0_i_bcwt_drv <= NOT((NOT(x_rsc_11_0_i_bcwt_drv OR x_rsc_11_0_i_biwt))
            OR x_rsc_11_0_i_bdwt);
        x_rsc_11_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_11_0_i_bcwt_1_drv OR x_rsc_11_0_i_biwt_1))
            OR x_rsc_11_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_11_0_i_biwt = '1' ) THEN
        x_rsc_11_0_i_s_din_bfwt <= x_rsc_11_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_11_0_i_oswt : IN STD_LOGIC;
    x_rsc_11_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_11_0_i_biwt : OUT STD_LOGIC;
    x_rsc_11_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_11_0_i_bcwt : IN STD_LOGIC;
    x_rsc_11_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_11_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_11_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_11_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_11_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_11_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_11_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_11_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_11_0_i_bdwt <= x_rsc_11_0_i_oswt AND core_wen;
  x_rsc_11_0_i_biwt <= x_rsc_11_0_i_ogwt AND x_rsc_11_0_i_s_rrdy;
  x_rsc_11_0_i_ogwt <= x_rsc_11_0_i_oswt AND (NOT x_rsc_11_0_i_bcwt);
  x_rsc_11_0_i_s_re_core_sct <= x_rsc_11_0_i_ogwt;
  x_rsc_11_0_i_bdwt_2 <= x_rsc_11_0_i_oswt_1 AND core_wen;
  x_rsc_11_0_i_biwt_1 <= x_rsc_11_0_i_ogwt_1 AND x_rsc_11_0_i_s_wrdy;
  x_rsc_11_0_i_ogwt_1 <= x_rsc_11_0_i_oswt_1 AND (NOT x_rsc_11_0_i_bcwt_1);
  x_rsc_11_0_i_s_we_core_sct <= x_rsc_11_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_10_0_i_oswt : IN STD_LOGIC;
    x_rsc_10_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_10_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_10_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_10_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_10_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_10_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_i_biwt : IN STD_LOGIC;
    x_rsc_10_0_i_bdwt : IN STD_LOGIC;
    x_rsc_10_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_10_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_10_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_10_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_10_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_10_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_10_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_10_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_10_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_10_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_10_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_10_0_i_bcwt <= x_rsc_10_0_i_bcwt_drv;
  x_rsc_10_0_i_bcwt_1 <= x_rsc_10_0_i_bcwt_1_drv;

  x_rsc_10_0_i_wen_comp <= (NOT x_rsc_10_0_i_oswt) OR x_rsc_10_0_i_biwt OR x_rsc_10_0_i_bcwt_drv;
  x_rsc_10_0_i_wen_comp_1 <= (NOT x_rsc_10_0_i_oswt_1) OR x_rsc_10_0_i_biwt_1 OR
      x_rsc_10_0_i_bcwt_1_drv;
  x_rsc_10_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_10_0_i_s_raddr_core,
      x_rsc_10_0_i_s_raddr_core_sct);
  x_rsc_10_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_10_0_i_s_waddr_core,
      x_rsc_10_0_i_s_waddr_core_sct);
  x_rsc_10_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_10_0_i_s_din, x_rsc_10_0_i_s_din_bfwt,
      x_rsc_10_0_i_bcwt_drv);
  x_rsc_10_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_10_0_i_s_dout_core, x_rsc_10_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_10_0_i_bcwt_drv <= '0';
        x_rsc_10_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_10_0_i_bcwt_drv <= NOT((NOT(x_rsc_10_0_i_bcwt_drv OR x_rsc_10_0_i_biwt))
            OR x_rsc_10_0_i_bdwt);
        x_rsc_10_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_10_0_i_bcwt_1_drv OR x_rsc_10_0_i_biwt_1))
            OR x_rsc_10_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_10_0_i_biwt = '1' ) THEN
        x_rsc_10_0_i_s_din_bfwt <= x_rsc_10_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_10_0_i_oswt : IN STD_LOGIC;
    x_rsc_10_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_10_0_i_biwt : OUT STD_LOGIC;
    x_rsc_10_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_10_0_i_bcwt : IN STD_LOGIC;
    x_rsc_10_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_10_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_10_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_10_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_10_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_10_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_10_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_10_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_10_0_i_bdwt <= x_rsc_10_0_i_oswt AND core_wen;
  x_rsc_10_0_i_biwt <= x_rsc_10_0_i_ogwt AND x_rsc_10_0_i_s_rrdy;
  x_rsc_10_0_i_ogwt <= x_rsc_10_0_i_oswt AND (NOT x_rsc_10_0_i_bcwt);
  x_rsc_10_0_i_s_re_core_sct <= x_rsc_10_0_i_ogwt;
  x_rsc_10_0_i_bdwt_2 <= x_rsc_10_0_i_oswt_1 AND core_wen;
  x_rsc_10_0_i_biwt_1 <= x_rsc_10_0_i_ogwt_1 AND x_rsc_10_0_i_s_wrdy;
  x_rsc_10_0_i_ogwt_1 <= x_rsc_10_0_i_oswt_1 AND (NOT x_rsc_10_0_i_bcwt_1);
  x_rsc_10_0_i_s_we_core_sct <= x_rsc_10_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_9_0_i_oswt : IN STD_LOGIC;
    x_rsc_9_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_9_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_9_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_9_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_9_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_9_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_i_biwt : IN STD_LOGIC;
    x_rsc_9_0_i_bdwt : IN STD_LOGIC;
    x_rsc_9_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_9_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_9_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_9_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_9_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_9_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_9_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_9_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_9_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_9_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_9_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_9_0_i_bcwt <= x_rsc_9_0_i_bcwt_drv;
  x_rsc_9_0_i_bcwt_1 <= x_rsc_9_0_i_bcwt_1_drv;

  x_rsc_9_0_i_wen_comp <= (NOT x_rsc_9_0_i_oswt) OR x_rsc_9_0_i_biwt OR x_rsc_9_0_i_bcwt_drv;
  x_rsc_9_0_i_wen_comp_1 <= (NOT x_rsc_9_0_i_oswt_1) OR x_rsc_9_0_i_biwt_1 OR x_rsc_9_0_i_bcwt_1_drv;
  x_rsc_9_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_9_0_i_s_raddr_core,
      x_rsc_9_0_i_s_raddr_core_sct);
  x_rsc_9_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_9_0_i_s_waddr_core,
      x_rsc_9_0_i_s_waddr_core_sct);
  x_rsc_9_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_9_0_i_s_din, x_rsc_9_0_i_s_din_bfwt,
      x_rsc_9_0_i_bcwt_drv);
  x_rsc_9_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_9_0_i_s_dout_core, x_rsc_9_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_9_0_i_bcwt_drv <= '0';
        x_rsc_9_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_9_0_i_bcwt_drv <= NOT((NOT(x_rsc_9_0_i_bcwt_drv OR x_rsc_9_0_i_biwt))
            OR x_rsc_9_0_i_bdwt);
        x_rsc_9_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_9_0_i_bcwt_1_drv OR x_rsc_9_0_i_biwt_1))
            OR x_rsc_9_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_9_0_i_biwt = '1' ) THEN
        x_rsc_9_0_i_s_din_bfwt <= x_rsc_9_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_9_0_i_oswt : IN STD_LOGIC;
    x_rsc_9_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_9_0_i_biwt : OUT STD_LOGIC;
    x_rsc_9_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_9_0_i_bcwt : IN STD_LOGIC;
    x_rsc_9_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_9_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_9_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_9_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_9_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_9_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_9_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_9_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_9_0_i_bdwt <= x_rsc_9_0_i_oswt AND core_wen;
  x_rsc_9_0_i_biwt <= x_rsc_9_0_i_ogwt AND x_rsc_9_0_i_s_rrdy;
  x_rsc_9_0_i_ogwt <= x_rsc_9_0_i_oswt AND (NOT x_rsc_9_0_i_bcwt);
  x_rsc_9_0_i_s_re_core_sct <= x_rsc_9_0_i_ogwt;
  x_rsc_9_0_i_bdwt_2 <= x_rsc_9_0_i_oswt_1 AND core_wen;
  x_rsc_9_0_i_biwt_1 <= x_rsc_9_0_i_ogwt_1 AND x_rsc_9_0_i_s_wrdy;
  x_rsc_9_0_i_ogwt_1 <= x_rsc_9_0_i_oswt_1 AND (NOT x_rsc_9_0_i_bcwt_1);
  x_rsc_9_0_i_s_we_core_sct <= x_rsc_9_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_8_0_i_oswt : IN STD_LOGIC;
    x_rsc_8_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_8_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_8_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_8_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_8_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_8_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_i_biwt : IN STD_LOGIC;
    x_rsc_8_0_i_bdwt : IN STD_LOGIC;
    x_rsc_8_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_8_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_8_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_8_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_8_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_8_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_8_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_8_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_8_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_8_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_8_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_8_0_i_bcwt <= x_rsc_8_0_i_bcwt_drv;
  x_rsc_8_0_i_bcwt_1 <= x_rsc_8_0_i_bcwt_1_drv;

  x_rsc_8_0_i_wen_comp <= (NOT x_rsc_8_0_i_oswt) OR x_rsc_8_0_i_biwt OR x_rsc_8_0_i_bcwt_drv;
  x_rsc_8_0_i_wen_comp_1 <= (NOT x_rsc_8_0_i_oswt_1) OR x_rsc_8_0_i_biwt_1 OR x_rsc_8_0_i_bcwt_1_drv;
  x_rsc_8_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_8_0_i_s_raddr_core,
      x_rsc_8_0_i_s_raddr_core_sct);
  x_rsc_8_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_8_0_i_s_waddr_core,
      x_rsc_8_0_i_s_waddr_core_sct);
  x_rsc_8_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_8_0_i_s_din, x_rsc_8_0_i_s_din_bfwt,
      x_rsc_8_0_i_bcwt_drv);
  x_rsc_8_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_8_0_i_s_dout_core, x_rsc_8_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_8_0_i_bcwt_drv <= '0';
        x_rsc_8_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_8_0_i_bcwt_drv <= NOT((NOT(x_rsc_8_0_i_bcwt_drv OR x_rsc_8_0_i_biwt))
            OR x_rsc_8_0_i_bdwt);
        x_rsc_8_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_8_0_i_bcwt_1_drv OR x_rsc_8_0_i_biwt_1))
            OR x_rsc_8_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_8_0_i_biwt = '1' ) THEN
        x_rsc_8_0_i_s_din_bfwt <= x_rsc_8_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_8_0_i_oswt : IN STD_LOGIC;
    x_rsc_8_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_8_0_i_biwt : OUT STD_LOGIC;
    x_rsc_8_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_8_0_i_bcwt : IN STD_LOGIC;
    x_rsc_8_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_8_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_8_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_8_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_8_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_8_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_8_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_8_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_8_0_i_bdwt <= x_rsc_8_0_i_oswt AND core_wen;
  x_rsc_8_0_i_biwt <= x_rsc_8_0_i_ogwt AND x_rsc_8_0_i_s_rrdy;
  x_rsc_8_0_i_ogwt <= x_rsc_8_0_i_oswt AND (NOT x_rsc_8_0_i_bcwt);
  x_rsc_8_0_i_s_re_core_sct <= x_rsc_8_0_i_ogwt;
  x_rsc_8_0_i_bdwt_2 <= x_rsc_8_0_i_oswt_1 AND core_wen;
  x_rsc_8_0_i_biwt_1 <= x_rsc_8_0_i_ogwt_1 AND x_rsc_8_0_i_s_wrdy;
  x_rsc_8_0_i_ogwt_1 <= x_rsc_8_0_i_oswt_1 AND (NOT x_rsc_8_0_i_bcwt_1);
  x_rsc_8_0_i_s_we_core_sct <= x_rsc_8_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_7_0_i_oswt : IN STD_LOGIC;
    x_rsc_7_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_7_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_7_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_7_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_7_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_7_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_i_biwt : IN STD_LOGIC;
    x_rsc_7_0_i_bdwt : IN STD_LOGIC;
    x_rsc_7_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_7_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_7_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_7_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_7_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_7_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_7_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_7_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_7_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_7_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_7_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_7_0_i_bcwt <= x_rsc_7_0_i_bcwt_drv;
  x_rsc_7_0_i_bcwt_1 <= x_rsc_7_0_i_bcwt_1_drv;

  x_rsc_7_0_i_wen_comp <= (NOT x_rsc_7_0_i_oswt) OR x_rsc_7_0_i_biwt OR x_rsc_7_0_i_bcwt_drv;
  x_rsc_7_0_i_wen_comp_1 <= (NOT x_rsc_7_0_i_oswt_1) OR x_rsc_7_0_i_biwt_1 OR x_rsc_7_0_i_bcwt_1_drv;
  x_rsc_7_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_7_0_i_s_raddr_core,
      x_rsc_7_0_i_s_raddr_core_sct);
  x_rsc_7_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_7_0_i_s_waddr_core,
      x_rsc_7_0_i_s_waddr_core_sct);
  x_rsc_7_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_7_0_i_s_din, x_rsc_7_0_i_s_din_bfwt,
      x_rsc_7_0_i_bcwt_drv);
  x_rsc_7_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_7_0_i_s_dout_core, x_rsc_7_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_7_0_i_bcwt_drv <= '0';
        x_rsc_7_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_7_0_i_bcwt_drv <= NOT((NOT(x_rsc_7_0_i_bcwt_drv OR x_rsc_7_0_i_biwt))
            OR x_rsc_7_0_i_bdwt);
        x_rsc_7_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_7_0_i_bcwt_1_drv OR x_rsc_7_0_i_biwt_1))
            OR x_rsc_7_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_7_0_i_biwt = '1' ) THEN
        x_rsc_7_0_i_s_din_bfwt <= x_rsc_7_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_7_0_i_oswt : IN STD_LOGIC;
    x_rsc_7_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_7_0_i_biwt : OUT STD_LOGIC;
    x_rsc_7_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_7_0_i_bcwt : IN STD_LOGIC;
    x_rsc_7_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_7_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_7_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_7_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_7_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_7_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_7_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_7_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_7_0_i_bdwt <= x_rsc_7_0_i_oswt AND core_wen;
  x_rsc_7_0_i_biwt <= x_rsc_7_0_i_ogwt AND x_rsc_7_0_i_s_rrdy;
  x_rsc_7_0_i_ogwt <= x_rsc_7_0_i_oswt AND (NOT x_rsc_7_0_i_bcwt);
  x_rsc_7_0_i_s_re_core_sct <= x_rsc_7_0_i_ogwt;
  x_rsc_7_0_i_bdwt_2 <= x_rsc_7_0_i_oswt_1 AND core_wen;
  x_rsc_7_0_i_biwt_1 <= x_rsc_7_0_i_ogwt_1 AND x_rsc_7_0_i_s_wrdy;
  x_rsc_7_0_i_ogwt_1 <= x_rsc_7_0_i_oswt_1 AND (NOT x_rsc_7_0_i_bcwt_1);
  x_rsc_7_0_i_s_we_core_sct <= x_rsc_7_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_6_0_i_oswt : IN STD_LOGIC;
    x_rsc_6_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_6_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_6_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_6_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_6_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_6_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_i_biwt : IN STD_LOGIC;
    x_rsc_6_0_i_bdwt : IN STD_LOGIC;
    x_rsc_6_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_6_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_6_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_6_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_6_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_6_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_6_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_6_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_6_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_6_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_6_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_6_0_i_bcwt <= x_rsc_6_0_i_bcwt_drv;
  x_rsc_6_0_i_bcwt_1 <= x_rsc_6_0_i_bcwt_1_drv;

  x_rsc_6_0_i_wen_comp <= (NOT x_rsc_6_0_i_oswt) OR x_rsc_6_0_i_biwt OR x_rsc_6_0_i_bcwt_drv;
  x_rsc_6_0_i_wen_comp_1 <= (NOT x_rsc_6_0_i_oswt_1) OR x_rsc_6_0_i_biwt_1 OR x_rsc_6_0_i_bcwt_1_drv;
  x_rsc_6_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_6_0_i_s_raddr_core,
      x_rsc_6_0_i_s_raddr_core_sct);
  x_rsc_6_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_6_0_i_s_waddr_core,
      x_rsc_6_0_i_s_waddr_core_sct);
  x_rsc_6_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_6_0_i_s_din, x_rsc_6_0_i_s_din_bfwt,
      x_rsc_6_0_i_bcwt_drv);
  x_rsc_6_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_6_0_i_s_dout_core, x_rsc_6_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_6_0_i_bcwt_drv <= '0';
        x_rsc_6_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_6_0_i_bcwt_drv <= NOT((NOT(x_rsc_6_0_i_bcwt_drv OR x_rsc_6_0_i_biwt))
            OR x_rsc_6_0_i_bdwt);
        x_rsc_6_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_6_0_i_bcwt_1_drv OR x_rsc_6_0_i_biwt_1))
            OR x_rsc_6_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_6_0_i_biwt = '1' ) THEN
        x_rsc_6_0_i_s_din_bfwt <= x_rsc_6_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_6_0_i_oswt : IN STD_LOGIC;
    x_rsc_6_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_6_0_i_biwt : OUT STD_LOGIC;
    x_rsc_6_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_6_0_i_bcwt : IN STD_LOGIC;
    x_rsc_6_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_6_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_6_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_6_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_6_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_6_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_6_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_6_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_6_0_i_bdwt <= x_rsc_6_0_i_oswt AND core_wen;
  x_rsc_6_0_i_biwt <= x_rsc_6_0_i_ogwt AND x_rsc_6_0_i_s_rrdy;
  x_rsc_6_0_i_ogwt <= x_rsc_6_0_i_oswt AND (NOT x_rsc_6_0_i_bcwt);
  x_rsc_6_0_i_s_re_core_sct <= x_rsc_6_0_i_ogwt;
  x_rsc_6_0_i_bdwt_2 <= x_rsc_6_0_i_oswt_1 AND core_wen;
  x_rsc_6_0_i_biwt_1 <= x_rsc_6_0_i_ogwt_1 AND x_rsc_6_0_i_s_wrdy;
  x_rsc_6_0_i_ogwt_1 <= x_rsc_6_0_i_oswt_1 AND (NOT x_rsc_6_0_i_bcwt_1);
  x_rsc_6_0_i_s_we_core_sct <= x_rsc_6_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_5_0_i_oswt : IN STD_LOGIC;
    x_rsc_5_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_5_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_5_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_5_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_5_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_5_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_i_biwt : IN STD_LOGIC;
    x_rsc_5_0_i_bdwt : IN STD_LOGIC;
    x_rsc_5_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_5_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_5_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_5_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_5_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_5_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_5_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_5_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_5_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_5_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_5_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_5_0_i_bcwt <= x_rsc_5_0_i_bcwt_drv;
  x_rsc_5_0_i_bcwt_1 <= x_rsc_5_0_i_bcwt_1_drv;

  x_rsc_5_0_i_wen_comp <= (NOT x_rsc_5_0_i_oswt) OR x_rsc_5_0_i_biwt OR x_rsc_5_0_i_bcwt_drv;
  x_rsc_5_0_i_wen_comp_1 <= (NOT x_rsc_5_0_i_oswt_1) OR x_rsc_5_0_i_biwt_1 OR x_rsc_5_0_i_bcwt_1_drv;
  x_rsc_5_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_5_0_i_s_raddr_core,
      x_rsc_5_0_i_s_raddr_core_sct);
  x_rsc_5_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_5_0_i_s_waddr_core,
      x_rsc_5_0_i_s_waddr_core_sct);
  x_rsc_5_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_5_0_i_s_din, x_rsc_5_0_i_s_din_bfwt,
      x_rsc_5_0_i_bcwt_drv);
  x_rsc_5_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_5_0_i_s_dout_core, x_rsc_5_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_5_0_i_bcwt_drv <= '0';
        x_rsc_5_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_5_0_i_bcwt_drv <= NOT((NOT(x_rsc_5_0_i_bcwt_drv OR x_rsc_5_0_i_biwt))
            OR x_rsc_5_0_i_bdwt);
        x_rsc_5_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_5_0_i_bcwt_1_drv OR x_rsc_5_0_i_biwt_1))
            OR x_rsc_5_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_5_0_i_biwt = '1' ) THEN
        x_rsc_5_0_i_s_din_bfwt <= x_rsc_5_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_5_0_i_oswt : IN STD_LOGIC;
    x_rsc_5_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_5_0_i_biwt : OUT STD_LOGIC;
    x_rsc_5_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_5_0_i_bcwt : IN STD_LOGIC;
    x_rsc_5_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_5_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_5_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_5_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_5_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_5_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_5_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_5_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_5_0_i_bdwt <= x_rsc_5_0_i_oswt AND core_wen;
  x_rsc_5_0_i_biwt <= x_rsc_5_0_i_ogwt AND x_rsc_5_0_i_s_rrdy;
  x_rsc_5_0_i_ogwt <= x_rsc_5_0_i_oswt AND (NOT x_rsc_5_0_i_bcwt);
  x_rsc_5_0_i_s_re_core_sct <= x_rsc_5_0_i_ogwt;
  x_rsc_5_0_i_bdwt_2 <= x_rsc_5_0_i_oswt_1 AND core_wen;
  x_rsc_5_0_i_biwt_1 <= x_rsc_5_0_i_ogwt_1 AND x_rsc_5_0_i_s_wrdy;
  x_rsc_5_0_i_ogwt_1 <= x_rsc_5_0_i_oswt_1 AND (NOT x_rsc_5_0_i_bcwt_1);
  x_rsc_5_0_i_s_we_core_sct <= x_rsc_5_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_4_0_i_oswt : IN STD_LOGIC;
    x_rsc_4_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_4_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_4_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_4_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_4_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_4_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_i_biwt : IN STD_LOGIC;
    x_rsc_4_0_i_bdwt : IN STD_LOGIC;
    x_rsc_4_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_4_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_4_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_4_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_4_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_4_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_4_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_4_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_4_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_4_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_4_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_4_0_i_bcwt <= x_rsc_4_0_i_bcwt_drv;
  x_rsc_4_0_i_bcwt_1 <= x_rsc_4_0_i_bcwt_1_drv;

  x_rsc_4_0_i_wen_comp <= (NOT x_rsc_4_0_i_oswt) OR x_rsc_4_0_i_biwt OR x_rsc_4_0_i_bcwt_drv;
  x_rsc_4_0_i_wen_comp_1 <= (NOT x_rsc_4_0_i_oswt_1) OR x_rsc_4_0_i_biwt_1 OR x_rsc_4_0_i_bcwt_1_drv;
  x_rsc_4_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_4_0_i_s_raddr_core,
      x_rsc_4_0_i_s_raddr_core_sct);
  x_rsc_4_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_4_0_i_s_waddr_core,
      x_rsc_4_0_i_s_waddr_core_sct);
  x_rsc_4_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_4_0_i_s_din, x_rsc_4_0_i_s_din_bfwt,
      x_rsc_4_0_i_bcwt_drv);
  x_rsc_4_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_4_0_i_s_dout_core, x_rsc_4_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_4_0_i_bcwt_drv <= '0';
        x_rsc_4_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_4_0_i_bcwt_drv <= NOT((NOT(x_rsc_4_0_i_bcwt_drv OR x_rsc_4_0_i_biwt))
            OR x_rsc_4_0_i_bdwt);
        x_rsc_4_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_4_0_i_bcwt_1_drv OR x_rsc_4_0_i_biwt_1))
            OR x_rsc_4_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_4_0_i_biwt = '1' ) THEN
        x_rsc_4_0_i_s_din_bfwt <= x_rsc_4_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_4_0_i_oswt : IN STD_LOGIC;
    x_rsc_4_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_4_0_i_biwt : OUT STD_LOGIC;
    x_rsc_4_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_4_0_i_bcwt : IN STD_LOGIC;
    x_rsc_4_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_4_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_4_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_4_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_4_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_4_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_4_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_4_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_4_0_i_bdwt <= x_rsc_4_0_i_oswt AND core_wen;
  x_rsc_4_0_i_biwt <= x_rsc_4_0_i_ogwt AND x_rsc_4_0_i_s_rrdy;
  x_rsc_4_0_i_ogwt <= x_rsc_4_0_i_oswt AND (NOT x_rsc_4_0_i_bcwt);
  x_rsc_4_0_i_s_re_core_sct <= x_rsc_4_0_i_ogwt;
  x_rsc_4_0_i_bdwt_2 <= x_rsc_4_0_i_oswt_1 AND core_wen;
  x_rsc_4_0_i_biwt_1 <= x_rsc_4_0_i_ogwt_1 AND x_rsc_4_0_i_s_wrdy;
  x_rsc_4_0_i_ogwt_1 <= x_rsc_4_0_i_oswt_1 AND (NOT x_rsc_4_0_i_bcwt_1);
  x_rsc_4_0_i_s_we_core_sct <= x_rsc_4_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_3_0_i_oswt : IN STD_LOGIC;
    x_rsc_3_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_3_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_3_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_3_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_3_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_3_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_i_biwt : IN STD_LOGIC;
    x_rsc_3_0_i_bdwt : IN STD_LOGIC;
    x_rsc_3_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_3_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_3_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_3_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_3_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_3_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_3_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_3_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_3_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_3_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_3_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_3_0_i_bcwt <= x_rsc_3_0_i_bcwt_drv;
  x_rsc_3_0_i_bcwt_1 <= x_rsc_3_0_i_bcwt_1_drv;

  x_rsc_3_0_i_wen_comp <= (NOT x_rsc_3_0_i_oswt) OR x_rsc_3_0_i_biwt OR x_rsc_3_0_i_bcwt_drv;
  x_rsc_3_0_i_wen_comp_1 <= (NOT x_rsc_3_0_i_oswt_1) OR x_rsc_3_0_i_biwt_1 OR x_rsc_3_0_i_bcwt_1_drv;
  x_rsc_3_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_3_0_i_s_raddr_core,
      x_rsc_3_0_i_s_raddr_core_sct);
  x_rsc_3_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_3_0_i_s_waddr_core,
      x_rsc_3_0_i_s_waddr_core_sct);
  x_rsc_3_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_3_0_i_s_din, x_rsc_3_0_i_s_din_bfwt,
      x_rsc_3_0_i_bcwt_drv);
  x_rsc_3_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_3_0_i_s_dout_core, x_rsc_3_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_3_0_i_bcwt_drv <= '0';
        x_rsc_3_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_3_0_i_bcwt_drv <= NOT((NOT(x_rsc_3_0_i_bcwt_drv OR x_rsc_3_0_i_biwt))
            OR x_rsc_3_0_i_bdwt);
        x_rsc_3_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_3_0_i_bcwt_1_drv OR x_rsc_3_0_i_biwt_1))
            OR x_rsc_3_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_3_0_i_biwt = '1' ) THEN
        x_rsc_3_0_i_s_din_bfwt <= x_rsc_3_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_3_0_i_oswt : IN STD_LOGIC;
    x_rsc_3_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_3_0_i_biwt : OUT STD_LOGIC;
    x_rsc_3_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_3_0_i_bcwt : IN STD_LOGIC;
    x_rsc_3_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_3_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_3_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_3_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_3_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_3_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_3_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_3_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_3_0_i_bdwt <= x_rsc_3_0_i_oswt AND core_wen;
  x_rsc_3_0_i_biwt <= x_rsc_3_0_i_ogwt AND x_rsc_3_0_i_s_rrdy;
  x_rsc_3_0_i_ogwt <= x_rsc_3_0_i_oswt AND (NOT x_rsc_3_0_i_bcwt);
  x_rsc_3_0_i_s_re_core_sct <= x_rsc_3_0_i_ogwt;
  x_rsc_3_0_i_bdwt_2 <= x_rsc_3_0_i_oswt_1 AND core_wen;
  x_rsc_3_0_i_biwt_1 <= x_rsc_3_0_i_ogwt_1 AND x_rsc_3_0_i_s_wrdy;
  x_rsc_3_0_i_ogwt_1 <= x_rsc_3_0_i_oswt_1 AND (NOT x_rsc_3_0_i_bcwt_1);
  x_rsc_3_0_i_s_we_core_sct <= x_rsc_3_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_2_0_i_oswt : IN STD_LOGIC;
    x_rsc_2_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_2_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_2_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_2_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_2_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_2_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_i_biwt : IN STD_LOGIC;
    x_rsc_2_0_i_bdwt : IN STD_LOGIC;
    x_rsc_2_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_2_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_2_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_2_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_2_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_2_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_2_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_2_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_2_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_2_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_2_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_2_0_i_bcwt <= x_rsc_2_0_i_bcwt_drv;
  x_rsc_2_0_i_bcwt_1 <= x_rsc_2_0_i_bcwt_1_drv;

  x_rsc_2_0_i_wen_comp <= (NOT x_rsc_2_0_i_oswt) OR x_rsc_2_0_i_biwt OR x_rsc_2_0_i_bcwt_drv;
  x_rsc_2_0_i_wen_comp_1 <= (NOT x_rsc_2_0_i_oswt_1) OR x_rsc_2_0_i_biwt_1 OR x_rsc_2_0_i_bcwt_1_drv;
  x_rsc_2_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_2_0_i_s_raddr_core,
      x_rsc_2_0_i_s_raddr_core_sct);
  x_rsc_2_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_2_0_i_s_waddr_core,
      x_rsc_2_0_i_s_waddr_core_sct);
  x_rsc_2_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_2_0_i_s_din, x_rsc_2_0_i_s_din_bfwt,
      x_rsc_2_0_i_bcwt_drv);
  x_rsc_2_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_2_0_i_s_dout_core, x_rsc_2_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_2_0_i_bcwt_drv <= '0';
        x_rsc_2_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_2_0_i_bcwt_drv <= NOT((NOT(x_rsc_2_0_i_bcwt_drv OR x_rsc_2_0_i_biwt))
            OR x_rsc_2_0_i_bdwt);
        x_rsc_2_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_2_0_i_bcwt_1_drv OR x_rsc_2_0_i_biwt_1))
            OR x_rsc_2_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_2_0_i_biwt = '1' ) THEN
        x_rsc_2_0_i_s_din_bfwt <= x_rsc_2_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_2_0_i_oswt : IN STD_LOGIC;
    x_rsc_2_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_2_0_i_biwt : OUT STD_LOGIC;
    x_rsc_2_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_2_0_i_bcwt : IN STD_LOGIC;
    x_rsc_2_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_2_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_2_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_2_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_2_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_2_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_2_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_2_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_2_0_i_bdwt <= x_rsc_2_0_i_oswt AND core_wen;
  x_rsc_2_0_i_biwt <= x_rsc_2_0_i_ogwt AND x_rsc_2_0_i_s_rrdy;
  x_rsc_2_0_i_ogwt <= x_rsc_2_0_i_oswt AND (NOT x_rsc_2_0_i_bcwt);
  x_rsc_2_0_i_s_re_core_sct <= x_rsc_2_0_i_ogwt;
  x_rsc_2_0_i_bdwt_2 <= x_rsc_2_0_i_oswt_1 AND core_wen;
  x_rsc_2_0_i_biwt_1 <= x_rsc_2_0_i_ogwt_1 AND x_rsc_2_0_i_s_wrdy;
  x_rsc_2_0_i_ogwt_1 <= x_rsc_2_0_i_oswt_1 AND (NOT x_rsc_2_0_i_bcwt_1);
  x_rsc_2_0_i_s_we_core_sct <= x_rsc_2_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_1_0_i_oswt : IN STD_LOGIC;
    x_rsc_1_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_1_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_1_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_1_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_1_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_i_biwt : IN STD_LOGIC;
    x_rsc_1_0_i_bdwt : IN STD_LOGIC;
    x_rsc_1_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_1_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_1_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_1_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_1_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_1_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_1_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_1_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_1_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_1_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_1_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_1_0_i_bcwt <= x_rsc_1_0_i_bcwt_drv;
  x_rsc_1_0_i_bcwt_1 <= x_rsc_1_0_i_bcwt_1_drv;

  x_rsc_1_0_i_wen_comp <= (NOT x_rsc_1_0_i_oswt) OR x_rsc_1_0_i_biwt OR x_rsc_1_0_i_bcwt_drv;
  x_rsc_1_0_i_wen_comp_1 <= (NOT x_rsc_1_0_i_oswt_1) OR x_rsc_1_0_i_biwt_1 OR x_rsc_1_0_i_bcwt_1_drv;
  x_rsc_1_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_1_0_i_s_raddr_core,
      x_rsc_1_0_i_s_raddr_core_sct);
  x_rsc_1_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_1_0_i_s_waddr_core,
      x_rsc_1_0_i_s_waddr_core_sct);
  x_rsc_1_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_1_0_i_s_din, x_rsc_1_0_i_s_din_bfwt,
      x_rsc_1_0_i_bcwt_drv);
  x_rsc_1_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_1_0_i_s_dout_core, x_rsc_1_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_1_0_i_bcwt_drv <= '0';
        x_rsc_1_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_1_0_i_bcwt_drv <= NOT((NOT(x_rsc_1_0_i_bcwt_drv OR x_rsc_1_0_i_biwt))
            OR x_rsc_1_0_i_bdwt);
        x_rsc_1_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_1_0_i_bcwt_1_drv OR x_rsc_1_0_i_biwt_1))
            OR x_rsc_1_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_1_0_i_biwt = '1' ) THEN
        x_rsc_1_0_i_s_din_bfwt <= x_rsc_1_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_1_0_i_oswt : IN STD_LOGIC;
    x_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_1_0_i_biwt : OUT STD_LOGIC;
    x_rsc_1_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_1_0_i_bcwt : IN STD_LOGIC;
    x_rsc_1_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_1_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_1_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_1_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_1_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_1_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_1_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_1_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_1_0_i_bdwt <= x_rsc_1_0_i_oswt AND core_wen;
  x_rsc_1_0_i_biwt <= x_rsc_1_0_i_ogwt AND x_rsc_1_0_i_s_rrdy;
  x_rsc_1_0_i_ogwt <= x_rsc_1_0_i_oswt AND (NOT x_rsc_1_0_i_bcwt);
  x_rsc_1_0_i_s_re_core_sct <= x_rsc_1_0_i_ogwt;
  x_rsc_1_0_i_bdwt_2 <= x_rsc_1_0_i_oswt_1 AND core_wen;
  x_rsc_1_0_i_biwt_1 <= x_rsc_1_0_i_ogwt_1 AND x_rsc_1_0_i_s_wrdy;
  x_rsc_1_0_i_ogwt_1 <= x_rsc_1_0_i_oswt_1 AND (NOT x_rsc_1_0_i_bcwt_1);
  x_rsc_1_0_i_s_we_core_sct <= x_rsc_1_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_0_0_i_oswt : IN STD_LOGIC;
    x_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_0_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_0_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_i_biwt : IN STD_LOGIC;
    x_rsc_0_0_i_bdwt : IN STD_LOGIC;
    x_rsc_0_0_i_bcwt : OUT STD_LOGIC;
    x_rsc_0_0_i_biwt_1 : IN STD_LOGIC;
    x_rsc_0_0_i_bdwt_2 : IN STD_LOGIC;
    x_rsc_0_0_i_bcwt_1 : OUT STD_LOGIC;
    x_rsc_0_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_0_0_i_s_raddr_core_sct : IN STD_LOGIC;
    x_rsc_0_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_0_0_i_s_waddr_core_sct : IN STD_LOGIC;
    x_rsc_0_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp;

ARCHITECTURE v14 OF hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL x_rsc_0_0_i_bcwt_drv : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_bcwt_1_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL x_rsc_0_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  x_rsc_0_0_i_bcwt <= x_rsc_0_0_i_bcwt_drv;
  x_rsc_0_0_i_bcwt_1 <= x_rsc_0_0_i_bcwt_1_drv;

  x_rsc_0_0_i_wen_comp <= (NOT x_rsc_0_0_i_oswt) OR x_rsc_0_0_i_biwt OR x_rsc_0_0_i_bcwt_drv;
  x_rsc_0_0_i_wen_comp_1 <= (NOT x_rsc_0_0_i_oswt_1) OR x_rsc_0_0_i_biwt_1 OR x_rsc_0_0_i_bcwt_1_drv;
  x_rsc_0_0_i_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_0_0_i_s_raddr_core,
      x_rsc_0_0_i_s_raddr_core_sct);
  x_rsc_0_0_i_s_waddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), x_rsc_0_0_i_s_waddr_core,
      x_rsc_0_0_i_s_waddr_core_sct);
  x_rsc_0_0_i_s_din_mxwt <= MUX_v_32_2_2(x_rsc_0_0_i_s_din, x_rsc_0_0_i_s_din_bfwt,
      x_rsc_0_0_i_bcwt_drv);
  x_rsc_0_0_i_s_dout <= MUX_v_32_2_2(STD_LOGIC_VECTOR'("00000000000000000000000000000000"),
      x_rsc_0_0_i_s_dout_core, x_rsc_0_0_i_s_waddr_core_sct);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_rsc_0_0_i_bcwt_drv <= '0';
        x_rsc_0_0_i_bcwt_1_drv <= '0';
      ELSE
        x_rsc_0_0_i_bcwt_drv <= NOT((NOT(x_rsc_0_0_i_bcwt_drv OR x_rsc_0_0_i_biwt))
            OR x_rsc_0_0_i_bdwt);
        x_rsc_0_0_i_bcwt_1_drv <= NOT((NOT(x_rsc_0_0_i_bcwt_1_drv OR x_rsc_0_0_i_biwt_1))
            OR x_rsc_0_0_i_bdwt_2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( x_rsc_0_0_i_biwt = '1' ) THEN
        x_rsc_0_0_i_s_din_bfwt <= x_rsc_0_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    x_rsc_0_0_i_oswt : IN STD_LOGIC;
    x_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_0_0_i_biwt : OUT STD_LOGIC;
    x_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    x_rsc_0_0_i_bcwt : IN STD_LOGIC;
    x_rsc_0_0_i_s_re_core_sct : OUT STD_LOGIC;
    x_rsc_0_0_i_biwt_1 : OUT STD_LOGIC;
    x_rsc_0_0_i_bdwt_2 : OUT STD_LOGIC;
    x_rsc_0_0_i_bcwt_1 : IN STD_LOGIC;
    x_rsc_0_0_i_s_we_core_sct : OUT STD_LOGIC;
    x_rsc_0_0_i_s_rrdy : IN STD_LOGIC;
    x_rsc_0_0_i_s_wrdy : IN STD_LOGIC
  );
END hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_0_0_i_ogwt : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_ogwt_1 : STD_LOGIC;

BEGIN
  x_rsc_0_0_i_bdwt <= x_rsc_0_0_i_oswt AND core_wen;
  x_rsc_0_0_i_biwt <= x_rsc_0_0_i_ogwt AND x_rsc_0_0_i_s_rrdy;
  x_rsc_0_0_i_ogwt <= x_rsc_0_0_i_oswt AND (NOT x_rsc_0_0_i_bcwt);
  x_rsc_0_0_i_s_re_core_sct <= x_rsc_0_0_i_ogwt;
  x_rsc_0_0_i_bdwt_2 <= x_rsc_0_0_i_oswt_1 AND core_wen;
  x_rsc_0_0_i_biwt_1 <= x_rsc_0_0_i_ogwt_1 AND x_rsc_0_0_i_s_wrdy;
  x_rsc_0_0_i_ogwt_1 <= x_rsc_0_0_i_oswt_1 AND (NOT x_rsc_0_0_i_bcwt_1);
  x_rsc_0_0_i_s_we_core_sct <= x_rsc_0_0_i_ogwt_1;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    tw_h_rsci_oswt : IN STD_LOGIC;
    tw_h_rsci_wen_comp : OUT STD_LOGIC;
    tw_h_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    tw_h_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
    tw_h_rsci_biwt : IN STD_LOGIC;
    tw_h_rsci_bdwt : IN STD_LOGIC;
    tw_h_rsci_bcwt : OUT STD_LOGIC;
    tw_h_rsci_s_raddr : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    tw_h_rsci_s_raddr_core_sct : IN STD_LOGIC;
    tw_h_rsci_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp;

ARCHITECTURE v14 OF hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL tw_h_rsci_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL tw_h_rsci_s_din_bfwt_19_0 : STD_LOGIC_VECTOR (19 DOWNTO 0);

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_20_2_2(input_0 : STD_LOGIC_VECTOR(19 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(19 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(19 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  tw_h_rsci_bcwt <= tw_h_rsci_bcwt_drv;

  tw_h_rsci_wen_comp <= (NOT tw_h_rsci_oswt) OR tw_h_rsci_biwt OR tw_h_rsci_bcwt_drv;
  tw_h_rsci_s_raddr <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"), tw_h_rsci_s_raddr_core,
      tw_h_rsci_s_raddr_core_sct);
  tw_h_rsci_s_din_mxwt <= MUX_v_20_2_2((tw_h_rsci_s_din(19 DOWNTO 0)), tw_h_rsci_s_din_bfwt_19_0,
      tw_h_rsci_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        tw_h_rsci_bcwt_drv <= '0';
      ELSE
        tw_h_rsci_bcwt_drv <= NOT((NOT(tw_h_rsci_bcwt_drv OR tw_h_rsci_biwt)) OR
            tw_h_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( tw_h_rsci_biwt = '1' ) THEN
        tw_h_rsci_s_din_bfwt_19_0 <= tw_h_rsci_s_din(19 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    tw_h_rsci_oswt : IN STD_LOGIC;
    tw_h_rsci_biwt : OUT STD_LOGIC;
    tw_h_rsci_bdwt : OUT STD_LOGIC;
    tw_h_rsci_bcwt : IN STD_LOGIC;
    tw_h_rsci_s_re_core_sct : OUT STD_LOGIC;
    tw_h_rsci_s_rrdy : IN STD_LOGIC
  );
END hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL tw_h_rsci_ogwt : STD_LOGIC;

BEGIN
  tw_h_rsci_bdwt <= tw_h_rsci_oswt AND core_wen;
  tw_h_rsci_biwt <= tw_h_rsci_ogwt AND tw_h_rsci_s_rrdy;
  tw_h_rsci_ogwt <= tw_h_rsci_oswt AND (NOT tw_h_rsci_bcwt);
  tw_h_rsci_s_re_core_sct <= tw_h_rsci_ogwt;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_rsci_tw_rsc_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_rsci_tw_rsc_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    tw_rsci_oswt : IN STD_LOGIC;
    tw_rsci_wen_comp : OUT STD_LOGIC;
    tw_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    tw_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
    tw_rsci_biwt : IN STD_LOGIC;
    tw_rsci_bdwt : IN STD_LOGIC;
    tw_rsci_bcwt : OUT STD_LOGIC;
    tw_rsci_s_raddr : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    tw_rsci_s_raddr_core_sct : IN STD_LOGIC;
    tw_rsci_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_tw_rsci_tw_rsc_wait_dp;

ARCHITECTURE v14 OF hybrid_core_tw_rsci_tw_rsc_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL tw_rsci_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL tw_rsci_s_din_bfwt_19_0 : STD_LOGIC_VECTOR (19 DOWNTO 0);

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_20_2_2(input_0 : STD_LOGIC_VECTOR(19 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(19 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(19 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  tw_rsci_bcwt <= tw_rsci_bcwt_drv;

  tw_rsci_wen_comp <= (NOT tw_rsci_oswt) OR tw_rsci_biwt OR tw_rsci_bcwt_drv;
  tw_rsci_s_raddr <= MUX_v_10_2_2(STD_LOGIC_VECTOR'("0000000000"), tw_rsci_s_raddr_core,
      tw_rsci_s_raddr_core_sct);
  tw_rsci_s_din_mxwt <= MUX_v_20_2_2((tw_rsci_s_din(19 DOWNTO 0)), tw_rsci_s_din_bfwt_19_0,
      tw_rsci_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        tw_rsci_bcwt_drv <= '0';
      ELSE
        tw_rsci_bcwt_drv <= NOT((NOT(tw_rsci_bcwt_drv OR tw_rsci_biwt)) OR tw_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( tw_rsci_biwt = '1' ) THEN
        tw_rsci_s_din_bfwt_19_0 <= tw_rsci_s_din(19 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_rsci_tw_rsc_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_rsci_tw_rsc_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    tw_rsci_oswt : IN STD_LOGIC;
    tw_rsci_biwt : OUT STD_LOGIC;
    tw_rsci_bdwt : OUT STD_LOGIC;
    tw_rsci_bcwt : IN STD_LOGIC;
    tw_rsci_s_re_core_sct : OUT STD_LOGIC;
    tw_rsci_s_rrdy : IN STD_LOGIC
  );
END hybrid_core_tw_rsci_tw_rsc_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_tw_rsci_tw_rsc_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL tw_rsci_ogwt : STD_LOGIC;

BEGIN
  tw_rsci_bdwt <= tw_rsci_oswt AND core_wen;
  tw_rsci_biwt <= tw_rsci_ogwt AND tw_rsci_s_rrdy;
  tw_rsci_ogwt <= tw_rsci_oswt AND (NOT tw_rsci_bcwt);
  tw_rsci_s_re_core_sct <= tw_rsci_ogwt;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_revArr_rsci_revArr_rsc_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_revArr_rsci_revArr_rsc_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    revArr_rsci_oswt : IN STD_LOGIC;
    revArr_rsci_wen_comp : OUT STD_LOGIC;
    revArr_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    revArr_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    revArr_rsci_biwt : IN STD_LOGIC;
    revArr_rsci_bdwt : IN STD_LOGIC;
    revArr_rsci_bcwt : OUT STD_LOGIC;
    revArr_rsci_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    revArr_rsci_s_raddr_core_sct : IN STD_LOGIC;
    revArr_rsci_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_revArr_rsci_revArr_rsc_wait_dp;

ARCHITECTURE v14 OF hybrid_core_revArr_rsci_revArr_rsc_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL revArr_rsci_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL revArr_rsci_s_din_bfwt_9_0 : STD_LOGIC_VECTOR (9 DOWNTO 0);

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  revArr_rsci_bcwt <= revArr_rsci_bcwt_drv;

  revArr_rsci_wen_comp <= (NOT revArr_rsci_oswt) OR revArr_rsci_biwt OR revArr_rsci_bcwt_drv;
  revArr_rsci_s_raddr <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), revArr_rsci_s_raddr_core,
      revArr_rsci_s_raddr_core_sct);
  revArr_rsci_s_din_mxwt <= MUX_v_10_2_2((revArr_rsci_s_din(9 DOWNTO 0)), revArr_rsci_s_din_bfwt_9_0,
      revArr_rsci_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        revArr_rsci_bcwt_drv <= '0';
      ELSE
        revArr_rsci_bcwt_drv <= NOT((NOT(revArr_rsci_bcwt_drv OR revArr_rsci_biwt))
            OR revArr_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( revArr_rsci_biwt = '1' ) THEN
        revArr_rsci_s_din_bfwt_9_0 <= revArr_rsci_s_din(9 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    revArr_rsci_oswt : IN STD_LOGIC;
    revArr_rsci_biwt : OUT STD_LOGIC;
    revArr_rsci_bdwt : OUT STD_LOGIC;
    revArr_rsci_bcwt : IN STD_LOGIC;
    revArr_rsci_s_re_core_sct : OUT STD_LOGIC;
    revArr_rsci_s_rrdy : IN STD_LOGIC
  );
END hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL revArr_rsci_ogwt : STD_LOGIC;

BEGIN
  revArr_rsci_bdwt <= revArr_rsci_oswt AND core_wen;
  revArr_rsci_biwt <= revArr_rsci_ogwt AND revArr_rsci_s_rrdy;
  revArr_rsci_ogwt <= revArr_rsci_oswt AND (NOT revArr_rsci_bcwt);
  revArr_rsci_s_re_core_sct <= revArr_rsci_ogwt;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_h_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_h_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsci_biwt : IN STD_LOGIC;
    twiddle_h_rsci_bdwt : IN STD_LOGIC;
    twiddle_h_rsci_adrb_d_core_sct : IN STD_LOGIC
  );
END hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp;

ARCHITECTURE v14 OF hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsci_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsci_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_h_rsci_qb_d_mxwt <= MUX_v_32_2_2(twiddle_h_rsci_qb_d, twiddle_h_rsci_qb_d_bfwt,
      twiddle_h_rsci_bcwt);
  twiddle_h_rsci_adrb_d <= (NOT twiddle_h_rsci_adrb_d_core_sct) & (twiddle_h_rsci_adrb_d_core(3
      DOWNTO 0));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsci_bcwt <= '0';
      ELSE
        twiddle_h_rsci_bcwt <= NOT((NOT(twiddle_h_rsci_bcwt OR twiddle_h_rsci_biwt))
            OR twiddle_h_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsci_biwt = '1' ) THEN
        twiddle_h_rsci_qb_d_bfwt <= twiddle_h_rsci_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsci_oswt : IN STD_LOGIC;
    twiddle_h_rsci_biwt : OUT STD_LOGIC;
    twiddle_h_rsci_bdwt : OUT STD_LOGIC;
    twiddle_h_rsci_adrb_d_core_sct_pff : OUT STD_LOGIC;
    twiddle_h_rsci_oswt_pff : IN STD_LOGIC
  );
END hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl IS
  -- Default Constants

BEGIN
  twiddle_h_rsci_bdwt <= twiddle_h_rsci_oswt AND core_wen;
  twiddle_h_rsci_biwt <= (NOT core_wten) AND twiddle_h_rsci_oswt;
  twiddle_h_rsci_adrb_d_core_sct_pff <= twiddle_h_rsci_oswt_pff AND core_wen;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    xx_rsc_0_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_1_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_2_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_3_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_4_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_5_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_6_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_7_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_8_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_9_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_10_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_11_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_12_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_13_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_14_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_15_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_16_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_17_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_18_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_19_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_20_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_21_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_22_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_23_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_24_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_25_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_26_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_27_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_28_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_29_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_30_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_31_0_cgo_iro : IN STD_LOGIC;
    xx_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_0_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_1_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_2_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_3_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_4_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_5_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_6_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_7_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_8_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_9_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_10_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_11_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_12_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_13_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_14_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_15_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_16_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_17_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_18_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_19_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_20_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_21_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_22_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_23_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_24_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_25_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_26_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_27_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_28_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_29_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_30_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_31_0_cgo_iro : IN STD_LOGIC;
    yy_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
    ensig_cgo_iro : IN STD_LOGIC;
    S34_OUTER_LOOP_for_tf_mul_cmp_z : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    ensig_cgo_iro_1 : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    xx_rsc_0_0_cgo : IN STD_LOGIC;
    xx_rsc_1_0_cgo : IN STD_LOGIC;
    xx_rsc_2_0_cgo : IN STD_LOGIC;
    xx_rsc_3_0_cgo : IN STD_LOGIC;
    xx_rsc_4_0_cgo : IN STD_LOGIC;
    xx_rsc_5_0_cgo : IN STD_LOGIC;
    xx_rsc_6_0_cgo : IN STD_LOGIC;
    xx_rsc_7_0_cgo : IN STD_LOGIC;
    xx_rsc_8_0_cgo : IN STD_LOGIC;
    xx_rsc_9_0_cgo : IN STD_LOGIC;
    xx_rsc_10_0_cgo : IN STD_LOGIC;
    xx_rsc_11_0_cgo : IN STD_LOGIC;
    xx_rsc_12_0_cgo : IN STD_LOGIC;
    xx_rsc_13_0_cgo : IN STD_LOGIC;
    xx_rsc_14_0_cgo : IN STD_LOGIC;
    xx_rsc_15_0_cgo : IN STD_LOGIC;
    xx_rsc_16_0_cgo : IN STD_LOGIC;
    xx_rsc_17_0_cgo : IN STD_LOGIC;
    xx_rsc_18_0_cgo : IN STD_LOGIC;
    xx_rsc_19_0_cgo : IN STD_LOGIC;
    xx_rsc_20_0_cgo : IN STD_LOGIC;
    xx_rsc_21_0_cgo : IN STD_LOGIC;
    xx_rsc_22_0_cgo : IN STD_LOGIC;
    xx_rsc_23_0_cgo : IN STD_LOGIC;
    xx_rsc_24_0_cgo : IN STD_LOGIC;
    xx_rsc_25_0_cgo : IN STD_LOGIC;
    xx_rsc_26_0_cgo : IN STD_LOGIC;
    xx_rsc_27_0_cgo : IN STD_LOGIC;
    xx_rsc_28_0_cgo : IN STD_LOGIC;
    xx_rsc_29_0_cgo : IN STD_LOGIC;
    xx_rsc_30_0_cgo : IN STD_LOGIC;
    xx_rsc_31_0_cgo : IN STD_LOGIC;
    yy_rsc_0_0_cgo : IN STD_LOGIC;
    yy_rsc_1_0_cgo : IN STD_LOGIC;
    yy_rsc_2_0_cgo : IN STD_LOGIC;
    yy_rsc_3_0_cgo : IN STD_LOGIC;
    yy_rsc_4_0_cgo : IN STD_LOGIC;
    yy_rsc_5_0_cgo : IN STD_LOGIC;
    yy_rsc_6_0_cgo : IN STD_LOGIC;
    yy_rsc_7_0_cgo : IN STD_LOGIC;
    yy_rsc_8_0_cgo : IN STD_LOGIC;
    yy_rsc_9_0_cgo : IN STD_LOGIC;
    yy_rsc_10_0_cgo : IN STD_LOGIC;
    yy_rsc_11_0_cgo : IN STD_LOGIC;
    yy_rsc_12_0_cgo : IN STD_LOGIC;
    yy_rsc_13_0_cgo : IN STD_LOGIC;
    yy_rsc_14_0_cgo : IN STD_LOGIC;
    yy_rsc_15_0_cgo : IN STD_LOGIC;
    yy_rsc_16_0_cgo : IN STD_LOGIC;
    yy_rsc_17_0_cgo : IN STD_LOGIC;
    yy_rsc_18_0_cgo : IN STD_LOGIC;
    yy_rsc_19_0_cgo : IN STD_LOGIC;
    yy_rsc_20_0_cgo : IN STD_LOGIC;
    yy_rsc_21_0_cgo : IN STD_LOGIC;
    yy_rsc_22_0_cgo : IN STD_LOGIC;
    yy_rsc_23_0_cgo : IN STD_LOGIC;
    yy_rsc_24_0_cgo : IN STD_LOGIC;
    yy_rsc_25_0_cgo : IN STD_LOGIC;
    yy_rsc_26_0_cgo : IN STD_LOGIC;
    yy_rsc_27_0_cgo : IN STD_LOGIC;
    yy_rsc_28_0_cgo : IN STD_LOGIC;
    yy_rsc_29_0_cgo : IN STD_LOGIC;
    yy_rsc_30_0_cgo : IN STD_LOGIC;
    yy_rsc_31_0_cgo : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    mult_12_z_mul_cmp_en : OUT STD_LOGIC;
    S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    ensig_cgo_1 : IN STD_LOGIC;
    mult_z_mul_cmp_en : OUT STD_LOGIC
  );
END hybrid_core_wait_dp;

ARCHITECTURE v14 OF hybrid_core_wait_dp IS
  -- Default Constants

BEGIN
  xx_rsc_0_0_i_clka_en_d <= core_wen AND (xx_rsc_0_0_cgo OR xx_rsc_0_0_cgo_iro);
  xx_rsc_1_0_i_clka_en_d <= core_wen AND (xx_rsc_1_0_cgo OR xx_rsc_1_0_cgo_iro);
  xx_rsc_2_0_i_clka_en_d <= core_wen AND (xx_rsc_2_0_cgo OR xx_rsc_2_0_cgo_iro);
  xx_rsc_3_0_i_clka_en_d <= core_wen AND (xx_rsc_3_0_cgo OR xx_rsc_3_0_cgo_iro);
  xx_rsc_4_0_i_clka_en_d <= core_wen AND (xx_rsc_4_0_cgo OR xx_rsc_4_0_cgo_iro);
  xx_rsc_5_0_i_clka_en_d <= core_wen AND (xx_rsc_5_0_cgo OR xx_rsc_5_0_cgo_iro);
  xx_rsc_6_0_i_clka_en_d <= core_wen AND (xx_rsc_6_0_cgo OR xx_rsc_6_0_cgo_iro);
  xx_rsc_7_0_i_clka_en_d <= core_wen AND (xx_rsc_7_0_cgo OR xx_rsc_7_0_cgo_iro);
  xx_rsc_8_0_i_clka_en_d <= core_wen AND (xx_rsc_8_0_cgo OR xx_rsc_8_0_cgo_iro);
  xx_rsc_9_0_i_clka_en_d <= core_wen AND (xx_rsc_9_0_cgo OR xx_rsc_9_0_cgo_iro);
  xx_rsc_10_0_i_clka_en_d <= core_wen AND (xx_rsc_10_0_cgo OR xx_rsc_10_0_cgo_iro);
  xx_rsc_11_0_i_clka_en_d <= core_wen AND (xx_rsc_11_0_cgo OR xx_rsc_11_0_cgo_iro);
  xx_rsc_12_0_i_clka_en_d <= core_wen AND (xx_rsc_12_0_cgo OR xx_rsc_12_0_cgo_iro);
  xx_rsc_13_0_i_clka_en_d <= core_wen AND (xx_rsc_13_0_cgo OR xx_rsc_13_0_cgo_iro);
  xx_rsc_14_0_i_clka_en_d <= core_wen AND (xx_rsc_14_0_cgo OR xx_rsc_14_0_cgo_iro);
  xx_rsc_15_0_i_clka_en_d <= core_wen AND (xx_rsc_15_0_cgo OR xx_rsc_15_0_cgo_iro);
  xx_rsc_16_0_i_clka_en_d <= core_wen AND (xx_rsc_16_0_cgo OR xx_rsc_16_0_cgo_iro);
  xx_rsc_17_0_i_clka_en_d <= core_wen AND (xx_rsc_17_0_cgo OR xx_rsc_17_0_cgo_iro);
  xx_rsc_18_0_i_clka_en_d <= core_wen AND (xx_rsc_18_0_cgo OR xx_rsc_18_0_cgo_iro);
  xx_rsc_19_0_i_clka_en_d <= core_wen AND (xx_rsc_19_0_cgo OR xx_rsc_19_0_cgo_iro);
  xx_rsc_20_0_i_clka_en_d <= core_wen AND (xx_rsc_20_0_cgo OR xx_rsc_20_0_cgo_iro);
  xx_rsc_21_0_i_clka_en_d <= core_wen AND (xx_rsc_21_0_cgo OR xx_rsc_21_0_cgo_iro);
  xx_rsc_22_0_i_clka_en_d <= core_wen AND (xx_rsc_22_0_cgo OR xx_rsc_22_0_cgo_iro);
  xx_rsc_23_0_i_clka_en_d <= core_wen AND (xx_rsc_23_0_cgo OR xx_rsc_23_0_cgo_iro);
  xx_rsc_24_0_i_clka_en_d <= core_wen AND (xx_rsc_24_0_cgo OR xx_rsc_24_0_cgo_iro);
  xx_rsc_25_0_i_clka_en_d <= core_wen AND (xx_rsc_25_0_cgo OR xx_rsc_25_0_cgo_iro);
  xx_rsc_26_0_i_clka_en_d <= core_wen AND (xx_rsc_26_0_cgo OR xx_rsc_26_0_cgo_iro);
  xx_rsc_27_0_i_clka_en_d <= core_wen AND (xx_rsc_27_0_cgo OR xx_rsc_27_0_cgo_iro);
  xx_rsc_28_0_i_clka_en_d <= core_wen AND (xx_rsc_28_0_cgo OR xx_rsc_28_0_cgo_iro);
  xx_rsc_29_0_i_clka_en_d <= core_wen AND (xx_rsc_29_0_cgo OR xx_rsc_29_0_cgo_iro);
  xx_rsc_30_0_i_clka_en_d <= core_wen AND (xx_rsc_30_0_cgo OR xx_rsc_30_0_cgo_iro);
  xx_rsc_31_0_i_clka_en_d <= core_wen AND (xx_rsc_31_0_cgo OR xx_rsc_31_0_cgo_iro);
  yy_rsc_0_0_i_clka_en_d <= core_wen AND (yy_rsc_0_0_cgo OR yy_rsc_0_0_cgo_iro);
  yy_rsc_1_0_i_clka_en_d <= core_wen AND (yy_rsc_1_0_cgo OR yy_rsc_1_0_cgo_iro);
  yy_rsc_2_0_i_clka_en_d <= core_wen AND (yy_rsc_2_0_cgo OR yy_rsc_2_0_cgo_iro);
  yy_rsc_3_0_i_clka_en_d <= core_wen AND (yy_rsc_3_0_cgo OR yy_rsc_3_0_cgo_iro);
  yy_rsc_4_0_i_clka_en_d <= core_wen AND (yy_rsc_4_0_cgo OR yy_rsc_4_0_cgo_iro);
  yy_rsc_5_0_i_clka_en_d <= core_wen AND (yy_rsc_5_0_cgo OR yy_rsc_5_0_cgo_iro);
  yy_rsc_6_0_i_clka_en_d <= core_wen AND (yy_rsc_6_0_cgo OR yy_rsc_6_0_cgo_iro);
  yy_rsc_7_0_i_clka_en_d <= core_wen AND (yy_rsc_7_0_cgo OR yy_rsc_7_0_cgo_iro);
  yy_rsc_8_0_i_clka_en_d <= core_wen AND (yy_rsc_8_0_cgo OR yy_rsc_8_0_cgo_iro);
  yy_rsc_9_0_i_clka_en_d <= core_wen AND (yy_rsc_9_0_cgo OR yy_rsc_9_0_cgo_iro);
  yy_rsc_10_0_i_clka_en_d <= core_wen AND (yy_rsc_10_0_cgo OR yy_rsc_10_0_cgo_iro);
  yy_rsc_11_0_i_clka_en_d <= core_wen AND (yy_rsc_11_0_cgo OR yy_rsc_11_0_cgo_iro);
  yy_rsc_12_0_i_clka_en_d <= core_wen AND (yy_rsc_12_0_cgo OR yy_rsc_12_0_cgo_iro);
  yy_rsc_13_0_i_clka_en_d <= core_wen AND (yy_rsc_13_0_cgo OR yy_rsc_13_0_cgo_iro);
  yy_rsc_14_0_i_clka_en_d <= core_wen AND (yy_rsc_14_0_cgo OR yy_rsc_14_0_cgo_iro);
  yy_rsc_15_0_i_clka_en_d <= core_wen AND (yy_rsc_15_0_cgo OR yy_rsc_15_0_cgo_iro);
  yy_rsc_16_0_i_clka_en_d <= core_wen AND (yy_rsc_16_0_cgo OR yy_rsc_16_0_cgo_iro);
  yy_rsc_17_0_i_clka_en_d <= core_wen AND (yy_rsc_17_0_cgo OR yy_rsc_17_0_cgo_iro);
  yy_rsc_18_0_i_clka_en_d <= core_wen AND (yy_rsc_18_0_cgo OR yy_rsc_18_0_cgo_iro);
  yy_rsc_19_0_i_clka_en_d <= core_wen AND (yy_rsc_19_0_cgo OR yy_rsc_19_0_cgo_iro);
  yy_rsc_20_0_i_clka_en_d <= core_wen AND (yy_rsc_20_0_cgo OR yy_rsc_20_0_cgo_iro);
  yy_rsc_21_0_i_clka_en_d <= core_wen AND (yy_rsc_21_0_cgo OR yy_rsc_21_0_cgo_iro);
  yy_rsc_22_0_i_clka_en_d <= core_wen AND (yy_rsc_22_0_cgo OR yy_rsc_22_0_cgo_iro);
  yy_rsc_23_0_i_clka_en_d <= core_wen AND (yy_rsc_23_0_cgo OR yy_rsc_23_0_cgo_iro);
  yy_rsc_24_0_i_clka_en_d <= core_wen AND (yy_rsc_24_0_cgo OR yy_rsc_24_0_cgo_iro);
  yy_rsc_25_0_i_clka_en_d <= core_wen AND (yy_rsc_25_0_cgo OR yy_rsc_25_0_cgo_iro);
  yy_rsc_26_0_i_clka_en_d <= core_wen AND (yy_rsc_26_0_cgo OR yy_rsc_26_0_cgo_iro);
  yy_rsc_27_0_i_clka_en_d <= core_wen AND (yy_rsc_27_0_cgo OR yy_rsc_27_0_cgo_iro);
  yy_rsc_28_0_i_clka_en_d <= core_wen AND (yy_rsc_28_0_cgo OR yy_rsc_28_0_cgo_iro);
  yy_rsc_29_0_i_clka_en_d <= core_wen AND (yy_rsc_29_0_cgo OR yy_rsc_29_0_cgo_iro);
  yy_rsc_30_0_i_clka_en_d <= core_wen AND (yy_rsc_30_0_cgo OR yy_rsc_30_0_cgo_iro);
  yy_rsc_31_0_i_clka_en_d <= core_wen AND (yy_rsc_31_0_cgo OR yy_rsc_31_0_cgo_iro);
  mult_12_z_mul_cmp_en <= core_wen AND (ensig_cgo OR ensig_cgo_iro);
  mult_z_mul_cmp_en <= core_wen AND (ensig_cgo_1 OR ensig_cgo_iro_1);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( core_wen = '1' ) THEN
        S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg <= S34_OUTER_LOOP_for_tf_mul_cmp_z;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsci_biwt : IN STD_LOGIC;
    twiddle_rsci_bdwt : IN STD_LOGIC;
    twiddle_rsci_adrb_d_core_sct : IN STD_LOGIC
  );
END hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp;

ARCHITECTURE v14 OF hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsci_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsci_qb_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  twiddle_rsci_qb_d_mxwt <= MUX_v_32_2_2(twiddle_rsci_qb_d, twiddle_rsci_qb_d_bfwt,
      twiddle_rsci_bcwt);
  twiddle_rsci_adrb_d <= (NOT twiddle_rsci_adrb_d_core_sct) & (twiddle_rsci_adrb_d_core(3
      DOWNTO 0));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsci_bcwt <= '0';
      ELSE
        twiddle_rsci_bcwt <= NOT((NOT(twiddle_rsci_bcwt OR twiddle_rsci_biwt)) OR
            twiddle_rsci_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsci_biwt = '1' ) THEN
        twiddle_rsci_qb_d_bfwt <= twiddle_rsci_qb_d;
      END IF;
    END IF;
  END PROCESS;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsci_oswt : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsci_biwt : OUT STD_LOGIC;
    twiddle_rsci_bdwt : OUT STD_LOGIC;
    twiddle_rsci_adrb_d_core_sct_pff : OUT STD_LOGIC;
    twiddle_rsci_oswt_pff : IN STD_LOGIC
  );
END hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl;

ARCHITECTURE v14 OF hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl IS
  -- Default Constants

BEGIN
  twiddle_rsci_bdwt <= twiddle_rsci_oswt AND core_wen;
  twiddle_rsci_biwt <= (NOT core_wten) AND twiddle_rsci_oswt;
  twiddle_rsci_adrb_d_core_sct_pff <= twiddle_rsci_oswt_pff AND core_wen;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_h_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_h_rsc_triosy_obj IS
  PORT(
    tw_h_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    tw_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_tw_h_rsc_triosy_obj;

ARCHITECTURE v14 OF hybrid_core_tw_h_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL tw_h_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      tw_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      tw_h_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  tw_h_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => tw_h_rsc_triosy_obj_ld_core_sct,
      lz => tw_h_rsc_triosy_lz
    );
  hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl_inst : hybrid_core_tw_h_rsc_triosy_obj_tw_h_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      tw_h_rsc_triosy_obj_iswt0 => tw_h_rsc_triosy_obj_iswt0,
      tw_h_rsc_triosy_obj_ld_core_sct => tw_h_rsc_triosy_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_rsc_triosy_obj IS
  PORT(
    tw_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    tw_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_tw_rsc_triosy_obj;

ARCHITECTURE v14 OF hybrid_core_tw_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL tw_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      tw_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      tw_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  tw_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => tw_rsc_triosy_obj_ld_core_sct,
      lz => tw_rsc_triosy_lz
    );
  hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl_inst : hybrid_core_tw_rsc_triosy_obj_tw_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      tw_rsc_triosy_obj_iswt0 => tw_rsc_triosy_obj_iswt0,
      tw_rsc_triosy_obj_ld_core_sct => tw_rsc_triosy_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_revArr_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_revArr_rsc_triosy_obj IS
  PORT(
    revArr_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    revArr_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_revArr_rsc_triosy_obj;

ARCHITECTURE v14 OF hybrid_core_revArr_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL revArr_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      revArr_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      revArr_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  revArr_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => revArr_rsc_triosy_obj_ld_core_sct,
      lz => revArr_rsc_triosy_lz
    );
  hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl_inst : hybrid_core_revArr_rsc_triosy_obj_revArr_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      revArr_rsc_triosy_obj_iswt0 => revArr_rsc_triosy_obj_iswt0,
      revArr_rsc_triosy_obj_ld_core_sct => revArr_rsc_triosy_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_h_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_h_rsc_triosy_obj IS
  PORT(
    twiddle_h_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_twiddle_h_rsc_triosy_obj;

ARCHITECTURE v14 OF hybrid_core_twiddle_h_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_lz
    );
  hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl_inst : hybrid_core_twiddle_h_rsc_triosy_obj_twiddle_h_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_obj_iswt0 => twiddle_h_rsc_triosy_obj_iswt0,
      twiddle_h_rsc_triosy_obj_ld_core_sct => twiddle_h_rsc_triosy_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_rsc_triosy_obj IS
  PORT(
    twiddle_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_twiddle_rsc_triosy_obj;

ARCHITECTURE v14 OF hybrid_core_twiddle_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_lz
    );
  hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl_inst : hybrid_core_twiddle_rsc_triosy_obj_twiddle_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_obj_iswt0 => twiddle_rsc_triosy_obj_iswt0,
      twiddle_rsc_triosy_obj_ld_core_sct => twiddle_rsc_triosy_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_m_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_m_rsc_triosy_obj IS
  PORT(
    m_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    m_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_m_rsc_triosy_obj;

ARCHITECTURE v14 OF hybrid_core_m_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL m_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      m_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      m_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  m_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => m_rsc_triosy_obj_ld_core_sct,
      lz => m_rsc_triosy_lz
    );
  hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl_inst : hybrid_core_m_rsc_triosy_obj_m_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      m_rsc_triosy_obj_iswt0 => m_rsc_triosy_obj_iswt0,
      m_rsc_triosy_obj_ld_core_sct => m_rsc_triosy_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_0_0_obj IS
  PORT(
    x_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_0_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_0_0_obj_ld_core_sct,
      lz => x_rsc_triosy_0_0_lz
    );
  hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_0_0_obj_x_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_0_0_obj_iswt0 => x_rsc_triosy_0_0_obj_iswt0,
      x_rsc_triosy_0_0_obj_ld_core_sct => x_rsc_triosy_0_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_1_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_1_0_obj IS
  PORT(
    x_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_1_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_1_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_1_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_1_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_1_0_obj_ld_core_sct,
      lz => x_rsc_triosy_1_0_lz
    );
  hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_1_0_obj_x_rsc_triosy_1_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_1_0_obj_iswt0 => x_rsc_triosy_1_0_obj_iswt0,
      x_rsc_triosy_1_0_obj_ld_core_sct => x_rsc_triosy_1_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_2_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_2_0_obj IS
  PORT(
    x_rsc_triosy_2_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_2_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_2_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_2_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_2_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_2_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_2_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_2_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_2_0_obj_ld_core_sct,
      lz => x_rsc_triosy_2_0_lz
    );
  hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_2_0_obj_x_rsc_triosy_2_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_2_0_obj_iswt0 => x_rsc_triosy_2_0_obj_iswt0,
      x_rsc_triosy_2_0_obj_ld_core_sct => x_rsc_triosy_2_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_3_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_3_0_obj IS
  PORT(
    x_rsc_triosy_3_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_3_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_3_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_3_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_3_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_3_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_3_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_3_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_3_0_obj_ld_core_sct,
      lz => x_rsc_triosy_3_0_lz
    );
  hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_3_0_obj_x_rsc_triosy_3_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_3_0_obj_iswt0 => x_rsc_triosy_3_0_obj_iswt0,
      x_rsc_triosy_3_0_obj_ld_core_sct => x_rsc_triosy_3_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_4_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_4_0_obj IS
  PORT(
    x_rsc_triosy_4_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_4_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_4_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_4_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_4_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_4_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_4_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_4_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_4_0_obj_ld_core_sct,
      lz => x_rsc_triosy_4_0_lz
    );
  hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_4_0_obj_x_rsc_triosy_4_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_4_0_obj_iswt0 => x_rsc_triosy_4_0_obj_iswt0,
      x_rsc_triosy_4_0_obj_ld_core_sct => x_rsc_triosy_4_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_5_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_5_0_obj IS
  PORT(
    x_rsc_triosy_5_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_5_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_5_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_5_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_5_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_5_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_5_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_5_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_5_0_obj_ld_core_sct,
      lz => x_rsc_triosy_5_0_lz
    );
  hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_5_0_obj_x_rsc_triosy_5_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_5_0_obj_iswt0 => x_rsc_triosy_5_0_obj_iswt0,
      x_rsc_triosy_5_0_obj_ld_core_sct => x_rsc_triosy_5_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_6_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_6_0_obj IS
  PORT(
    x_rsc_triosy_6_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_6_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_6_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_6_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_6_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_6_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_6_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_6_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_6_0_obj_ld_core_sct,
      lz => x_rsc_triosy_6_0_lz
    );
  hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_6_0_obj_x_rsc_triosy_6_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_6_0_obj_iswt0 => x_rsc_triosy_6_0_obj_iswt0,
      x_rsc_triosy_6_0_obj_ld_core_sct => x_rsc_triosy_6_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_7_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_7_0_obj IS
  PORT(
    x_rsc_triosy_7_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_7_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_7_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_7_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_7_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_7_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_7_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_7_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_7_0_obj_ld_core_sct,
      lz => x_rsc_triosy_7_0_lz
    );
  hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_7_0_obj_x_rsc_triosy_7_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_7_0_obj_iswt0 => x_rsc_triosy_7_0_obj_iswt0,
      x_rsc_triosy_7_0_obj_ld_core_sct => x_rsc_triosy_7_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_8_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_8_0_obj IS
  PORT(
    x_rsc_triosy_8_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_8_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_8_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_8_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_8_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_8_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_8_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_8_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_8_0_obj_ld_core_sct,
      lz => x_rsc_triosy_8_0_lz
    );
  hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_8_0_obj_x_rsc_triosy_8_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_8_0_obj_iswt0 => x_rsc_triosy_8_0_obj_iswt0,
      x_rsc_triosy_8_0_obj_ld_core_sct => x_rsc_triosy_8_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_9_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_9_0_obj IS
  PORT(
    x_rsc_triosy_9_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_9_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_9_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_9_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_9_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_9_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_9_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_9_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_9_0_obj_ld_core_sct,
      lz => x_rsc_triosy_9_0_lz
    );
  hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_9_0_obj_x_rsc_triosy_9_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_9_0_obj_iswt0 => x_rsc_triosy_9_0_obj_iswt0,
      x_rsc_triosy_9_0_obj_ld_core_sct => x_rsc_triosy_9_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_10_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_10_0_obj IS
  PORT(
    x_rsc_triosy_10_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_10_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_10_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_10_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_10_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_10_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_10_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_10_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_10_0_obj_ld_core_sct,
      lz => x_rsc_triosy_10_0_lz
    );
  hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_10_0_obj_x_rsc_triosy_10_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_10_0_obj_iswt0 => x_rsc_triosy_10_0_obj_iswt0,
      x_rsc_triosy_10_0_obj_ld_core_sct => x_rsc_triosy_10_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_11_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_11_0_obj IS
  PORT(
    x_rsc_triosy_11_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_11_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_11_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_11_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_11_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_11_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_11_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_11_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_11_0_obj_ld_core_sct,
      lz => x_rsc_triosy_11_0_lz
    );
  hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_11_0_obj_x_rsc_triosy_11_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_11_0_obj_iswt0 => x_rsc_triosy_11_0_obj_iswt0,
      x_rsc_triosy_11_0_obj_ld_core_sct => x_rsc_triosy_11_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_12_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_12_0_obj IS
  PORT(
    x_rsc_triosy_12_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_12_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_12_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_12_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_12_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_12_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_12_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_12_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_12_0_obj_ld_core_sct,
      lz => x_rsc_triosy_12_0_lz
    );
  hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_12_0_obj_x_rsc_triosy_12_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_12_0_obj_iswt0 => x_rsc_triosy_12_0_obj_iswt0,
      x_rsc_triosy_12_0_obj_ld_core_sct => x_rsc_triosy_12_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_13_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_13_0_obj IS
  PORT(
    x_rsc_triosy_13_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_13_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_13_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_13_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_13_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_13_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_13_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_13_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_13_0_obj_ld_core_sct,
      lz => x_rsc_triosy_13_0_lz
    );
  hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_13_0_obj_x_rsc_triosy_13_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_13_0_obj_iswt0 => x_rsc_triosy_13_0_obj_iswt0,
      x_rsc_triosy_13_0_obj_ld_core_sct => x_rsc_triosy_13_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_14_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_14_0_obj IS
  PORT(
    x_rsc_triosy_14_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_14_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_14_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_14_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_14_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_14_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_14_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_14_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_14_0_obj_ld_core_sct,
      lz => x_rsc_triosy_14_0_lz
    );
  hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_14_0_obj_x_rsc_triosy_14_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_14_0_obj_iswt0 => x_rsc_triosy_14_0_obj_iswt0,
      x_rsc_triosy_14_0_obj_ld_core_sct => x_rsc_triosy_14_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_15_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_15_0_obj IS
  PORT(
    x_rsc_triosy_15_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_15_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_15_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_15_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_15_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_15_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_15_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_15_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_15_0_obj_ld_core_sct,
      lz => x_rsc_triosy_15_0_lz
    );
  hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_15_0_obj_x_rsc_triosy_15_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_15_0_obj_iswt0 => x_rsc_triosy_15_0_obj_iswt0,
      x_rsc_triosy_15_0_obj_ld_core_sct => x_rsc_triosy_15_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_16_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_16_0_obj IS
  PORT(
    x_rsc_triosy_16_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_16_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_16_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_16_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_16_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_16_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_16_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_16_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_16_0_obj_ld_core_sct,
      lz => x_rsc_triosy_16_0_lz
    );
  hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_16_0_obj_x_rsc_triosy_16_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_16_0_obj_iswt0 => x_rsc_triosy_16_0_obj_iswt0,
      x_rsc_triosy_16_0_obj_ld_core_sct => x_rsc_triosy_16_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_17_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_17_0_obj IS
  PORT(
    x_rsc_triosy_17_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_17_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_17_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_17_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_17_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_17_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_17_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_17_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_17_0_obj_ld_core_sct,
      lz => x_rsc_triosy_17_0_lz
    );
  hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_17_0_obj_x_rsc_triosy_17_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_17_0_obj_iswt0 => x_rsc_triosy_17_0_obj_iswt0,
      x_rsc_triosy_17_0_obj_ld_core_sct => x_rsc_triosy_17_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_18_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_18_0_obj IS
  PORT(
    x_rsc_triosy_18_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_18_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_18_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_18_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_18_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_18_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_18_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_18_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_18_0_obj_ld_core_sct,
      lz => x_rsc_triosy_18_0_lz
    );
  hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_18_0_obj_x_rsc_triosy_18_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_18_0_obj_iswt0 => x_rsc_triosy_18_0_obj_iswt0,
      x_rsc_triosy_18_0_obj_ld_core_sct => x_rsc_triosy_18_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_19_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_19_0_obj IS
  PORT(
    x_rsc_triosy_19_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_19_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_19_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_19_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_19_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_19_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_19_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_19_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_19_0_obj_ld_core_sct,
      lz => x_rsc_triosy_19_0_lz
    );
  hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_19_0_obj_x_rsc_triosy_19_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_19_0_obj_iswt0 => x_rsc_triosy_19_0_obj_iswt0,
      x_rsc_triosy_19_0_obj_ld_core_sct => x_rsc_triosy_19_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_20_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_20_0_obj IS
  PORT(
    x_rsc_triosy_20_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_20_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_20_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_20_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_20_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_20_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_20_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_20_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_20_0_obj_ld_core_sct,
      lz => x_rsc_triosy_20_0_lz
    );
  hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_20_0_obj_x_rsc_triosy_20_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_20_0_obj_iswt0 => x_rsc_triosy_20_0_obj_iswt0,
      x_rsc_triosy_20_0_obj_ld_core_sct => x_rsc_triosy_20_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_21_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_21_0_obj IS
  PORT(
    x_rsc_triosy_21_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_21_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_21_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_21_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_21_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_21_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_21_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_21_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_21_0_obj_ld_core_sct,
      lz => x_rsc_triosy_21_0_lz
    );
  hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_21_0_obj_x_rsc_triosy_21_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_21_0_obj_iswt0 => x_rsc_triosy_21_0_obj_iswt0,
      x_rsc_triosy_21_0_obj_ld_core_sct => x_rsc_triosy_21_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_22_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_22_0_obj IS
  PORT(
    x_rsc_triosy_22_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_22_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_22_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_22_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_22_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_22_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_22_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_22_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_22_0_obj_ld_core_sct,
      lz => x_rsc_triosy_22_0_lz
    );
  hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_22_0_obj_x_rsc_triosy_22_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_22_0_obj_iswt0 => x_rsc_triosy_22_0_obj_iswt0,
      x_rsc_triosy_22_0_obj_ld_core_sct => x_rsc_triosy_22_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_23_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_23_0_obj IS
  PORT(
    x_rsc_triosy_23_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_23_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_23_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_23_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_23_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_23_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_23_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_23_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_23_0_obj_ld_core_sct,
      lz => x_rsc_triosy_23_0_lz
    );
  hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_23_0_obj_x_rsc_triosy_23_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_23_0_obj_iswt0 => x_rsc_triosy_23_0_obj_iswt0,
      x_rsc_triosy_23_0_obj_ld_core_sct => x_rsc_triosy_23_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_24_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_24_0_obj IS
  PORT(
    x_rsc_triosy_24_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_24_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_24_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_24_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_24_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_24_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_24_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_24_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_24_0_obj_ld_core_sct,
      lz => x_rsc_triosy_24_0_lz
    );
  hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_24_0_obj_x_rsc_triosy_24_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_24_0_obj_iswt0 => x_rsc_triosy_24_0_obj_iswt0,
      x_rsc_triosy_24_0_obj_ld_core_sct => x_rsc_triosy_24_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_25_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_25_0_obj IS
  PORT(
    x_rsc_triosy_25_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_25_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_25_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_25_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_25_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_25_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_25_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_25_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_25_0_obj_ld_core_sct,
      lz => x_rsc_triosy_25_0_lz
    );
  hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_25_0_obj_x_rsc_triosy_25_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_25_0_obj_iswt0 => x_rsc_triosy_25_0_obj_iswt0,
      x_rsc_triosy_25_0_obj_ld_core_sct => x_rsc_triosy_25_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_26_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_26_0_obj IS
  PORT(
    x_rsc_triosy_26_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_26_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_26_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_26_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_26_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_26_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_26_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_26_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_26_0_obj_ld_core_sct,
      lz => x_rsc_triosy_26_0_lz
    );
  hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_26_0_obj_x_rsc_triosy_26_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_26_0_obj_iswt0 => x_rsc_triosy_26_0_obj_iswt0,
      x_rsc_triosy_26_0_obj_ld_core_sct => x_rsc_triosy_26_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_27_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_27_0_obj IS
  PORT(
    x_rsc_triosy_27_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_27_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_27_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_27_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_27_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_27_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_27_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_27_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_27_0_obj_ld_core_sct,
      lz => x_rsc_triosy_27_0_lz
    );
  hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_27_0_obj_x_rsc_triosy_27_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_27_0_obj_iswt0 => x_rsc_triosy_27_0_obj_iswt0,
      x_rsc_triosy_27_0_obj_ld_core_sct => x_rsc_triosy_27_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_28_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_28_0_obj IS
  PORT(
    x_rsc_triosy_28_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_28_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_28_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_28_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_28_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_28_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_28_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_28_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_28_0_obj_ld_core_sct,
      lz => x_rsc_triosy_28_0_lz
    );
  hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_28_0_obj_x_rsc_triosy_28_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_28_0_obj_iswt0 => x_rsc_triosy_28_0_obj_iswt0,
      x_rsc_triosy_28_0_obj_ld_core_sct => x_rsc_triosy_28_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_29_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_29_0_obj IS
  PORT(
    x_rsc_triosy_29_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_29_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_29_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_29_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_29_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_29_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_29_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_29_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_29_0_obj_ld_core_sct,
      lz => x_rsc_triosy_29_0_lz
    );
  hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_29_0_obj_x_rsc_triosy_29_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_29_0_obj_iswt0 => x_rsc_triosy_29_0_obj_iswt0,
      x_rsc_triosy_29_0_obj_ld_core_sct => x_rsc_triosy_29_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_30_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_30_0_obj IS
  PORT(
    x_rsc_triosy_30_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_30_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_30_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_30_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_30_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_30_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_30_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_30_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_30_0_obj_ld_core_sct,
      lz => x_rsc_triosy_30_0_lz
    );
  hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_30_0_obj_x_rsc_triosy_30_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_30_0_obj_iswt0 => x_rsc_triosy_30_0_obj_iswt0,
      x_rsc_triosy_30_0_obj_ld_core_sct => x_rsc_triosy_30_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_triosy_31_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_triosy_31_0_obj IS
  PORT(
    x_rsc_triosy_31_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    x_rsc_triosy_31_0_obj_iswt0 : IN STD_LOGIC
  );
END hybrid_core_x_rsc_triosy_31_0_obj;

ARCHITECTURE v14 OF hybrid_core_x_rsc_triosy_31_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL x_rsc_triosy_31_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_31_0_obj_iswt0 : IN STD_LOGIC;
      x_rsc_triosy_31_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  x_rsc_triosy_31_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => x_rsc_triosy_31_0_obj_ld_core_sct,
      lz => x_rsc_triosy_31_0_lz
    );
  hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl_inst : hybrid_core_x_rsc_triosy_31_0_obj_x_rsc_triosy_31_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      x_rsc_triosy_31_0_obj_iswt0 => x_rsc_triosy_31_0_obj_iswt0,
      x_rsc_triosy_31_0_obj_ld_core_sct => x_rsc_triosy_31_0_obj_ld_core_sct
    );
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_31_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_31_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_31_0_s_tdone : IN STD_LOGIC;
    x_rsc_31_0_tr_write_done : IN STD_LOGIC;
    x_rsc_31_0_RREADY : IN STD_LOGIC;
    x_rsc_31_0_RVALID : OUT STD_LOGIC;
    x_rsc_31_0_RUSER : OUT STD_LOGIC;
    x_rsc_31_0_RLAST : OUT STD_LOGIC;
    x_rsc_31_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_RID : OUT STD_LOGIC;
    x_rsc_31_0_ARREADY : OUT STD_LOGIC;
    x_rsc_31_0_ARVALID : IN STD_LOGIC;
    x_rsc_31_0_ARUSER : IN STD_LOGIC;
    x_rsc_31_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARLOCK : IN STD_LOGIC;
    x_rsc_31_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_31_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_31_0_ARID : IN STD_LOGIC;
    x_rsc_31_0_BREADY : IN STD_LOGIC;
    x_rsc_31_0_BVALID : OUT STD_LOGIC;
    x_rsc_31_0_BUSER : OUT STD_LOGIC;
    x_rsc_31_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_BID : OUT STD_LOGIC;
    x_rsc_31_0_WREADY : OUT STD_LOGIC;
    x_rsc_31_0_WVALID : IN STD_LOGIC;
    x_rsc_31_0_WUSER : IN STD_LOGIC;
    x_rsc_31_0_WLAST : IN STD_LOGIC;
    x_rsc_31_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_AWREADY : OUT STD_LOGIC;
    x_rsc_31_0_AWVALID : IN STD_LOGIC;
    x_rsc_31_0_AWUSER : IN STD_LOGIC;
    x_rsc_31_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWLOCK : IN STD_LOGIC;
    x_rsc_31_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_31_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_31_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_31_0_i_oswt : IN STD_LOGIC;
    x_rsc_31_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_31_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_31_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_31_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_31_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_31_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_31_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_31_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_31_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_31_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_31_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_31_0_i_oswt : IN STD_LOGIC;
      x_rsc_31_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_31_0_i_biwt : OUT STD_LOGIC;
      x_rsc_31_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_31_0_i_bcwt : IN STD_LOGIC;
      x_rsc_31_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_31_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_31_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_31_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_31_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_31_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_31_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_31_0_i_oswt : IN STD_LOGIC;
      x_rsc_31_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_31_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_31_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_31_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_31_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_31_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_i_biwt : IN STD_LOGIC;
      x_rsc_31_0_i_bdwt : IN STD_LOGIC;
      x_rsc_31_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_31_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_31_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_31_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_31_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_31_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_31_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_31_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_31_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_31_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_31_0_i_AWID,
      AWADDR => x_rsc_31_0_i_AWADDR,
      AWLEN => x_rsc_31_0_i_AWLEN,
      AWSIZE => x_rsc_31_0_i_AWSIZE,
      AWBURST => x_rsc_31_0_i_AWBURST,
      AWLOCK => x_rsc_31_0_AWLOCK,
      AWCACHE => x_rsc_31_0_i_AWCACHE,
      AWPROT => x_rsc_31_0_i_AWPROT,
      AWQOS => x_rsc_31_0_i_AWQOS,
      AWREGION => x_rsc_31_0_i_AWREGION,
      AWUSER => x_rsc_31_0_i_AWUSER,
      AWVALID => x_rsc_31_0_AWVALID,
      AWREADY => x_rsc_31_0_AWREADY,
      WDATA => x_rsc_31_0_i_WDATA,
      WSTRB => x_rsc_31_0_i_WSTRB,
      WLAST => x_rsc_31_0_WLAST,
      WUSER => x_rsc_31_0_i_WUSER,
      WVALID => x_rsc_31_0_WVALID,
      WREADY => x_rsc_31_0_WREADY,
      BID => x_rsc_31_0_i_BID,
      BRESP => x_rsc_31_0_i_BRESP,
      BUSER => x_rsc_31_0_i_BUSER,
      BVALID => x_rsc_31_0_BVALID,
      BREADY => x_rsc_31_0_BREADY,
      ARID => x_rsc_31_0_i_ARID,
      ARADDR => x_rsc_31_0_i_ARADDR,
      ARLEN => x_rsc_31_0_i_ARLEN,
      ARSIZE => x_rsc_31_0_i_ARSIZE,
      ARBURST => x_rsc_31_0_i_ARBURST,
      ARLOCK => x_rsc_31_0_ARLOCK,
      ARCACHE => x_rsc_31_0_i_ARCACHE,
      ARPROT => x_rsc_31_0_i_ARPROT,
      ARQOS => x_rsc_31_0_i_ARQOS,
      ARREGION => x_rsc_31_0_i_ARREGION,
      ARUSER => x_rsc_31_0_i_ARUSER,
      ARVALID => x_rsc_31_0_ARVALID,
      ARREADY => x_rsc_31_0_ARREADY,
      RID => x_rsc_31_0_i_RID,
      RDATA => x_rsc_31_0_i_RDATA,
      RRESP => x_rsc_31_0_i_RRESP,
      RLAST => x_rsc_31_0_RLAST,
      RUSER => x_rsc_31_0_i_RUSER,
      RVALID => x_rsc_31_0_RVALID,
      RREADY => x_rsc_31_0_RREADY,
      s_re => x_rsc_31_0_i_s_re_core_sct,
      s_we => x_rsc_31_0_i_s_we_core_sct,
      s_raddr => x_rsc_31_0_i_s_raddr_1,
      s_waddr => x_rsc_31_0_i_s_waddr_1,
      s_din => x_rsc_31_0_i_s_din_1,
      s_dout => x_rsc_31_0_i_s_dout_1,
      s_rrdy => x_rsc_31_0_i_s_rrdy,
      s_wrdy => x_rsc_31_0_i_s_wrdy,
      is_idle => x_rsc_31_0_is_idle_1,
      tr_write_done => x_rsc_31_0_tr_write_done,
      s_tdone => x_rsc_31_0_s_tdone
    );
  x_rsc_31_0_i_AWID(0) <= x_rsc_31_0_AWID;
  x_rsc_31_0_i_AWADDR <= x_rsc_31_0_AWADDR;
  x_rsc_31_0_i_AWLEN <= x_rsc_31_0_AWLEN;
  x_rsc_31_0_i_AWSIZE <= x_rsc_31_0_AWSIZE;
  x_rsc_31_0_i_AWBURST <= x_rsc_31_0_AWBURST;
  x_rsc_31_0_i_AWCACHE <= x_rsc_31_0_AWCACHE;
  x_rsc_31_0_i_AWPROT <= x_rsc_31_0_AWPROT;
  x_rsc_31_0_i_AWQOS <= x_rsc_31_0_AWQOS;
  x_rsc_31_0_i_AWREGION <= x_rsc_31_0_AWREGION;
  x_rsc_31_0_i_AWUSER(0) <= x_rsc_31_0_AWUSER;
  x_rsc_31_0_i_WDATA <= x_rsc_31_0_WDATA;
  x_rsc_31_0_i_WSTRB <= x_rsc_31_0_WSTRB;
  x_rsc_31_0_i_WUSER(0) <= x_rsc_31_0_WUSER;
  x_rsc_31_0_BID <= x_rsc_31_0_i_BID(0);
  x_rsc_31_0_BRESP <= x_rsc_31_0_i_BRESP;
  x_rsc_31_0_BUSER <= x_rsc_31_0_i_BUSER(0);
  x_rsc_31_0_i_ARID(0) <= x_rsc_31_0_ARID;
  x_rsc_31_0_i_ARADDR <= x_rsc_31_0_ARADDR;
  x_rsc_31_0_i_ARLEN <= x_rsc_31_0_ARLEN;
  x_rsc_31_0_i_ARSIZE <= x_rsc_31_0_ARSIZE;
  x_rsc_31_0_i_ARBURST <= x_rsc_31_0_ARBURST;
  x_rsc_31_0_i_ARCACHE <= x_rsc_31_0_ARCACHE;
  x_rsc_31_0_i_ARPROT <= x_rsc_31_0_ARPROT;
  x_rsc_31_0_i_ARQOS <= x_rsc_31_0_ARQOS;
  x_rsc_31_0_i_ARREGION <= x_rsc_31_0_ARREGION;
  x_rsc_31_0_i_ARUSER(0) <= x_rsc_31_0_ARUSER;
  x_rsc_31_0_RID <= x_rsc_31_0_i_RID(0);
  x_rsc_31_0_RDATA <= x_rsc_31_0_i_RDATA;
  x_rsc_31_0_RRESP <= x_rsc_31_0_i_RRESP;
  x_rsc_31_0_RUSER <= x_rsc_31_0_i_RUSER(0);
  x_rsc_31_0_i_s_raddr_1 <= x_rsc_31_0_i_s_raddr;
  x_rsc_31_0_i_s_waddr_1 <= x_rsc_31_0_i_s_waddr;
  x_rsc_31_0_i_s_din <= x_rsc_31_0_i_s_din_1;
  x_rsc_31_0_i_s_dout_1 <= x_rsc_31_0_i_s_dout;

  hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl_inst : hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_31_0_i_oswt => x_rsc_31_0_i_oswt,
      x_rsc_31_0_i_oswt_1 => x_rsc_31_0_i_oswt_1,
      x_rsc_31_0_i_biwt => x_rsc_31_0_i_biwt,
      x_rsc_31_0_i_bdwt => x_rsc_31_0_i_bdwt,
      x_rsc_31_0_i_bcwt => x_rsc_31_0_i_bcwt,
      x_rsc_31_0_i_s_re_core_sct => x_rsc_31_0_i_s_re_core_sct,
      x_rsc_31_0_i_biwt_1 => x_rsc_31_0_i_biwt_1,
      x_rsc_31_0_i_bdwt_2 => x_rsc_31_0_i_bdwt_2,
      x_rsc_31_0_i_bcwt_1 => x_rsc_31_0_i_bcwt_1,
      x_rsc_31_0_i_s_we_core_sct => x_rsc_31_0_i_s_we_core_sct,
      x_rsc_31_0_i_s_rrdy => x_rsc_31_0_i_s_rrdy,
      x_rsc_31_0_i_s_wrdy => x_rsc_31_0_i_s_wrdy
    );
  hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst : hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_31_0_i_oswt => x_rsc_31_0_i_oswt,
      x_rsc_31_0_i_wen_comp => x_rsc_31_0_i_wen_comp,
      x_rsc_31_0_i_oswt_1 => x_rsc_31_0_i_oswt_1,
      x_rsc_31_0_i_wen_comp_1 => x_rsc_31_0_i_wen_comp_1,
      x_rsc_31_0_i_s_raddr_core => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_raddr_core,
      x_rsc_31_0_i_s_waddr_core => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_waddr_core,
      x_rsc_31_0_i_s_din_mxwt => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_din_mxwt,
      x_rsc_31_0_i_s_dout_core => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_dout_core,
      x_rsc_31_0_i_biwt => x_rsc_31_0_i_biwt,
      x_rsc_31_0_i_bdwt => x_rsc_31_0_i_bdwt,
      x_rsc_31_0_i_bcwt => x_rsc_31_0_i_bcwt,
      x_rsc_31_0_i_biwt_1 => x_rsc_31_0_i_biwt_1,
      x_rsc_31_0_i_bdwt_2 => x_rsc_31_0_i_bdwt_2,
      x_rsc_31_0_i_bcwt_1 => x_rsc_31_0_i_bcwt_1,
      x_rsc_31_0_i_s_raddr => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_raddr,
      x_rsc_31_0_i_s_raddr_core_sct => x_rsc_31_0_i_s_re_core_sct,
      x_rsc_31_0_i_s_waddr => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_waddr,
      x_rsc_31_0_i_s_waddr_core_sct => x_rsc_31_0_i_s_we_core_sct,
      x_rsc_31_0_i_s_din => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_din,
      x_rsc_31_0_i_s_dout => hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_dout
    );
  hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_raddr_core <= x_rsc_31_0_i_s_raddr_core;
  hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_waddr_core <= x_rsc_31_0_i_s_waddr_core;
  x_rsc_31_0_i_s_din_mxwt <= hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_din_mxwt;
  hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_dout_core <= x_rsc_31_0_i_s_dout_core;
  x_rsc_31_0_i_s_raddr <= hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_raddr;
  x_rsc_31_0_i_s_waddr <= hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_waddr;
  hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_din <= x_rsc_31_0_i_s_din;
  x_rsc_31_0_i_s_dout <= hybrid_core_x_rsc_31_0_i_x_rsc_31_0_wait_dp_inst_x_rsc_31_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_30_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_30_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_30_0_s_tdone : IN STD_LOGIC;
    x_rsc_30_0_tr_write_done : IN STD_LOGIC;
    x_rsc_30_0_RREADY : IN STD_LOGIC;
    x_rsc_30_0_RVALID : OUT STD_LOGIC;
    x_rsc_30_0_RUSER : OUT STD_LOGIC;
    x_rsc_30_0_RLAST : OUT STD_LOGIC;
    x_rsc_30_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_RID : OUT STD_LOGIC;
    x_rsc_30_0_ARREADY : OUT STD_LOGIC;
    x_rsc_30_0_ARVALID : IN STD_LOGIC;
    x_rsc_30_0_ARUSER : IN STD_LOGIC;
    x_rsc_30_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARLOCK : IN STD_LOGIC;
    x_rsc_30_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_30_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_30_0_ARID : IN STD_LOGIC;
    x_rsc_30_0_BREADY : IN STD_LOGIC;
    x_rsc_30_0_BVALID : OUT STD_LOGIC;
    x_rsc_30_0_BUSER : OUT STD_LOGIC;
    x_rsc_30_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_BID : OUT STD_LOGIC;
    x_rsc_30_0_WREADY : OUT STD_LOGIC;
    x_rsc_30_0_WVALID : IN STD_LOGIC;
    x_rsc_30_0_WUSER : IN STD_LOGIC;
    x_rsc_30_0_WLAST : IN STD_LOGIC;
    x_rsc_30_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_AWREADY : OUT STD_LOGIC;
    x_rsc_30_0_AWVALID : IN STD_LOGIC;
    x_rsc_30_0_AWUSER : IN STD_LOGIC;
    x_rsc_30_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWLOCK : IN STD_LOGIC;
    x_rsc_30_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_30_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_30_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_30_0_i_oswt : IN STD_LOGIC;
    x_rsc_30_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_30_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_30_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_30_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_30_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_30_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_30_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_30_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_30_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_30_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_30_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_30_0_i_oswt : IN STD_LOGIC;
      x_rsc_30_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_30_0_i_biwt : OUT STD_LOGIC;
      x_rsc_30_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_30_0_i_bcwt : IN STD_LOGIC;
      x_rsc_30_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_30_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_30_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_30_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_30_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_30_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_30_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_30_0_i_oswt : IN STD_LOGIC;
      x_rsc_30_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_30_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_30_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_30_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_30_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_30_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_i_biwt : IN STD_LOGIC;
      x_rsc_30_0_i_bdwt : IN STD_LOGIC;
      x_rsc_30_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_30_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_30_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_30_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_30_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_30_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_30_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_30_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_30_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_30_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_30_0_i_AWID,
      AWADDR => x_rsc_30_0_i_AWADDR,
      AWLEN => x_rsc_30_0_i_AWLEN,
      AWSIZE => x_rsc_30_0_i_AWSIZE,
      AWBURST => x_rsc_30_0_i_AWBURST,
      AWLOCK => x_rsc_30_0_AWLOCK,
      AWCACHE => x_rsc_30_0_i_AWCACHE,
      AWPROT => x_rsc_30_0_i_AWPROT,
      AWQOS => x_rsc_30_0_i_AWQOS,
      AWREGION => x_rsc_30_0_i_AWREGION,
      AWUSER => x_rsc_30_0_i_AWUSER,
      AWVALID => x_rsc_30_0_AWVALID,
      AWREADY => x_rsc_30_0_AWREADY,
      WDATA => x_rsc_30_0_i_WDATA,
      WSTRB => x_rsc_30_0_i_WSTRB,
      WLAST => x_rsc_30_0_WLAST,
      WUSER => x_rsc_30_0_i_WUSER,
      WVALID => x_rsc_30_0_WVALID,
      WREADY => x_rsc_30_0_WREADY,
      BID => x_rsc_30_0_i_BID,
      BRESP => x_rsc_30_0_i_BRESP,
      BUSER => x_rsc_30_0_i_BUSER,
      BVALID => x_rsc_30_0_BVALID,
      BREADY => x_rsc_30_0_BREADY,
      ARID => x_rsc_30_0_i_ARID,
      ARADDR => x_rsc_30_0_i_ARADDR,
      ARLEN => x_rsc_30_0_i_ARLEN,
      ARSIZE => x_rsc_30_0_i_ARSIZE,
      ARBURST => x_rsc_30_0_i_ARBURST,
      ARLOCK => x_rsc_30_0_ARLOCK,
      ARCACHE => x_rsc_30_0_i_ARCACHE,
      ARPROT => x_rsc_30_0_i_ARPROT,
      ARQOS => x_rsc_30_0_i_ARQOS,
      ARREGION => x_rsc_30_0_i_ARREGION,
      ARUSER => x_rsc_30_0_i_ARUSER,
      ARVALID => x_rsc_30_0_ARVALID,
      ARREADY => x_rsc_30_0_ARREADY,
      RID => x_rsc_30_0_i_RID,
      RDATA => x_rsc_30_0_i_RDATA,
      RRESP => x_rsc_30_0_i_RRESP,
      RLAST => x_rsc_30_0_RLAST,
      RUSER => x_rsc_30_0_i_RUSER,
      RVALID => x_rsc_30_0_RVALID,
      RREADY => x_rsc_30_0_RREADY,
      s_re => x_rsc_30_0_i_s_re_core_sct,
      s_we => x_rsc_30_0_i_s_we_core_sct,
      s_raddr => x_rsc_30_0_i_s_raddr_1,
      s_waddr => x_rsc_30_0_i_s_waddr_1,
      s_din => x_rsc_30_0_i_s_din_1,
      s_dout => x_rsc_30_0_i_s_dout_1,
      s_rrdy => x_rsc_30_0_i_s_rrdy,
      s_wrdy => x_rsc_30_0_i_s_wrdy,
      is_idle => x_rsc_30_0_is_idle_1,
      tr_write_done => x_rsc_30_0_tr_write_done,
      s_tdone => x_rsc_30_0_s_tdone
    );
  x_rsc_30_0_i_AWID(0) <= x_rsc_30_0_AWID;
  x_rsc_30_0_i_AWADDR <= x_rsc_30_0_AWADDR;
  x_rsc_30_0_i_AWLEN <= x_rsc_30_0_AWLEN;
  x_rsc_30_0_i_AWSIZE <= x_rsc_30_0_AWSIZE;
  x_rsc_30_0_i_AWBURST <= x_rsc_30_0_AWBURST;
  x_rsc_30_0_i_AWCACHE <= x_rsc_30_0_AWCACHE;
  x_rsc_30_0_i_AWPROT <= x_rsc_30_0_AWPROT;
  x_rsc_30_0_i_AWQOS <= x_rsc_30_0_AWQOS;
  x_rsc_30_0_i_AWREGION <= x_rsc_30_0_AWREGION;
  x_rsc_30_0_i_AWUSER(0) <= x_rsc_30_0_AWUSER;
  x_rsc_30_0_i_WDATA <= x_rsc_30_0_WDATA;
  x_rsc_30_0_i_WSTRB <= x_rsc_30_0_WSTRB;
  x_rsc_30_0_i_WUSER(0) <= x_rsc_30_0_WUSER;
  x_rsc_30_0_BID <= x_rsc_30_0_i_BID(0);
  x_rsc_30_0_BRESP <= x_rsc_30_0_i_BRESP;
  x_rsc_30_0_BUSER <= x_rsc_30_0_i_BUSER(0);
  x_rsc_30_0_i_ARID(0) <= x_rsc_30_0_ARID;
  x_rsc_30_0_i_ARADDR <= x_rsc_30_0_ARADDR;
  x_rsc_30_0_i_ARLEN <= x_rsc_30_0_ARLEN;
  x_rsc_30_0_i_ARSIZE <= x_rsc_30_0_ARSIZE;
  x_rsc_30_0_i_ARBURST <= x_rsc_30_0_ARBURST;
  x_rsc_30_0_i_ARCACHE <= x_rsc_30_0_ARCACHE;
  x_rsc_30_0_i_ARPROT <= x_rsc_30_0_ARPROT;
  x_rsc_30_0_i_ARQOS <= x_rsc_30_0_ARQOS;
  x_rsc_30_0_i_ARREGION <= x_rsc_30_0_ARREGION;
  x_rsc_30_0_i_ARUSER(0) <= x_rsc_30_0_ARUSER;
  x_rsc_30_0_RID <= x_rsc_30_0_i_RID(0);
  x_rsc_30_0_RDATA <= x_rsc_30_0_i_RDATA;
  x_rsc_30_0_RRESP <= x_rsc_30_0_i_RRESP;
  x_rsc_30_0_RUSER <= x_rsc_30_0_i_RUSER(0);
  x_rsc_30_0_i_s_raddr_1 <= x_rsc_30_0_i_s_raddr;
  x_rsc_30_0_i_s_waddr_1 <= x_rsc_30_0_i_s_waddr;
  x_rsc_30_0_i_s_din <= x_rsc_30_0_i_s_din_1;
  x_rsc_30_0_i_s_dout_1 <= x_rsc_30_0_i_s_dout;

  hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl_inst : hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_30_0_i_oswt => x_rsc_30_0_i_oswt,
      x_rsc_30_0_i_oswt_1 => x_rsc_30_0_i_oswt_1,
      x_rsc_30_0_i_biwt => x_rsc_30_0_i_biwt,
      x_rsc_30_0_i_bdwt => x_rsc_30_0_i_bdwt,
      x_rsc_30_0_i_bcwt => x_rsc_30_0_i_bcwt,
      x_rsc_30_0_i_s_re_core_sct => x_rsc_30_0_i_s_re_core_sct,
      x_rsc_30_0_i_biwt_1 => x_rsc_30_0_i_biwt_1,
      x_rsc_30_0_i_bdwt_2 => x_rsc_30_0_i_bdwt_2,
      x_rsc_30_0_i_bcwt_1 => x_rsc_30_0_i_bcwt_1,
      x_rsc_30_0_i_s_we_core_sct => x_rsc_30_0_i_s_we_core_sct,
      x_rsc_30_0_i_s_rrdy => x_rsc_30_0_i_s_rrdy,
      x_rsc_30_0_i_s_wrdy => x_rsc_30_0_i_s_wrdy
    );
  hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst : hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_30_0_i_oswt => x_rsc_30_0_i_oswt,
      x_rsc_30_0_i_wen_comp => x_rsc_30_0_i_wen_comp,
      x_rsc_30_0_i_oswt_1 => x_rsc_30_0_i_oswt_1,
      x_rsc_30_0_i_wen_comp_1 => x_rsc_30_0_i_wen_comp_1,
      x_rsc_30_0_i_s_raddr_core => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_raddr_core,
      x_rsc_30_0_i_s_waddr_core => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_waddr_core,
      x_rsc_30_0_i_s_din_mxwt => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_din_mxwt,
      x_rsc_30_0_i_s_dout_core => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_dout_core,
      x_rsc_30_0_i_biwt => x_rsc_30_0_i_biwt,
      x_rsc_30_0_i_bdwt => x_rsc_30_0_i_bdwt,
      x_rsc_30_0_i_bcwt => x_rsc_30_0_i_bcwt,
      x_rsc_30_0_i_biwt_1 => x_rsc_30_0_i_biwt_1,
      x_rsc_30_0_i_bdwt_2 => x_rsc_30_0_i_bdwt_2,
      x_rsc_30_0_i_bcwt_1 => x_rsc_30_0_i_bcwt_1,
      x_rsc_30_0_i_s_raddr => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_raddr,
      x_rsc_30_0_i_s_raddr_core_sct => x_rsc_30_0_i_s_re_core_sct,
      x_rsc_30_0_i_s_waddr => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_waddr,
      x_rsc_30_0_i_s_waddr_core_sct => x_rsc_30_0_i_s_we_core_sct,
      x_rsc_30_0_i_s_din => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_din,
      x_rsc_30_0_i_s_dout => hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_dout
    );
  hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_raddr_core <= x_rsc_30_0_i_s_raddr_core;
  hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_waddr_core <= x_rsc_30_0_i_s_waddr_core;
  x_rsc_30_0_i_s_din_mxwt <= hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_din_mxwt;
  hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_dout_core <= x_rsc_30_0_i_s_dout_core;
  x_rsc_30_0_i_s_raddr <= hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_raddr;
  x_rsc_30_0_i_s_waddr <= hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_waddr;
  hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_din <= x_rsc_30_0_i_s_din;
  x_rsc_30_0_i_s_dout <= hybrid_core_x_rsc_30_0_i_x_rsc_30_0_wait_dp_inst_x_rsc_30_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_29_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_29_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_29_0_s_tdone : IN STD_LOGIC;
    x_rsc_29_0_tr_write_done : IN STD_LOGIC;
    x_rsc_29_0_RREADY : IN STD_LOGIC;
    x_rsc_29_0_RVALID : OUT STD_LOGIC;
    x_rsc_29_0_RUSER : OUT STD_LOGIC;
    x_rsc_29_0_RLAST : OUT STD_LOGIC;
    x_rsc_29_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_RID : OUT STD_LOGIC;
    x_rsc_29_0_ARREADY : OUT STD_LOGIC;
    x_rsc_29_0_ARVALID : IN STD_LOGIC;
    x_rsc_29_0_ARUSER : IN STD_LOGIC;
    x_rsc_29_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARLOCK : IN STD_LOGIC;
    x_rsc_29_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_29_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_29_0_ARID : IN STD_LOGIC;
    x_rsc_29_0_BREADY : IN STD_LOGIC;
    x_rsc_29_0_BVALID : OUT STD_LOGIC;
    x_rsc_29_0_BUSER : OUT STD_LOGIC;
    x_rsc_29_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_BID : OUT STD_LOGIC;
    x_rsc_29_0_WREADY : OUT STD_LOGIC;
    x_rsc_29_0_WVALID : IN STD_LOGIC;
    x_rsc_29_0_WUSER : IN STD_LOGIC;
    x_rsc_29_0_WLAST : IN STD_LOGIC;
    x_rsc_29_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_AWREADY : OUT STD_LOGIC;
    x_rsc_29_0_AWVALID : IN STD_LOGIC;
    x_rsc_29_0_AWUSER : IN STD_LOGIC;
    x_rsc_29_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWLOCK : IN STD_LOGIC;
    x_rsc_29_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_29_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_29_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_29_0_i_oswt : IN STD_LOGIC;
    x_rsc_29_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_29_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_29_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_29_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_29_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_29_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_29_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_29_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_29_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_29_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_29_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_29_0_i_oswt : IN STD_LOGIC;
      x_rsc_29_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_29_0_i_biwt : OUT STD_LOGIC;
      x_rsc_29_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_29_0_i_bcwt : IN STD_LOGIC;
      x_rsc_29_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_29_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_29_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_29_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_29_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_29_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_29_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_29_0_i_oswt : IN STD_LOGIC;
      x_rsc_29_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_29_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_29_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_29_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_29_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_29_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_i_biwt : IN STD_LOGIC;
      x_rsc_29_0_i_bdwt : IN STD_LOGIC;
      x_rsc_29_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_29_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_29_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_29_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_29_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_29_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_29_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_29_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_29_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_29_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_29_0_i_AWID,
      AWADDR => x_rsc_29_0_i_AWADDR,
      AWLEN => x_rsc_29_0_i_AWLEN,
      AWSIZE => x_rsc_29_0_i_AWSIZE,
      AWBURST => x_rsc_29_0_i_AWBURST,
      AWLOCK => x_rsc_29_0_AWLOCK,
      AWCACHE => x_rsc_29_0_i_AWCACHE,
      AWPROT => x_rsc_29_0_i_AWPROT,
      AWQOS => x_rsc_29_0_i_AWQOS,
      AWREGION => x_rsc_29_0_i_AWREGION,
      AWUSER => x_rsc_29_0_i_AWUSER,
      AWVALID => x_rsc_29_0_AWVALID,
      AWREADY => x_rsc_29_0_AWREADY,
      WDATA => x_rsc_29_0_i_WDATA,
      WSTRB => x_rsc_29_0_i_WSTRB,
      WLAST => x_rsc_29_0_WLAST,
      WUSER => x_rsc_29_0_i_WUSER,
      WVALID => x_rsc_29_0_WVALID,
      WREADY => x_rsc_29_0_WREADY,
      BID => x_rsc_29_0_i_BID,
      BRESP => x_rsc_29_0_i_BRESP,
      BUSER => x_rsc_29_0_i_BUSER,
      BVALID => x_rsc_29_0_BVALID,
      BREADY => x_rsc_29_0_BREADY,
      ARID => x_rsc_29_0_i_ARID,
      ARADDR => x_rsc_29_0_i_ARADDR,
      ARLEN => x_rsc_29_0_i_ARLEN,
      ARSIZE => x_rsc_29_0_i_ARSIZE,
      ARBURST => x_rsc_29_0_i_ARBURST,
      ARLOCK => x_rsc_29_0_ARLOCK,
      ARCACHE => x_rsc_29_0_i_ARCACHE,
      ARPROT => x_rsc_29_0_i_ARPROT,
      ARQOS => x_rsc_29_0_i_ARQOS,
      ARREGION => x_rsc_29_0_i_ARREGION,
      ARUSER => x_rsc_29_0_i_ARUSER,
      ARVALID => x_rsc_29_0_ARVALID,
      ARREADY => x_rsc_29_0_ARREADY,
      RID => x_rsc_29_0_i_RID,
      RDATA => x_rsc_29_0_i_RDATA,
      RRESP => x_rsc_29_0_i_RRESP,
      RLAST => x_rsc_29_0_RLAST,
      RUSER => x_rsc_29_0_i_RUSER,
      RVALID => x_rsc_29_0_RVALID,
      RREADY => x_rsc_29_0_RREADY,
      s_re => x_rsc_29_0_i_s_re_core_sct,
      s_we => x_rsc_29_0_i_s_we_core_sct,
      s_raddr => x_rsc_29_0_i_s_raddr_1,
      s_waddr => x_rsc_29_0_i_s_waddr_1,
      s_din => x_rsc_29_0_i_s_din_1,
      s_dout => x_rsc_29_0_i_s_dout_1,
      s_rrdy => x_rsc_29_0_i_s_rrdy,
      s_wrdy => x_rsc_29_0_i_s_wrdy,
      is_idle => x_rsc_29_0_is_idle_1,
      tr_write_done => x_rsc_29_0_tr_write_done,
      s_tdone => x_rsc_29_0_s_tdone
    );
  x_rsc_29_0_i_AWID(0) <= x_rsc_29_0_AWID;
  x_rsc_29_0_i_AWADDR <= x_rsc_29_0_AWADDR;
  x_rsc_29_0_i_AWLEN <= x_rsc_29_0_AWLEN;
  x_rsc_29_0_i_AWSIZE <= x_rsc_29_0_AWSIZE;
  x_rsc_29_0_i_AWBURST <= x_rsc_29_0_AWBURST;
  x_rsc_29_0_i_AWCACHE <= x_rsc_29_0_AWCACHE;
  x_rsc_29_0_i_AWPROT <= x_rsc_29_0_AWPROT;
  x_rsc_29_0_i_AWQOS <= x_rsc_29_0_AWQOS;
  x_rsc_29_0_i_AWREGION <= x_rsc_29_0_AWREGION;
  x_rsc_29_0_i_AWUSER(0) <= x_rsc_29_0_AWUSER;
  x_rsc_29_0_i_WDATA <= x_rsc_29_0_WDATA;
  x_rsc_29_0_i_WSTRB <= x_rsc_29_0_WSTRB;
  x_rsc_29_0_i_WUSER(0) <= x_rsc_29_0_WUSER;
  x_rsc_29_0_BID <= x_rsc_29_0_i_BID(0);
  x_rsc_29_0_BRESP <= x_rsc_29_0_i_BRESP;
  x_rsc_29_0_BUSER <= x_rsc_29_0_i_BUSER(0);
  x_rsc_29_0_i_ARID(0) <= x_rsc_29_0_ARID;
  x_rsc_29_0_i_ARADDR <= x_rsc_29_0_ARADDR;
  x_rsc_29_0_i_ARLEN <= x_rsc_29_0_ARLEN;
  x_rsc_29_0_i_ARSIZE <= x_rsc_29_0_ARSIZE;
  x_rsc_29_0_i_ARBURST <= x_rsc_29_0_ARBURST;
  x_rsc_29_0_i_ARCACHE <= x_rsc_29_0_ARCACHE;
  x_rsc_29_0_i_ARPROT <= x_rsc_29_0_ARPROT;
  x_rsc_29_0_i_ARQOS <= x_rsc_29_0_ARQOS;
  x_rsc_29_0_i_ARREGION <= x_rsc_29_0_ARREGION;
  x_rsc_29_0_i_ARUSER(0) <= x_rsc_29_0_ARUSER;
  x_rsc_29_0_RID <= x_rsc_29_0_i_RID(0);
  x_rsc_29_0_RDATA <= x_rsc_29_0_i_RDATA;
  x_rsc_29_0_RRESP <= x_rsc_29_0_i_RRESP;
  x_rsc_29_0_RUSER <= x_rsc_29_0_i_RUSER(0);
  x_rsc_29_0_i_s_raddr_1 <= x_rsc_29_0_i_s_raddr;
  x_rsc_29_0_i_s_waddr_1 <= x_rsc_29_0_i_s_waddr;
  x_rsc_29_0_i_s_din <= x_rsc_29_0_i_s_din_1;
  x_rsc_29_0_i_s_dout_1 <= x_rsc_29_0_i_s_dout;

  hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl_inst : hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_29_0_i_oswt => x_rsc_29_0_i_oswt,
      x_rsc_29_0_i_oswt_1 => x_rsc_29_0_i_oswt_1,
      x_rsc_29_0_i_biwt => x_rsc_29_0_i_biwt,
      x_rsc_29_0_i_bdwt => x_rsc_29_0_i_bdwt,
      x_rsc_29_0_i_bcwt => x_rsc_29_0_i_bcwt,
      x_rsc_29_0_i_s_re_core_sct => x_rsc_29_0_i_s_re_core_sct,
      x_rsc_29_0_i_biwt_1 => x_rsc_29_0_i_biwt_1,
      x_rsc_29_0_i_bdwt_2 => x_rsc_29_0_i_bdwt_2,
      x_rsc_29_0_i_bcwt_1 => x_rsc_29_0_i_bcwt_1,
      x_rsc_29_0_i_s_we_core_sct => x_rsc_29_0_i_s_we_core_sct,
      x_rsc_29_0_i_s_rrdy => x_rsc_29_0_i_s_rrdy,
      x_rsc_29_0_i_s_wrdy => x_rsc_29_0_i_s_wrdy
    );
  hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst : hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_29_0_i_oswt => x_rsc_29_0_i_oswt,
      x_rsc_29_0_i_wen_comp => x_rsc_29_0_i_wen_comp,
      x_rsc_29_0_i_oswt_1 => x_rsc_29_0_i_oswt_1,
      x_rsc_29_0_i_wen_comp_1 => x_rsc_29_0_i_wen_comp_1,
      x_rsc_29_0_i_s_raddr_core => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_raddr_core,
      x_rsc_29_0_i_s_waddr_core => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_waddr_core,
      x_rsc_29_0_i_s_din_mxwt => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_din_mxwt,
      x_rsc_29_0_i_s_dout_core => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_dout_core,
      x_rsc_29_0_i_biwt => x_rsc_29_0_i_biwt,
      x_rsc_29_0_i_bdwt => x_rsc_29_0_i_bdwt,
      x_rsc_29_0_i_bcwt => x_rsc_29_0_i_bcwt,
      x_rsc_29_0_i_biwt_1 => x_rsc_29_0_i_biwt_1,
      x_rsc_29_0_i_bdwt_2 => x_rsc_29_0_i_bdwt_2,
      x_rsc_29_0_i_bcwt_1 => x_rsc_29_0_i_bcwt_1,
      x_rsc_29_0_i_s_raddr => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_raddr,
      x_rsc_29_0_i_s_raddr_core_sct => x_rsc_29_0_i_s_re_core_sct,
      x_rsc_29_0_i_s_waddr => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_waddr,
      x_rsc_29_0_i_s_waddr_core_sct => x_rsc_29_0_i_s_we_core_sct,
      x_rsc_29_0_i_s_din => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_din,
      x_rsc_29_0_i_s_dout => hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_dout
    );
  hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_raddr_core <= x_rsc_29_0_i_s_raddr_core;
  hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_waddr_core <= x_rsc_29_0_i_s_waddr_core;
  x_rsc_29_0_i_s_din_mxwt <= hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_din_mxwt;
  hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_dout_core <= x_rsc_29_0_i_s_dout_core;
  x_rsc_29_0_i_s_raddr <= hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_raddr;
  x_rsc_29_0_i_s_waddr <= hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_waddr;
  hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_din <= x_rsc_29_0_i_s_din;
  x_rsc_29_0_i_s_dout <= hybrid_core_x_rsc_29_0_i_x_rsc_29_0_wait_dp_inst_x_rsc_29_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_28_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_28_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_28_0_s_tdone : IN STD_LOGIC;
    x_rsc_28_0_tr_write_done : IN STD_LOGIC;
    x_rsc_28_0_RREADY : IN STD_LOGIC;
    x_rsc_28_0_RVALID : OUT STD_LOGIC;
    x_rsc_28_0_RUSER : OUT STD_LOGIC;
    x_rsc_28_0_RLAST : OUT STD_LOGIC;
    x_rsc_28_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_RID : OUT STD_LOGIC;
    x_rsc_28_0_ARREADY : OUT STD_LOGIC;
    x_rsc_28_0_ARVALID : IN STD_LOGIC;
    x_rsc_28_0_ARUSER : IN STD_LOGIC;
    x_rsc_28_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARLOCK : IN STD_LOGIC;
    x_rsc_28_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_28_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_28_0_ARID : IN STD_LOGIC;
    x_rsc_28_0_BREADY : IN STD_LOGIC;
    x_rsc_28_0_BVALID : OUT STD_LOGIC;
    x_rsc_28_0_BUSER : OUT STD_LOGIC;
    x_rsc_28_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_BID : OUT STD_LOGIC;
    x_rsc_28_0_WREADY : OUT STD_LOGIC;
    x_rsc_28_0_WVALID : IN STD_LOGIC;
    x_rsc_28_0_WUSER : IN STD_LOGIC;
    x_rsc_28_0_WLAST : IN STD_LOGIC;
    x_rsc_28_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_AWREADY : OUT STD_LOGIC;
    x_rsc_28_0_AWVALID : IN STD_LOGIC;
    x_rsc_28_0_AWUSER : IN STD_LOGIC;
    x_rsc_28_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWLOCK : IN STD_LOGIC;
    x_rsc_28_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_28_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_28_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_28_0_i_oswt : IN STD_LOGIC;
    x_rsc_28_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_28_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_28_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_28_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_28_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_28_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_28_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_28_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_28_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_28_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_28_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_28_0_i_oswt : IN STD_LOGIC;
      x_rsc_28_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_28_0_i_biwt : OUT STD_LOGIC;
      x_rsc_28_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_28_0_i_bcwt : IN STD_LOGIC;
      x_rsc_28_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_28_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_28_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_28_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_28_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_28_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_28_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_28_0_i_oswt : IN STD_LOGIC;
      x_rsc_28_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_28_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_28_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_28_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_28_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_28_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_i_biwt : IN STD_LOGIC;
      x_rsc_28_0_i_bdwt : IN STD_LOGIC;
      x_rsc_28_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_28_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_28_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_28_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_28_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_28_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_28_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_28_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_28_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_28_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_28_0_i_AWID,
      AWADDR => x_rsc_28_0_i_AWADDR,
      AWLEN => x_rsc_28_0_i_AWLEN,
      AWSIZE => x_rsc_28_0_i_AWSIZE,
      AWBURST => x_rsc_28_0_i_AWBURST,
      AWLOCK => x_rsc_28_0_AWLOCK,
      AWCACHE => x_rsc_28_0_i_AWCACHE,
      AWPROT => x_rsc_28_0_i_AWPROT,
      AWQOS => x_rsc_28_0_i_AWQOS,
      AWREGION => x_rsc_28_0_i_AWREGION,
      AWUSER => x_rsc_28_0_i_AWUSER,
      AWVALID => x_rsc_28_0_AWVALID,
      AWREADY => x_rsc_28_0_AWREADY,
      WDATA => x_rsc_28_0_i_WDATA,
      WSTRB => x_rsc_28_0_i_WSTRB,
      WLAST => x_rsc_28_0_WLAST,
      WUSER => x_rsc_28_0_i_WUSER,
      WVALID => x_rsc_28_0_WVALID,
      WREADY => x_rsc_28_0_WREADY,
      BID => x_rsc_28_0_i_BID,
      BRESP => x_rsc_28_0_i_BRESP,
      BUSER => x_rsc_28_0_i_BUSER,
      BVALID => x_rsc_28_0_BVALID,
      BREADY => x_rsc_28_0_BREADY,
      ARID => x_rsc_28_0_i_ARID,
      ARADDR => x_rsc_28_0_i_ARADDR,
      ARLEN => x_rsc_28_0_i_ARLEN,
      ARSIZE => x_rsc_28_0_i_ARSIZE,
      ARBURST => x_rsc_28_0_i_ARBURST,
      ARLOCK => x_rsc_28_0_ARLOCK,
      ARCACHE => x_rsc_28_0_i_ARCACHE,
      ARPROT => x_rsc_28_0_i_ARPROT,
      ARQOS => x_rsc_28_0_i_ARQOS,
      ARREGION => x_rsc_28_0_i_ARREGION,
      ARUSER => x_rsc_28_0_i_ARUSER,
      ARVALID => x_rsc_28_0_ARVALID,
      ARREADY => x_rsc_28_0_ARREADY,
      RID => x_rsc_28_0_i_RID,
      RDATA => x_rsc_28_0_i_RDATA,
      RRESP => x_rsc_28_0_i_RRESP,
      RLAST => x_rsc_28_0_RLAST,
      RUSER => x_rsc_28_0_i_RUSER,
      RVALID => x_rsc_28_0_RVALID,
      RREADY => x_rsc_28_0_RREADY,
      s_re => x_rsc_28_0_i_s_re_core_sct,
      s_we => x_rsc_28_0_i_s_we_core_sct,
      s_raddr => x_rsc_28_0_i_s_raddr_1,
      s_waddr => x_rsc_28_0_i_s_waddr_1,
      s_din => x_rsc_28_0_i_s_din_1,
      s_dout => x_rsc_28_0_i_s_dout_1,
      s_rrdy => x_rsc_28_0_i_s_rrdy,
      s_wrdy => x_rsc_28_0_i_s_wrdy,
      is_idle => x_rsc_28_0_is_idle_1,
      tr_write_done => x_rsc_28_0_tr_write_done,
      s_tdone => x_rsc_28_0_s_tdone
    );
  x_rsc_28_0_i_AWID(0) <= x_rsc_28_0_AWID;
  x_rsc_28_0_i_AWADDR <= x_rsc_28_0_AWADDR;
  x_rsc_28_0_i_AWLEN <= x_rsc_28_0_AWLEN;
  x_rsc_28_0_i_AWSIZE <= x_rsc_28_0_AWSIZE;
  x_rsc_28_0_i_AWBURST <= x_rsc_28_0_AWBURST;
  x_rsc_28_0_i_AWCACHE <= x_rsc_28_0_AWCACHE;
  x_rsc_28_0_i_AWPROT <= x_rsc_28_0_AWPROT;
  x_rsc_28_0_i_AWQOS <= x_rsc_28_0_AWQOS;
  x_rsc_28_0_i_AWREGION <= x_rsc_28_0_AWREGION;
  x_rsc_28_0_i_AWUSER(0) <= x_rsc_28_0_AWUSER;
  x_rsc_28_0_i_WDATA <= x_rsc_28_0_WDATA;
  x_rsc_28_0_i_WSTRB <= x_rsc_28_0_WSTRB;
  x_rsc_28_0_i_WUSER(0) <= x_rsc_28_0_WUSER;
  x_rsc_28_0_BID <= x_rsc_28_0_i_BID(0);
  x_rsc_28_0_BRESP <= x_rsc_28_0_i_BRESP;
  x_rsc_28_0_BUSER <= x_rsc_28_0_i_BUSER(0);
  x_rsc_28_0_i_ARID(0) <= x_rsc_28_0_ARID;
  x_rsc_28_0_i_ARADDR <= x_rsc_28_0_ARADDR;
  x_rsc_28_0_i_ARLEN <= x_rsc_28_0_ARLEN;
  x_rsc_28_0_i_ARSIZE <= x_rsc_28_0_ARSIZE;
  x_rsc_28_0_i_ARBURST <= x_rsc_28_0_ARBURST;
  x_rsc_28_0_i_ARCACHE <= x_rsc_28_0_ARCACHE;
  x_rsc_28_0_i_ARPROT <= x_rsc_28_0_ARPROT;
  x_rsc_28_0_i_ARQOS <= x_rsc_28_0_ARQOS;
  x_rsc_28_0_i_ARREGION <= x_rsc_28_0_ARREGION;
  x_rsc_28_0_i_ARUSER(0) <= x_rsc_28_0_ARUSER;
  x_rsc_28_0_RID <= x_rsc_28_0_i_RID(0);
  x_rsc_28_0_RDATA <= x_rsc_28_0_i_RDATA;
  x_rsc_28_0_RRESP <= x_rsc_28_0_i_RRESP;
  x_rsc_28_0_RUSER <= x_rsc_28_0_i_RUSER(0);
  x_rsc_28_0_i_s_raddr_1 <= x_rsc_28_0_i_s_raddr;
  x_rsc_28_0_i_s_waddr_1 <= x_rsc_28_0_i_s_waddr;
  x_rsc_28_0_i_s_din <= x_rsc_28_0_i_s_din_1;
  x_rsc_28_0_i_s_dout_1 <= x_rsc_28_0_i_s_dout;

  hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl_inst : hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_28_0_i_oswt => x_rsc_28_0_i_oswt,
      x_rsc_28_0_i_oswt_1 => x_rsc_28_0_i_oswt_1,
      x_rsc_28_0_i_biwt => x_rsc_28_0_i_biwt,
      x_rsc_28_0_i_bdwt => x_rsc_28_0_i_bdwt,
      x_rsc_28_0_i_bcwt => x_rsc_28_0_i_bcwt,
      x_rsc_28_0_i_s_re_core_sct => x_rsc_28_0_i_s_re_core_sct,
      x_rsc_28_0_i_biwt_1 => x_rsc_28_0_i_biwt_1,
      x_rsc_28_0_i_bdwt_2 => x_rsc_28_0_i_bdwt_2,
      x_rsc_28_0_i_bcwt_1 => x_rsc_28_0_i_bcwt_1,
      x_rsc_28_0_i_s_we_core_sct => x_rsc_28_0_i_s_we_core_sct,
      x_rsc_28_0_i_s_rrdy => x_rsc_28_0_i_s_rrdy,
      x_rsc_28_0_i_s_wrdy => x_rsc_28_0_i_s_wrdy
    );
  hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst : hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_28_0_i_oswt => x_rsc_28_0_i_oswt,
      x_rsc_28_0_i_wen_comp => x_rsc_28_0_i_wen_comp,
      x_rsc_28_0_i_oswt_1 => x_rsc_28_0_i_oswt_1,
      x_rsc_28_0_i_wen_comp_1 => x_rsc_28_0_i_wen_comp_1,
      x_rsc_28_0_i_s_raddr_core => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_raddr_core,
      x_rsc_28_0_i_s_waddr_core => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_waddr_core,
      x_rsc_28_0_i_s_din_mxwt => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_din_mxwt,
      x_rsc_28_0_i_s_dout_core => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_dout_core,
      x_rsc_28_0_i_biwt => x_rsc_28_0_i_biwt,
      x_rsc_28_0_i_bdwt => x_rsc_28_0_i_bdwt,
      x_rsc_28_0_i_bcwt => x_rsc_28_0_i_bcwt,
      x_rsc_28_0_i_biwt_1 => x_rsc_28_0_i_biwt_1,
      x_rsc_28_0_i_bdwt_2 => x_rsc_28_0_i_bdwt_2,
      x_rsc_28_0_i_bcwt_1 => x_rsc_28_0_i_bcwt_1,
      x_rsc_28_0_i_s_raddr => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_raddr,
      x_rsc_28_0_i_s_raddr_core_sct => x_rsc_28_0_i_s_re_core_sct,
      x_rsc_28_0_i_s_waddr => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_waddr,
      x_rsc_28_0_i_s_waddr_core_sct => x_rsc_28_0_i_s_we_core_sct,
      x_rsc_28_0_i_s_din => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_din,
      x_rsc_28_0_i_s_dout => hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_dout
    );
  hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_raddr_core <= x_rsc_28_0_i_s_raddr_core;
  hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_waddr_core <= x_rsc_28_0_i_s_waddr_core;
  x_rsc_28_0_i_s_din_mxwt <= hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_din_mxwt;
  hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_dout_core <= x_rsc_28_0_i_s_dout_core;
  x_rsc_28_0_i_s_raddr <= hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_raddr;
  x_rsc_28_0_i_s_waddr <= hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_waddr;
  hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_din <= x_rsc_28_0_i_s_din;
  x_rsc_28_0_i_s_dout <= hybrid_core_x_rsc_28_0_i_x_rsc_28_0_wait_dp_inst_x_rsc_28_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_27_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_27_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_27_0_s_tdone : IN STD_LOGIC;
    x_rsc_27_0_tr_write_done : IN STD_LOGIC;
    x_rsc_27_0_RREADY : IN STD_LOGIC;
    x_rsc_27_0_RVALID : OUT STD_LOGIC;
    x_rsc_27_0_RUSER : OUT STD_LOGIC;
    x_rsc_27_0_RLAST : OUT STD_LOGIC;
    x_rsc_27_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_RID : OUT STD_LOGIC;
    x_rsc_27_0_ARREADY : OUT STD_LOGIC;
    x_rsc_27_0_ARVALID : IN STD_LOGIC;
    x_rsc_27_0_ARUSER : IN STD_LOGIC;
    x_rsc_27_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARLOCK : IN STD_LOGIC;
    x_rsc_27_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_27_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_27_0_ARID : IN STD_LOGIC;
    x_rsc_27_0_BREADY : IN STD_LOGIC;
    x_rsc_27_0_BVALID : OUT STD_LOGIC;
    x_rsc_27_0_BUSER : OUT STD_LOGIC;
    x_rsc_27_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_BID : OUT STD_LOGIC;
    x_rsc_27_0_WREADY : OUT STD_LOGIC;
    x_rsc_27_0_WVALID : IN STD_LOGIC;
    x_rsc_27_0_WUSER : IN STD_LOGIC;
    x_rsc_27_0_WLAST : IN STD_LOGIC;
    x_rsc_27_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_AWREADY : OUT STD_LOGIC;
    x_rsc_27_0_AWVALID : IN STD_LOGIC;
    x_rsc_27_0_AWUSER : IN STD_LOGIC;
    x_rsc_27_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWLOCK : IN STD_LOGIC;
    x_rsc_27_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_27_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_27_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_27_0_i_oswt : IN STD_LOGIC;
    x_rsc_27_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_27_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_27_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_27_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_27_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_27_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_27_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_27_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_27_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_27_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_27_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_27_0_i_oswt : IN STD_LOGIC;
      x_rsc_27_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_27_0_i_biwt : OUT STD_LOGIC;
      x_rsc_27_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_27_0_i_bcwt : IN STD_LOGIC;
      x_rsc_27_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_27_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_27_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_27_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_27_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_27_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_27_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_27_0_i_oswt : IN STD_LOGIC;
      x_rsc_27_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_27_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_27_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_27_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_27_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_27_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_i_biwt : IN STD_LOGIC;
      x_rsc_27_0_i_bdwt : IN STD_LOGIC;
      x_rsc_27_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_27_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_27_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_27_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_27_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_27_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_27_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_27_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_27_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_27_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_27_0_i_AWID,
      AWADDR => x_rsc_27_0_i_AWADDR,
      AWLEN => x_rsc_27_0_i_AWLEN,
      AWSIZE => x_rsc_27_0_i_AWSIZE,
      AWBURST => x_rsc_27_0_i_AWBURST,
      AWLOCK => x_rsc_27_0_AWLOCK,
      AWCACHE => x_rsc_27_0_i_AWCACHE,
      AWPROT => x_rsc_27_0_i_AWPROT,
      AWQOS => x_rsc_27_0_i_AWQOS,
      AWREGION => x_rsc_27_0_i_AWREGION,
      AWUSER => x_rsc_27_0_i_AWUSER,
      AWVALID => x_rsc_27_0_AWVALID,
      AWREADY => x_rsc_27_0_AWREADY,
      WDATA => x_rsc_27_0_i_WDATA,
      WSTRB => x_rsc_27_0_i_WSTRB,
      WLAST => x_rsc_27_0_WLAST,
      WUSER => x_rsc_27_0_i_WUSER,
      WVALID => x_rsc_27_0_WVALID,
      WREADY => x_rsc_27_0_WREADY,
      BID => x_rsc_27_0_i_BID,
      BRESP => x_rsc_27_0_i_BRESP,
      BUSER => x_rsc_27_0_i_BUSER,
      BVALID => x_rsc_27_0_BVALID,
      BREADY => x_rsc_27_0_BREADY,
      ARID => x_rsc_27_0_i_ARID,
      ARADDR => x_rsc_27_0_i_ARADDR,
      ARLEN => x_rsc_27_0_i_ARLEN,
      ARSIZE => x_rsc_27_0_i_ARSIZE,
      ARBURST => x_rsc_27_0_i_ARBURST,
      ARLOCK => x_rsc_27_0_ARLOCK,
      ARCACHE => x_rsc_27_0_i_ARCACHE,
      ARPROT => x_rsc_27_0_i_ARPROT,
      ARQOS => x_rsc_27_0_i_ARQOS,
      ARREGION => x_rsc_27_0_i_ARREGION,
      ARUSER => x_rsc_27_0_i_ARUSER,
      ARVALID => x_rsc_27_0_ARVALID,
      ARREADY => x_rsc_27_0_ARREADY,
      RID => x_rsc_27_0_i_RID,
      RDATA => x_rsc_27_0_i_RDATA,
      RRESP => x_rsc_27_0_i_RRESP,
      RLAST => x_rsc_27_0_RLAST,
      RUSER => x_rsc_27_0_i_RUSER,
      RVALID => x_rsc_27_0_RVALID,
      RREADY => x_rsc_27_0_RREADY,
      s_re => x_rsc_27_0_i_s_re_core_sct,
      s_we => x_rsc_27_0_i_s_we_core_sct,
      s_raddr => x_rsc_27_0_i_s_raddr_1,
      s_waddr => x_rsc_27_0_i_s_waddr_1,
      s_din => x_rsc_27_0_i_s_din_1,
      s_dout => x_rsc_27_0_i_s_dout_1,
      s_rrdy => x_rsc_27_0_i_s_rrdy,
      s_wrdy => x_rsc_27_0_i_s_wrdy,
      is_idle => x_rsc_27_0_is_idle_1,
      tr_write_done => x_rsc_27_0_tr_write_done,
      s_tdone => x_rsc_27_0_s_tdone
    );
  x_rsc_27_0_i_AWID(0) <= x_rsc_27_0_AWID;
  x_rsc_27_0_i_AWADDR <= x_rsc_27_0_AWADDR;
  x_rsc_27_0_i_AWLEN <= x_rsc_27_0_AWLEN;
  x_rsc_27_0_i_AWSIZE <= x_rsc_27_0_AWSIZE;
  x_rsc_27_0_i_AWBURST <= x_rsc_27_0_AWBURST;
  x_rsc_27_0_i_AWCACHE <= x_rsc_27_0_AWCACHE;
  x_rsc_27_0_i_AWPROT <= x_rsc_27_0_AWPROT;
  x_rsc_27_0_i_AWQOS <= x_rsc_27_0_AWQOS;
  x_rsc_27_0_i_AWREGION <= x_rsc_27_0_AWREGION;
  x_rsc_27_0_i_AWUSER(0) <= x_rsc_27_0_AWUSER;
  x_rsc_27_0_i_WDATA <= x_rsc_27_0_WDATA;
  x_rsc_27_0_i_WSTRB <= x_rsc_27_0_WSTRB;
  x_rsc_27_0_i_WUSER(0) <= x_rsc_27_0_WUSER;
  x_rsc_27_0_BID <= x_rsc_27_0_i_BID(0);
  x_rsc_27_0_BRESP <= x_rsc_27_0_i_BRESP;
  x_rsc_27_0_BUSER <= x_rsc_27_0_i_BUSER(0);
  x_rsc_27_0_i_ARID(0) <= x_rsc_27_0_ARID;
  x_rsc_27_0_i_ARADDR <= x_rsc_27_0_ARADDR;
  x_rsc_27_0_i_ARLEN <= x_rsc_27_0_ARLEN;
  x_rsc_27_0_i_ARSIZE <= x_rsc_27_0_ARSIZE;
  x_rsc_27_0_i_ARBURST <= x_rsc_27_0_ARBURST;
  x_rsc_27_0_i_ARCACHE <= x_rsc_27_0_ARCACHE;
  x_rsc_27_0_i_ARPROT <= x_rsc_27_0_ARPROT;
  x_rsc_27_0_i_ARQOS <= x_rsc_27_0_ARQOS;
  x_rsc_27_0_i_ARREGION <= x_rsc_27_0_ARREGION;
  x_rsc_27_0_i_ARUSER(0) <= x_rsc_27_0_ARUSER;
  x_rsc_27_0_RID <= x_rsc_27_0_i_RID(0);
  x_rsc_27_0_RDATA <= x_rsc_27_0_i_RDATA;
  x_rsc_27_0_RRESP <= x_rsc_27_0_i_RRESP;
  x_rsc_27_0_RUSER <= x_rsc_27_0_i_RUSER(0);
  x_rsc_27_0_i_s_raddr_1 <= x_rsc_27_0_i_s_raddr;
  x_rsc_27_0_i_s_waddr_1 <= x_rsc_27_0_i_s_waddr;
  x_rsc_27_0_i_s_din <= x_rsc_27_0_i_s_din_1;
  x_rsc_27_0_i_s_dout_1 <= x_rsc_27_0_i_s_dout;

  hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl_inst : hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_27_0_i_oswt => x_rsc_27_0_i_oswt,
      x_rsc_27_0_i_oswt_1 => x_rsc_27_0_i_oswt_1,
      x_rsc_27_0_i_biwt => x_rsc_27_0_i_biwt,
      x_rsc_27_0_i_bdwt => x_rsc_27_0_i_bdwt,
      x_rsc_27_0_i_bcwt => x_rsc_27_0_i_bcwt,
      x_rsc_27_0_i_s_re_core_sct => x_rsc_27_0_i_s_re_core_sct,
      x_rsc_27_0_i_biwt_1 => x_rsc_27_0_i_biwt_1,
      x_rsc_27_0_i_bdwt_2 => x_rsc_27_0_i_bdwt_2,
      x_rsc_27_0_i_bcwt_1 => x_rsc_27_0_i_bcwt_1,
      x_rsc_27_0_i_s_we_core_sct => x_rsc_27_0_i_s_we_core_sct,
      x_rsc_27_0_i_s_rrdy => x_rsc_27_0_i_s_rrdy,
      x_rsc_27_0_i_s_wrdy => x_rsc_27_0_i_s_wrdy
    );
  hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst : hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_27_0_i_oswt => x_rsc_27_0_i_oswt,
      x_rsc_27_0_i_wen_comp => x_rsc_27_0_i_wen_comp,
      x_rsc_27_0_i_oswt_1 => x_rsc_27_0_i_oswt_1,
      x_rsc_27_0_i_wen_comp_1 => x_rsc_27_0_i_wen_comp_1,
      x_rsc_27_0_i_s_raddr_core => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_raddr_core,
      x_rsc_27_0_i_s_waddr_core => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_waddr_core,
      x_rsc_27_0_i_s_din_mxwt => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_din_mxwt,
      x_rsc_27_0_i_s_dout_core => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_dout_core,
      x_rsc_27_0_i_biwt => x_rsc_27_0_i_biwt,
      x_rsc_27_0_i_bdwt => x_rsc_27_0_i_bdwt,
      x_rsc_27_0_i_bcwt => x_rsc_27_0_i_bcwt,
      x_rsc_27_0_i_biwt_1 => x_rsc_27_0_i_biwt_1,
      x_rsc_27_0_i_bdwt_2 => x_rsc_27_0_i_bdwt_2,
      x_rsc_27_0_i_bcwt_1 => x_rsc_27_0_i_bcwt_1,
      x_rsc_27_0_i_s_raddr => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_raddr,
      x_rsc_27_0_i_s_raddr_core_sct => x_rsc_27_0_i_s_re_core_sct,
      x_rsc_27_0_i_s_waddr => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_waddr,
      x_rsc_27_0_i_s_waddr_core_sct => x_rsc_27_0_i_s_we_core_sct,
      x_rsc_27_0_i_s_din => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_din,
      x_rsc_27_0_i_s_dout => hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_dout
    );
  hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_raddr_core <= x_rsc_27_0_i_s_raddr_core;
  hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_waddr_core <= x_rsc_27_0_i_s_waddr_core;
  x_rsc_27_0_i_s_din_mxwt <= hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_din_mxwt;
  hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_dout_core <= x_rsc_27_0_i_s_dout_core;
  x_rsc_27_0_i_s_raddr <= hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_raddr;
  x_rsc_27_0_i_s_waddr <= hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_waddr;
  hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_din <= x_rsc_27_0_i_s_din;
  x_rsc_27_0_i_s_dout <= hybrid_core_x_rsc_27_0_i_x_rsc_27_0_wait_dp_inst_x_rsc_27_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_26_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_26_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_26_0_s_tdone : IN STD_LOGIC;
    x_rsc_26_0_tr_write_done : IN STD_LOGIC;
    x_rsc_26_0_RREADY : IN STD_LOGIC;
    x_rsc_26_0_RVALID : OUT STD_LOGIC;
    x_rsc_26_0_RUSER : OUT STD_LOGIC;
    x_rsc_26_0_RLAST : OUT STD_LOGIC;
    x_rsc_26_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_RID : OUT STD_LOGIC;
    x_rsc_26_0_ARREADY : OUT STD_LOGIC;
    x_rsc_26_0_ARVALID : IN STD_LOGIC;
    x_rsc_26_0_ARUSER : IN STD_LOGIC;
    x_rsc_26_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARLOCK : IN STD_LOGIC;
    x_rsc_26_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_26_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_26_0_ARID : IN STD_LOGIC;
    x_rsc_26_0_BREADY : IN STD_LOGIC;
    x_rsc_26_0_BVALID : OUT STD_LOGIC;
    x_rsc_26_0_BUSER : OUT STD_LOGIC;
    x_rsc_26_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_BID : OUT STD_LOGIC;
    x_rsc_26_0_WREADY : OUT STD_LOGIC;
    x_rsc_26_0_WVALID : IN STD_LOGIC;
    x_rsc_26_0_WUSER : IN STD_LOGIC;
    x_rsc_26_0_WLAST : IN STD_LOGIC;
    x_rsc_26_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_AWREADY : OUT STD_LOGIC;
    x_rsc_26_0_AWVALID : IN STD_LOGIC;
    x_rsc_26_0_AWUSER : IN STD_LOGIC;
    x_rsc_26_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWLOCK : IN STD_LOGIC;
    x_rsc_26_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_26_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_26_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_26_0_i_oswt : IN STD_LOGIC;
    x_rsc_26_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_26_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_26_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_26_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_26_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_26_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_26_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_26_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_26_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_26_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_26_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_26_0_i_oswt : IN STD_LOGIC;
      x_rsc_26_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_26_0_i_biwt : OUT STD_LOGIC;
      x_rsc_26_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_26_0_i_bcwt : IN STD_LOGIC;
      x_rsc_26_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_26_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_26_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_26_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_26_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_26_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_26_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_26_0_i_oswt : IN STD_LOGIC;
      x_rsc_26_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_26_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_26_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_26_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_26_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_26_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_i_biwt : IN STD_LOGIC;
      x_rsc_26_0_i_bdwt : IN STD_LOGIC;
      x_rsc_26_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_26_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_26_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_26_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_26_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_26_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_26_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_26_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_26_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_26_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_26_0_i_AWID,
      AWADDR => x_rsc_26_0_i_AWADDR,
      AWLEN => x_rsc_26_0_i_AWLEN,
      AWSIZE => x_rsc_26_0_i_AWSIZE,
      AWBURST => x_rsc_26_0_i_AWBURST,
      AWLOCK => x_rsc_26_0_AWLOCK,
      AWCACHE => x_rsc_26_0_i_AWCACHE,
      AWPROT => x_rsc_26_0_i_AWPROT,
      AWQOS => x_rsc_26_0_i_AWQOS,
      AWREGION => x_rsc_26_0_i_AWREGION,
      AWUSER => x_rsc_26_0_i_AWUSER,
      AWVALID => x_rsc_26_0_AWVALID,
      AWREADY => x_rsc_26_0_AWREADY,
      WDATA => x_rsc_26_0_i_WDATA,
      WSTRB => x_rsc_26_0_i_WSTRB,
      WLAST => x_rsc_26_0_WLAST,
      WUSER => x_rsc_26_0_i_WUSER,
      WVALID => x_rsc_26_0_WVALID,
      WREADY => x_rsc_26_0_WREADY,
      BID => x_rsc_26_0_i_BID,
      BRESP => x_rsc_26_0_i_BRESP,
      BUSER => x_rsc_26_0_i_BUSER,
      BVALID => x_rsc_26_0_BVALID,
      BREADY => x_rsc_26_0_BREADY,
      ARID => x_rsc_26_0_i_ARID,
      ARADDR => x_rsc_26_0_i_ARADDR,
      ARLEN => x_rsc_26_0_i_ARLEN,
      ARSIZE => x_rsc_26_0_i_ARSIZE,
      ARBURST => x_rsc_26_0_i_ARBURST,
      ARLOCK => x_rsc_26_0_ARLOCK,
      ARCACHE => x_rsc_26_0_i_ARCACHE,
      ARPROT => x_rsc_26_0_i_ARPROT,
      ARQOS => x_rsc_26_0_i_ARQOS,
      ARREGION => x_rsc_26_0_i_ARREGION,
      ARUSER => x_rsc_26_0_i_ARUSER,
      ARVALID => x_rsc_26_0_ARVALID,
      ARREADY => x_rsc_26_0_ARREADY,
      RID => x_rsc_26_0_i_RID,
      RDATA => x_rsc_26_0_i_RDATA,
      RRESP => x_rsc_26_0_i_RRESP,
      RLAST => x_rsc_26_0_RLAST,
      RUSER => x_rsc_26_0_i_RUSER,
      RVALID => x_rsc_26_0_RVALID,
      RREADY => x_rsc_26_0_RREADY,
      s_re => x_rsc_26_0_i_s_re_core_sct,
      s_we => x_rsc_26_0_i_s_we_core_sct,
      s_raddr => x_rsc_26_0_i_s_raddr_1,
      s_waddr => x_rsc_26_0_i_s_waddr_1,
      s_din => x_rsc_26_0_i_s_din_1,
      s_dout => x_rsc_26_0_i_s_dout_1,
      s_rrdy => x_rsc_26_0_i_s_rrdy,
      s_wrdy => x_rsc_26_0_i_s_wrdy,
      is_idle => x_rsc_26_0_is_idle_1,
      tr_write_done => x_rsc_26_0_tr_write_done,
      s_tdone => x_rsc_26_0_s_tdone
    );
  x_rsc_26_0_i_AWID(0) <= x_rsc_26_0_AWID;
  x_rsc_26_0_i_AWADDR <= x_rsc_26_0_AWADDR;
  x_rsc_26_0_i_AWLEN <= x_rsc_26_0_AWLEN;
  x_rsc_26_0_i_AWSIZE <= x_rsc_26_0_AWSIZE;
  x_rsc_26_0_i_AWBURST <= x_rsc_26_0_AWBURST;
  x_rsc_26_0_i_AWCACHE <= x_rsc_26_0_AWCACHE;
  x_rsc_26_0_i_AWPROT <= x_rsc_26_0_AWPROT;
  x_rsc_26_0_i_AWQOS <= x_rsc_26_0_AWQOS;
  x_rsc_26_0_i_AWREGION <= x_rsc_26_0_AWREGION;
  x_rsc_26_0_i_AWUSER(0) <= x_rsc_26_0_AWUSER;
  x_rsc_26_0_i_WDATA <= x_rsc_26_0_WDATA;
  x_rsc_26_0_i_WSTRB <= x_rsc_26_0_WSTRB;
  x_rsc_26_0_i_WUSER(0) <= x_rsc_26_0_WUSER;
  x_rsc_26_0_BID <= x_rsc_26_0_i_BID(0);
  x_rsc_26_0_BRESP <= x_rsc_26_0_i_BRESP;
  x_rsc_26_0_BUSER <= x_rsc_26_0_i_BUSER(0);
  x_rsc_26_0_i_ARID(0) <= x_rsc_26_0_ARID;
  x_rsc_26_0_i_ARADDR <= x_rsc_26_0_ARADDR;
  x_rsc_26_0_i_ARLEN <= x_rsc_26_0_ARLEN;
  x_rsc_26_0_i_ARSIZE <= x_rsc_26_0_ARSIZE;
  x_rsc_26_0_i_ARBURST <= x_rsc_26_0_ARBURST;
  x_rsc_26_0_i_ARCACHE <= x_rsc_26_0_ARCACHE;
  x_rsc_26_0_i_ARPROT <= x_rsc_26_0_ARPROT;
  x_rsc_26_0_i_ARQOS <= x_rsc_26_0_ARQOS;
  x_rsc_26_0_i_ARREGION <= x_rsc_26_0_ARREGION;
  x_rsc_26_0_i_ARUSER(0) <= x_rsc_26_0_ARUSER;
  x_rsc_26_0_RID <= x_rsc_26_0_i_RID(0);
  x_rsc_26_0_RDATA <= x_rsc_26_0_i_RDATA;
  x_rsc_26_0_RRESP <= x_rsc_26_0_i_RRESP;
  x_rsc_26_0_RUSER <= x_rsc_26_0_i_RUSER(0);
  x_rsc_26_0_i_s_raddr_1 <= x_rsc_26_0_i_s_raddr;
  x_rsc_26_0_i_s_waddr_1 <= x_rsc_26_0_i_s_waddr;
  x_rsc_26_0_i_s_din <= x_rsc_26_0_i_s_din_1;
  x_rsc_26_0_i_s_dout_1 <= x_rsc_26_0_i_s_dout;

  hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl_inst : hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_26_0_i_oswt => x_rsc_26_0_i_oswt,
      x_rsc_26_0_i_oswt_1 => x_rsc_26_0_i_oswt_1,
      x_rsc_26_0_i_biwt => x_rsc_26_0_i_biwt,
      x_rsc_26_0_i_bdwt => x_rsc_26_0_i_bdwt,
      x_rsc_26_0_i_bcwt => x_rsc_26_0_i_bcwt,
      x_rsc_26_0_i_s_re_core_sct => x_rsc_26_0_i_s_re_core_sct,
      x_rsc_26_0_i_biwt_1 => x_rsc_26_0_i_biwt_1,
      x_rsc_26_0_i_bdwt_2 => x_rsc_26_0_i_bdwt_2,
      x_rsc_26_0_i_bcwt_1 => x_rsc_26_0_i_bcwt_1,
      x_rsc_26_0_i_s_we_core_sct => x_rsc_26_0_i_s_we_core_sct,
      x_rsc_26_0_i_s_rrdy => x_rsc_26_0_i_s_rrdy,
      x_rsc_26_0_i_s_wrdy => x_rsc_26_0_i_s_wrdy
    );
  hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst : hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_26_0_i_oswt => x_rsc_26_0_i_oswt,
      x_rsc_26_0_i_wen_comp => x_rsc_26_0_i_wen_comp,
      x_rsc_26_0_i_oswt_1 => x_rsc_26_0_i_oswt_1,
      x_rsc_26_0_i_wen_comp_1 => x_rsc_26_0_i_wen_comp_1,
      x_rsc_26_0_i_s_raddr_core => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_raddr_core,
      x_rsc_26_0_i_s_waddr_core => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_waddr_core,
      x_rsc_26_0_i_s_din_mxwt => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_din_mxwt,
      x_rsc_26_0_i_s_dout_core => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_dout_core,
      x_rsc_26_0_i_biwt => x_rsc_26_0_i_biwt,
      x_rsc_26_0_i_bdwt => x_rsc_26_0_i_bdwt,
      x_rsc_26_0_i_bcwt => x_rsc_26_0_i_bcwt,
      x_rsc_26_0_i_biwt_1 => x_rsc_26_0_i_biwt_1,
      x_rsc_26_0_i_bdwt_2 => x_rsc_26_0_i_bdwt_2,
      x_rsc_26_0_i_bcwt_1 => x_rsc_26_0_i_bcwt_1,
      x_rsc_26_0_i_s_raddr => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_raddr,
      x_rsc_26_0_i_s_raddr_core_sct => x_rsc_26_0_i_s_re_core_sct,
      x_rsc_26_0_i_s_waddr => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_waddr,
      x_rsc_26_0_i_s_waddr_core_sct => x_rsc_26_0_i_s_we_core_sct,
      x_rsc_26_0_i_s_din => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_din,
      x_rsc_26_0_i_s_dout => hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_dout
    );
  hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_raddr_core <= x_rsc_26_0_i_s_raddr_core;
  hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_waddr_core <= x_rsc_26_0_i_s_waddr_core;
  x_rsc_26_0_i_s_din_mxwt <= hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_din_mxwt;
  hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_dout_core <= x_rsc_26_0_i_s_dout_core;
  x_rsc_26_0_i_s_raddr <= hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_raddr;
  x_rsc_26_0_i_s_waddr <= hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_waddr;
  hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_din <= x_rsc_26_0_i_s_din;
  x_rsc_26_0_i_s_dout <= hybrid_core_x_rsc_26_0_i_x_rsc_26_0_wait_dp_inst_x_rsc_26_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_25_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_25_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_25_0_s_tdone : IN STD_LOGIC;
    x_rsc_25_0_tr_write_done : IN STD_LOGIC;
    x_rsc_25_0_RREADY : IN STD_LOGIC;
    x_rsc_25_0_RVALID : OUT STD_LOGIC;
    x_rsc_25_0_RUSER : OUT STD_LOGIC;
    x_rsc_25_0_RLAST : OUT STD_LOGIC;
    x_rsc_25_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_RID : OUT STD_LOGIC;
    x_rsc_25_0_ARREADY : OUT STD_LOGIC;
    x_rsc_25_0_ARVALID : IN STD_LOGIC;
    x_rsc_25_0_ARUSER : IN STD_LOGIC;
    x_rsc_25_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARLOCK : IN STD_LOGIC;
    x_rsc_25_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_25_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_25_0_ARID : IN STD_LOGIC;
    x_rsc_25_0_BREADY : IN STD_LOGIC;
    x_rsc_25_0_BVALID : OUT STD_LOGIC;
    x_rsc_25_0_BUSER : OUT STD_LOGIC;
    x_rsc_25_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_BID : OUT STD_LOGIC;
    x_rsc_25_0_WREADY : OUT STD_LOGIC;
    x_rsc_25_0_WVALID : IN STD_LOGIC;
    x_rsc_25_0_WUSER : IN STD_LOGIC;
    x_rsc_25_0_WLAST : IN STD_LOGIC;
    x_rsc_25_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_AWREADY : OUT STD_LOGIC;
    x_rsc_25_0_AWVALID : IN STD_LOGIC;
    x_rsc_25_0_AWUSER : IN STD_LOGIC;
    x_rsc_25_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWLOCK : IN STD_LOGIC;
    x_rsc_25_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_25_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_25_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_25_0_i_oswt : IN STD_LOGIC;
    x_rsc_25_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_25_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_25_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_25_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_25_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_25_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_25_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_25_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_25_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_25_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_25_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_25_0_i_oswt : IN STD_LOGIC;
      x_rsc_25_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_25_0_i_biwt : OUT STD_LOGIC;
      x_rsc_25_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_25_0_i_bcwt : IN STD_LOGIC;
      x_rsc_25_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_25_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_25_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_25_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_25_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_25_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_25_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_25_0_i_oswt : IN STD_LOGIC;
      x_rsc_25_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_25_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_25_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_25_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_25_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_25_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_i_biwt : IN STD_LOGIC;
      x_rsc_25_0_i_bdwt : IN STD_LOGIC;
      x_rsc_25_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_25_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_25_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_25_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_25_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_25_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_25_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_25_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_25_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_25_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_25_0_i_AWID,
      AWADDR => x_rsc_25_0_i_AWADDR,
      AWLEN => x_rsc_25_0_i_AWLEN,
      AWSIZE => x_rsc_25_0_i_AWSIZE,
      AWBURST => x_rsc_25_0_i_AWBURST,
      AWLOCK => x_rsc_25_0_AWLOCK,
      AWCACHE => x_rsc_25_0_i_AWCACHE,
      AWPROT => x_rsc_25_0_i_AWPROT,
      AWQOS => x_rsc_25_0_i_AWQOS,
      AWREGION => x_rsc_25_0_i_AWREGION,
      AWUSER => x_rsc_25_0_i_AWUSER,
      AWVALID => x_rsc_25_0_AWVALID,
      AWREADY => x_rsc_25_0_AWREADY,
      WDATA => x_rsc_25_0_i_WDATA,
      WSTRB => x_rsc_25_0_i_WSTRB,
      WLAST => x_rsc_25_0_WLAST,
      WUSER => x_rsc_25_0_i_WUSER,
      WVALID => x_rsc_25_0_WVALID,
      WREADY => x_rsc_25_0_WREADY,
      BID => x_rsc_25_0_i_BID,
      BRESP => x_rsc_25_0_i_BRESP,
      BUSER => x_rsc_25_0_i_BUSER,
      BVALID => x_rsc_25_0_BVALID,
      BREADY => x_rsc_25_0_BREADY,
      ARID => x_rsc_25_0_i_ARID,
      ARADDR => x_rsc_25_0_i_ARADDR,
      ARLEN => x_rsc_25_0_i_ARLEN,
      ARSIZE => x_rsc_25_0_i_ARSIZE,
      ARBURST => x_rsc_25_0_i_ARBURST,
      ARLOCK => x_rsc_25_0_ARLOCK,
      ARCACHE => x_rsc_25_0_i_ARCACHE,
      ARPROT => x_rsc_25_0_i_ARPROT,
      ARQOS => x_rsc_25_0_i_ARQOS,
      ARREGION => x_rsc_25_0_i_ARREGION,
      ARUSER => x_rsc_25_0_i_ARUSER,
      ARVALID => x_rsc_25_0_ARVALID,
      ARREADY => x_rsc_25_0_ARREADY,
      RID => x_rsc_25_0_i_RID,
      RDATA => x_rsc_25_0_i_RDATA,
      RRESP => x_rsc_25_0_i_RRESP,
      RLAST => x_rsc_25_0_RLAST,
      RUSER => x_rsc_25_0_i_RUSER,
      RVALID => x_rsc_25_0_RVALID,
      RREADY => x_rsc_25_0_RREADY,
      s_re => x_rsc_25_0_i_s_re_core_sct,
      s_we => x_rsc_25_0_i_s_we_core_sct,
      s_raddr => x_rsc_25_0_i_s_raddr_1,
      s_waddr => x_rsc_25_0_i_s_waddr_1,
      s_din => x_rsc_25_0_i_s_din_1,
      s_dout => x_rsc_25_0_i_s_dout_1,
      s_rrdy => x_rsc_25_0_i_s_rrdy,
      s_wrdy => x_rsc_25_0_i_s_wrdy,
      is_idle => x_rsc_25_0_is_idle_1,
      tr_write_done => x_rsc_25_0_tr_write_done,
      s_tdone => x_rsc_25_0_s_tdone
    );
  x_rsc_25_0_i_AWID(0) <= x_rsc_25_0_AWID;
  x_rsc_25_0_i_AWADDR <= x_rsc_25_0_AWADDR;
  x_rsc_25_0_i_AWLEN <= x_rsc_25_0_AWLEN;
  x_rsc_25_0_i_AWSIZE <= x_rsc_25_0_AWSIZE;
  x_rsc_25_0_i_AWBURST <= x_rsc_25_0_AWBURST;
  x_rsc_25_0_i_AWCACHE <= x_rsc_25_0_AWCACHE;
  x_rsc_25_0_i_AWPROT <= x_rsc_25_0_AWPROT;
  x_rsc_25_0_i_AWQOS <= x_rsc_25_0_AWQOS;
  x_rsc_25_0_i_AWREGION <= x_rsc_25_0_AWREGION;
  x_rsc_25_0_i_AWUSER(0) <= x_rsc_25_0_AWUSER;
  x_rsc_25_0_i_WDATA <= x_rsc_25_0_WDATA;
  x_rsc_25_0_i_WSTRB <= x_rsc_25_0_WSTRB;
  x_rsc_25_0_i_WUSER(0) <= x_rsc_25_0_WUSER;
  x_rsc_25_0_BID <= x_rsc_25_0_i_BID(0);
  x_rsc_25_0_BRESP <= x_rsc_25_0_i_BRESP;
  x_rsc_25_0_BUSER <= x_rsc_25_0_i_BUSER(0);
  x_rsc_25_0_i_ARID(0) <= x_rsc_25_0_ARID;
  x_rsc_25_0_i_ARADDR <= x_rsc_25_0_ARADDR;
  x_rsc_25_0_i_ARLEN <= x_rsc_25_0_ARLEN;
  x_rsc_25_0_i_ARSIZE <= x_rsc_25_0_ARSIZE;
  x_rsc_25_0_i_ARBURST <= x_rsc_25_0_ARBURST;
  x_rsc_25_0_i_ARCACHE <= x_rsc_25_0_ARCACHE;
  x_rsc_25_0_i_ARPROT <= x_rsc_25_0_ARPROT;
  x_rsc_25_0_i_ARQOS <= x_rsc_25_0_ARQOS;
  x_rsc_25_0_i_ARREGION <= x_rsc_25_0_ARREGION;
  x_rsc_25_0_i_ARUSER(0) <= x_rsc_25_0_ARUSER;
  x_rsc_25_0_RID <= x_rsc_25_0_i_RID(0);
  x_rsc_25_0_RDATA <= x_rsc_25_0_i_RDATA;
  x_rsc_25_0_RRESP <= x_rsc_25_0_i_RRESP;
  x_rsc_25_0_RUSER <= x_rsc_25_0_i_RUSER(0);
  x_rsc_25_0_i_s_raddr_1 <= x_rsc_25_0_i_s_raddr;
  x_rsc_25_0_i_s_waddr_1 <= x_rsc_25_0_i_s_waddr;
  x_rsc_25_0_i_s_din <= x_rsc_25_0_i_s_din_1;
  x_rsc_25_0_i_s_dout_1 <= x_rsc_25_0_i_s_dout;

  hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl_inst : hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_25_0_i_oswt => x_rsc_25_0_i_oswt,
      x_rsc_25_0_i_oswt_1 => x_rsc_25_0_i_oswt_1,
      x_rsc_25_0_i_biwt => x_rsc_25_0_i_biwt,
      x_rsc_25_0_i_bdwt => x_rsc_25_0_i_bdwt,
      x_rsc_25_0_i_bcwt => x_rsc_25_0_i_bcwt,
      x_rsc_25_0_i_s_re_core_sct => x_rsc_25_0_i_s_re_core_sct,
      x_rsc_25_0_i_biwt_1 => x_rsc_25_0_i_biwt_1,
      x_rsc_25_0_i_bdwt_2 => x_rsc_25_0_i_bdwt_2,
      x_rsc_25_0_i_bcwt_1 => x_rsc_25_0_i_bcwt_1,
      x_rsc_25_0_i_s_we_core_sct => x_rsc_25_0_i_s_we_core_sct,
      x_rsc_25_0_i_s_rrdy => x_rsc_25_0_i_s_rrdy,
      x_rsc_25_0_i_s_wrdy => x_rsc_25_0_i_s_wrdy
    );
  hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst : hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_25_0_i_oswt => x_rsc_25_0_i_oswt,
      x_rsc_25_0_i_wen_comp => x_rsc_25_0_i_wen_comp,
      x_rsc_25_0_i_oswt_1 => x_rsc_25_0_i_oswt_1,
      x_rsc_25_0_i_wen_comp_1 => x_rsc_25_0_i_wen_comp_1,
      x_rsc_25_0_i_s_raddr_core => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_raddr_core,
      x_rsc_25_0_i_s_waddr_core => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_waddr_core,
      x_rsc_25_0_i_s_din_mxwt => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_din_mxwt,
      x_rsc_25_0_i_s_dout_core => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_dout_core,
      x_rsc_25_0_i_biwt => x_rsc_25_0_i_biwt,
      x_rsc_25_0_i_bdwt => x_rsc_25_0_i_bdwt,
      x_rsc_25_0_i_bcwt => x_rsc_25_0_i_bcwt,
      x_rsc_25_0_i_biwt_1 => x_rsc_25_0_i_biwt_1,
      x_rsc_25_0_i_bdwt_2 => x_rsc_25_0_i_bdwt_2,
      x_rsc_25_0_i_bcwt_1 => x_rsc_25_0_i_bcwt_1,
      x_rsc_25_0_i_s_raddr => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_raddr,
      x_rsc_25_0_i_s_raddr_core_sct => x_rsc_25_0_i_s_re_core_sct,
      x_rsc_25_0_i_s_waddr => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_waddr,
      x_rsc_25_0_i_s_waddr_core_sct => x_rsc_25_0_i_s_we_core_sct,
      x_rsc_25_0_i_s_din => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_din,
      x_rsc_25_0_i_s_dout => hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_dout
    );
  hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_raddr_core <= x_rsc_25_0_i_s_raddr_core;
  hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_waddr_core <= x_rsc_25_0_i_s_waddr_core;
  x_rsc_25_0_i_s_din_mxwt <= hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_din_mxwt;
  hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_dout_core <= x_rsc_25_0_i_s_dout_core;
  x_rsc_25_0_i_s_raddr <= hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_raddr;
  x_rsc_25_0_i_s_waddr <= hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_waddr;
  hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_din <= x_rsc_25_0_i_s_din;
  x_rsc_25_0_i_s_dout <= hybrid_core_x_rsc_25_0_i_x_rsc_25_0_wait_dp_inst_x_rsc_25_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_24_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_24_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_24_0_s_tdone : IN STD_LOGIC;
    x_rsc_24_0_tr_write_done : IN STD_LOGIC;
    x_rsc_24_0_RREADY : IN STD_LOGIC;
    x_rsc_24_0_RVALID : OUT STD_LOGIC;
    x_rsc_24_0_RUSER : OUT STD_LOGIC;
    x_rsc_24_0_RLAST : OUT STD_LOGIC;
    x_rsc_24_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_RID : OUT STD_LOGIC;
    x_rsc_24_0_ARREADY : OUT STD_LOGIC;
    x_rsc_24_0_ARVALID : IN STD_LOGIC;
    x_rsc_24_0_ARUSER : IN STD_LOGIC;
    x_rsc_24_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARLOCK : IN STD_LOGIC;
    x_rsc_24_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_24_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_24_0_ARID : IN STD_LOGIC;
    x_rsc_24_0_BREADY : IN STD_LOGIC;
    x_rsc_24_0_BVALID : OUT STD_LOGIC;
    x_rsc_24_0_BUSER : OUT STD_LOGIC;
    x_rsc_24_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_BID : OUT STD_LOGIC;
    x_rsc_24_0_WREADY : OUT STD_LOGIC;
    x_rsc_24_0_WVALID : IN STD_LOGIC;
    x_rsc_24_0_WUSER : IN STD_LOGIC;
    x_rsc_24_0_WLAST : IN STD_LOGIC;
    x_rsc_24_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_AWREADY : OUT STD_LOGIC;
    x_rsc_24_0_AWVALID : IN STD_LOGIC;
    x_rsc_24_0_AWUSER : IN STD_LOGIC;
    x_rsc_24_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWLOCK : IN STD_LOGIC;
    x_rsc_24_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_24_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_24_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_24_0_i_oswt : IN STD_LOGIC;
    x_rsc_24_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_24_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_24_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_24_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_24_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_24_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_24_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_24_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_24_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_24_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_24_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_24_0_i_oswt : IN STD_LOGIC;
      x_rsc_24_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_24_0_i_biwt : OUT STD_LOGIC;
      x_rsc_24_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_24_0_i_bcwt : IN STD_LOGIC;
      x_rsc_24_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_24_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_24_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_24_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_24_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_24_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_24_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_24_0_i_oswt : IN STD_LOGIC;
      x_rsc_24_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_24_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_24_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_24_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_24_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_24_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_i_biwt : IN STD_LOGIC;
      x_rsc_24_0_i_bdwt : IN STD_LOGIC;
      x_rsc_24_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_24_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_24_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_24_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_24_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_24_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_24_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_24_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_24_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_24_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_24_0_i_AWID,
      AWADDR => x_rsc_24_0_i_AWADDR,
      AWLEN => x_rsc_24_0_i_AWLEN,
      AWSIZE => x_rsc_24_0_i_AWSIZE,
      AWBURST => x_rsc_24_0_i_AWBURST,
      AWLOCK => x_rsc_24_0_AWLOCK,
      AWCACHE => x_rsc_24_0_i_AWCACHE,
      AWPROT => x_rsc_24_0_i_AWPROT,
      AWQOS => x_rsc_24_0_i_AWQOS,
      AWREGION => x_rsc_24_0_i_AWREGION,
      AWUSER => x_rsc_24_0_i_AWUSER,
      AWVALID => x_rsc_24_0_AWVALID,
      AWREADY => x_rsc_24_0_AWREADY,
      WDATA => x_rsc_24_0_i_WDATA,
      WSTRB => x_rsc_24_0_i_WSTRB,
      WLAST => x_rsc_24_0_WLAST,
      WUSER => x_rsc_24_0_i_WUSER,
      WVALID => x_rsc_24_0_WVALID,
      WREADY => x_rsc_24_0_WREADY,
      BID => x_rsc_24_0_i_BID,
      BRESP => x_rsc_24_0_i_BRESP,
      BUSER => x_rsc_24_0_i_BUSER,
      BVALID => x_rsc_24_0_BVALID,
      BREADY => x_rsc_24_0_BREADY,
      ARID => x_rsc_24_0_i_ARID,
      ARADDR => x_rsc_24_0_i_ARADDR,
      ARLEN => x_rsc_24_0_i_ARLEN,
      ARSIZE => x_rsc_24_0_i_ARSIZE,
      ARBURST => x_rsc_24_0_i_ARBURST,
      ARLOCK => x_rsc_24_0_ARLOCK,
      ARCACHE => x_rsc_24_0_i_ARCACHE,
      ARPROT => x_rsc_24_0_i_ARPROT,
      ARQOS => x_rsc_24_0_i_ARQOS,
      ARREGION => x_rsc_24_0_i_ARREGION,
      ARUSER => x_rsc_24_0_i_ARUSER,
      ARVALID => x_rsc_24_0_ARVALID,
      ARREADY => x_rsc_24_0_ARREADY,
      RID => x_rsc_24_0_i_RID,
      RDATA => x_rsc_24_0_i_RDATA,
      RRESP => x_rsc_24_0_i_RRESP,
      RLAST => x_rsc_24_0_RLAST,
      RUSER => x_rsc_24_0_i_RUSER,
      RVALID => x_rsc_24_0_RVALID,
      RREADY => x_rsc_24_0_RREADY,
      s_re => x_rsc_24_0_i_s_re_core_sct,
      s_we => x_rsc_24_0_i_s_we_core_sct,
      s_raddr => x_rsc_24_0_i_s_raddr_1,
      s_waddr => x_rsc_24_0_i_s_waddr_1,
      s_din => x_rsc_24_0_i_s_din_1,
      s_dout => x_rsc_24_0_i_s_dout_1,
      s_rrdy => x_rsc_24_0_i_s_rrdy,
      s_wrdy => x_rsc_24_0_i_s_wrdy,
      is_idle => x_rsc_24_0_is_idle_1,
      tr_write_done => x_rsc_24_0_tr_write_done,
      s_tdone => x_rsc_24_0_s_tdone
    );
  x_rsc_24_0_i_AWID(0) <= x_rsc_24_0_AWID;
  x_rsc_24_0_i_AWADDR <= x_rsc_24_0_AWADDR;
  x_rsc_24_0_i_AWLEN <= x_rsc_24_0_AWLEN;
  x_rsc_24_0_i_AWSIZE <= x_rsc_24_0_AWSIZE;
  x_rsc_24_0_i_AWBURST <= x_rsc_24_0_AWBURST;
  x_rsc_24_0_i_AWCACHE <= x_rsc_24_0_AWCACHE;
  x_rsc_24_0_i_AWPROT <= x_rsc_24_0_AWPROT;
  x_rsc_24_0_i_AWQOS <= x_rsc_24_0_AWQOS;
  x_rsc_24_0_i_AWREGION <= x_rsc_24_0_AWREGION;
  x_rsc_24_0_i_AWUSER(0) <= x_rsc_24_0_AWUSER;
  x_rsc_24_0_i_WDATA <= x_rsc_24_0_WDATA;
  x_rsc_24_0_i_WSTRB <= x_rsc_24_0_WSTRB;
  x_rsc_24_0_i_WUSER(0) <= x_rsc_24_0_WUSER;
  x_rsc_24_0_BID <= x_rsc_24_0_i_BID(0);
  x_rsc_24_0_BRESP <= x_rsc_24_0_i_BRESP;
  x_rsc_24_0_BUSER <= x_rsc_24_0_i_BUSER(0);
  x_rsc_24_0_i_ARID(0) <= x_rsc_24_0_ARID;
  x_rsc_24_0_i_ARADDR <= x_rsc_24_0_ARADDR;
  x_rsc_24_0_i_ARLEN <= x_rsc_24_0_ARLEN;
  x_rsc_24_0_i_ARSIZE <= x_rsc_24_0_ARSIZE;
  x_rsc_24_0_i_ARBURST <= x_rsc_24_0_ARBURST;
  x_rsc_24_0_i_ARCACHE <= x_rsc_24_0_ARCACHE;
  x_rsc_24_0_i_ARPROT <= x_rsc_24_0_ARPROT;
  x_rsc_24_0_i_ARQOS <= x_rsc_24_0_ARQOS;
  x_rsc_24_0_i_ARREGION <= x_rsc_24_0_ARREGION;
  x_rsc_24_0_i_ARUSER(0) <= x_rsc_24_0_ARUSER;
  x_rsc_24_0_RID <= x_rsc_24_0_i_RID(0);
  x_rsc_24_0_RDATA <= x_rsc_24_0_i_RDATA;
  x_rsc_24_0_RRESP <= x_rsc_24_0_i_RRESP;
  x_rsc_24_0_RUSER <= x_rsc_24_0_i_RUSER(0);
  x_rsc_24_0_i_s_raddr_1 <= x_rsc_24_0_i_s_raddr;
  x_rsc_24_0_i_s_waddr_1 <= x_rsc_24_0_i_s_waddr;
  x_rsc_24_0_i_s_din <= x_rsc_24_0_i_s_din_1;
  x_rsc_24_0_i_s_dout_1 <= x_rsc_24_0_i_s_dout;

  hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl_inst : hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_24_0_i_oswt => x_rsc_24_0_i_oswt,
      x_rsc_24_0_i_oswt_1 => x_rsc_24_0_i_oswt_1,
      x_rsc_24_0_i_biwt => x_rsc_24_0_i_biwt,
      x_rsc_24_0_i_bdwt => x_rsc_24_0_i_bdwt,
      x_rsc_24_0_i_bcwt => x_rsc_24_0_i_bcwt,
      x_rsc_24_0_i_s_re_core_sct => x_rsc_24_0_i_s_re_core_sct,
      x_rsc_24_0_i_biwt_1 => x_rsc_24_0_i_biwt_1,
      x_rsc_24_0_i_bdwt_2 => x_rsc_24_0_i_bdwt_2,
      x_rsc_24_0_i_bcwt_1 => x_rsc_24_0_i_bcwt_1,
      x_rsc_24_0_i_s_we_core_sct => x_rsc_24_0_i_s_we_core_sct,
      x_rsc_24_0_i_s_rrdy => x_rsc_24_0_i_s_rrdy,
      x_rsc_24_0_i_s_wrdy => x_rsc_24_0_i_s_wrdy
    );
  hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst : hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_24_0_i_oswt => x_rsc_24_0_i_oswt,
      x_rsc_24_0_i_wen_comp => x_rsc_24_0_i_wen_comp,
      x_rsc_24_0_i_oswt_1 => x_rsc_24_0_i_oswt_1,
      x_rsc_24_0_i_wen_comp_1 => x_rsc_24_0_i_wen_comp_1,
      x_rsc_24_0_i_s_raddr_core => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_raddr_core,
      x_rsc_24_0_i_s_waddr_core => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_waddr_core,
      x_rsc_24_0_i_s_din_mxwt => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_din_mxwt,
      x_rsc_24_0_i_s_dout_core => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_dout_core,
      x_rsc_24_0_i_biwt => x_rsc_24_0_i_biwt,
      x_rsc_24_0_i_bdwt => x_rsc_24_0_i_bdwt,
      x_rsc_24_0_i_bcwt => x_rsc_24_0_i_bcwt,
      x_rsc_24_0_i_biwt_1 => x_rsc_24_0_i_biwt_1,
      x_rsc_24_0_i_bdwt_2 => x_rsc_24_0_i_bdwt_2,
      x_rsc_24_0_i_bcwt_1 => x_rsc_24_0_i_bcwt_1,
      x_rsc_24_0_i_s_raddr => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_raddr,
      x_rsc_24_0_i_s_raddr_core_sct => x_rsc_24_0_i_s_re_core_sct,
      x_rsc_24_0_i_s_waddr => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_waddr,
      x_rsc_24_0_i_s_waddr_core_sct => x_rsc_24_0_i_s_we_core_sct,
      x_rsc_24_0_i_s_din => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_din,
      x_rsc_24_0_i_s_dout => hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_dout
    );
  hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_raddr_core <= x_rsc_24_0_i_s_raddr_core;
  hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_waddr_core <= x_rsc_24_0_i_s_waddr_core;
  x_rsc_24_0_i_s_din_mxwt <= hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_din_mxwt;
  hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_dout_core <= x_rsc_24_0_i_s_dout_core;
  x_rsc_24_0_i_s_raddr <= hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_raddr;
  x_rsc_24_0_i_s_waddr <= hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_waddr;
  hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_din <= x_rsc_24_0_i_s_din;
  x_rsc_24_0_i_s_dout <= hybrid_core_x_rsc_24_0_i_x_rsc_24_0_wait_dp_inst_x_rsc_24_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_23_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_23_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_23_0_s_tdone : IN STD_LOGIC;
    x_rsc_23_0_tr_write_done : IN STD_LOGIC;
    x_rsc_23_0_RREADY : IN STD_LOGIC;
    x_rsc_23_0_RVALID : OUT STD_LOGIC;
    x_rsc_23_0_RUSER : OUT STD_LOGIC;
    x_rsc_23_0_RLAST : OUT STD_LOGIC;
    x_rsc_23_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_RID : OUT STD_LOGIC;
    x_rsc_23_0_ARREADY : OUT STD_LOGIC;
    x_rsc_23_0_ARVALID : IN STD_LOGIC;
    x_rsc_23_0_ARUSER : IN STD_LOGIC;
    x_rsc_23_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARLOCK : IN STD_LOGIC;
    x_rsc_23_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_23_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_23_0_ARID : IN STD_LOGIC;
    x_rsc_23_0_BREADY : IN STD_LOGIC;
    x_rsc_23_0_BVALID : OUT STD_LOGIC;
    x_rsc_23_0_BUSER : OUT STD_LOGIC;
    x_rsc_23_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_BID : OUT STD_LOGIC;
    x_rsc_23_0_WREADY : OUT STD_LOGIC;
    x_rsc_23_0_WVALID : IN STD_LOGIC;
    x_rsc_23_0_WUSER : IN STD_LOGIC;
    x_rsc_23_0_WLAST : IN STD_LOGIC;
    x_rsc_23_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_AWREADY : OUT STD_LOGIC;
    x_rsc_23_0_AWVALID : IN STD_LOGIC;
    x_rsc_23_0_AWUSER : IN STD_LOGIC;
    x_rsc_23_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWLOCK : IN STD_LOGIC;
    x_rsc_23_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_23_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_23_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_23_0_i_oswt : IN STD_LOGIC;
    x_rsc_23_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_23_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_23_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_23_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_23_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_23_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_23_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_23_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_23_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_23_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_23_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_23_0_i_oswt : IN STD_LOGIC;
      x_rsc_23_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_23_0_i_biwt : OUT STD_LOGIC;
      x_rsc_23_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_23_0_i_bcwt : IN STD_LOGIC;
      x_rsc_23_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_23_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_23_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_23_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_23_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_23_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_23_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_23_0_i_oswt : IN STD_LOGIC;
      x_rsc_23_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_23_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_23_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_23_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_23_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_23_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_i_biwt : IN STD_LOGIC;
      x_rsc_23_0_i_bdwt : IN STD_LOGIC;
      x_rsc_23_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_23_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_23_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_23_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_23_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_23_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_23_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_23_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_23_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_23_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_23_0_i_AWID,
      AWADDR => x_rsc_23_0_i_AWADDR,
      AWLEN => x_rsc_23_0_i_AWLEN,
      AWSIZE => x_rsc_23_0_i_AWSIZE,
      AWBURST => x_rsc_23_0_i_AWBURST,
      AWLOCK => x_rsc_23_0_AWLOCK,
      AWCACHE => x_rsc_23_0_i_AWCACHE,
      AWPROT => x_rsc_23_0_i_AWPROT,
      AWQOS => x_rsc_23_0_i_AWQOS,
      AWREGION => x_rsc_23_0_i_AWREGION,
      AWUSER => x_rsc_23_0_i_AWUSER,
      AWVALID => x_rsc_23_0_AWVALID,
      AWREADY => x_rsc_23_0_AWREADY,
      WDATA => x_rsc_23_0_i_WDATA,
      WSTRB => x_rsc_23_0_i_WSTRB,
      WLAST => x_rsc_23_0_WLAST,
      WUSER => x_rsc_23_0_i_WUSER,
      WVALID => x_rsc_23_0_WVALID,
      WREADY => x_rsc_23_0_WREADY,
      BID => x_rsc_23_0_i_BID,
      BRESP => x_rsc_23_0_i_BRESP,
      BUSER => x_rsc_23_0_i_BUSER,
      BVALID => x_rsc_23_0_BVALID,
      BREADY => x_rsc_23_0_BREADY,
      ARID => x_rsc_23_0_i_ARID,
      ARADDR => x_rsc_23_0_i_ARADDR,
      ARLEN => x_rsc_23_0_i_ARLEN,
      ARSIZE => x_rsc_23_0_i_ARSIZE,
      ARBURST => x_rsc_23_0_i_ARBURST,
      ARLOCK => x_rsc_23_0_ARLOCK,
      ARCACHE => x_rsc_23_0_i_ARCACHE,
      ARPROT => x_rsc_23_0_i_ARPROT,
      ARQOS => x_rsc_23_0_i_ARQOS,
      ARREGION => x_rsc_23_0_i_ARREGION,
      ARUSER => x_rsc_23_0_i_ARUSER,
      ARVALID => x_rsc_23_0_ARVALID,
      ARREADY => x_rsc_23_0_ARREADY,
      RID => x_rsc_23_0_i_RID,
      RDATA => x_rsc_23_0_i_RDATA,
      RRESP => x_rsc_23_0_i_RRESP,
      RLAST => x_rsc_23_0_RLAST,
      RUSER => x_rsc_23_0_i_RUSER,
      RVALID => x_rsc_23_0_RVALID,
      RREADY => x_rsc_23_0_RREADY,
      s_re => x_rsc_23_0_i_s_re_core_sct,
      s_we => x_rsc_23_0_i_s_we_core_sct,
      s_raddr => x_rsc_23_0_i_s_raddr_1,
      s_waddr => x_rsc_23_0_i_s_waddr_1,
      s_din => x_rsc_23_0_i_s_din_1,
      s_dout => x_rsc_23_0_i_s_dout_1,
      s_rrdy => x_rsc_23_0_i_s_rrdy,
      s_wrdy => x_rsc_23_0_i_s_wrdy,
      is_idle => x_rsc_23_0_is_idle_1,
      tr_write_done => x_rsc_23_0_tr_write_done,
      s_tdone => x_rsc_23_0_s_tdone
    );
  x_rsc_23_0_i_AWID(0) <= x_rsc_23_0_AWID;
  x_rsc_23_0_i_AWADDR <= x_rsc_23_0_AWADDR;
  x_rsc_23_0_i_AWLEN <= x_rsc_23_0_AWLEN;
  x_rsc_23_0_i_AWSIZE <= x_rsc_23_0_AWSIZE;
  x_rsc_23_0_i_AWBURST <= x_rsc_23_0_AWBURST;
  x_rsc_23_0_i_AWCACHE <= x_rsc_23_0_AWCACHE;
  x_rsc_23_0_i_AWPROT <= x_rsc_23_0_AWPROT;
  x_rsc_23_0_i_AWQOS <= x_rsc_23_0_AWQOS;
  x_rsc_23_0_i_AWREGION <= x_rsc_23_0_AWREGION;
  x_rsc_23_0_i_AWUSER(0) <= x_rsc_23_0_AWUSER;
  x_rsc_23_0_i_WDATA <= x_rsc_23_0_WDATA;
  x_rsc_23_0_i_WSTRB <= x_rsc_23_0_WSTRB;
  x_rsc_23_0_i_WUSER(0) <= x_rsc_23_0_WUSER;
  x_rsc_23_0_BID <= x_rsc_23_0_i_BID(0);
  x_rsc_23_0_BRESP <= x_rsc_23_0_i_BRESP;
  x_rsc_23_0_BUSER <= x_rsc_23_0_i_BUSER(0);
  x_rsc_23_0_i_ARID(0) <= x_rsc_23_0_ARID;
  x_rsc_23_0_i_ARADDR <= x_rsc_23_0_ARADDR;
  x_rsc_23_0_i_ARLEN <= x_rsc_23_0_ARLEN;
  x_rsc_23_0_i_ARSIZE <= x_rsc_23_0_ARSIZE;
  x_rsc_23_0_i_ARBURST <= x_rsc_23_0_ARBURST;
  x_rsc_23_0_i_ARCACHE <= x_rsc_23_0_ARCACHE;
  x_rsc_23_0_i_ARPROT <= x_rsc_23_0_ARPROT;
  x_rsc_23_0_i_ARQOS <= x_rsc_23_0_ARQOS;
  x_rsc_23_0_i_ARREGION <= x_rsc_23_0_ARREGION;
  x_rsc_23_0_i_ARUSER(0) <= x_rsc_23_0_ARUSER;
  x_rsc_23_0_RID <= x_rsc_23_0_i_RID(0);
  x_rsc_23_0_RDATA <= x_rsc_23_0_i_RDATA;
  x_rsc_23_0_RRESP <= x_rsc_23_0_i_RRESP;
  x_rsc_23_0_RUSER <= x_rsc_23_0_i_RUSER(0);
  x_rsc_23_0_i_s_raddr_1 <= x_rsc_23_0_i_s_raddr;
  x_rsc_23_0_i_s_waddr_1 <= x_rsc_23_0_i_s_waddr;
  x_rsc_23_0_i_s_din <= x_rsc_23_0_i_s_din_1;
  x_rsc_23_0_i_s_dout_1 <= x_rsc_23_0_i_s_dout;

  hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl_inst : hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_23_0_i_oswt => x_rsc_23_0_i_oswt,
      x_rsc_23_0_i_oswt_1 => x_rsc_23_0_i_oswt_1,
      x_rsc_23_0_i_biwt => x_rsc_23_0_i_biwt,
      x_rsc_23_0_i_bdwt => x_rsc_23_0_i_bdwt,
      x_rsc_23_0_i_bcwt => x_rsc_23_0_i_bcwt,
      x_rsc_23_0_i_s_re_core_sct => x_rsc_23_0_i_s_re_core_sct,
      x_rsc_23_0_i_biwt_1 => x_rsc_23_0_i_biwt_1,
      x_rsc_23_0_i_bdwt_2 => x_rsc_23_0_i_bdwt_2,
      x_rsc_23_0_i_bcwt_1 => x_rsc_23_0_i_bcwt_1,
      x_rsc_23_0_i_s_we_core_sct => x_rsc_23_0_i_s_we_core_sct,
      x_rsc_23_0_i_s_rrdy => x_rsc_23_0_i_s_rrdy,
      x_rsc_23_0_i_s_wrdy => x_rsc_23_0_i_s_wrdy
    );
  hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst : hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_23_0_i_oswt => x_rsc_23_0_i_oswt,
      x_rsc_23_0_i_wen_comp => x_rsc_23_0_i_wen_comp,
      x_rsc_23_0_i_oswt_1 => x_rsc_23_0_i_oswt_1,
      x_rsc_23_0_i_wen_comp_1 => x_rsc_23_0_i_wen_comp_1,
      x_rsc_23_0_i_s_raddr_core => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_raddr_core,
      x_rsc_23_0_i_s_waddr_core => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_waddr_core,
      x_rsc_23_0_i_s_din_mxwt => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_din_mxwt,
      x_rsc_23_0_i_s_dout_core => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_dout_core,
      x_rsc_23_0_i_biwt => x_rsc_23_0_i_biwt,
      x_rsc_23_0_i_bdwt => x_rsc_23_0_i_bdwt,
      x_rsc_23_0_i_bcwt => x_rsc_23_0_i_bcwt,
      x_rsc_23_0_i_biwt_1 => x_rsc_23_0_i_biwt_1,
      x_rsc_23_0_i_bdwt_2 => x_rsc_23_0_i_bdwt_2,
      x_rsc_23_0_i_bcwt_1 => x_rsc_23_0_i_bcwt_1,
      x_rsc_23_0_i_s_raddr => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_raddr,
      x_rsc_23_0_i_s_raddr_core_sct => x_rsc_23_0_i_s_re_core_sct,
      x_rsc_23_0_i_s_waddr => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_waddr,
      x_rsc_23_0_i_s_waddr_core_sct => x_rsc_23_0_i_s_we_core_sct,
      x_rsc_23_0_i_s_din => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_din,
      x_rsc_23_0_i_s_dout => hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_dout
    );
  hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_raddr_core <= x_rsc_23_0_i_s_raddr_core;
  hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_waddr_core <= x_rsc_23_0_i_s_waddr_core;
  x_rsc_23_0_i_s_din_mxwt <= hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_din_mxwt;
  hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_dout_core <= x_rsc_23_0_i_s_dout_core;
  x_rsc_23_0_i_s_raddr <= hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_raddr;
  x_rsc_23_0_i_s_waddr <= hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_waddr;
  hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_din <= x_rsc_23_0_i_s_din;
  x_rsc_23_0_i_s_dout <= hybrid_core_x_rsc_23_0_i_x_rsc_23_0_wait_dp_inst_x_rsc_23_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_22_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_22_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_22_0_s_tdone : IN STD_LOGIC;
    x_rsc_22_0_tr_write_done : IN STD_LOGIC;
    x_rsc_22_0_RREADY : IN STD_LOGIC;
    x_rsc_22_0_RVALID : OUT STD_LOGIC;
    x_rsc_22_0_RUSER : OUT STD_LOGIC;
    x_rsc_22_0_RLAST : OUT STD_LOGIC;
    x_rsc_22_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_RID : OUT STD_LOGIC;
    x_rsc_22_0_ARREADY : OUT STD_LOGIC;
    x_rsc_22_0_ARVALID : IN STD_LOGIC;
    x_rsc_22_0_ARUSER : IN STD_LOGIC;
    x_rsc_22_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARLOCK : IN STD_LOGIC;
    x_rsc_22_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_22_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_22_0_ARID : IN STD_LOGIC;
    x_rsc_22_0_BREADY : IN STD_LOGIC;
    x_rsc_22_0_BVALID : OUT STD_LOGIC;
    x_rsc_22_0_BUSER : OUT STD_LOGIC;
    x_rsc_22_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_BID : OUT STD_LOGIC;
    x_rsc_22_0_WREADY : OUT STD_LOGIC;
    x_rsc_22_0_WVALID : IN STD_LOGIC;
    x_rsc_22_0_WUSER : IN STD_LOGIC;
    x_rsc_22_0_WLAST : IN STD_LOGIC;
    x_rsc_22_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_AWREADY : OUT STD_LOGIC;
    x_rsc_22_0_AWVALID : IN STD_LOGIC;
    x_rsc_22_0_AWUSER : IN STD_LOGIC;
    x_rsc_22_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWLOCK : IN STD_LOGIC;
    x_rsc_22_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_22_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_22_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_22_0_i_oswt : IN STD_LOGIC;
    x_rsc_22_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_22_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_22_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_22_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_22_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_22_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_22_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_22_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_22_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_22_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_22_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_22_0_i_oswt : IN STD_LOGIC;
      x_rsc_22_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_22_0_i_biwt : OUT STD_LOGIC;
      x_rsc_22_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_22_0_i_bcwt : IN STD_LOGIC;
      x_rsc_22_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_22_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_22_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_22_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_22_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_22_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_22_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_22_0_i_oswt : IN STD_LOGIC;
      x_rsc_22_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_22_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_22_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_22_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_22_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_22_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_i_biwt : IN STD_LOGIC;
      x_rsc_22_0_i_bdwt : IN STD_LOGIC;
      x_rsc_22_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_22_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_22_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_22_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_22_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_22_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_22_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_22_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_22_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_22_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_22_0_i_AWID,
      AWADDR => x_rsc_22_0_i_AWADDR,
      AWLEN => x_rsc_22_0_i_AWLEN,
      AWSIZE => x_rsc_22_0_i_AWSIZE,
      AWBURST => x_rsc_22_0_i_AWBURST,
      AWLOCK => x_rsc_22_0_AWLOCK,
      AWCACHE => x_rsc_22_0_i_AWCACHE,
      AWPROT => x_rsc_22_0_i_AWPROT,
      AWQOS => x_rsc_22_0_i_AWQOS,
      AWREGION => x_rsc_22_0_i_AWREGION,
      AWUSER => x_rsc_22_0_i_AWUSER,
      AWVALID => x_rsc_22_0_AWVALID,
      AWREADY => x_rsc_22_0_AWREADY,
      WDATA => x_rsc_22_0_i_WDATA,
      WSTRB => x_rsc_22_0_i_WSTRB,
      WLAST => x_rsc_22_0_WLAST,
      WUSER => x_rsc_22_0_i_WUSER,
      WVALID => x_rsc_22_0_WVALID,
      WREADY => x_rsc_22_0_WREADY,
      BID => x_rsc_22_0_i_BID,
      BRESP => x_rsc_22_0_i_BRESP,
      BUSER => x_rsc_22_0_i_BUSER,
      BVALID => x_rsc_22_0_BVALID,
      BREADY => x_rsc_22_0_BREADY,
      ARID => x_rsc_22_0_i_ARID,
      ARADDR => x_rsc_22_0_i_ARADDR,
      ARLEN => x_rsc_22_0_i_ARLEN,
      ARSIZE => x_rsc_22_0_i_ARSIZE,
      ARBURST => x_rsc_22_0_i_ARBURST,
      ARLOCK => x_rsc_22_0_ARLOCK,
      ARCACHE => x_rsc_22_0_i_ARCACHE,
      ARPROT => x_rsc_22_0_i_ARPROT,
      ARQOS => x_rsc_22_0_i_ARQOS,
      ARREGION => x_rsc_22_0_i_ARREGION,
      ARUSER => x_rsc_22_0_i_ARUSER,
      ARVALID => x_rsc_22_0_ARVALID,
      ARREADY => x_rsc_22_0_ARREADY,
      RID => x_rsc_22_0_i_RID,
      RDATA => x_rsc_22_0_i_RDATA,
      RRESP => x_rsc_22_0_i_RRESP,
      RLAST => x_rsc_22_0_RLAST,
      RUSER => x_rsc_22_0_i_RUSER,
      RVALID => x_rsc_22_0_RVALID,
      RREADY => x_rsc_22_0_RREADY,
      s_re => x_rsc_22_0_i_s_re_core_sct,
      s_we => x_rsc_22_0_i_s_we_core_sct,
      s_raddr => x_rsc_22_0_i_s_raddr_1,
      s_waddr => x_rsc_22_0_i_s_waddr_1,
      s_din => x_rsc_22_0_i_s_din_1,
      s_dout => x_rsc_22_0_i_s_dout_1,
      s_rrdy => x_rsc_22_0_i_s_rrdy,
      s_wrdy => x_rsc_22_0_i_s_wrdy,
      is_idle => x_rsc_22_0_is_idle_1,
      tr_write_done => x_rsc_22_0_tr_write_done,
      s_tdone => x_rsc_22_0_s_tdone
    );
  x_rsc_22_0_i_AWID(0) <= x_rsc_22_0_AWID;
  x_rsc_22_0_i_AWADDR <= x_rsc_22_0_AWADDR;
  x_rsc_22_0_i_AWLEN <= x_rsc_22_0_AWLEN;
  x_rsc_22_0_i_AWSIZE <= x_rsc_22_0_AWSIZE;
  x_rsc_22_0_i_AWBURST <= x_rsc_22_0_AWBURST;
  x_rsc_22_0_i_AWCACHE <= x_rsc_22_0_AWCACHE;
  x_rsc_22_0_i_AWPROT <= x_rsc_22_0_AWPROT;
  x_rsc_22_0_i_AWQOS <= x_rsc_22_0_AWQOS;
  x_rsc_22_0_i_AWREGION <= x_rsc_22_0_AWREGION;
  x_rsc_22_0_i_AWUSER(0) <= x_rsc_22_0_AWUSER;
  x_rsc_22_0_i_WDATA <= x_rsc_22_0_WDATA;
  x_rsc_22_0_i_WSTRB <= x_rsc_22_0_WSTRB;
  x_rsc_22_0_i_WUSER(0) <= x_rsc_22_0_WUSER;
  x_rsc_22_0_BID <= x_rsc_22_0_i_BID(0);
  x_rsc_22_0_BRESP <= x_rsc_22_0_i_BRESP;
  x_rsc_22_0_BUSER <= x_rsc_22_0_i_BUSER(0);
  x_rsc_22_0_i_ARID(0) <= x_rsc_22_0_ARID;
  x_rsc_22_0_i_ARADDR <= x_rsc_22_0_ARADDR;
  x_rsc_22_0_i_ARLEN <= x_rsc_22_0_ARLEN;
  x_rsc_22_0_i_ARSIZE <= x_rsc_22_0_ARSIZE;
  x_rsc_22_0_i_ARBURST <= x_rsc_22_0_ARBURST;
  x_rsc_22_0_i_ARCACHE <= x_rsc_22_0_ARCACHE;
  x_rsc_22_0_i_ARPROT <= x_rsc_22_0_ARPROT;
  x_rsc_22_0_i_ARQOS <= x_rsc_22_0_ARQOS;
  x_rsc_22_0_i_ARREGION <= x_rsc_22_0_ARREGION;
  x_rsc_22_0_i_ARUSER(0) <= x_rsc_22_0_ARUSER;
  x_rsc_22_0_RID <= x_rsc_22_0_i_RID(0);
  x_rsc_22_0_RDATA <= x_rsc_22_0_i_RDATA;
  x_rsc_22_0_RRESP <= x_rsc_22_0_i_RRESP;
  x_rsc_22_0_RUSER <= x_rsc_22_0_i_RUSER(0);
  x_rsc_22_0_i_s_raddr_1 <= x_rsc_22_0_i_s_raddr;
  x_rsc_22_0_i_s_waddr_1 <= x_rsc_22_0_i_s_waddr;
  x_rsc_22_0_i_s_din <= x_rsc_22_0_i_s_din_1;
  x_rsc_22_0_i_s_dout_1 <= x_rsc_22_0_i_s_dout;

  hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl_inst : hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_22_0_i_oswt => x_rsc_22_0_i_oswt,
      x_rsc_22_0_i_oswt_1 => x_rsc_22_0_i_oswt_1,
      x_rsc_22_0_i_biwt => x_rsc_22_0_i_biwt,
      x_rsc_22_0_i_bdwt => x_rsc_22_0_i_bdwt,
      x_rsc_22_0_i_bcwt => x_rsc_22_0_i_bcwt,
      x_rsc_22_0_i_s_re_core_sct => x_rsc_22_0_i_s_re_core_sct,
      x_rsc_22_0_i_biwt_1 => x_rsc_22_0_i_biwt_1,
      x_rsc_22_0_i_bdwt_2 => x_rsc_22_0_i_bdwt_2,
      x_rsc_22_0_i_bcwt_1 => x_rsc_22_0_i_bcwt_1,
      x_rsc_22_0_i_s_we_core_sct => x_rsc_22_0_i_s_we_core_sct,
      x_rsc_22_0_i_s_rrdy => x_rsc_22_0_i_s_rrdy,
      x_rsc_22_0_i_s_wrdy => x_rsc_22_0_i_s_wrdy
    );
  hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst : hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_22_0_i_oswt => x_rsc_22_0_i_oswt,
      x_rsc_22_0_i_wen_comp => x_rsc_22_0_i_wen_comp,
      x_rsc_22_0_i_oswt_1 => x_rsc_22_0_i_oswt_1,
      x_rsc_22_0_i_wen_comp_1 => x_rsc_22_0_i_wen_comp_1,
      x_rsc_22_0_i_s_raddr_core => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_raddr_core,
      x_rsc_22_0_i_s_waddr_core => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_waddr_core,
      x_rsc_22_0_i_s_din_mxwt => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_din_mxwt,
      x_rsc_22_0_i_s_dout_core => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_dout_core,
      x_rsc_22_0_i_biwt => x_rsc_22_0_i_biwt,
      x_rsc_22_0_i_bdwt => x_rsc_22_0_i_bdwt,
      x_rsc_22_0_i_bcwt => x_rsc_22_0_i_bcwt,
      x_rsc_22_0_i_biwt_1 => x_rsc_22_0_i_biwt_1,
      x_rsc_22_0_i_bdwt_2 => x_rsc_22_0_i_bdwt_2,
      x_rsc_22_0_i_bcwt_1 => x_rsc_22_0_i_bcwt_1,
      x_rsc_22_0_i_s_raddr => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_raddr,
      x_rsc_22_0_i_s_raddr_core_sct => x_rsc_22_0_i_s_re_core_sct,
      x_rsc_22_0_i_s_waddr => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_waddr,
      x_rsc_22_0_i_s_waddr_core_sct => x_rsc_22_0_i_s_we_core_sct,
      x_rsc_22_0_i_s_din => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_din,
      x_rsc_22_0_i_s_dout => hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_dout
    );
  hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_raddr_core <= x_rsc_22_0_i_s_raddr_core;
  hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_waddr_core <= x_rsc_22_0_i_s_waddr_core;
  x_rsc_22_0_i_s_din_mxwt <= hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_din_mxwt;
  hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_dout_core <= x_rsc_22_0_i_s_dout_core;
  x_rsc_22_0_i_s_raddr <= hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_raddr;
  x_rsc_22_0_i_s_waddr <= hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_waddr;
  hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_din <= x_rsc_22_0_i_s_din;
  x_rsc_22_0_i_s_dout <= hybrid_core_x_rsc_22_0_i_x_rsc_22_0_wait_dp_inst_x_rsc_22_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_21_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_21_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_21_0_s_tdone : IN STD_LOGIC;
    x_rsc_21_0_tr_write_done : IN STD_LOGIC;
    x_rsc_21_0_RREADY : IN STD_LOGIC;
    x_rsc_21_0_RVALID : OUT STD_LOGIC;
    x_rsc_21_0_RUSER : OUT STD_LOGIC;
    x_rsc_21_0_RLAST : OUT STD_LOGIC;
    x_rsc_21_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_RID : OUT STD_LOGIC;
    x_rsc_21_0_ARREADY : OUT STD_LOGIC;
    x_rsc_21_0_ARVALID : IN STD_LOGIC;
    x_rsc_21_0_ARUSER : IN STD_LOGIC;
    x_rsc_21_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARLOCK : IN STD_LOGIC;
    x_rsc_21_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_21_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_21_0_ARID : IN STD_LOGIC;
    x_rsc_21_0_BREADY : IN STD_LOGIC;
    x_rsc_21_0_BVALID : OUT STD_LOGIC;
    x_rsc_21_0_BUSER : OUT STD_LOGIC;
    x_rsc_21_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_BID : OUT STD_LOGIC;
    x_rsc_21_0_WREADY : OUT STD_LOGIC;
    x_rsc_21_0_WVALID : IN STD_LOGIC;
    x_rsc_21_0_WUSER : IN STD_LOGIC;
    x_rsc_21_0_WLAST : IN STD_LOGIC;
    x_rsc_21_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_AWREADY : OUT STD_LOGIC;
    x_rsc_21_0_AWVALID : IN STD_LOGIC;
    x_rsc_21_0_AWUSER : IN STD_LOGIC;
    x_rsc_21_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWLOCK : IN STD_LOGIC;
    x_rsc_21_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_21_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_21_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_21_0_i_oswt : IN STD_LOGIC;
    x_rsc_21_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_21_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_21_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_21_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_21_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_21_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_21_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_21_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_21_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_21_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_21_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_21_0_i_oswt : IN STD_LOGIC;
      x_rsc_21_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_21_0_i_biwt : OUT STD_LOGIC;
      x_rsc_21_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_21_0_i_bcwt : IN STD_LOGIC;
      x_rsc_21_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_21_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_21_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_21_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_21_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_21_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_21_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_21_0_i_oswt : IN STD_LOGIC;
      x_rsc_21_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_21_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_21_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_21_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_21_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_21_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_i_biwt : IN STD_LOGIC;
      x_rsc_21_0_i_bdwt : IN STD_LOGIC;
      x_rsc_21_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_21_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_21_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_21_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_21_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_21_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_21_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_21_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_21_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_21_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_21_0_i_AWID,
      AWADDR => x_rsc_21_0_i_AWADDR,
      AWLEN => x_rsc_21_0_i_AWLEN,
      AWSIZE => x_rsc_21_0_i_AWSIZE,
      AWBURST => x_rsc_21_0_i_AWBURST,
      AWLOCK => x_rsc_21_0_AWLOCK,
      AWCACHE => x_rsc_21_0_i_AWCACHE,
      AWPROT => x_rsc_21_0_i_AWPROT,
      AWQOS => x_rsc_21_0_i_AWQOS,
      AWREGION => x_rsc_21_0_i_AWREGION,
      AWUSER => x_rsc_21_0_i_AWUSER,
      AWVALID => x_rsc_21_0_AWVALID,
      AWREADY => x_rsc_21_0_AWREADY,
      WDATA => x_rsc_21_0_i_WDATA,
      WSTRB => x_rsc_21_0_i_WSTRB,
      WLAST => x_rsc_21_0_WLAST,
      WUSER => x_rsc_21_0_i_WUSER,
      WVALID => x_rsc_21_0_WVALID,
      WREADY => x_rsc_21_0_WREADY,
      BID => x_rsc_21_0_i_BID,
      BRESP => x_rsc_21_0_i_BRESP,
      BUSER => x_rsc_21_0_i_BUSER,
      BVALID => x_rsc_21_0_BVALID,
      BREADY => x_rsc_21_0_BREADY,
      ARID => x_rsc_21_0_i_ARID,
      ARADDR => x_rsc_21_0_i_ARADDR,
      ARLEN => x_rsc_21_0_i_ARLEN,
      ARSIZE => x_rsc_21_0_i_ARSIZE,
      ARBURST => x_rsc_21_0_i_ARBURST,
      ARLOCK => x_rsc_21_0_ARLOCK,
      ARCACHE => x_rsc_21_0_i_ARCACHE,
      ARPROT => x_rsc_21_0_i_ARPROT,
      ARQOS => x_rsc_21_0_i_ARQOS,
      ARREGION => x_rsc_21_0_i_ARREGION,
      ARUSER => x_rsc_21_0_i_ARUSER,
      ARVALID => x_rsc_21_0_ARVALID,
      ARREADY => x_rsc_21_0_ARREADY,
      RID => x_rsc_21_0_i_RID,
      RDATA => x_rsc_21_0_i_RDATA,
      RRESP => x_rsc_21_0_i_RRESP,
      RLAST => x_rsc_21_0_RLAST,
      RUSER => x_rsc_21_0_i_RUSER,
      RVALID => x_rsc_21_0_RVALID,
      RREADY => x_rsc_21_0_RREADY,
      s_re => x_rsc_21_0_i_s_re_core_sct,
      s_we => x_rsc_21_0_i_s_we_core_sct,
      s_raddr => x_rsc_21_0_i_s_raddr_1,
      s_waddr => x_rsc_21_0_i_s_waddr_1,
      s_din => x_rsc_21_0_i_s_din_1,
      s_dout => x_rsc_21_0_i_s_dout_1,
      s_rrdy => x_rsc_21_0_i_s_rrdy,
      s_wrdy => x_rsc_21_0_i_s_wrdy,
      is_idle => x_rsc_21_0_is_idle_1,
      tr_write_done => x_rsc_21_0_tr_write_done,
      s_tdone => x_rsc_21_0_s_tdone
    );
  x_rsc_21_0_i_AWID(0) <= x_rsc_21_0_AWID;
  x_rsc_21_0_i_AWADDR <= x_rsc_21_0_AWADDR;
  x_rsc_21_0_i_AWLEN <= x_rsc_21_0_AWLEN;
  x_rsc_21_0_i_AWSIZE <= x_rsc_21_0_AWSIZE;
  x_rsc_21_0_i_AWBURST <= x_rsc_21_0_AWBURST;
  x_rsc_21_0_i_AWCACHE <= x_rsc_21_0_AWCACHE;
  x_rsc_21_0_i_AWPROT <= x_rsc_21_0_AWPROT;
  x_rsc_21_0_i_AWQOS <= x_rsc_21_0_AWQOS;
  x_rsc_21_0_i_AWREGION <= x_rsc_21_0_AWREGION;
  x_rsc_21_0_i_AWUSER(0) <= x_rsc_21_0_AWUSER;
  x_rsc_21_0_i_WDATA <= x_rsc_21_0_WDATA;
  x_rsc_21_0_i_WSTRB <= x_rsc_21_0_WSTRB;
  x_rsc_21_0_i_WUSER(0) <= x_rsc_21_0_WUSER;
  x_rsc_21_0_BID <= x_rsc_21_0_i_BID(0);
  x_rsc_21_0_BRESP <= x_rsc_21_0_i_BRESP;
  x_rsc_21_0_BUSER <= x_rsc_21_0_i_BUSER(0);
  x_rsc_21_0_i_ARID(0) <= x_rsc_21_0_ARID;
  x_rsc_21_0_i_ARADDR <= x_rsc_21_0_ARADDR;
  x_rsc_21_0_i_ARLEN <= x_rsc_21_0_ARLEN;
  x_rsc_21_0_i_ARSIZE <= x_rsc_21_0_ARSIZE;
  x_rsc_21_0_i_ARBURST <= x_rsc_21_0_ARBURST;
  x_rsc_21_0_i_ARCACHE <= x_rsc_21_0_ARCACHE;
  x_rsc_21_0_i_ARPROT <= x_rsc_21_0_ARPROT;
  x_rsc_21_0_i_ARQOS <= x_rsc_21_0_ARQOS;
  x_rsc_21_0_i_ARREGION <= x_rsc_21_0_ARREGION;
  x_rsc_21_0_i_ARUSER(0) <= x_rsc_21_0_ARUSER;
  x_rsc_21_0_RID <= x_rsc_21_0_i_RID(0);
  x_rsc_21_0_RDATA <= x_rsc_21_0_i_RDATA;
  x_rsc_21_0_RRESP <= x_rsc_21_0_i_RRESP;
  x_rsc_21_0_RUSER <= x_rsc_21_0_i_RUSER(0);
  x_rsc_21_0_i_s_raddr_1 <= x_rsc_21_0_i_s_raddr;
  x_rsc_21_0_i_s_waddr_1 <= x_rsc_21_0_i_s_waddr;
  x_rsc_21_0_i_s_din <= x_rsc_21_0_i_s_din_1;
  x_rsc_21_0_i_s_dout_1 <= x_rsc_21_0_i_s_dout;

  hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl_inst : hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_21_0_i_oswt => x_rsc_21_0_i_oswt,
      x_rsc_21_0_i_oswt_1 => x_rsc_21_0_i_oswt_1,
      x_rsc_21_0_i_biwt => x_rsc_21_0_i_biwt,
      x_rsc_21_0_i_bdwt => x_rsc_21_0_i_bdwt,
      x_rsc_21_0_i_bcwt => x_rsc_21_0_i_bcwt,
      x_rsc_21_0_i_s_re_core_sct => x_rsc_21_0_i_s_re_core_sct,
      x_rsc_21_0_i_biwt_1 => x_rsc_21_0_i_biwt_1,
      x_rsc_21_0_i_bdwt_2 => x_rsc_21_0_i_bdwt_2,
      x_rsc_21_0_i_bcwt_1 => x_rsc_21_0_i_bcwt_1,
      x_rsc_21_0_i_s_we_core_sct => x_rsc_21_0_i_s_we_core_sct,
      x_rsc_21_0_i_s_rrdy => x_rsc_21_0_i_s_rrdy,
      x_rsc_21_0_i_s_wrdy => x_rsc_21_0_i_s_wrdy
    );
  hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst : hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_21_0_i_oswt => x_rsc_21_0_i_oswt,
      x_rsc_21_0_i_wen_comp => x_rsc_21_0_i_wen_comp,
      x_rsc_21_0_i_oswt_1 => x_rsc_21_0_i_oswt_1,
      x_rsc_21_0_i_wen_comp_1 => x_rsc_21_0_i_wen_comp_1,
      x_rsc_21_0_i_s_raddr_core => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_raddr_core,
      x_rsc_21_0_i_s_waddr_core => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_waddr_core,
      x_rsc_21_0_i_s_din_mxwt => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_din_mxwt,
      x_rsc_21_0_i_s_dout_core => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_dout_core,
      x_rsc_21_0_i_biwt => x_rsc_21_0_i_biwt,
      x_rsc_21_0_i_bdwt => x_rsc_21_0_i_bdwt,
      x_rsc_21_0_i_bcwt => x_rsc_21_0_i_bcwt,
      x_rsc_21_0_i_biwt_1 => x_rsc_21_0_i_biwt_1,
      x_rsc_21_0_i_bdwt_2 => x_rsc_21_0_i_bdwt_2,
      x_rsc_21_0_i_bcwt_1 => x_rsc_21_0_i_bcwt_1,
      x_rsc_21_0_i_s_raddr => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_raddr,
      x_rsc_21_0_i_s_raddr_core_sct => x_rsc_21_0_i_s_re_core_sct,
      x_rsc_21_0_i_s_waddr => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_waddr,
      x_rsc_21_0_i_s_waddr_core_sct => x_rsc_21_0_i_s_we_core_sct,
      x_rsc_21_0_i_s_din => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_din,
      x_rsc_21_0_i_s_dout => hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_dout
    );
  hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_raddr_core <= x_rsc_21_0_i_s_raddr_core;
  hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_waddr_core <= x_rsc_21_0_i_s_waddr_core;
  x_rsc_21_0_i_s_din_mxwt <= hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_din_mxwt;
  hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_dout_core <= x_rsc_21_0_i_s_dout_core;
  x_rsc_21_0_i_s_raddr <= hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_raddr;
  x_rsc_21_0_i_s_waddr <= hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_waddr;
  hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_din <= x_rsc_21_0_i_s_din;
  x_rsc_21_0_i_s_dout <= hybrid_core_x_rsc_21_0_i_x_rsc_21_0_wait_dp_inst_x_rsc_21_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_20_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_20_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_20_0_s_tdone : IN STD_LOGIC;
    x_rsc_20_0_tr_write_done : IN STD_LOGIC;
    x_rsc_20_0_RREADY : IN STD_LOGIC;
    x_rsc_20_0_RVALID : OUT STD_LOGIC;
    x_rsc_20_0_RUSER : OUT STD_LOGIC;
    x_rsc_20_0_RLAST : OUT STD_LOGIC;
    x_rsc_20_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_RID : OUT STD_LOGIC;
    x_rsc_20_0_ARREADY : OUT STD_LOGIC;
    x_rsc_20_0_ARVALID : IN STD_LOGIC;
    x_rsc_20_0_ARUSER : IN STD_LOGIC;
    x_rsc_20_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARLOCK : IN STD_LOGIC;
    x_rsc_20_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_20_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_20_0_ARID : IN STD_LOGIC;
    x_rsc_20_0_BREADY : IN STD_LOGIC;
    x_rsc_20_0_BVALID : OUT STD_LOGIC;
    x_rsc_20_0_BUSER : OUT STD_LOGIC;
    x_rsc_20_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_BID : OUT STD_LOGIC;
    x_rsc_20_0_WREADY : OUT STD_LOGIC;
    x_rsc_20_0_WVALID : IN STD_LOGIC;
    x_rsc_20_0_WUSER : IN STD_LOGIC;
    x_rsc_20_0_WLAST : IN STD_LOGIC;
    x_rsc_20_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_AWREADY : OUT STD_LOGIC;
    x_rsc_20_0_AWVALID : IN STD_LOGIC;
    x_rsc_20_0_AWUSER : IN STD_LOGIC;
    x_rsc_20_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWLOCK : IN STD_LOGIC;
    x_rsc_20_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_20_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_20_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_20_0_i_oswt : IN STD_LOGIC;
    x_rsc_20_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_20_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_20_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_20_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_20_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_20_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_20_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_20_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_20_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_20_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_20_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_20_0_i_oswt : IN STD_LOGIC;
      x_rsc_20_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_20_0_i_biwt : OUT STD_LOGIC;
      x_rsc_20_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_20_0_i_bcwt : IN STD_LOGIC;
      x_rsc_20_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_20_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_20_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_20_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_20_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_20_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_20_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_20_0_i_oswt : IN STD_LOGIC;
      x_rsc_20_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_20_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_20_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_20_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_20_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_20_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_i_biwt : IN STD_LOGIC;
      x_rsc_20_0_i_bdwt : IN STD_LOGIC;
      x_rsc_20_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_20_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_20_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_20_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_20_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_20_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_20_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_20_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_20_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_20_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_20_0_i_AWID,
      AWADDR => x_rsc_20_0_i_AWADDR,
      AWLEN => x_rsc_20_0_i_AWLEN,
      AWSIZE => x_rsc_20_0_i_AWSIZE,
      AWBURST => x_rsc_20_0_i_AWBURST,
      AWLOCK => x_rsc_20_0_AWLOCK,
      AWCACHE => x_rsc_20_0_i_AWCACHE,
      AWPROT => x_rsc_20_0_i_AWPROT,
      AWQOS => x_rsc_20_0_i_AWQOS,
      AWREGION => x_rsc_20_0_i_AWREGION,
      AWUSER => x_rsc_20_0_i_AWUSER,
      AWVALID => x_rsc_20_0_AWVALID,
      AWREADY => x_rsc_20_0_AWREADY,
      WDATA => x_rsc_20_0_i_WDATA,
      WSTRB => x_rsc_20_0_i_WSTRB,
      WLAST => x_rsc_20_0_WLAST,
      WUSER => x_rsc_20_0_i_WUSER,
      WVALID => x_rsc_20_0_WVALID,
      WREADY => x_rsc_20_0_WREADY,
      BID => x_rsc_20_0_i_BID,
      BRESP => x_rsc_20_0_i_BRESP,
      BUSER => x_rsc_20_0_i_BUSER,
      BVALID => x_rsc_20_0_BVALID,
      BREADY => x_rsc_20_0_BREADY,
      ARID => x_rsc_20_0_i_ARID,
      ARADDR => x_rsc_20_0_i_ARADDR,
      ARLEN => x_rsc_20_0_i_ARLEN,
      ARSIZE => x_rsc_20_0_i_ARSIZE,
      ARBURST => x_rsc_20_0_i_ARBURST,
      ARLOCK => x_rsc_20_0_ARLOCK,
      ARCACHE => x_rsc_20_0_i_ARCACHE,
      ARPROT => x_rsc_20_0_i_ARPROT,
      ARQOS => x_rsc_20_0_i_ARQOS,
      ARREGION => x_rsc_20_0_i_ARREGION,
      ARUSER => x_rsc_20_0_i_ARUSER,
      ARVALID => x_rsc_20_0_ARVALID,
      ARREADY => x_rsc_20_0_ARREADY,
      RID => x_rsc_20_0_i_RID,
      RDATA => x_rsc_20_0_i_RDATA,
      RRESP => x_rsc_20_0_i_RRESP,
      RLAST => x_rsc_20_0_RLAST,
      RUSER => x_rsc_20_0_i_RUSER,
      RVALID => x_rsc_20_0_RVALID,
      RREADY => x_rsc_20_0_RREADY,
      s_re => x_rsc_20_0_i_s_re_core_sct,
      s_we => x_rsc_20_0_i_s_we_core_sct,
      s_raddr => x_rsc_20_0_i_s_raddr_1,
      s_waddr => x_rsc_20_0_i_s_waddr_1,
      s_din => x_rsc_20_0_i_s_din_1,
      s_dout => x_rsc_20_0_i_s_dout_1,
      s_rrdy => x_rsc_20_0_i_s_rrdy,
      s_wrdy => x_rsc_20_0_i_s_wrdy,
      is_idle => x_rsc_20_0_is_idle_1,
      tr_write_done => x_rsc_20_0_tr_write_done,
      s_tdone => x_rsc_20_0_s_tdone
    );
  x_rsc_20_0_i_AWID(0) <= x_rsc_20_0_AWID;
  x_rsc_20_0_i_AWADDR <= x_rsc_20_0_AWADDR;
  x_rsc_20_0_i_AWLEN <= x_rsc_20_0_AWLEN;
  x_rsc_20_0_i_AWSIZE <= x_rsc_20_0_AWSIZE;
  x_rsc_20_0_i_AWBURST <= x_rsc_20_0_AWBURST;
  x_rsc_20_0_i_AWCACHE <= x_rsc_20_0_AWCACHE;
  x_rsc_20_0_i_AWPROT <= x_rsc_20_0_AWPROT;
  x_rsc_20_0_i_AWQOS <= x_rsc_20_0_AWQOS;
  x_rsc_20_0_i_AWREGION <= x_rsc_20_0_AWREGION;
  x_rsc_20_0_i_AWUSER(0) <= x_rsc_20_0_AWUSER;
  x_rsc_20_0_i_WDATA <= x_rsc_20_0_WDATA;
  x_rsc_20_0_i_WSTRB <= x_rsc_20_0_WSTRB;
  x_rsc_20_0_i_WUSER(0) <= x_rsc_20_0_WUSER;
  x_rsc_20_0_BID <= x_rsc_20_0_i_BID(0);
  x_rsc_20_0_BRESP <= x_rsc_20_0_i_BRESP;
  x_rsc_20_0_BUSER <= x_rsc_20_0_i_BUSER(0);
  x_rsc_20_0_i_ARID(0) <= x_rsc_20_0_ARID;
  x_rsc_20_0_i_ARADDR <= x_rsc_20_0_ARADDR;
  x_rsc_20_0_i_ARLEN <= x_rsc_20_0_ARLEN;
  x_rsc_20_0_i_ARSIZE <= x_rsc_20_0_ARSIZE;
  x_rsc_20_0_i_ARBURST <= x_rsc_20_0_ARBURST;
  x_rsc_20_0_i_ARCACHE <= x_rsc_20_0_ARCACHE;
  x_rsc_20_0_i_ARPROT <= x_rsc_20_0_ARPROT;
  x_rsc_20_0_i_ARQOS <= x_rsc_20_0_ARQOS;
  x_rsc_20_0_i_ARREGION <= x_rsc_20_0_ARREGION;
  x_rsc_20_0_i_ARUSER(0) <= x_rsc_20_0_ARUSER;
  x_rsc_20_0_RID <= x_rsc_20_0_i_RID(0);
  x_rsc_20_0_RDATA <= x_rsc_20_0_i_RDATA;
  x_rsc_20_0_RRESP <= x_rsc_20_0_i_RRESP;
  x_rsc_20_0_RUSER <= x_rsc_20_0_i_RUSER(0);
  x_rsc_20_0_i_s_raddr_1 <= x_rsc_20_0_i_s_raddr;
  x_rsc_20_0_i_s_waddr_1 <= x_rsc_20_0_i_s_waddr;
  x_rsc_20_0_i_s_din <= x_rsc_20_0_i_s_din_1;
  x_rsc_20_0_i_s_dout_1 <= x_rsc_20_0_i_s_dout;

  hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl_inst : hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_20_0_i_oswt => x_rsc_20_0_i_oswt,
      x_rsc_20_0_i_oswt_1 => x_rsc_20_0_i_oswt_1,
      x_rsc_20_0_i_biwt => x_rsc_20_0_i_biwt,
      x_rsc_20_0_i_bdwt => x_rsc_20_0_i_bdwt,
      x_rsc_20_0_i_bcwt => x_rsc_20_0_i_bcwt,
      x_rsc_20_0_i_s_re_core_sct => x_rsc_20_0_i_s_re_core_sct,
      x_rsc_20_0_i_biwt_1 => x_rsc_20_0_i_biwt_1,
      x_rsc_20_0_i_bdwt_2 => x_rsc_20_0_i_bdwt_2,
      x_rsc_20_0_i_bcwt_1 => x_rsc_20_0_i_bcwt_1,
      x_rsc_20_0_i_s_we_core_sct => x_rsc_20_0_i_s_we_core_sct,
      x_rsc_20_0_i_s_rrdy => x_rsc_20_0_i_s_rrdy,
      x_rsc_20_0_i_s_wrdy => x_rsc_20_0_i_s_wrdy
    );
  hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst : hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_20_0_i_oswt => x_rsc_20_0_i_oswt,
      x_rsc_20_0_i_wen_comp => x_rsc_20_0_i_wen_comp,
      x_rsc_20_0_i_oswt_1 => x_rsc_20_0_i_oswt_1,
      x_rsc_20_0_i_wen_comp_1 => x_rsc_20_0_i_wen_comp_1,
      x_rsc_20_0_i_s_raddr_core => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_raddr_core,
      x_rsc_20_0_i_s_waddr_core => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_waddr_core,
      x_rsc_20_0_i_s_din_mxwt => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_din_mxwt,
      x_rsc_20_0_i_s_dout_core => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_dout_core,
      x_rsc_20_0_i_biwt => x_rsc_20_0_i_biwt,
      x_rsc_20_0_i_bdwt => x_rsc_20_0_i_bdwt,
      x_rsc_20_0_i_bcwt => x_rsc_20_0_i_bcwt,
      x_rsc_20_0_i_biwt_1 => x_rsc_20_0_i_biwt_1,
      x_rsc_20_0_i_bdwt_2 => x_rsc_20_0_i_bdwt_2,
      x_rsc_20_0_i_bcwt_1 => x_rsc_20_0_i_bcwt_1,
      x_rsc_20_0_i_s_raddr => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_raddr,
      x_rsc_20_0_i_s_raddr_core_sct => x_rsc_20_0_i_s_re_core_sct,
      x_rsc_20_0_i_s_waddr => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_waddr,
      x_rsc_20_0_i_s_waddr_core_sct => x_rsc_20_0_i_s_we_core_sct,
      x_rsc_20_0_i_s_din => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_din,
      x_rsc_20_0_i_s_dout => hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_dout
    );
  hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_raddr_core <= x_rsc_20_0_i_s_raddr_core;
  hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_waddr_core <= x_rsc_20_0_i_s_waddr_core;
  x_rsc_20_0_i_s_din_mxwt <= hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_din_mxwt;
  hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_dout_core <= x_rsc_20_0_i_s_dout_core;
  x_rsc_20_0_i_s_raddr <= hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_raddr;
  x_rsc_20_0_i_s_waddr <= hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_waddr;
  hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_din <= x_rsc_20_0_i_s_din;
  x_rsc_20_0_i_s_dout <= hybrid_core_x_rsc_20_0_i_x_rsc_20_0_wait_dp_inst_x_rsc_20_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_19_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_19_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_19_0_s_tdone : IN STD_LOGIC;
    x_rsc_19_0_tr_write_done : IN STD_LOGIC;
    x_rsc_19_0_RREADY : IN STD_LOGIC;
    x_rsc_19_0_RVALID : OUT STD_LOGIC;
    x_rsc_19_0_RUSER : OUT STD_LOGIC;
    x_rsc_19_0_RLAST : OUT STD_LOGIC;
    x_rsc_19_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_RID : OUT STD_LOGIC;
    x_rsc_19_0_ARREADY : OUT STD_LOGIC;
    x_rsc_19_0_ARVALID : IN STD_LOGIC;
    x_rsc_19_0_ARUSER : IN STD_LOGIC;
    x_rsc_19_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARLOCK : IN STD_LOGIC;
    x_rsc_19_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_19_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_19_0_ARID : IN STD_LOGIC;
    x_rsc_19_0_BREADY : IN STD_LOGIC;
    x_rsc_19_0_BVALID : OUT STD_LOGIC;
    x_rsc_19_0_BUSER : OUT STD_LOGIC;
    x_rsc_19_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_BID : OUT STD_LOGIC;
    x_rsc_19_0_WREADY : OUT STD_LOGIC;
    x_rsc_19_0_WVALID : IN STD_LOGIC;
    x_rsc_19_0_WUSER : IN STD_LOGIC;
    x_rsc_19_0_WLAST : IN STD_LOGIC;
    x_rsc_19_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_AWREADY : OUT STD_LOGIC;
    x_rsc_19_0_AWVALID : IN STD_LOGIC;
    x_rsc_19_0_AWUSER : IN STD_LOGIC;
    x_rsc_19_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWLOCK : IN STD_LOGIC;
    x_rsc_19_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_19_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_19_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_19_0_i_oswt : IN STD_LOGIC;
    x_rsc_19_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_19_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_19_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_19_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_19_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_19_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_19_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_19_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_19_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_19_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_19_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_19_0_i_oswt : IN STD_LOGIC;
      x_rsc_19_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_19_0_i_biwt : OUT STD_LOGIC;
      x_rsc_19_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_19_0_i_bcwt : IN STD_LOGIC;
      x_rsc_19_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_19_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_19_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_19_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_19_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_19_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_19_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_19_0_i_oswt : IN STD_LOGIC;
      x_rsc_19_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_19_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_19_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_19_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_19_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_19_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_i_biwt : IN STD_LOGIC;
      x_rsc_19_0_i_bdwt : IN STD_LOGIC;
      x_rsc_19_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_19_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_19_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_19_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_19_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_19_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_19_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_19_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_19_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_19_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_19_0_i_AWID,
      AWADDR => x_rsc_19_0_i_AWADDR,
      AWLEN => x_rsc_19_0_i_AWLEN,
      AWSIZE => x_rsc_19_0_i_AWSIZE,
      AWBURST => x_rsc_19_0_i_AWBURST,
      AWLOCK => x_rsc_19_0_AWLOCK,
      AWCACHE => x_rsc_19_0_i_AWCACHE,
      AWPROT => x_rsc_19_0_i_AWPROT,
      AWQOS => x_rsc_19_0_i_AWQOS,
      AWREGION => x_rsc_19_0_i_AWREGION,
      AWUSER => x_rsc_19_0_i_AWUSER,
      AWVALID => x_rsc_19_0_AWVALID,
      AWREADY => x_rsc_19_0_AWREADY,
      WDATA => x_rsc_19_0_i_WDATA,
      WSTRB => x_rsc_19_0_i_WSTRB,
      WLAST => x_rsc_19_0_WLAST,
      WUSER => x_rsc_19_0_i_WUSER,
      WVALID => x_rsc_19_0_WVALID,
      WREADY => x_rsc_19_0_WREADY,
      BID => x_rsc_19_0_i_BID,
      BRESP => x_rsc_19_0_i_BRESP,
      BUSER => x_rsc_19_0_i_BUSER,
      BVALID => x_rsc_19_0_BVALID,
      BREADY => x_rsc_19_0_BREADY,
      ARID => x_rsc_19_0_i_ARID,
      ARADDR => x_rsc_19_0_i_ARADDR,
      ARLEN => x_rsc_19_0_i_ARLEN,
      ARSIZE => x_rsc_19_0_i_ARSIZE,
      ARBURST => x_rsc_19_0_i_ARBURST,
      ARLOCK => x_rsc_19_0_ARLOCK,
      ARCACHE => x_rsc_19_0_i_ARCACHE,
      ARPROT => x_rsc_19_0_i_ARPROT,
      ARQOS => x_rsc_19_0_i_ARQOS,
      ARREGION => x_rsc_19_0_i_ARREGION,
      ARUSER => x_rsc_19_0_i_ARUSER,
      ARVALID => x_rsc_19_0_ARVALID,
      ARREADY => x_rsc_19_0_ARREADY,
      RID => x_rsc_19_0_i_RID,
      RDATA => x_rsc_19_0_i_RDATA,
      RRESP => x_rsc_19_0_i_RRESP,
      RLAST => x_rsc_19_0_RLAST,
      RUSER => x_rsc_19_0_i_RUSER,
      RVALID => x_rsc_19_0_RVALID,
      RREADY => x_rsc_19_0_RREADY,
      s_re => x_rsc_19_0_i_s_re_core_sct,
      s_we => x_rsc_19_0_i_s_we_core_sct,
      s_raddr => x_rsc_19_0_i_s_raddr_1,
      s_waddr => x_rsc_19_0_i_s_waddr_1,
      s_din => x_rsc_19_0_i_s_din_1,
      s_dout => x_rsc_19_0_i_s_dout_1,
      s_rrdy => x_rsc_19_0_i_s_rrdy,
      s_wrdy => x_rsc_19_0_i_s_wrdy,
      is_idle => x_rsc_19_0_is_idle_1,
      tr_write_done => x_rsc_19_0_tr_write_done,
      s_tdone => x_rsc_19_0_s_tdone
    );
  x_rsc_19_0_i_AWID(0) <= x_rsc_19_0_AWID;
  x_rsc_19_0_i_AWADDR <= x_rsc_19_0_AWADDR;
  x_rsc_19_0_i_AWLEN <= x_rsc_19_0_AWLEN;
  x_rsc_19_0_i_AWSIZE <= x_rsc_19_0_AWSIZE;
  x_rsc_19_0_i_AWBURST <= x_rsc_19_0_AWBURST;
  x_rsc_19_0_i_AWCACHE <= x_rsc_19_0_AWCACHE;
  x_rsc_19_0_i_AWPROT <= x_rsc_19_0_AWPROT;
  x_rsc_19_0_i_AWQOS <= x_rsc_19_0_AWQOS;
  x_rsc_19_0_i_AWREGION <= x_rsc_19_0_AWREGION;
  x_rsc_19_0_i_AWUSER(0) <= x_rsc_19_0_AWUSER;
  x_rsc_19_0_i_WDATA <= x_rsc_19_0_WDATA;
  x_rsc_19_0_i_WSTRB <= x_rsc_19_0_WSTRB;
  x_rsc_19_0_i_WUSER(0) <= x_rsc_19_0_WUSER;
  x_rsc_19_0_BID <= x_rsc_19_0_i_BID(0);
  x_rsc_19_0_BRESP <= x_rsc_19_0_i_BRESP;
  x_rsc_19_0_BUSER <= x_rsc_19_0_i_BUSER(0);
  x_rsc_19_0_i_ARID(0) <= x_rsc_19_0_ARID;
  x_rsc_19_0_i_ARADDR <= x_rsc_19_0_ARADDR;
  x_rsc_19_0_i_ARLEN <= x_rsc_19_0_ARLEN;
  x_rsc_19_0_i_ARSIZE <= x_rsc_19_0_ARSIZE;
  x_rsc_19_0_i_ARBURST <= x_rsc_19_0_ARBURST;
  x_rsc_19_0_i_ARCACHE <= x_rsc_19_0_ARCACHE;
  x_rsc_19_0_i_ARPROT <= x_rsc_19_0_ARPROT;
  x_rsc_19_0_i_ARQOS <= x_rsc_19_0_ARQOS;
  x_rsc_19_0_i_ARREGION <= x_rsc_19_0_ARREGION;
  x_rsc_19_0_i_ARUSER(0) <= x_rsc_19_0_ARUSER;
  x_rsc_19_0_RID <= x_rsc_19_0_i_RID(0);
  x_rsc_19_0_RDATA <= x_rsc_19_0_i_RDATA;
  x_rsc_19_0_RRESP <= x_rsc_19_0_i_RRESP;
  x_rsc_19_0_RUSER <= x_rsc_19_0_i_RUSER(0);
  x_rsc_19_0_i_s_raddr_1 <= x_rsc_19_0_i_s_raddr;
  x_rsc_19_0_i_s_waddr_1 <= x_rsc_19_0_i_s_waddr;
  x_rsc_19_0_i_s_din <= x_rsc_19_0_i_s_din_1;
  x_rsc_19_0_i_s_dout_1 <= x_rsc_19_0_i_s_dout;

  hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl_inst : hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_19_0_i_oswt => x_rsc_19_0_i_oswt,
      x_rsc_19_0_i_oswt_1 => x_rsc_19_0_i_oswt_1,
      x_rsc_19_0_i_biwt => x_rsc_19_0_i_biwt,
      x_rsc_19_0_i_bdwt => x_rsc_19_0_i_bdwt,
      x_rsc_19_0_i_bcwt => x_rsc_19_0_i_bcwt,
      x_rsc_19_0_i_s_re_core_sct => x_rsc_19_0_i_s_re_core_sct,
      x_rsc_19_0_i_biwt_1 => x_rsc_19_0_i_biwt_1,
      x_rsc_19_0_i_bdwt_2 => x_rsc_19_0_i_bdwt_2,
      x_rsc_19_0_i_bcwt_1 => x_rsc_19_0_i_bcwt_1,
      x_rsc_19_0_i_s_we_core_sct => x_rsc_19_0_i_s_we_core_sct,
      x_rsc_19_0_i_s_rrdy => x_rsc_19_0_i_s_rrdy,
      x_rsc_19_0_i_s_wrdy => x_rsc_19_0_i_s_wrdy
    );
  hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst : hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_19_0_i_oswt => x_rsc_19_0_i_oswt,
      x_rsc_19_0_i_wen_comp => x_rsc_19_0_i_wen_comp,
      x_rsc_19_0_i_oswt_1 => x_rsc_19_0_i_oswt_1,
      x_rsc_19_0_i_wen_comp_1 => x_rsc_19_0_i_wen_comp_1,
      x_rsc_19_0_i_s_raddr_core => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_raddr_core,
      x_rsc_19_0_i_s_waddr_core => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_waddr_core,
      x_rsc_19_0_i_s_din_mxwt => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_din_mxwt,
      x_rsc_19_0_i_s_dout_core => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_dout_core,
      x_rsc_19_0_i_biwt => x_rsc_19_0_i_biwt,
      x_rsc_19_0_i_bdwt => x_rsc_19_0_i_bdwt,
      x_rsc_19_0_i_bcwt => x_rsc_19_0_i_bcwt,
      x_rsc_19_0_i_biwt_1 => x_rsc_19_0_i_biwt_1,
      x_rsc_19_0_i_bdwt_2 => x_rsc_19_0_i_bdwt_2,
      x_rsc_19_0_i_bcwt_1 => x_rsc_19_0_i_bcwt_1,
      x_rsc_19_0_i_s_raddr => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_raddr,
      x_rsc_19_0_i_s_raddr_core_sct => x_rsc_19_0_i_s_re_core_sct,
      x_rsc_19_0_i_s_waddr => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_waddr,
      x_rsc_19_0_i_s_waddr_core_sct => x_rsc_19_0_i_s_we_core_sct,
      x_rsc_19_0_i_s_din => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_din,
      x_rsc_19_0_i_s_dout => hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_dout
    );
  hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_raddr_core <= x_rsc_19_0_i_s_raddr_core;
  hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_waddr_core <= x_rsc_19_0_i_s_waddr_core;
  x_rsc_19_0_i_s_din_mxwt <= hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_din_mxwt;
  hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_dout_core <= x_rsc_19_0_i_s_dout_core;
  x_rsc_19_0_i_s_raddr <= hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_raddr;
  x_rsc_19_0_i_s_waddr <= hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_waddr;
  hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_din <= x_rsc_19_0_i_s_din;
  x_rsc_19_0_i_s_dout <= hybrid_core_x_rsc_19_0_i_x_rsc_19_0_wait_dp_inst_x_rsc_19_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_18_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_18_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_18_0_s_tdone : IN STD_LOGIC;
    x_rsc_18_0_tr_write_done : IN STD_LOGIC;
    x_rsc_18_0_RREADY : IN STD_LOGIC;
    x_rsc_18_0_RVALID : OUT STD_LOGIC;
    x_rsc_18_0_RUSER : OUT STD_LOGIC;
    x_rsc_18_0_RLAST : OUT STD_LOGIC;
    x_rsc_18_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_RID : OUT STD_LOGIC;
    x_rsc_18_0_ARREADY : OUT STD_LOGIC;
    x_rsc_18_0_ARVALID : IN STD_LOGIC;
    x_rsc_18_0_ARUSER : IN STD_LOGIC;
    x_rsc_18_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARLOCK : IN STD_LOGIC;
    x_rsc_18_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_18_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_18_0_ARID : IN STD_LOGIC;
    x_rsc_18_0_BREADY : IN STD_LOGIC;
    x_rsc_18_0_BVALID : OUT STD_LOGIC;
    x_rsc_18_0_BUSER : OUT STD_LOGIC;
    x_rsc_18_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_BID : OUT STD_LOGIC;
    x_rsc_18_0_WREADY : OUT STD_LOGIC;
    x_rsc_18_0_WVALID : IN STD_LOGIC;
    x_rsc_18_0_WUSER : IN STD_LOGIC;
    x_rsc_18_0_WLAST : IN STD_LOGIC;
    x_rsc_18_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_AWREADY : OUT STD_LOGIC;
    x_rsc_18_0_AWVALID : IN STD_LOGIC;
    x_rsc_18_0_AWUSER : IN STD_LOGIC;
    x_rsc_18_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWLOCK : IN STD_LOGIC;
    x_rsc_18_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_18_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_18_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_18_0_i_oswt : IN STD_LOGIC;
    x_rsc_18_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_18_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_18_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_18_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_18_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_18_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_18_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_18_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_18_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_18_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_18_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_18_0_i_oswt : IN STD_LOGIC;
      x_rsc_18_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_18_0_i_biwt : OUT STD_LOGIC;
      x_rsc_18_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_18_0_i_bcwt : IN STD_LOGIC;
      x_rsc_18_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_18_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_18_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_18_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_18_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_18_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_18_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_18_0_i_oswt : IN STD_LOGIC;
      x_rsc_18_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_18_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_18_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_18_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_18_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_18_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_i_biwt : IN STD_LOGIC;
      x_rsc_18_0_i_bdwt : IN STD_LOGIC;
      x_rsc_18_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_18_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_18_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_18_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_18_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_18_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_18_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_18_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_18_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_18_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_18_0_i_AWID,
      AWADDR => x_rsc_18_0_i_AWADDR,
      AWLEN => x_rsc_18_0_i_AWLEN,
      AWSIZE => x_rsc_18_0_i_AWSIZE,
      AWBURST => x_rsc_18_0_i_AWBURST,
      AWLOCK => x_rsc_18_0_AWLOCK,
      AWCACHE => x_rsc_18_0_i_AWCACHE,
      AWPROT => x_rsc_18_0_i_AWPROT,
      AWQOS => x_rsc_18_0_i_AWQOS,
      AWREGION => x_rsc_18_0_i_AWREGION,
      AWUSER => x_rsc_18_0_i_AWUSER,
      AWVALID => x_rsc_18_0_AWVALID,
      AWREADY => x_rsc_18_0_AWREADY,
      WDATA => x_rsc_18_0_i_WDATA,
      WSTRB => x_rsc_18_0_i_WSTRB,
      WLAST => x_rsc_18_0_WLAST,
      WUSER => x_rsc_18_0_i_WUSER,
      WVALID => x_rsc_18_0_WVALID,
      WREADY => x_rsc_18_0_WREADY,
      BID => x_rsc_18_0_i_BID,
      BRESP => x_rsc_18_0_i_BRESP,
      BUSER => x_rsc_18_0_i_BUSER,
      BVALID => x_rsc_18_0_BVALID,
      BREADY => x_rsc_18_0_BREADY,
      ARID => x_rsc_18_0_i_ARID,
      ARADDR => x_rsc_18_0_i_ARADDR,
      ARLEN => x_rsc_18_0_i_ARLEN,
      ARSIZE => x_rsc_18_0_i_ARSIZE,
      ARBURST => x_rsc_18_0_i_ARBURST,
      ARLOCK => x_rsc_18_0_ARLOCK,
      ARCACHE => x_rsc_18_0_i_ARCACHE,
      ARPROT => x_rsc_18_0_i_ARPROT,
      ARQOS => x_rsc_18_0_i_ARQOS,
      ARREGION => x_rsc_18_0_i_ARREGION,
      ARUSER => x_rsc_18_0_i_ARUSER,
      ARVALID => x_rsc_18_0_ARVALID,
      ARREADY => x_rsc_18_0_ARREADY,
      RID => x_rsc_18_0_i_RID,
      RDATA => x_rsc_18_0_i_RDATA,
      RRESP => x_rsc_18_0_i_RRESP,
      RLAST => x_rsc_18_0_RLAST,
      RUSER => x_rsc_18_0_i_RUSER,
      RVALID => x_rsc_18_0_RVALID,
      RREADY => x_rsc_18_0_RREADY,
      s_re => x_rsc_18_0_i_s_re_core_sct,
      s_we => x_rsc_18_0_i_s_we_core_sct,
      s_raddr => x_rsc_18_0_i_s_raddr_1,
      s_waddr => x_rsc_18_0_i_s_waddr_1,
      s_din => x_rsc_18_0_i_s_din_1,
      s_dout => x_rsc_18_0_i_s_dout_1,
      s_rrdy => x_rsc_18_0_i_s_rrdy,
      s_wrdy => x_rsc_18_0_i_s_wrdy,
      is_idle => x_rsc_18_0_is_idle_1,
      tr_write_done => x_rsc_18_0_tr_write_done,
      s_tdone => x_rsc_18_0_s_tdone
    );
  x_rsc_18_0_i_AWID(0) <= x_rsc_18_0_AWID;
  x_rsc_18_0_i_AWADDR <= x_rsc_18_0_AWADDR;
  x_rsc_18_0_i_AWLEN <= x_rsc_18_0_AWLEN;
  x_rsc_18_0_i_AWSIZE <= x_rsc_18_0_AWSIZE;
  x_rsc_18_0_i_AWBURST <= x_rsc_18_0_AWBURST;
  x_rsc_18_0_i_AWCACHE <= x_rsc_18_0_AWCACHE;
  x_rsc_18_0_i_AWPROT <= x_rsc_18_0_AWPROT;
  x_rsc_18_0_i_AWQOS <= x_rsc_18_0_AWQOS;
  x_rsc_18_0_i_AWREGION <= x_rsc_18_0_AWREGION;
  x_rsc_18_0_i_AWUSER(0) <= x_rsc_18_0_AWUSER;
  x_rsc_18_0_i_WDATA <= x_rsc_18_0_WDATA;
  x_rsc_18_0_i_WSTRB <= x_rsc_18_0_WSTRB;
  x_rsc_18_0_i_WUSER(0) <= x_rsc_18_0_WUSER;
  x_rsc_18_0_BID <= x_rsc_18_0_i_BID(0);
  x_rsc_18_0_BRESP <= x_rsc_18_0_i_BRESP;
  x_rsc_18_0_BUSER <= x_rsc_18_0_i_BUSER(0);
  x_rsc_18_0_i_ARID(0) <= x_rsc_18_0_ARID;
  x_rsc_18_0_i_ARADDR <= x_rsc_18_0_ARADDR;
  x_rsc_18_0_i_ARLEN <= x_rsc_18_0_ARLEN;
  x_rsc_18_0_i_ARSIZE <= x_rsc_18_0_ARSIZE;
  x_rsc_18_0_i_ARBURST <= x_rsc_18_0_ARBURST;
  x_rsc_18_0_i_ARCACHE <= x_rsc_18_0_ARCACHE;
  x_rsc_18_0_i_ARPROT <= x_rsc_18_0_ARPROT;
  x_rsc_18_0_i_ARQOS <= x_rsc_18_0_ARQOS;
  x_rsc_18_0_i_ARREGION <= x_rsc_18_0_ARREGION;
  x_rsc_18_0_i_ARUSER(0) <= x_rsc_18_0_ARUSER;
  x_rsc_18_0_RID <= x_rsc_18_0_i_RID(0);
  x_rsc_18_0_RDATA <= x_rsc_18_0_i_RDATA;
  x_rsc_18_0_RRESP <= x_rsc_18_0_i_RRESP;
  x_rsc_18_0_RUSER <= x_rsc_18_0_i_RUSER(0);
  x_rsc_18_0_i_s_raddr_1 <= x_rsc_18_0_i_s_raddr;
  x_rsc_18_0_i_s_waddr_1 <= x_rsc_18_0_i_s_waddr;
  x_rsc_18_0_i_s_din <= x_rsc_18_0_i_s_din_1;
  x_rsc_18_0_i_s_dout_1 <= x_rsc_18_0_i_s_dout;

  hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl_inst : hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_18_0_i_oswt => x_rsc_18_0_i_oswt,
      x_rsc_18_0_i_oswt_1 => x_rsc_18_0_i_oswt_1,
      x_rsc_18_0_i_biwt => x_rsc_18_0_i_biwt,
      x_rsc_18_0_i_bdwt => x_rsc_18_0_i_bdwt,
      x_rsc_18_0_i_bcwt => x_rsc_18_0_i_bcwt,
      x_rsc_18_0_i_s_re_core_sct => x_rsc_18_0_i_s_re_core_sct,
      x_rsc_18_0_i_biwt_1 => x_rsc_18_0_i_biwt_1,
      x_rsc_18_0_i_bdwt_2 => x_rsc_18_0_i_bdwt_2,
      x_rsc_18_0_i_bcwt_1 => x_rsc_18_0_i_bcwt_1,
      x_rsc_18_0_i_s_we_core_sct => x_rsc_18_0_i_s_we_core_sct,
      x_rsc_18_0_i_s_rrdy => x_rsc_18_0_i_s_rrdy,
      x_rsc_18_0_i_s_wrdy => x_rsc_18_0_i_s_wrdy
    );
  hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst : hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_18_0_i_oswt => x_rsc_18_0_i_oswt,
      x_rsc_18_0_i_wen_comp => x_rsc_18_0_i_wen_comp,
      x_rsc_18_0_i_oswt_1 => x_rsc_18_0_i_oswt_1,
      x_rsc_18_0_i_wen_comp_1 => x_rsc_18_0_i_wen_comp_1,
      x_rsc_18_0_i_s_raddr_core => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_raddr_core,
      x_rsc_18_0_i_s_waddr_core => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_waddr_core,
      x_rsc_18_0_i_s_din_mxwt => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_din_mxwt,
      x_rsc_18_0_i_s_dout_core => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_dout_core,
      x_rsc_18_0_i_biwt => x_rsc_18_0_i_biwt,
      x_rsc_18_0_i_bdwt => x_rsc_18_0_i_bdwt,
      x_rsc_18_0_i_bcwt => x_rsc_18_0_i_bcwt,
      x_rsc_18_0_i_biwt_1 => x_rsc_18_0_i_biwt_1,
      x_rsc_18_0_i_bdwt_2 => x_rsc_18_0_i_bdwt_2,
      x_rsc_18_0_i_bcwt_1 => x_rsc_18_0_i_bcwt_1,
      x_rsc_18_0_i_s_raddr => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_raddr,
      x_rsc_18_0_i_s_raddr_core_sct => x_rsc_18_0_i_s_re_core_sct,
      x_rsc_18_0_i_s_waddr => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_waddr,
      x_rsc_18_0_i_s_waddr_core_sct => x_rsc_18_0_i_s_we_core_sct,
      x_rsc_18_0_i_s_din => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_din,
      x_rsc_18_0_i_s_dout => hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_dout
    );
  hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_raddr_core <= x_rsc_18_0_i_s_raddr_core;
  hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_waddr_core <= x_rsc_18_0_i_s_waddr_core;
  x_rsc_18_0_i_s_din_mxwt <= hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_din_mxwt;
  hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_dout_core <= x_rsc_18_0_i_s_dout_core;
  x_rsc_18_0_i_s_raddr <= hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_raddr;
  x_rsc_18_0_i_s_waddr <= hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_waddr;
  hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_din <= x_rsc_18_0_i_s_din;
  x_rsc_18_0_i_s_dout <= hybrid_core_x_rsc_18_0_i_x_rsc_18_0_wait_dp_inst_x_rsc_18_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_17_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_17_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_17_0_s_tdone : IN STD_LOGIC;
    x_rsc_17_0_tr_write_done : IN STD_LOGIC;
    x_rsc_17_0_RREADY : IN STD_LOGIC;
    x_rsc_17_0_RVALID : OUT STD_LOGIC;
    x_rsc_17_0_RUSER : OUT STD_LOGIC;
    x_rsc_17_0_RLAST : OUT STD_LOGIC;
    x_rsc_17_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_RID : OUT STD_LOGIC;
    x_rsc_17_0_ARREADY : OUT STD_LOGIC;
    x_rsc_17_0_ARVALID : IN STD_LOGIC;
    x_rsc_17_0_ARUSER : IN STD_LOGIC;
    x_rsc_17_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARLOCK : IN STD_LOGIC;
    x_rsc_17_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_17_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_17_0_ARID : IN STD_LOGIC;
    x_rsc_17_0_BREADY : IN STD_LOGIC;
    x_rsc_17_0_BVALID : OUT STD_LOGIC;
    x_rsc_17_0_BUSER : OUT STD_LOGIC;
    x_rsc_17_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_BID : OUT STD_LOGIC;
    x_rsc_17_0_WREADY : OUT STD_LOGIC;
    x_rsc_17_0_WVALID : IN STD_LOGIC;
    x_rsc_17_0_WUSER : IN STD_LOGIC;
    x_rsc_17_0_WLAST : IN STD_LOGIC;
    x_rsc_17_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_AWREADY : OUT STD_LOGIC;
    x_rsc_17_0_AWVALID : IN STD_LOGIC;
    x_rsc_17_0_AWUSER : IN STD_LOGIC;
    x_rsc_17_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWLOCK : IN STD_LOGIC;
    x_rsc_17_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_17_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_17_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_17_0_i_oswt : IN STD_LOGIC;
    x_rsc_17_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_17_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_17_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_17_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_17_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_17_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_17_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_17_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_17_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_17_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_17_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_17_0_i_oswt : IN STD_LOGIC;
      x_rsc_17_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_17_0_i_biwt : OUT STD_LOGIC;
      x_rsc_17_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_17_0_i_bcwt : IN STD_LOGIC;
      x_rsc_17_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_17_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_17_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_17_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_17_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_17_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_17_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_17_0_i_oswt : IN STD_LOGIC;
      x_rsc_17_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_17_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_17_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_17_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_17_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_17_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_i_biwt : IN STD_LOGIC;
      x_rsc_17_0_i_bdwt : IN STD_LOGIC;
      x_rsc_17_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_17_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_17_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_17_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_17_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_17_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_17_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_17_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_17_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_17_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_17_0_i_AWID,
      AWADDR => x_rsc_17_0_i_AWADDR,
      AWLEN => x_rsc_17_0_i_AWLEN,
      AWSIZE => x_rsc_17_0_i_AWSIZE,
      AWBURST => x_rsc_17_0_i_AWBURST,
      AWLOCK => x_rsc_17_0_AWLOCK,
      AWCACHE => x_rsc_17_0_i_AWCACHE,
      AWPROT => x_rsc_17_0_i_AWPROT,
      AWQOS => x_rsc_17_0_i_AWQOS,
      AWREGION => x_rsc_17_0_i_AWREGION,
      AWUSER => x_rsc_17_0_i_AWUSER,
      AWVALID => x_rsc_17_0_AWVALID,
      AWREADY => x_rsc_17_0_AWREADY,
      WDATA => x_rsc_17_0_i_WDATA,
      WSTRB => x_rsc_17_0_i_WSTRB,
      WLAST => x_rsc_17_0_WLAST,
      WUSER => x_rsc_17_0_i_WUSER,
      WVALID => x_rsc_17_0_WVALID,
      WREADY => x_rsc_17_0_WREADY,
      BID => x_rsc_17_0_i_BID,
      BRESP => x_rsc_17_0_i_BRESP,
      BUSER => x_rsc_17_0_i_BUSER,
      BVALID => x_rsc_17_0_BVALID,
      BREADY => x_rsc_17_0_BREADY,
      ARID => x_rsc_17_0_i_ARID,
      ARADDR => x_rsc_17_0_i_ARADDR,
      ARLEN => x_rsc_17_0_i_ARLEN,
      ARSIZE => x_rsc_17_0_i_ARSIZE,
      ARBURST => x_rsc_17_0_i_ARBURST,
      ARLOCK => x_rsc_17_0_ARLOCK,
      ARCACHE => x_rsc_17_0_i_ARCACHE,
      ARPROT => x_rsc_17_0_i_ARPROT,
      ARQOS => x_rsc_17_0_i_ARQOS,
      ARREGION => x_rsc_17_0_i_ARREGION,
      ARUSER => x_rsc_17_0_i_ARUSER,
      ARVALID => x_rsc_17_0_ARVALID,
      ARREADY => x_rsc_17_0_ARREADY,
      RID => x_rsc_17_0_i_RID,
      RDATA => x_rsc_17_0_i_RDATA,
      RRESP => x_rsc_17_0_i_RRESP,
      RLAST => x_rsc_17_0_RLAST,
      RUSER => x_rsc_17_0_i_RUSER,
      RVALID => x_rsc_17_0_RVALID,
      RREADY => x_rsc_17_0_RREADY,
      s_re => x_rsc_17_0_i_s_re_core_sct,
      s_we => x_rsc_17_0_i_s_we_core_sct,
      s_raddr => x_rsc_17_0_i_s_raddr_1,
      s_waddr => x_rsc_17_0_i_s_waddr_1,
      s_din => x_rsc_17_0_i_s_din_1,
      s_dout => x_rsc_17_0_i_s_dout_1,
      s_rrdy => x_rsc_17_0_i_s_rrdy,
      s_wrdy => x_rsc_17_0_i_s_wrdy,
      is_idle => x_rsc_17_0_is_idle_1,
      tr_write_done => x_rsc_17_0_tr_write_done,
      s_tdone => x_rsc_17_0_s_tdone
    );
  x_rsc_17_0_i_AWID(0) <= x_rsc_17_0_AWID;
  x_rsc_17_0_i_AWADDR <= x_rsc_17_0_AWADDR;
  x_rsc_17_0_i_AWLEN <= x_rsc_17_0_AWLEN;
  x_rsc_17_0_i_AWSIZE <= x_rsc_17_0_AWSIZE;
  x_rsc_17_0_i_AWBURST <= x_rsc_17_0_AWBURST;
  x_rsc_17_0_i_AWCACHE <= x_rsc_17_0_AWCACHE;
  x_rsc_17_0_i_AWPROT <= x_rsc_17_0_AWPROT;
  x_rsc_17_0_i_AWQOS <= x_rsc_17_0_AWQOS;
  x_rsc_17_0_i_AWREGION <= x_rsc_17_0_AWREGION;
  x_rsc_17_0_i_AWUSER(0) <= x_rsc_17_0_AWUSER;
  x_rsc_17_0_i_WDATA <= x_rsc_17_0_WDATA;
  x_rsc_17_0_i_WSTRB <= x_rsc_17_0_WSTRB;
  x_rsc_17_0_i_WUSER(0) <= x_rsc_17_0_WUSER;
  x_rsc_17_0_BID <= x_rsc_17_0_i_BID(0);
  x_rsc_17_0_BRESP <= x_rsc_17_0_i_BRESP;
  x_rsc_17_0_BUSER <= x_rsc_17_0_i_BUSER(0);
  x_rsc_17_0_i_ARID(0) <= x_rsc_17_0_ARID;
  x_rsc_17_0_i_ARADDR <= x_rsc_17_0_ARADDR;
  x_rsc_17_0_i_ARLEN <= x_rsc_17_0_ARLEN;
  x_rsc_17_0_i_ARSIZE <= x_rsc_17_0_ARSIZE;
  x_rsc_17_0_i_ARBURST <= x_rsc_17_0_ARBURST;
  x_rsc_17_0_i_ARCACHE <= x_rsc_17_0_ARCACHE;
  x_rsc_17_0_i_ARPROT <= x_rsc_17_0_ARPROT;
  x_rsc_17_0_i_ARQOS <= x_rsc_17_0_ARQOS;
  x_rsc_17_0_i_ARREGION <= x_rsc_17_0_ARREGION;
  x_rsc_17_0_i_ARUSER(0) <= x_rsc_17_0_ARUSER;
  x_rsc_17_0_RID <= x_rsc_17_0_i_RID(0);
  x_rsc_17_0_RDATA <= x_rsc_17_0_i_RDATA;
  x_rsc_17_0_RRESP <= x_rsc_17_0_i_RRESP;
  x_rsc_17_0_RUSER <= x_rsc_17_0_i_RUSER(0);
  x_rsc_17_0_i_s_raddr_1 <= x_rsc_17_0_i_s_raddr;
  x_rsc_17_0_i_s_waddr_1 <= x_rsc_17_0_i_s_waddr;
  x_rsc_17_0_i_s_din <= x_rsc_17_0_i_s_din_1;
  x_rsc_17_0_i_s_dout_1 <= x_rsc_17_0_i_s_dout;

  hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl_inst : hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_17_0_i_oswt => x_rsc_17_0_i_oswt,
      x_rsc_17_0_i_oswt_1 => x_rsc_17_0_i_oswt_1,
      x_rsc_17_0_i_biwt => x_rsc_17_0_i_biwt,
      x_rsc_17_0_i_bdwt => x_rsc_17_0_i_bdwt,
      x_rsc_17_0_i_bcwt => x_rsc_17_0_i_bcwt,
      x_rsc_17_0_i_s_re_core_sct => x_rsc_17_0_i_s_re_core_sct,
      x_rsc_17_0_i_biwt_1 => x_rsc_17_0_i_biwt_1,
      x_rsc_17_0_i_bdwt_2 => x_rsc_17_0_i_bdwt_2,
      x_rsc_17_0_i_bcwt_1 => x_rsc_17_0_i_bcwt_1,
      x_rsc_17_0_i_s_we_core_sct => x_rsc_17_0_i_s_we_core_sct,
      x_rsc_17_0_i_s_rrdy => x_rsc_17_0_i_s_rrdy,
      x_rsc_17_0_i_s_wrdy => x_rsc_17_0_i_s_wrdy
    );
  hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst : hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_17_0_i_oswt => x_rsc_17_0_i_oswt,
      x_rsc_17_0_i_wen_comp => x_rsc_17_0_i_wen_comp,
      x_rsc_17_0_i_oswt_1 => x_rsc_17_0_i_oswt_1,
      x_rsc_17_0_i_wen_comp_1 => x_rsc_17_0_i_wen_comp_1,
      x_rsc_17_0_i_s_raddr_core => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_raddr_core,
      x_rsc_17_0_i_s_waddr_core => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_waddr_core,
      x_rsc_17_0_i_s_din_mxwt => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_din_mxwt,
      x_rsc_17_0_i_s_dout_core => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_dout_core,
      x_rsc_17_0_i_biwt => x_rsc_17_0_i_biwt,
      x_rsc_17_0_i_bdwt => x_rsc_17_0_i_bdwt,
      x_rsc_17_0_i_bcwt => x_rsc_17_0_i_bcwt,
      x_rsc_17_0_i_biwt_1 => x_rsc_17_0_i_biwt_1,
      x_rsc_17_0_i_bdwt_2 => x_rsc_17_0_i_bdwt_2,
      x_rsc_17_0_i_bcwt_1 => x_rsc_17_0_i_bcwt_1,
      x_rsc_17_0_i_s_raddr => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_raddr,
      x_rsc_17_0_i_s_raddr_core_sct => x_rsc_17_0_i_s_re_core_sct,
      x_rsc_17_0_i_s_waddr => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_waddr,
      x_rsc_17_0_i_s_waddr_core_sct => x_rsc_17_0_i_s_we_core_sct,
      x_rsc_17_0_i_s_din => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_din,
      x_rsc_17_0_i_s_dout => hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_dout
    );
  hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_raddr_core <= x_rsc_17_0_i_s_raddr_core;
  hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_waddr_core <= x_rsc_17_0_i_s_waddr_core;
  x_rsc_17_0_i_s_din_mxwt <= hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_din_mxwt;
  hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_dout_core <= x_rsc_17_0_i_s_dout_core;
  x_rsc_17_0_i_s_raddr <= hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_raddr;
  x_rsc_17_0_i_s_waddr <= hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_waddr;
  hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_din <= x_rsc_17_0_i_s_din;
  x_rsc_17_0_i_s_dout <= hybrid_core_x_rsc_17_0_i_x_rsc_17_0_wait_dp_inst_x_rsc_17_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_16_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_16_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_16_0_s_tdone : IN STD_LOGIC;
    x_rsc_16_0_tr_write_done : IN STD_LOGIC;
    x_rsc_16_0_RREADY : IN STD_LOGIC;
    x_rsc_16_0_RVALID : OUT STD_LOGIC;
    x_rsc_16_0_RUSER : OUT STD_LOGIC;
    x_rsc_16_0_RLAST : OUT STD_LOGIC;
    x_rsc_16_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_RID : OUT STD_LOGIC;
    x_rsc_16_0_ARREADY : OUT STD_LOGIC;
    x_rsc_16_0_ARVALID : IN STD_LOGIC;
    x_rsc_16_0_ARUSER : IN STD_LOGIC;
    x_rsc_16_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARLOCK : IN STD_LOGIC;
    x_rsc_16_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_16_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_16_0_ARID : IN STD_LOGIC;
    x_rsc_16_0_BREADY : IN STD_LOGIC;
    x_rsc_16_0_BVALID : OUT STD_LOGIC;
    x_rsc_16_0_BUSER : OUT STD_LOGIC;
    x_rsc_16_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_BID : OUT STD_LOGIC;
    x_rsc_16_0_WREADY : OUT STD_LOGIC;
    x_rsc_16_0_WVALID : IN STD_LOGIC;
    x_rsc_16_0_WUSER : IN STD_LOGIC;
    x_rsc_16_0_WLAST : IN STD_LOGIC;
    x_rsc_16_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_AWREADY : OUT STD_LOGIC;
    x_rsc_16_0_AWVALID : IN STD_LOGIC;
    x_rsc_16_0_AWUSER : IN STD_LOGIC;
    x_rsc_16_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWLOCK : IN STD_LOGIC;
    x_rsc_16_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_16_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_16_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_16_0_i_oswt : IN STD_LOGIC;
    x_rsc_16_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_16_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_16_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_16_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_16_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_16_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_16_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_16_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_16_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_16_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_16_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_16_0_i_oswt : IN STD_LOGIC;
      x_rsc_16_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_16_0_i_biwt : OUT STD_LOGIC;
      x_rsc_16_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_16_0_i_bcwt : IN STD_LOGIC;
      x_rsc_16_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_16_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_16_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_16_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_16_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_16_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_16_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_16_0_i_oswt : IN STD_LOGIC;
      x_rsc_16_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_16_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_16_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_16_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_16_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_16_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_i_biwt : IN STD_LOGIC;
      x_rsc_16_0_i_bdwt : IN STD_LOGIC;
      x_rsc_16_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_16_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_16_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_16_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_16_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_16_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_16_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_16_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_16_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_16_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_16_0_i_AWID,
      AWADDR => x_rsc_16_0_i_AWADDR,
      AWLEN => x_rsc_16_0_i_AWLEN,
      AWSIZE => x_rsc_16_0_i_AWSIZE,
      AWBURST => x_rsc_16_0_i_AWBURST,
      AWLOCK => x_rsc_16_0_AWLOCK,
      AWCACHE => x_rsc_16_0_i_AWCACHE,
      AWPROT => x_rsc_16_0_i_AWPROT,
      AWQOS => x_rsc_16_0_i_AWQOS,
      AWREGION => x_rsc_16_0_i_AWREGION,
      AWUSER => x_rsc_16_0_i_AWUSER,
      AWVALID => x_rsc_16_0_AWVALID,
      AWREADY => x_rsc_16_0_AWREADY,
      WDATA => x_rsc_16_0_i_WDATA,
      WSTRB => x_rsc_16_0_i_WSTRB,
      WLAST => x_rsc_16_0_WLAST,
      WUSER => x_rsc_16_0_i_WUSER,
      WVALID => x_rsc_16_0_WVALID,
      WREADY => x_rsc_16_0_WREADY,
      BID => x_rsc_16_0_i_BID,
      BRESP => x_rsc_16_0_i_BRESP,
      BUSER => x_rsc_16_0_i_BUSER,
      BVALID => x_rsc_16_0_BVALID,
      BREADY => x_rsc_16_0_BREADY,
      ARID => x_rsc_16_0_i_ARID,
      ARADDR => x_rsc_16_0_i_ARADDR,
      ARLEN => x_rsc_16_0_i_ARLEN,
      ARSIZE => x_rsc_16_0_i_ARSIZE,
      ARBURST => x_rsc_16_0_i_ARBURST,
      ARLOCK => x_rsc_16_0_ARLOCK,
      ARCACHE => x_rsc_16_0_i_ARCACHE,
      ARPROT => x_rsc_16_0_i_ARPROT,
      ARQOS => x_rsc_16_0_i_ARQOS,
      ARREGION => x_rsc_16_0_i_ARREGION,
      ARUSER => x_rsc_16_0_i_ARUSER,
      ARVALID => x_rsc_16_0_ARVALID,
      ARREADY => x_rsc_16_0_ARREADY,
      RID => x_rsc_16_0_i_RID,
      RDATA => x_rsc_16_0_i_RDATA,
      RRESP => x_rsc_16_0_i_RRESP,
      RLAST => x_rsc_16_0_RLAST,
      RUSER => x_rsc_16_0_i_RUSER,
      RVALID => x_rsc_16_0_RVALID,
      RREADY => x_rsc_16_0_RREADY,
      s_re => x_rsc_16_0_i_s_re_core_sct,
      s_we => x_rsc_16_0_i_s_we_core_sct,
      s_raddr => x_rsc_16_0_i_s_raddr_1,
      s_waddr => x_rsc_16_0_i_s_waddr_1,
      s_din => x_rsc_16_0_i_s_din_1,
      s_dout => x_rsc_16_0_i_s_dout_1,
      s_rrdy => x_rsc_16_0_i_s_rrdy,
      s_wrdy => x_rsc_16_0_i_s_wrdy,
      is_idle => x_rsc_16_0_is_idle_1,
      tr_write_done => x_rsc_16_0_tr_write_done,
      s_tdone => x_rsc_16_0_s_tdone
    );
  x_rsc_16_0_i_AWID(0) <= x_rsc_16_0_AWID;
  x_rsc_16_0_i_AWADDR <= x_rsc_16_0_AWADDR;
  x_rsc_16_0_i_AWLEN <= x_rsc_16_0_AWLEN;
  x_rsc_16_0_i_AWSIZE <= x_rsc_16_0_AWSIZE;
  x_rsc_16_0_i_AWBURST <= x_rsc_16_0_AWBURST;
  x_rsc_16_0_i_AWCACHE <= x_rsc_16_0_AWCACHE;
  x_rsc_16_0_i_AWPROT <= x_rsc_16_0_AWPROT;
  x_rsc_16_0_i_AWQOS <= x_rsc_16_0_AWQOS;
  x_rsc_16_0_i_AWREGION <= x_rsc_16_0_AWREGION;
  x_rsc_16_0_i_AWUSER(0) <= x_rsc_16_0_AWUSER;
  x_rsc_16_0_i_WDATA <= x_rsc_16_0_WDATA;
  x_rsc_16_0_i_WSTRB <= x_rsc_16_0_WSTRB;
  x_rsc_16_0_i_WUSER(0) <= x_rsc_16_0_WUSER;
  x_rsc_16_0_BID <= x_rsc_16_0_i_BID(0);
  x_rsc_16_0_BRESP <= x_rsc_16_0_i_BRESP;
  x_rsc_16_0_BUSER <= x_rsc_16_0_i_BUSER(0);
  x_rsc_16_0_i_ARID(0) <= x_rsc_16_0_ARID;
  x_rsc_16_0_i_ARADDR <= x_rsc_16_0_ARADDR;
  x_rsc_16_0_i_ARLEN <= x_rsc_16_0_ARLEN;
  x_rsc_16_0_i_ARSIZE <= x_rsc_16_0_ARSIZE;
  x_rsc_16_0_i_ARBURST <= x_rsc_16_0_ARBURST;
  x_rsc_16_0_i_ARCACHE <= x_rsc_16_0_ARCACHE;
  x_rsc_16_0_i_ARPROT <= x_rsc_16_0_ARPROT;
  x_rsc_16_0_i_ARQOS <= x_rsc_16_0_ARQOS;
  x_rsc_16_0_i_ARREGION <= x_rsc_16_0_ARREGION;
  x_rsc_16_0_i_ARUSER(0) <= x_rsc_16_0_ARUSER;
  x_rsc_16_0_RID <= x_rsc_16_0_i_RID(0);
  x_rsc_16_0_RDATA <= x_rsc_16_0_i_RDATA;
  x_rsc_16_0_RRESP <= x_rsc_16_0_i_RRESP;
  x_rsc_16_0_RUSER <= x_rsc_16_0_i_RUSER(0);
  x_rsc_16_0_i_s_raddr_1 <= x_rsc_16_0_i_s_raddr;
  x_rsc_16_0_i_s_waddr_1 <= x_rsc_16_0_i_s_waddr;
  x_rsc_16_0_i_s_din <= x_rsc_16_0_i_s_din_1;
  x_rsc_16_0_i_s_dout_1 <= x_rsc_16_0_i_s_dout;

  hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl_inst : hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_16_0_i_oswt => x_rsc_16_0_i_oswt,
      x_rsc_16_0_i_oswt_1 => x_rsc_16_0_i_oswt_1,
      x_rsc_16_0_i_biwt => x_rsc_16_0_i_biwt,
      x_rsc_16_0_i_bdwt => x_rsc_16_0_i_bdwt,
      x_rsc_16_0_i_bcwt => x_rsc_16_0_i_bcwt,
      x_rsc_16_0_i_s_re_core_sct => x_rsc_16_0_i_s_re_core_sct,
      x_rsc_16_0_i_biwt_1 => x_rsc_16_0_i_biwt_1,
      x_rsc_16_0_i_bdwt_2 => x_rsc_16_0_i_bdwt_2,
      x_rsc_16_0_i_bcwt_1 => x_rsc_16_0_i_bcwt_1,
      x_rsc_16_0_i_s_we_core_sct => x_rsc_16_0_i_s_we_core_sct,
      x_rsc_16_0_i_s_rrdy => x_rsc_16_0_i_s_rrdy,
      x_rsc_16_0_i_s_wrdy => x_rsc_16_0_i_s_wrdy
    );
  hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst : hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_16_0_i_oswt => x_rsc_16_0_i_oswt,
      x_rsc_16_0_i_wen_comp => x_rsc_16_0_i_wen_comp,
      x_rsc_16_0_i_oswt_1 => x_rsc_16_0_i_oswt_1,
      x_rsc_16_0_i_wen_comp_1 => x_rsc_16_0_i_wen_comp_1,
      x_rsc_16_0_i_s_raddr_core => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_raddr_core,
      x_rsc_16_0_i_s_waddr_core => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_waddr_core,
      x_rsc_16_0_i_s_din_mxwt => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_din_mxwt,
      x_rsc_16_0_i_s_dout_core => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_dout_core,
      x_rsc_16_0_i_biwt => x_rsc_16_0_i_biwt,
      x_rsc_16_0_i_bdwt => x_rsc_16_0_i_bdwt,
      x_rsc_16_0_i_bcwt => x_rsc_16_0_i_bcwt,
      x_rsc_16_0_i_biwt_1 => x_rsc_16_0_i_biwt_1,
      x_rsc_16_0_i_bdwt_2 => x_rsc_16_0_i_bdwt_2,
      x_rsc_16_0_i_bcwt_1 => x_rsc_16_0_i_bcwt_1,
      x_rsc_16_0_i_s_raddr => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_raddr,
      x_rsc_16_0_i_s_raddr_core_sct => x_rsc_16_0_i_s_re_core_sct,
      x_rsc_16_0_i_s_waddr => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_waddr,
      x_rsc_16_0_i_s_waddr_core_sct => x_rsc_16_0_i_s_we_core_sct,
      x_rsc_16_0_i_s_din => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_din,
      x_rsc_16_0_i_s_dout => hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_dout
    );
  hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_raddr_core <= x_rsc_16_0_i_s_raddr_core;
  hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_waddr_core <= x_rsc_16_0_i_s_waddr_core;
  x_rsc_16_0_i_s_din_mxwt <= hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_din_mxwt;
  hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_dout_core <= x_rsc_16_0_i_s_dout_core;
  x_rsc_16_0_i_s_raddr <= hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_raddr;
  x_rsc_16_0_i_s_waddr <= hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_waddr;
  hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_din <= x_rsc_16_0_i_s_din;
  x_rsc_16_0_i_s_dout <= hybrid_core_x_rsc_16_0_i_x_rsc_16_0_wait_dp_inst_x_rsc_16_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_15_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_15_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_15_0_s_tdone : IN STD_LOGIC;
    x_rsc_15_0_tr_write_done : IN STD_LOGIC;
    x_rsc_15_0_RREADY : IN STD_LOGIC;
    x_rsc_15_0_RVALID : OUT STD_LOGIC;
    x_rsc_15_0_RUSER : OUT STD_LOGIC;
    x_rsc_15_0_RLAST : OUT STD_LOGIC;
    x_rsc_15_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_RID : OUT STD_LOGIC;
    x_rsc_15_0_ARREADY : OUT STD_LOGIC;
    x_rsc_15_0_ARVALID : IN STD_LOGIC;
    x_rsc_15_0_ARUSER : IN STD_LOGIC;
    x_rsc_15_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARLOCK : IN STD_LOGIC;
    x_rsc_15_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_15_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_15_0_ARID : IN STD_LOGIC;
    x_rsc_15_0_BREADY : IN STD_LOGIC;
    x_rsc_15_0_BVALID : OUT STD_LOGIC;
    x_rsc_15_0_BUSER : OUT STD_LOGIC;
    x_rsc_15_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_BID : OUT STD_LOGIC;
    x_rsc_15_0_WREADY : OUT STD_LOGIC;
    x_rsc_15_0_WVALID : IN STD_LOGIC;
    x_rsc_15_0_WUSER : IN STD_LOGIC;
    x_rsc_15_0_WLAST : IN STD_LOGIC;
    x_rsc_15_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_AWREADY : OUT STD_LOGIC;
    x_rsc_15_0_AWVALID : IN STD_LOGIC;
    x_rsc_15_0_AWUSER : IN STD_LOGIC;
    x_rsc_15_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWLOCK : IN STD_LOGIC;
    x_rsc_15_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_15_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_15_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_15_0_i_oswt : IN STD_LOGIC;
    x_rsc_15_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_15_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_15_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_15_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_15_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_15_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_15_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_15_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_15_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_15_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_15_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_15_0_i_oswt : IN STD_LOGIC;
      x_rsc_15_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_15_0_i_biwt : OUT STD_LOGIC;
      x_rsc_15_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_15_0_i_bcwt : IN STD_LOGIC;
      x_rsc_15_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_15_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_15_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_15_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_15_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_15_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_15_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_15_0_i_oswt : IN STD_LOGIC;
      x_rsc_15_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_15_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_15_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_15_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_15_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_15_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_i_biwt : IN STD_LOGIC;
      x_rsc_15_0_i_bdwt : IN STD_LOGIC;
      x_rsc_15_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_15_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_15_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_15_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_15_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_15_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_15_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_15_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_15_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_15_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_15_0_i_AWID,
      AWADDR => x_rsc_15_0_i_AWADDR,
      AWLEN => x_rsc_15_0_i_AWLEN,
      AWSIZE => x_rsc_15_0_i_AWSIZE,
      AWBURST => x_rsc_15_0_i_AWBURST,
      AWLOCK => x_rsc_15_0_AWLOCK,
      AWCACHE => x_rsc_15_0_i_AWCACHE,
      AWPROT => x_rsc_15_0_i_AWPROT,
      AWQOS => x_rsc_15_0_i_AWQOS,
      AWREGION => x_rsc_15_0_i_AWREGION,
      AWUSER => x_rsc_15_0_i_AWUSER,
      AWVALID => x_rsc_15_0_AWVALID,
      AWREADY => x_rsc_15_0_AWREADY,
      WDATA => x_rsc_15_0_i_WDATA,
      WSTRB => x_rsc_15_0_i_WSTRB,
      WLAST => x_rsc_15_0_WLAST,
      WUSER => x_rsc_15_0_i_WUSER,
      WVALID => x_rsc_15_0_WVALID,
      WREADY => x_rsc_15_0_WREADY,
      BID => x_rsc_15_0_i_BID,
      BRESP => x_rsc_15_0_i_BRESP,
      BUSER => x_rsc_15_0_i_BUSER,
      BVALID => x_rsc_15_0_BVALID,
      BREADY => x_rsc_15_0_BREADY,
      ARID => x_rsc_15_0_i_ARID,
      ARADDR => x_rsc_15_0_i_ARADDR,
      ARLEN => x_rsc_15_0_i_ARLEN,
      ARSIZE => x_rsc_15_0_i_ARSIZE,
      ARBURST => x_rsc_15_0_i_ARBURST,
      ARLOCK => x_rsc_15_0_ARLOCK,
      ARCACHE => x_rsc_15_0_i_ARCACHE,
      ARPROT => x_rsc_15_0_i_ARPROT,
      ARQOS => x_rsc_15_0_i_ARQOS,
      ARREGION => x_rsc_15_0_i_ARREGION,
      ARUSER => x_rsc_15_0_i_ARUSER,
      ARVALID => x_rsc_15_0_ARVALID,
      ARREADY => x_rsc_15_0_ARREADY,
      RID => x_rsc_15_0_i_RID,
      RDATA => x_rsc_15_0_i_RDATA,
      RRESP => x_rsc_15_0_i_RRESP,
      RLAST => x_rsc_15_0_RLAST,
      RUSER => x_rsc_15_0_i_RUSER,
      RVALID => x_rsc_15_0_RVALID,
      RREADY => x_rsc_15_0_RREADY,
      s_re => x_rsc_15_0_i_s_re_core_sct,
      s_we => x_rsc_15_0_i_s_we_core_sct,
      s_raddr => x_rsc_15_0_i_s_raddr_1,
      s_waddr => x_rsc_15_0_i_s_waddr_1,
      s_din => x_rsc_15_0_i_s_din_1,
      s_dout => x_rsc_15_0_i_s_dout_1,
      s_rrdy => x_rsc_15_0_i_s_rrdy,
      s_wrdy => x_rsc_15_0_i_s_wrdy,
      is_idle => x_rsc_15_0_is_idle_1,
      tr_write_done => x_rsc_15_0_tr_write_done,
      s_tdone => x_rsc_15_0_s_tdone
    );
  x_rsc_15_0_i_AWID(0) <= x_rsc_15_0_AWID;
  x_rsc_15_0_i_AWADDR <= x_rsc_15_0_AWADDR;
  x_rsc_15_0_i_AWLEN <= x_rsc_15_0_AWLEN;
  x_rsc_15_0_i_AWSIZE <= x_rsc_15_0_AWSIZE;
  x_rsc_15_0_i_AWBURST <= x_rsc_15_0_AWBURST;
  x_rsc_15_0_i_AWCACHE <= x_rsc_15_0_AWCACHE;
  x_rsc_15_0_i_AWPROT <= x_rsc_15_0_AWPROT;
  x_rsc_15_0_i_AWQOS <= x_rsc_15_0_AWQOS;
  x_rsc_15_0_i_AWREGION <= x_rsc_15_0_AWREGION;
  x_rsc_15_0_i_AWUSER(0) <= x_rsc_15_0_AWUSER;
  x_rsc_15_0_i_WDATA <= x_rsc_15_0_WDATA;
  x_rsc_15_0_i_WSTRB <= x_rsc_15_0_WSTRB;
  x_rsc_15_0_i_WUSER(0) <= x_rsc_15_0_WUSER;
  x_rsc_15_0_BID <= x_rsc_15_0_i_BID(0);
  x_rsc_15_0_BRESP <= x_rsc_15_0_i_BRESP;
  x_rsc_15_0_BUSER <= x_rsc_15_0_i_BUSER(0);
  x_rsc_15_0_i_ARID(0) <= x_rsc_15_0_ARID;
  x_rsc_15_0_i_ARADDR <= x_rsc_15_0_ARADDR;
  x_rsc_15_0_i_ARLEN <= x_rsc_15_0_ARLEN;
  x_rsc_15_0_i_ARSIZE <= x_rsc_15_0_ARSIZE;
  x_rsc_15_0_i_ARBURST <= x_rsc_15_0_ARBURST;
  x_rsc_15_0_i_ARCACHE <= x_rsc_15_0_ARCACHE;
  x_rsc_15_0_i_ARPROT <= x_rsc_15_0_ARPROT;
  x_rsc_15_0_i_ARQOS <= x_rsc_15_0_ARQOS;
  x_rsc_15_0_i_ARREGION <= x_rsc_15_0_ARREGION;
  x_rsc_15_0_i_ARUSER(0) <= x_rsc_15_0_ARUSER;
  x_rsc_15_0_RID <= x_rsc_15_0_i_RID(0);
  x_rsc_15_0_RDATA <= x_rsc_15_0_i_RDATA;
  x_rsc_15_0_RRESP <= x_rsc_15_0_i_RRESP;
  x_rsc_15_0_RUSER <= x_rsc_15_0_i_RUSER(0);
  x_rsc_15_0_i_s_raddr_1 <= x_rsc_15_0_i_s_raddr;
  x_rsc_15_0_i_s_waddr_1 <= x_rsc_15_0_i_s_waddr;
  x_rsc_15_0_i_s_din <= x_rsc_15_0_i_s_din_1;
  x_rsc_15_0_i_s_dout_1 <= x_rsc_15_0_i_s_dout;

  hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl_inst : hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_15_0_i_oswt => x_rsc_15_0_i_oswt,
      x_rsc_15_0_i_oswt_1 => x_rsc_15_0_i_oswt_1,
      x_rsc_15_0_i_biwt => x_rsc_15_0_i_biwt,
      x_rsc_15_0_i_bdwt => x_rsc_15_0_i_bdwt,
      x_rsc_15_0_i_bcwt => x_rsc_15_0_i_bcwt,
      x_rsc_15_0_i_s_re_core_sct => x_rsc_15_0_i_s_re_core_sct,
      x_rsc_15_0_i_biwt_1 => x_rsc_15_0_i_biwt_1,
      x_rsc_15_0_i_bdwt_2 => x_rsc_15_0_i_bdwt_2,
      x_rsc_15_0_i_bcwt_1 => x_rsc_15_0_i_bcwt_1,
      x_rsc_15_0_i_s_we_core_sct => x_rsc_15_0_i_s_we_core_sct,
      x_rsc_15_0_i_s_rrdy => x_rsc_15_0_i_s_rrdy,
      x_rsc_15_0_i_s_wrdy => x_rsc_15_0_i_s_wrdy
    );
  hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst : hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_15_0_i_oswt => x_rsc_15_0_i_oswt,
      x_rsc_15_0_i_wen_comp => x_rsc_15_0_i_wen_comp,
      x_rsc_15_0_i_oswt_1 => x_rsc_15_0_i_oswt_1,
      x_rsc_15_0_i_wen_comp_1 => x_rsc_15_0_i_wen_comp_1,
      x_rsc_15_0_i_s_raddr_core => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_raddr_core,
      x_rsc_15_0_i_s_waddr_core => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_waddr_core,
      x_rsc_15_0_i_s_din_mxwt => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_din_mxwt,
      x_rsc_15_0_i_s_dout_core => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_dout_core,
      x_rsc_15_0_i_biwt => x_rsc_15_0_i_biwt,
      x_rsc_15_0_i_bdwt => x_rsc_15_0_i_bdwt,
      x_rsc_15_0_i_bcwt => x_rsc_15_0_i_bcwt,
      x_rsc_15_0_i_biwt_1 => x_rsc_15_0_i_biwt_1,
      x_rsc_15_0_i_bdwt_2 => x_rsc_15_0_i_bdwt_2,
      x_rsc_15_0_i_bcwt_1 => x_rsc_15_0_i_bcwt_1,
      x_rsc_15_0_i_s_raddr => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_raddr,
      x_rsc_15_0_i_s_raddr_core_sct => x_rsc_15_0_i_s_re_core_sct,
      x_rsc_15_0_i_s_waddr => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_waddr,
      x_rsc_15_0_i_s_waddr_core_sct => x_rsc_15_0_i_s_we_core_sct,
      x_rsc_15_0_i_s_din => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_din,
      x_rsc_15_0_i_s_dout => hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_dout
    );
  hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_raddr_core <= x_rsc_15_0_i_s_raddr_core;
  hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_waddr_core <= x_rsc_15_0_i_s_waddr_core;
  x_rsc_15_0_i_s_din_mxwt <= hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_din_mxwt;
  hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_dout_core <= x_rsc_15_0_i_s_dout_core;
  x_rsc_15_0_i_s_raddr <= hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_raddr;
  x_rsc_15_0_i_s_waddr <= hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_waddr;
  hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_din <= x_rsc_15_0_i_s_din;
  x_rsc_15_0_i_s_dout <= hybrid_core_x_rsc_15_0_i_x_rsc_15_0_wait_dp_inst_x_rsc_15_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_14_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_14_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_14_0_s_tdone : IN STD_LOGIC;
    x_rsc_14_0_tr_write_done : IN STD_LOGIC;
    x_rsc_14_0_RREADY : IN STD_LOGIC;
    x_rsc_14_0_RVALID : OUT STD_LOGIC;
    x_rsc_14_0_RUSER : OUT STD_LOGIC;
    x_rsc_14_0_RLAST : OUT STD_LOGIC;
    x_rsc_14_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_RID : OUT STD_LOGIC;
    x_rsc_14_0_ARREADY : OUT STD_LOGIC;
    x_rsc_14_0_ARVALID : IN STD_LOGIC;
    x_rsc_14_0_ARUSER : IN STD_LOGIC;
    x_rsc_14_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARLOCK : IN STD_LOGIC;
    x_rsc_14_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_14_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_14_0_ARID : IN STD_LOGIC;
    x_rsc_14_0_BREADY : IN STD_LOGIC;
    x_rsc_14_0_BVALID : OUT STD_LOGIC;
    x_rsc_14_0_BUSER : OUT STD_LOGIC;
    x_rsc_14_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_BID : OUT STD_LOGIC;
    x_rsc_14_0_WREADY : OUT STD_LOGIC;
    x_rsc_14_0_WVALID : IN STD_LOGIC;
    x_rsc_14_0_WUSER : IN STD_LOGIC;
    x_rsc_14_0_WLAST : IN STD_LOGIC;
    x_rsc_14_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_AWREADY : OUT STD_LOGIC;
    x_rsc_14_0_AWVALID : IN STD_LOGIC;
    x_rsc_14_0_AWUSER : IN STD_LOGIC;
    x_rsc_14_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWLOCK : IN STD_LOGIC;
    x_rsc_14_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_14_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_14_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_14_0_i_oswt : IN STD_LOGIC;
    x_rsc_14_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_14_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_14_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_14_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_14_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_14_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_14_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_14_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_14_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_14_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_14_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_14_0_i_oswt : IN STD_LOGIC;
      x_rsc_14_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_14_0_i_biwt : OUT STD_LOGIC;
      x_rsc_14_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_14_0_i_bcwt : IN STD_LOGIC;
      x_rsc_14_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_14_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_14_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_14_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_14_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_14_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_14_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_14_0_i_oswt : IN STD_LOGIC;
      x_rsc_14_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_14_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_14_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_14_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_14_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_14_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_i_biwt : IN STD_LOGIC;
      x_rsc_14_0_i_bdwt : IN STD_LOGIC;
      x_rsc_14_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_14_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_14_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_14_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_14_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_14_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_14_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_14_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_14_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_14_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_14_0_i_AWID,
      AWADDR => x_rsc_14_0_i_AWADDR,
      AWLEN => x_rsc_14_0_i_AWLEN,
      AWSIZE => x_rsc_14_0_i_AWSIZE,
      AWBURST => x_rsc_14_0_i_AWBURST,
      AWLOCK => x_rsc_14_0_AWLOCK,
      AWCACHE => x_rsc_14_0_i_AWCACHE,
      AWPROT => x_rsc_14_0_i_AWPROT,
      AWQOS => x_rsc_14_0_i_AWQOS,
      AWREGION => x_rsc_14_0_i_AWREGION,
      AWUSER => x_rsc_14_0_i_AWUSER,
      AWVALID => x_rsc_14_0_AWVALID,
      AWREADY => x_rsc_14_0_AWREADY,
      WDATA => x_rsc_14_0_i_WDATA,
      WSTRB => x_rsc_14_0_i_WSTRB,
      WLAST => x_rsc_14_0_WLAST,
      WUSER => x_rsc_14_0_i_WUSER,
      WVALID => x_rsc_14_0_WVALID,
      WREADY => x_rsc_14_0_WREADY,
      BID => x_rsc_14_0_i_BID,
      BRESP => x_rsc_14_0_i_BRESP,
      BUSER => x_rsc_14_0_i_BUSER,
      BVALID => x_rsc_14_0_BVALID,
      BREADY => x_rsc_14_0_BREADY,
      ARID => x_rsc_14_0_i_ARID,
      ARADDR => x_rsc_14_0_i_ARADDR,
      ARLEN => x_rsc_14_0_i_ARLEN,
      ARSIZE => x_rsc_14_0_i_ARSIZE,
      ARBURST => x_rsc_14_0_i_ARBURST,
      ARLOCK => x_rsc_14_0_ARLOCK,
      ARCACHE => x_rsc_14_0_i_ARCACHE,
      ARPROT => x_rsc_14_0_i_ARPROT,
      ARQOS => x_rsc_14_0_i_ARQOS,
      ARREGION => x_rsc_14_0_i_ARREGION,
      ARUSER => x_rsc_14_0_i_ARUSER,
      ARVALID => x_rsc_14_0_ARVALID,
      ARREADY => x_rsc_14_0_ARREADY,
      RID => x_rsc_14_0_i_RID,
      RDATA => x_rsc_14_0_i_RDATA,
      RRESP => x_rsc_14_0_i_RRESP,
      RLAST => x_rsc_14_0_RLAST,
      RUSER => x_rsc_14_0_i_RUSER,
      RVALID => x_rsc_14_0_RVALID,
      RREADY => x_rsc_14_0_RREADY,
      s_re => x_rsc_14_0_i_s_re_core_sct,
      s_we => x_rsc_14_0_i_s_we_core_sct,
      s_raddr => x_rsc_14_0_i_s_raddr_1,
      s_waddr => x_rsc_14_0_i_s_waddr_1,
      s_din => x_rsc_14_0_i_s_din_1,
      s_dout => x_rsc_14_0_i_s_dout_1,
      s_rrdy => x_rsc_14_0_i_s_rrdy,
      s_wrdy => x_rsc_14_0_i_s_wrdy,
      is_idle => x_rsc_14_0_is_idle_1,
      tr_write_done => x_rsc_14_0_tr_write_done,
      s_tdone => x_rsc_14_0_s_tdone
    );
  x_rsc_14_0_i_AWID(0) <= x_rsc_14_0_AWID;
  x_rsc_14_0_i_AWADDR <= x_rsc_14_0_AWADDR;
  x_rsc_14_0_i_AWLEN <= x_rsc_14_0_AWLEN;
  x_rsc_14_0_i_AWSIZE <= x_rsc_14_0_AWSIZE;
  x_rsc_14_0_i_AWBURST <= x_rsc_14_0_AWBURST;
  x_rsc_14_0_i_AWCACHE <= x_rsc_14_0_AWCACHE;
  x_rsc_14_0_i_AWPROT <= x_rsc_14_0_AWPROT;
  x_rsc_14_0_i_AWQOS <= x_rsc_14_0_AWQOS;
  x_rsc_14_0_i_AWREGION <= x_rsc_14_0_AWREGION;
  x_rsc_14_0_i_AWUSER(0) <= x_rsc_14_0_AWUSER;
  x_rsc_14_0_i_WDATA <= x_rsc_14_0_WDATA;
  x_rsc_14_0_i_WSTRB <= x_rsc_14_0_WSTRB;
  x_rsc_14_0_i_WUSER(0) <= x_rsc_14_0_WUSER;
  x_rsc_14_0_BID <= x_rsc_14_0_i_BID(0);
  x_rsc_14_0_BRESP <= x_rsc_14_0_i_BRESP;
  x_rsc_14_0_BUSER <= x_rsc_14_0_i_BUSER(0);
  x_rsc_14_0_i_ARID(0) <= x_rsc_14_0_ARID;
  x_rsc_14_0_i_ARADDR <= x_rsc_14_0_ARADDR;
  x_rsc_14_0_i_ARLEN <= x_rsc_14_0_ARLEN;
  x_rsc_14_0_i_ARSIZE <= x_rsc_14_0_ARSIZE;
  x_rsc_14_0_i_ARBURST <= x_rsc_14_0_ARBURST;
  x_rsc_14_0_i_ARCACHE <= x_rsc_14_0_ARCACHE;
  x_rsc_14_0_i_ARPROT <= x_rsc_14_0_ARPROT;
  x_rsc_14_0_i_ARQOS <= x_rsc_14_0_ARQOS;
  x_rsc_14_0_i_ARREGION <= x_rsc_14_0_ARREGION;
  x_rsc_14_0_i_ARUSER(0) <= x_rsc_14_0_ARUSER;
  x_rsc_14_0_RID <= x_rsc_14_0_i_RID(0);
  x_rsc_14_0_RDATA <= x_rsc_14_0_i_RDATA;
  x_rsc_14_0_RRESP <= x_rsc_14_0_i_RRESP;
  x_rsc_14_0_RUSER <= x_rsc_14_0_i_RUSER(0);
  x_rsc_14_0_i_s_raddr_1 <= x_rsc_14_0_i_s_raddr;
  x_rsc_14_0_i_s_waddr_1 <= x_rsc_14_0_i_s_waddr;
  x_rsc_14_0_i_s_din <= x_rsc_14_0_i_s_din_1;
  x_rsc_14_0_i_s_dout_1 <= x_rsc_14_0_i_s_dout;

  hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl_inst : hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_14_0_i_oswt => x_rsc_14_0_i_oswt,
      x_rsc_14_0_i_oswt_1 => x_rsc_14_0_i_oswt_1,
      x_rsc_14_0_i_biwt => x_rsc_14_0_i_biwt,
      x_rsc_14_0_i_bdwt => x_rsc_14_0_i_bdwt,
      x_rsc_14_0_i_bcwt => x_rsc_14_0_i_bcwt,
      x_rsc_14_0_i_s_re_core_sct => x_rsc_14_0_i_s_re_core_sct,
      x_rsc_14_0_i_biwt_1 => x_rsc_14_0_i_biwt_1,
      x_rsc_14_0_i_bdwt_2 => x_rsc_14_0_i_bdwt_2,
      x_rsc_14_0_i_bcwt_1 => x_rsc_14_0_i_bcwt_1,
      x_rsc_14_0_i_s_we_core_sct => x_rsc_14_0_i_s_we_core_sct,
      x_rsc_14_0_i_s_rrdy => x_rsc_14_0_i_s_rrdy,
      x_rsc_14_0_i_s_wrdy => x_rsc_14_0_i_s_wrdy
    );
  hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst : hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_14_0_i_oswt => x_rsc_14_0_i_oswt,
      x_rsc_14_0_i_wen_comp => x_rsc_14_0_i_wen_comp,
      x_rsc_14_0_i_oswt_1 => x_rsc_14_0_i_oswt_1,
      x_rsc_14_0_i_wen_comp_1 => x_rsc_14_0_i_wen_comp_1,
      x_rsc_14_0_i_s_raddr_core => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_raddr_core,
      x_rsc_14_0_i_s_waddr_core => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_waddr_core,
      x_rsc_14_0_i_s_din_mxwt => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_din_mxwt,
      x_rsc_14_0_i_s_dout_core => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_dout_core,
      x_rsc_14_0_i_biwt => x_rsc_14_0_i_biwt,
      x_rsc_14_0_i_bdwt => x_rsc_14_0_i_bdwt,
      x_rsc_14_0_i_bcwt => x_rsc_14_0_i_bcwt,
      x_rsc_14_0_i_biwt_1 => x_rsc_14_0_i_biwt_1,
      x_rsc_14_0_i_bdwt_2 => x_rsc_14_0_i_bdwt_2,
      x_rsc_14_0_i_bcwt_1 => x_rsc_14_0_i_bcwt_1,
      x_rsc_14_0_i_s_raddr => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_raddr,
      x_rsc_14_0_i_s_raddr_core_sct => x_rsc_14_0_i_s_re_core_sct,
      x_rsc_14_0_i_s_waddr => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_waddr,
      x_rsc_14_0_i_s_waddr_core_sct => x_rsc_14_0_i_s_we_core_sct,
      x_rsc_14_0_i_s_din => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_din,
      x_rsc_14_0_i_s_dout => hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_dout
    );
  hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_raddr_core <= x_rsc_14_0_i_s_raddr_core;
  hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_waddr_core <= x_rsc_14_0_i_s_waddr_core;
  x_rsc_14_0_i_s_din_mxwt <= hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_din_mxwt;
  hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_dout_core <= x_rsc_14_0_i_s_dout_core;
  x_rsc_14_0_i_s_raddr <= hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_raddr;
  x_rsc_14_0_i_s_waddr <= hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_waddr;
  hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_din <= x_rsc_14_0_i_s_din;
  x_rsc_14_0_i_s_dout <= hybrid_core_x_rsc_14_0_i_x_rsc_14_0_wait_dp_inst_x_rsc_14_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_13_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_13_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_13_0_s_tdone : IN STD_LOGIC;
    x_rsc_13_0_tr_write_done : IN STD_LOGIC;
    x_rsc_13_0_RREADY : IN STD_LOGIC;
    x_rsc_13_0_RVALID : OUT STD_LOGIC;
    x_rsc_13_0_RUSER : OUT STD_LOGIC;
    x_rsc_13_0_RLAST : OUT STD_LOGIC;
    x_rsc_13_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_RID : OUT STD_LOGIC;
    x_rsc_13_0_ARREADY : OUT STD_LOGIC;
    x_rsc_13_0_ARVALID : IN STD_LOGIC;
    x_rsc_13_0_ARUSER : IN STD_LOGIC;
    x_rsc_13_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARLOCK : IN STD_LOGIC;
    x_rsc_13_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_13_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_13_0_ARID : IN STD_LOGIC;
    x_rsc_13_0_BREADY : IN STD_LOGIC;
    x_rsc_13_0_BVALID : OUT STD_LOGIC;
    x_rsc_13_0_BUSER : OUT STD_LOGIC;
    x_rsc_13_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_BID : OUT STD_LOGIC;
    x_rsc_13_0_WREADY : OUT STD_LOGIC;
    x_rsc_13_0_WVALID : IN STD_LOGIC;
    x_rsc_13_0_WUSER : IN STD_LOGIC;
    x_rsc_13_0_WLAST : IN STD_LOGIC;
    x_rsc_13_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_AWREADY : OUT STD_LOGIC;
    x_rsc_13_0_AWVALID : IN STD_LOGIC;
    x_rsc_13_0_AWUSER : IN STD_LOGIC;
    x_rsc_13_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWLOCK : IN STD_LOGIC;
    x_rsc_13_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_13_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_13_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_13_0_i_oswt : IN STD_LOGIC;
    x_rsc_13_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_13_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_13_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_13_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_13_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_13_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_13_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_13_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_13_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_13_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_13_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_13_0_i_oswt : IN STD_LOGIC;
      x_rsc_13_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_13_0_i_biwt : OUT STD_LOGIC;
      x_rsc_13_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_13_0_i_bcwt : IN STD_LOGIC;
      x_rsc_13_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_13_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_13_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_13_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_13_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_13_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_13_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_13_0_i_oswt : IN STD_LOGIC;
      x_rsc_13_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_13_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_13_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_13_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_13_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_13_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_i_biwt : IN STD_LOGIC;
      x_rsc_13_0_i_bdwt : IN STD_LOGIC;
      x_rsc_13_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_13_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_13_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_13_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_13_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_13_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_13_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_13_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_13_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_13_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_13_0_i_AWID,
      AWADDR => x_rsc_13_0_i_AWADDR,
      AWLEN => x_rsc_13_0_i_AWLEN,
      AWSIZE => x_rsc_13_0_i_AWSIZE,
      AWBURST => x_rsc_13_0_i_AWBURST,
      AWLOCK => x_rsc_13_0_AWLOCK,
      AWCACHE => x_rsc_13_0_i_AWCACHE,
      AWPROT => x_rsc_13_0_i_AWPROT,
      AWQOS => x_rsc_13_0_i_AWQOS,
      AWREGION => x_rsc_13_0_i_AWREGION,
      AWUSER => x_rsc_13_0_i_AWUSER,
      AWVALID => x_rsc_13_0_AWVALID,
      AWREADY => x_rsc_13_0_AWREADY,
      WDATA => x_rsc_13_0_i_WDATA,
      WSTRB => x_rsc_13_0_i_WSTRB,
      WLAST => x_rsc_13_0_WLAST,
      WUSER => x_rsc_13_0_i_WUSER,
      WVALID => x_rsc_13_0_WVALID,
      WREADY => x_rsc_13_0_WREADY,
      BID => x_rsc_13_0_i_BID,
      BRESP => x_rsc_13_0_i_BRESP,
      BUSER => x_rsc_13_0_i_BUSER,
      BVALID => x_rsc_13_0_BVALID,
      BREADY => x_rsc_13_0_BREADY,
      ARID => x_rsc_13_0_i_ARID,
      ARADDR => x_rsc_13_0_i_ARADDR,
      ARLEN => x_rsc_13_0_i_ARLEN,
      ARSIZE => x_rsc_13_0_i_ARSIZE,
      ARBURST => x_rsc_13_0_i_ARBURST,
      ARLOCK => x_rsc_13_0_ARLOCK,
      ARCACHE => x_rsc_13_0_i_ARCACHE,
      ARPROT => x_rsc_13_0_i_ARPROT,
      ARQOS => x_rsc_13_0_i_ARQOS,
      ARREGION => x_rsc_13_0_i_ARREGION,
      ARUSER => x_rsc_13_0_i_ARUSER,
      ARVALID => x_rsc_13_0_ARVALID,
      ARREADY => x_rsc_13_0_ARREADY,
      RID => x_rsc_13_0_i_RID,
      RDATA => x_rsc_13_0_i_RDATA,
      RRESP => x_rsc_13_0_i_RRESP,
      RLAST => x_rsc_13_0_RLAST,
      RUSER => x_rsc_13_0_i_RUSER,
      RVALID => x_rsc_13_0_RVALID,
      RREADY => x_rsc_13_0_RREADY,
      s_re => x_rsc_13_0_i_s_re_core_sct,
      s_we => x_rsc_13_0_i_s_we_core_sct,
      s_raddr => x_rsc_13_0_i_s_raddr_1,
      s_waddr => x_rsc_13_0_i_s_waddr_1,
      s_din => x_rsc_13_0_i_s_din_1,
      s_dout => x_rsc_13_0_i_s_dout_1,
      s_rrdy => x_rsc_13_0_i_s_rrdy,
      s_wrdy => x_rsc_13_0_i_s_wrdy,
      is_idle => x_rsc_13_0_is_idle_1,
      tr_write_done => x_rsc_13_0_tr_write_done,
      s_tdone => x_rsc_13_0_s_tdone
    );
  x_rsc_13_0_i_AWID(0) <= x_rsc_13_0_AWID;
  x_rsc_13_0_i_AWADDR <= x_rsc_13_0_AWADDR;
  x_rsc_13_0_i_AWLEN <= x_rsc_13_0_AWLEN;
  x_rsc_13_0_i_AWSIZE <= x_rsc_13_0_AWSIZE;
  x_rsc_13_0_i_AWBURST <= x_rsc_13_0_AWBURST;
  x_rsc_13_0_i_AWCACHE <= x_rsc_13_0_AWCACHE;
  x_rsc_13_0_i_AWPROT <= x_rsc_13_0_AWPROT;
  x_rsc_13_0_i_AWQOS <= x_rsc_13_0_AWQOS;
  x_rsc_13_0_i_AWREGION <= x_rsc_13_0_AWREGION;
  x_rsc_13_0_i_AWUSER(0) <= x_rsc_13_0_AWUSER;
  x_rsc_13_0_i_WDATA <= x_rsc_13_0_WDATA;
  x_rsc_13_0_i_WSTRB <= x_rsc_13_0_WSTRB;
  x_rsc_13_0_i_WUSER(0) <= x_rsc_13_0_WUSER;
  x_rsc_13_0_BID <= x_rsc_13_0_i_BID(0);
  x_rsc_13_0_BRESP <= x_rsc_13_0_i_BRESP;
  x_rsc_13_0_BUSER <= x_rsc_13_0_i_BUSER(0);
  x_rsc_13_0_i_ARID(0) <= x_rsc_13_0_ARID;
  x_rsc_13_0_i_ARADDR <= x_rsc_13_0_ARADDR;
  x_rsc_13_0_i_ARLEN <= x_rsc_13_0_ARLEN;
  x_rsc_13_0_i_ARSIZE <= x_rsc_13_0_ARSIZE;
  x_rsc_13_0_i_ARBURST <= x_rsc_13_0_ARBURST;
  x_rsc_13_0_i_ARCACHE <= x_rsc_13_0_ARCACHE;
  x_rsc_13_0_i_ARPROT <= x_rsc_13_0_ARPROT;
  x_rsc_13_0_i_ARQOS <= x_rsc_13_0_ARQOS;
  x_rsc_13_0_i_ARREGION <= x_rsc_13_0_ARREGION;
  x_rsc_13_0_i_ARUSER(0) <= x_rsc_13_0_ARUSER;
  x_rsc_13_0_RID <= x_rsc_13_0_i_RID(0);
  x_rsc_13_0_RDATA <= x_rsc_13_0_i_RDATA;
  x_rsc_13_0_RRESP <= x_rsc_13_0_i_RRESP;
  x_rsc_13_0_RUSER <= x_rsc_13_0_i_RUSER(0);
  x_rsc_13_0_i_s_raddr_1 <= x_rsc_13_0_i_s_raddr;
  x_rsc_13_0_i_s_waddr_1 <= x_rsc_13_0_i_s_waddr;
  x_rsc_13_0_i_s_din <= x_rsc_13_0_i_s_din_1;
  x_rsc_13_0_i_s_dout_1 <= x_rsc_13_0_i_s_dout;

  hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl_inst : hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_13_0_i_oswt => x_rsc_13_0_i_oswt,
      x_rsc_13_0_i_oswt_1 => x_rsc_13_0_i_oswt_1,
      x_rsc_13_0_i_biwt => x_rsc_13_0_i_biwt,
      x_rsc_13_0_i_bdwt => x_rsc_13_0_i_bdwt,
      x_rsc_13_0_i_bcwt => x_rsc_13_0_i_bcwt,
      x_rsc_13_0_i_s_re_core_sct => x_rsc_13_0_i_s_re_core_sct,
      x_rsc_13_0_i_biwt_1 => x_rsc_13_0_i_biwt_1,
      x_rsc_13_0_i_bdwt_2 => x_rsc_13_0_i_bdwt_2,
      x_rsc_13_0_i_bcwt_1 => x_rsc_13_0_i_bcwt_1,
      x_rsc_13_0_i_s_we_core_sct => x_rsc_13_0_i_s_we_core_sct,
      x_rsc_13_0_i_s_rrdy => x_rsc_13_0_i_s_rrdy,
      x_rsc_13_0_i_s_wrdy => x_rsc_13_0_i_s_wrdy
    );
  hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst : hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_13_0_i_oswt => x_rsc_13_0_i_oswt,
      x_rsc_13_0_i_wen_comp => x_rsc_13_0_i_wen_comp,
      x_rsc_13_0_i_oswt_1 => x_rsc_13_0_i_oswt_1,
      x_rsc_13_0_i_wen_comp_1 => x_rsc_13_0_i_wen_comp_1,
      x_rsc_13_0_i_s_raddr_core => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_raddr_core,
      x_rsc_13_0_i_s_waddr_core => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_waddr_core,
      x_rsc_13_0_i_s_din_mxwt => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_din_mxwt,
      x_rsc_13_0_i_s_dout_core => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_dout_core,
      x_rsc_13_0_i_biwt => x_rsc_13_0_i_biwt,
      x_rsc_13_0_i_bdwt => x_rsc_13_0_i_bdwt,
      x_rsc_13_0_i_bcwt => x_rsc_13_0_i_bcwt,
      x_rsc_13_0_i_biwt_1 => x_rsc_13_0_i_biwt_1,
      x_rsc_13_0_i_bdwt_2 => x_rsc_13_0_i_bdwt_2,
      x_rsc_13_0_i_bcwt_1 => x_rsc_13_0_i_bcwt_1,
      x_rsc_13_0_i_s_raddr => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_raddr,
      x_rsc_13_0_i_s_raddr_core_sct => x_rsc_13_0_i_s_re_core_sct,
      x_rsc_13_0_i_s_waddr => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_waddr,
      x_rsc_13_0_i_s_waddr_core_sct => x_rsc_13_0_i_s_we_core_sct,
      x_rsc_13_0_i_s_din => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_din,
      x_rsc_13_0_i_s_dout => hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_dout
    );
  hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_raddr_core <= x_rsc_13_0_i_s_raddr_core;
  hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_waddr_core <= x_rsc_13_0_i_s_waddr_core;
  x_rsc_13_0_i_s_din_mxwt <= hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_din_mxwt;
  hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_dout_core <= x_rsc_13_0_i_s_dout_core;
  x_rsc_13_0_i_s_raddr <= hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_raddr;
  x_rsc_13_0_i_s_waddr <= hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_waddr;
  hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_din <= x_rsc_13_0_i_s_din;
  x_rsc_13_0_i_s_dout <= hybrid_core_x_rsc_13_0_i_x_rsc_13_0_wait_dp_inst_x_rsc_13_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_12_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_12_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_12_0_s_tdone : IN STD_LOGIC;
    x_rsc_12_0_tr_write_done : IN STD_LOGIC;
    x_rsc_12_0_RREADY : IN STD_LOGIC;
    x_rsc_12_0_RVALID : OUT STD_LOGIC;
    x_rsc_12_0_RUSER : OUT STD_LOGIC;
    x_rsc_12_0_RLAST : OUT STD_LOGIC;
    x_rsc_12_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_RID : OUT STD_LOGIC;
    x_rsc_12_0_ARREADY : OUT STD_LOGIC;
    x_rsc_12_0_ARVALID : IN STD_LOGIC;
    x_rsc_12_0_ARUSER : IN STD_LOGIC;
    x_rsc_12_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARLOCK : IN STD_LOGIC;
    x_rsc_12_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_12_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_12_0_ARID : IN STD_LOGIC;
    x_rsc_12_0_BREADY : IN STD_LOGIC;
    x_rsc_12_0_BVALID : OUT STD_LOGIC;
    x_rsc_12_0_BUSER : OUT STD_LOGIC;
    x_rsc_12_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_BID : OUT STD_LOGIC;
    x_rsc_12_0_WREADY : OUT STD_LOGIC;
    x_rsc_12_0_WVALID : IN STD_LOGIC;
    x_rsc_12_0_WUSER : IN STD_LOGIC;
    x_rsc_12_0_WLAST : IN STD_LOGIC;
    x_rsc_12_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_AWREADY : OUT STD_LOGIC;
    x_rsc_12_0_AWVALID : IN STD_LOGIC;
    x_rsc_12_0_AWUSER : IN STD_LOGIC;
    x_rsc_12_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWLOCK : IN STD_LOGIC;
    x_rsc_12_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_12_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_12_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_12_0_i_oswt : IN STD_LOGIC;
    x_rsc_12_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_12_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_12_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_12_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_12_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_12_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_12_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_12_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_12_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_12_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_12_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_12_0_i_oswt : IN STD_LOGIC;
      x_rsc_12_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_12_0_i_biwt : OUT STD_LOGIC;
      x_rsc_12_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_12_0_i_bcwt : IN STD_LOGIC;
      x_rsc_12_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_12_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_12_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_12_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_12_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_12_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_12_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_12_0_i_oswt : IN STD_LOGIC;
      x_rsc_12_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_12_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_12_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_12_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_12_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_12_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_i_biwt : IN STD_LOGIC;
      x_rsc_12_0_i_bdwt : IN STD_LOGIC;
      x_rsc_12_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_12_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_12_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_12_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_12_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_12_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_12_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_12_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_12_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_12_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_12_0_i_AWID,
      AWADDR => x_rsc_12_0_i_AWADDR,
      AWLEN => x_rsc_12_0_i_AWLEN,
      AWSIZE => x_rsc_12_0_i_AWSIZE,
      AWBURST => x_rsc_12_0_i_AWBURST,
      AWLOCK => x_rsc_12_0_AWLOCK,
      AWCACHE => x_rsc_12_0_i_AWCACHE,
      AWPROT => x_rsc_12_0_i_AWPROT,
      AWQOS => x_rsc_12_0_i_AWQOS,
      AWREGION => x_rsc_12_0_i_AWREGION,
      AWUSER => x_rsc_12_0_i_AWUSER,
      AWVALID => x_rsc_12_0_AWVALID,
      AWREADY => x_rsc_12_0_AWREADY,
      WDATA => x_rsc_12_0_i_WDATA,
      WSTRB => x_rsc_12_0_i_WSTRB,
      WLAST => x_rsc_12_0_WLAST,
      WUSER => x_rsc_12_0_i_WUSER,
      WVALID => x_rsc_12_0_WVALID,
      WREADY => x_rsc_12_0_WREADY,
      BID => x_rsc_12_0_i_BID,
      BRESP => x_rsc_12_0_i_BRESP,
      BUSER => x_rsc_12_0_i_BUSER,
      BVALID => x_rsc_12_0_BVALID,
      BREADY => x_rsc_12_0_BREADY,
      ARID => x_rsc_12_0_i_ARID,
      ARADDR => x_rsc_12_0_i_ARADDR,
      ARLEN => x_rsc_12_0_i_ARLEN,
      ARSIZE => x_rsc_12_0_i_ARSIZE,
      ARBURST => x_rsc_12_0_i_ARBURST,
      ARLOCK => x_rsc_12_0_ARLOCK,
      ARCACHE => x_rsc_12_0_i_ARCACHE,
      ARPROT => x_rsc_12_0_i_ARPROT,
      ARQOS => x_rsc_12_0_i_ARQOS,
      ARREGION => x_rsc_12_0_i_ARREGION,
      ARUSER => x_rsc_12_0_i_ARUSER,
      ARVALID => x_rsc_12_0_ARVALID,
      ARREADY => x_rsc_12_0_ARREADY,
      RID => x_rsc_12_0_i_RID,
      RDATA => x_rsc_12_0_i_RDATA,
      RRESP => x_rsc_12_0_i_RRESP,
      RLAST => x_rsc_12_0_RLAST,
      RUSER => x_rsc_12_0_i_RUSER,
      RVALID => x_rsc_12_0_RVALID,
      RREADY => x_rsc_12_0_RREADY,
      s_re => x_rsc_12_0_i_s_re_core_sct,
      s_we => x_rsc_12_0_i_s_we_core_sct,
      s_raddr => x_rsc_12_0_i_s_raddr_1,
      s_waddr => x_rsc_12_0_i_s_waddr_1,
      s_din => x_rsc_12_0_i_s_din_1,
      s_dout => x_rsc_12_0_i_s_dout_1,
      s_rrdy => x_rsc_12_0_i_s_rrdy,
      s_wrdy => x_rsc_12_0_i_s_wrdy,
      is_idle => x_rsc_12_0_is_idle_1,
      tr_write_done => x_rsc_12_0_tr_write_done,
      s_tdone => x_rsc_12_0_s_tdone
    );
  x_rsc_12_0_i_AWID(0) <= x_rsc_12_0_AWID;
  x_rsc_12_0_i_AWADDR <= x_rsc_12_0_AWADDR;
  x_rsc_12_0_i_AWLEN <= x_rsc_12_0_AWLEN;
  x_rsc_12_0_i_AWSIZE <= x_rsc_12_0_AWSIZE;
  x_rsc_12_0_i_AWBURST <= x_rsc_12_0_AWBURST;
  x_rsc_12_0_i_AWCACHE <= x_rsc_12_0_AWCACHE;
  x_rsc_12_0_i_AWPROT <= x_rsc_12_0_AWPROT;
  x_rsc_12_0_i_AWQOS <= x_rsc_12_0_AWQOS;
  x_rsc_12_0_i_AWREGION <= x_rsc_12_0_AWREGION;
  x_rsc_12_0_i_AWUSER(0) <= x_rsc_12_0_AWUSER;
  x_rsc_12_0_i_WDATA <= x_rsc_12_0_WDATA;
  x_rsc_12_0_i_WSTRB <= x_rsc_12_0_WSTRB;
  x_rsc_12_0_i_WUSER(0) <= x_rsc_12_0_WUSER;
  x_rsc_12_0_BID <= x_rsc_12_0_i_BID(0);
  x_rsc_12_0_BRESP <= x_rsc_12_0_i_BRESP;
  x_rsc_12_0_BUSER <= x_rsc_12_0_i_BUSER(0);
  x_rsc_12_0_i_ARID(0) <= x_rsc_12_0_ARID;
  x_rsc_12_0_i_ARADDR <= x_rsc_12_0_ARADDR;
  x_rsc_12_0_i_ARLEN <= x_rsc_12_0_ARLEN;
  x_rsc_12_0_i_ARSIZE <= x_rsc_12_0_ARSIZE;
  x_rsc_12_0_i_ARBURST <= x_rsc_12_0_ARBURST;
  x_rsc_12_0_i_ARCACHE <= x_rsc_12_0_ARCACHE;
  x_rsc_12_0_i_ARPROT <= x_rsc_12_0_ARPROT;
  x_rsc_12_0_i_ARQOS <= x_rsc_12_0_ARQOS;
  x_rsc_12_0_i_ARREGION <= x_rsc_12_0_ARREGION;
  x_rsc_12_0_i_ARUSER(0) <= x_rsc_12_0_ARUSER;
  x_rsc_12_0_RID <= x_rsc_12_0_i_RID(0);
  x_rsc_12_0_RDATA <= x_rsc_12_0_i_RDATA;
  x_rsc_12_0_RRESP <= x_rsc_12_0_i_RRESP;
  x_rsc_12_0_RUSER <= x_rsc_12_0_i_RUSER(0);
  x_rsc_12_0_i_s_raddr_1 <= x_rsc_12_0_i_s_raddr;
  x_rsc_12_0_i_s_waddr_1 <= x_rsc_12_0_i_s_waddr;
  x_rsc_12_0_i_s_din <= x_rsc_12_0_i_s_din_1;
  x_rsc_12_0_i_s_dout_1 <= x_rsc_12_0_i_s_dout;

  hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl_inst : hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_12_0_i_oswt => x_rsc_12_0_i_oswt,
      x_rsc_12_0_i_oswt_1 => x_rsc_12_0_i_oswt_1,
      x_rsc_12_0_i_biwt => x_rsc_12_0_i_biwt,
      x_rsc_12_0_i_bdwt => x_rsc_12_0_i_bdwt,
      x_rsc_12_0_i_bcwt => x_rsc_12_0_i_bcwt,
      x_rsc_12_0_i_s_re_core_sct => x_rsc_12_0_i_s_re_core_sct,
      x_rsc_12_0_i_biwt_1 => x_rsc_12_0_i_biwt_1,
      x_rsc_12_0_i_bdwt_2 => x_rsc_12_0_i_bdwt_2,
      x_rsc_12_0_i_bcwt_1 => x_rsc_12_0_i_bcwt_1,
      x_rsc_12_0_i_s_we_core_sct => x_rsc_12_0_i_s_we_core_sct,
      x_rsc_12_0_i_s_rrdy => x_rsc_12_0_i_s_rrdy,
      x_rsc_12_0_i_s_wrdy => x_rsc_12_0_i_s_wrdy
    );
  hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst : hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_12_0_i_oswt => x_rsc_12_0_i_oswt,
      x_rsc_12_0_i_wen_comp => x_rsc_12_0_i_wen_comp,
      x_rsc_12_0_i_oswt_1 => x_rsc_12_0_i_oswt_1,
      x_rsc_12_0_i_wen_comp_1 => x_rsc_12_0_i_wen_comp_1,
      x_rsc_12_0_i_s_raddr_core => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_raddr_core,
      x_rsc_12_0_i_s_waddr_core => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_waddr_core,
      x_rsc_12_0_i_s_din_mxwt => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_din_mxwt,
      x_rsc_12_0_i_s_dout_core => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_dout_core,
      x_rsc_12_0_i_biwt => x_rsc_12_0_i_biwt,
      x_rsc_12_0_i_bdwt => x_rsc_12_0_i_bdwt,
      x_rsc_12_0_i_bcwt => x_rsc_12_0_i_bcwt,
      x_rsc_12_0_i_biwt_1 => x_rsc_12_0_i_biwt_1,
      x_rsc_12_0_i_bdwt_2 => x_rsc_12_0_i_bdwt_2,
      x_rsc_12_0_i_bcwt_1 => x_rsc_12_0_i_bcwt_1,
      x_rsc_12_0_i_s_raddr => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_raddr,
      x_rsc_12_0_i_s_raddr_core_sct => x_rsc_12_0_i_s_re_core_sct,
      x_rsc_12_0_i_s_waddr => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_waddr,
      x_rsc_12_0_i_s_waddr_core_sct => x_rsc_12_0_i_s_we_core_sct,
      x_rsc_12_0_i_s_din => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_din,
      x_rsc_12_0_i_s_dout => hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_dout
    );
  hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_raddr_core <= x_rsc_12_0_i_s_raddr_core;
  hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_waddr_core <= x_rsc_12_0_i_s_waddr_core;
  x_rsc_12_0_i_s_din_mxwt <= hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_din_mxwt;
  hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_dout_core <= x_rsc_12_0_i_s_dout_core;
  x_rsc_12_0_i_s_raddr <= hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_raddr;
  x_rsc_12_0_i_s_waddr <= hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_waddr;
  hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_din <= x_rsc_12_0_i_s_din;
  x_rsc_12_0_i_s_dout <= hybrid_core_x_rsc_12_0_i_x_rsc_12_0_wait_dp_inst_x_rsc_12_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_11_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_11_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_11_0_s_tdone : IN STD_LOGIC;
    x_rsc_11_0_tr_write_done : IN STD_LOGIC;
    x_rsc_11_0_RREADY : IN STD_LOGIC;
    x_rsc_11_0_RVALID : OUT STD_LOGIC;
    x_rsc_11_0_RUSER : OUT STD_LOGIC;
    x_rsc_11_0_RLAST : OUT STD_LOGIC;
    x_rsc_11_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_RID : OUT STD_LOGIC;
    x_rsc_11_0_ARREADY : OUT STD_LOGIC;
    x_rsc_11_0_ARVALID : IN STD_LOGIC;
    x_rsc_11_0_ARUSER : IN STD_LOGIC;
    x_rsc_11_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARLOCK : IN STD_LOGIC;
    x_rsc_11_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_11_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_11_0_ARID : IN STD_LOGIC;
    x_rsc_11_0_BREADY : IN STD_LOGIC;
    x_rsc_11_0_BVALID : OUT STD_LOGIC;
    x_rsc_11_0_BUSER : OUT STD_LOGIC;
    x_rsc_11_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_BID : OUT STD_LOGIC;
    x_rsc_11_0_WREADY : OUT STD_LOGIC;
    x_rsc_11_0_WVALID : IN STD_LOGIC;
    x_rsc_11_0_WUSER : IN STD_LOGIC;
    x_rsc_11_0_WLAST : IN STD_LOGIC;
    x_rsc_11_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_AWREADY : OUT STD_LOGIC;
    x_rsc_11_0_AWVALID : IN STD_LOGIC;
    x_rsc_11_0_AWUSER : IN STD_LOGIC;
    x_rsc_11_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWLOCK : IN STD_LOGIC;
    x_rsc_11_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_11_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_11_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_11_0_i_oswt : IN STD_LOGIC;
    x_rsc_11_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_11_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_11_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_11_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_11_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_11_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_11_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_11_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_11_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_11_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_11_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_11_0_i_oswt : IN STD_LOGIC;
      x_rsc_11_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_11_0_i_biwt : OUT STD_LOGIC;
      x_rsc_11_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_11_0_i_bcwt : IN STD_LOGIC;
      x_rsc_11_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_11_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_11_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_11_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_11_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_11_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_11_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_11_0_i_oswt : IN STD_LOGIC;
      x_rsc_11_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_11_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_11_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_11_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_11_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_11_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_i_biwt : IN STD_LOGIC;
      x_rsc_11_0_i_bdwt : IN STD_LOGIC;
      x_rsc_11_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_11_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_11_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_11_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_11_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_11_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_11_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_11_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_11_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_11_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_11_0_i_AWID,
      AWADDR => x_rsc_11_0_i_AWADDR,
      AWLEN => x_rsc_11_0_i_AWLEN,
      AWSIZE => x_rsc_11_0_i_AWSIZE,
      AWBURST => x_rsc_11_0_i_AWBURST,
      AWLOCK => x_rsc_11_0_AWLOCK,
      AWCACHE => x_rsc_11_0_i_AWCACHE,
      AWPROT => x_rsc_11_0_i_AWPROT,
      AWQOS => x_rsc_11_0_i_AWQOS,
      AWREGION => x_rsc_11_0_i_AWREGION,
      AWUSER => x_rsc_11_0_i_AWUSER,
      AWVALID => x_rsc_11_0_AWVALID,
      AWREADY => x_rsc_11_0_AWREADY,
      WDATA => x_rsc_11_0_i_WDATA,
      WSTRB => x_rsc_11_0_i_WSTRB,
      WLAST => x_rsc_11_0_WLAST,
      WUSER => x_rsc_11_0_i_WUSER,
      WVALID => x_rsc_11_0_WVALID,
      WREADY => x_rsc_11_0_WREADY,
      BID => x_rsc_11_0_i_BID,
      BRESP => x_rsc_11_0_i_BRESP,
      BUSER => x_rsc_11_0_i_BUSER,
      BVALID => x_rsc_11_0_BVALID,
      BREADY => x_rsc_11_0_BREADY,
      ARID => x_rsc_11_0_i_ARID,
      ARADDR => x_rsc_11_0_i_ARADDR,
      ARLEN => x_rsc_11_0_i_ARLEN,
      ARSIZE => x_rsc_11_0_i_ARSIZE,
      ARBURST => x_rsc_11_0_i_ARBURST,
      ARLOCK => x_rsc_11_0_ARLOCK,
      ARCACHE => x_rsc_11_0_i_ARCACHE,
      ARPROT => x_rsc_11_0_i_ARPROT,
      ARQOS => x_rsc_11_0_i_ARQOS,
      ARREGION => x_rsc_11_0_i_ARREGION,
      ARUSER => x_rsc_11_0_i_ARUSER,
      ARVALID => x_rsc_11_0_ARVALID,
      ARREADY => x_rsc_11_0_ARREADY,
      RID => x_rsc_11_0_i_RID,
      RDATA => x_rsc_11_0_i_RDATA,
      RRESP => x_rsc_11_0_i_RRESP,
      RLAST => x_rsc_11_0_RLAST,
      RUSER => x_rsc_11_0_i_RUSER,
      RVALID => x_rsc_11_0_RVALID,
      RREADY => x_rsc_11_0_RREADY,
      s_re => x_rsc_11_0_i_s_re_core_sct,
      s_we => x_rsc_11_0_i_s_we_core_sct,
      s_raddr => x_rsc_11_0_i_s_raddr_1,
      s_waddr => x_rsc_11_0_i_s_waddr_1,
      s_din => x_rsc_11_0_i_s_din_1,
      s_dout => x_rsc_11_0_i_s_dout_1,
      s_rrdy => x_rsc_11_0_i_s_rrdy,
      s_wrdy => x_rsc_11_0_i_s_wrdy,
      is_idle => x_rsc_11_0_is_idle_1,
      tr_write_done => x_rsc_11_0_tr_write_done,
      s_tdone => x_rsc_11_0_s_tdone
    );
  x_rsc_11_0_i_AWID(0) <= x_rsc_11_0_AWID;
  x_rsc_11_0_i_AWADDR <= x_rsc_11_0_AWADDR;
  x_rsc_11_0_i_AWLEN <= x_rsc_11_0_AWLEN;
  x_rsc_11_0_i_AWSIZE <= x_rsc_11_0_AWSIZE;
  x_rsc_11_0_i_AWBURST <= x_rsc_11_0_AWBURST;
  x_rsc_11_0_i_AWCACHE <= x_rsc_11_0_AWCACHE;
  x_rsc_11_0_i_AWPROT <= x_rsc_11_0_AWPROT;
  x_rsc_11_0_i_AWQOS <= x_rsc_11_0_AWQOS;
  x_rsc_11_0_i_AWREGION <= x_rsc_11_0_AWREGION;
  x_rsc_11_0_i_AWUSER(0) <= x_rsc_11_0_AWUSER;
  x_rsc_11_0_i_WDATA <= x_rsc_11_0_WDATA;
  x_rsc_11_0_i_WSTRB <= x_rsc_11_0_WSTRB;
  x_rsc_11_0_i_WUSER(0) <= x_rsc_11_0_WUSER;
  x_rsc_11_0_BID <= x_rsc_11_0_i_BID(0);
  x_rsc_11_0_BRESP <= x_rsc_11_0_i_BRESP;
  x_rsc_11_0_BUSER <= x_rsc_11_0_i_BUSER(0);
  x_rsc_11_0_i_ARID(0) <= x_rsc_11_0_ARID;
  x_rsc_11_0_i_ARADDR <= x_rsc_11_0_ARADDR;
  x_rsc_11_0_i_ARLEN <= x_rsc_11_0_ARLEN;
  x_rsc_11_0_i_ARSIZE <= x_rsc_11_0_ARSIZE;
  x_rsc_11_0_i_ARBURST <= x_rsc_11_0_ARBURST;
  x_rsc_11_0_i_ARCACHE <= x_rsc_11_0_ARCACHE;
  x_rsc_11_0_i_ARPROT <= x_rsc_11_0_ARPROT;
  x_rsc_11_0_i_ARQOS <= x_rsc_11_0_ARQOS;
  x_rsc_11_0_i_ARREGION <= x_rsc_11_0_ARREGION;
  x_rsc_11_0_i_ARUSER(0) <= x_rsc_11_0_ARUSER;
  x_rsc_11_0_RID <= x_rsc_11_0_i_RID(0);
  x_rsc_11_0_RDATA <= x_rsc_11_0_i_RDATA;
  x_rsc_11_0_RRESP <= x_rsc_11_0_i_RRESP;
  x_rsc_11_0_RUSER <= x_rsc_11_0_i_RUSER(0);
  x_rsc_11_0_i_s_raddr_1 <= x_rsc_11_0_i_s_raddr;
  x_rsc_11_0_i_s_waddr_1 <= x_rsc_11_0_i_s_waddr;
  x_rsc_11_0_i_s_din <= x_rsc_11_0_i_s_din_1;
  x_rsc_11_0_i_s_dout_1 <= x_rsc_11_0_i_s_dout;

  hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl_inst : hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_11_0_i_oswt => x_rsc_11_0_i_oswt,
      x_rsc_11_0_i_oswt_1 => x_rsc_11_0_i_oswt_1,
      x_rsc_11_0_i_biwt => x_rsc_11_0_i_biwt,
      x_rsc_11_0_i_bdwt => x_rsc_11_0_i_bdwt,
      x_rsc_11_0_i_bcwt => x_rsc_11_0_i_bcwt,
      x_rsc_11_0_i_s_re_core_sct => x_rsc_11_0_i_s_re_core_sct,
      x_rsc_11_0_i_biwt_1 => x_rsc_11_0_i_biwt_1,
      x_rsc_11_0_i_bdwt_2 => x_rsc_11_0_i_bdwt_2,
      x_rsc_11_0_i_bcwt_1 => x_rsc_11_0_i_bcwt_1,
      x_rsc_11_0_i_s_we_core_sct => x_rsc_11_0_i_s_we_core_sct,
      x_rsc_11_0_i_s_rrdy => x_rsc_11_0_i_s_rrdy,
      x_rsc_11_0_i_s_wrdy => x_rsc_11_0_i_s_wrdy
    );
  hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst : hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_11_0_i_oswt => x_rsc_11_0_i_oswt,
      x_rsc_11_0_i_wen_comp => x_rsc_11_0_i_wen_comp,
      x_rsc_11_0_i_oswt_1 => x_rsc_11_0_i_oswt_1,
      x_rsc_11_0_i_wen_comp_1 => x_rsc_11_0_i_wen_comp_1,
      x_rsc_11_0_i_s_raddr_core => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_raddr_core,
      x_rsc_11_0_i_s_waddr_core => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_waddr_core,
      x_rsc_11_0_i_s_din_mxwt => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_din_mxwt,
      x_rsc_11_0_i_s_dout_core => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_dout_core,
      x_rsc_11_0_i_biwt => x_rsc_11_0_i_biwt,
      x_rsc_11_0_i_bdwt => x_rsc_11_0_i_bdwt,
      x_rsc_11_0_i_bcwt => x_rsc_11_0_i_bcwt,
      x_rsc_11_0_i_biwt_1 => x_rsc_11_0_i_biwt_1,
      x_rsc_11_0_i_bdwt_2 => x_rsc_11_0_i_bdwt_2,
      x_rsc_11_0_i_bcwt_1 => x_rsc_11_0_i_bcwt_1,
      x_rsc_11_0_i_s_raddr => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_raddr,
      x_rsc_11_0_i_s_raddr_core_sct => x_rsc_11_0_i_s_re_core_sct,
      x_rsc_11_0_i_s_waddr => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_waddr,
      x_rsc_11_0_i_s_waddr_core_sct => x_rsc_11_0_i_s_we_core_sct,
      x_rsc_11_0_i_s_din => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_din,
      x_rsc_11_0_i_s_dout => hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_dout
    );
  hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_raddr_core <= x_rsc_11_0_i_s_raddr_core;
  hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_waddr_core <= x_rsc_11_0_i_s_waddr_core;
  x_rsc_11_0_i_s_din_mxwt <= hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_din_mxwt;
  hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_dout_core <= x_rsc_11_0_i_s_dout_core;
  x_rsc_11_0_i_s_raddr <= hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_raddr;
  x_rsc_11_0_i_s_waddr <= hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_waddr;
  hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_din <= x_rsc_11_0_i_s_din;
  x_rsc_11_0_i_s_dout <= hybrid_core_x_rsc_11_0_i_x_rsc_11_0_wait_dp_inst_x_rsc_11_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_10_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_10_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_10_0_s_tdone : IN STD_LOGIC;
    x_rsc_10_0_tr_write_done : IN STD_LOGIC;
    x_rsc_10_0_RREADY : IN STD_LOGIC;
    x_rsc_10_0_RVALID : OUT STD_LOGIC;
    x_rsc_10_0_RUSER : OUT STD_LOGIC;
    x_rsc_10_0_RLAST : OUT STD_LOGIC;
    x_rsc_10_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_RID : OUT STD_LOGIC;
    x_rsc_10_0_ARREADY : OUT STD_LOGIC;
    x_rsc_10_0_ARVALID : IN STD_LOGIC;
    x_rsc_10_0_ARUSER : IN STD_LOGIC;
    x_rsc_10_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARLOCK : IN STD_LOGIC;
    x_rsc_10_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_10_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_10_0_ARID : IN STD_LOGIC;
    x_rsc_10_0_BREADY : IN STD_LOGIC;
    x_rsc_10_0_BVALID : OUT STD_LOGIC;
    x_rsc_10_0_BUSER : OUT STD_LOGIC;
    x_rsc_10_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_BID : OUT STD_LOGIC;
    x_rsc_10_0_WREADY : OUT STD_LOGIC;
    x_rsc_10_0_WVALID : IN STD_LOGIC;
    x_rsc_10_0_WUSER : IN STD_LOGIC;
    x_rsc_10_0_WLAST : IN STD_LOGIC;
    x_rsc_10_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_AWREADY : OUT STD_LOGIC;
    x_rsc_10_0_AWVALID : IN STD_LOGIC;
    x_rsc_10_0_AWUSER : IN STD_LOGIC;
    x_rsc_10_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWLOCK : IN STD_LOGIC;
    x_rsc_10_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_10_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_10_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_10_0_i_oswt : IN STD_LOGIC;
    x_rsc_10_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_10_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_10_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_10_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_10_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_10_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_10_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_10_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_10_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_10_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_10_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_10_0_i_oswt : IN STD_LOGIC;
      x_rsc_10_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_10_0_i_biwt : OUT STD_LOGIC;
      x_rsc_10_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_10_0_i_bcwt : IN STD_LOGIC;
      x_rsc_10_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_10_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_10_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_10_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_10_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_10_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_10_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_10_0_i_oswt : IN STD_LOGIC;
      x_rsc_10_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_10_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_10_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_10_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_10_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_10_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_i_biwt : IN STD_LOGIC;
      x_rsc_10_0_i_bdwt : IN STD_LOGIC;
      x_rsc_10_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_10_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_10_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_10_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_10_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_10_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_10_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_10_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_10_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_dout_core
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_raddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_waddr :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_10_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_10_0_i_AWID,
      AWADDR => x_rsc_10_0_i_AWADDR,
      AWLEN => x_rsc_10_0_i_AWLEN,
      AWSIZE => x_rsc_10_0_i_AWSIZE,
      AWBURST => x_rsc_10_0_i_AWBURST,
      AWLOCK => x_rsc_10_0_AWLOCK,
      AWCACHE => x_rsc_10_0_i_AWCACHE,
      AWPROT => x_rsc_10_0_i_AWPROT,
      AWQOS => x_rsc_10_0_i_AWQOS,
      AWREGION => x_rsc_10_0_i_AWREGION,
      AWUSER => x_rsc_10_0_i_AWUSER,
      AWVALID => x_rsc_10_0_AWVALID,
      AWREADY => x_rsc_10_0_AWREADY,
      WDATA => x_rsc_10_0_i_WDATA,
      WSTRB => x_rsc_10_0_i_WSTRB,
      WLAST => x_rsc_10_0_WLAST,
      WUSER => x_rsc_10_0_i_WUSER,
      WVALID => x_rsc_10_0_WVALID,
      WREADY => x_rsc_10_0_WREADY,
      BID => x_rsc_10_0_i_BID,
      BRESP => x_rsc_10_0_i_BRESP,
      BUSER => x_rsc_10_0_i_BUSER,
      BVALID => x_rsc_10_0_BVALID,
      BREADY => x_rsc_10_0_BREADY,
      ARID => x_rsc_10_0_i_ARID,
      ARADDR => x_rsc_10_0_i_ARADDR,
      ARLEN => x_rsc_10_0_i_ARLEN,
      ARSIZE => x_rsc_10_0_i_ARSIZE,
      ARBURST => x_rsc_10_0_i_ARBURST,
      ARLOCK => x_rsc_10_0_ARLOCK,
      ARCACHE => x_rsc_10_0_i_ARCACHE,
      ARPROT => x_rsc_10_0_i_ARPROT,
      ARQOS => x_rsc_10_0_i_ARQOS,
      ARREGION => x_rsc_10_0_i_ARREGION,
      ARUSER => x_rsc_10_0_i_ARUSER,
      ARVALID => x_rsc_10_0_ARVALID,
      ARREADY => x_rsc_10_0_ARREADY,
      RID => x_rsc_10_0_i_RID,
      RDATA => x_rsc_10_0_i_RDATA,
      RRESP => x_rsc_10_0_i_RRESP,
      RLAST => x_rsc_10_0_RLAST,
      RUSER => x_rsc_10_0_i_RUSER,
      RVALID => x_rsc_10_0_RVALID,
      RREADY => x_rsc_10_0_RREADY,
      s_re => x_rsc_10_0_i_s_re_core_sct,
      s_we => x_rsc_10_0_i_s_we_core_sct,
      s_raddr => x_rsc_10_0_i_s_raddr_1,
      s_waddr => x_rsc_10_0_i_s_waddr_1,
      s_din => x_rsc_10_0_i_s_din_1,
      s_dout => x_rsc_10_0_i_s_dout_1,
      s_rrdy => x_rsc_10_0_i_s_rrdy,
      s_wrdy => x_rsc_10_0_i_s_wrdy,
      is_idle => x_rsc_10_0_is_idle_1,
      tr_write_done => x_rsc_10_0_tr_write_done,
      s_tdone => x_rsc_10_0_s_tdone
    );
  x_rsc_10_0_i_AWID(0) <= x_rsc_10_0_AWID;
  x_rsc_10_0_i_AWADDR <= x_rsc_10_0_AWADDR;
  x_rsc_10_0_i_AWLEN <= x_rsc_10_0_AWLEN;
  x_rsc_10_0_i_AWSIZE <= x_rsc_10_0_AWSIZE;
  x_rsc_10_0_i_AWBURST <= x_rsc_10_0_AWBURST;
  x_rsc_10_0_i_AWCACHE <= x_rsc_10_0_AWCACHE;
  x_rsc_10_0_i_AWPROT <= x_rsc_10_0_AWPROT;
  x_rsc_10_0_i_AWQOS <= x_rsc_10_0_AWQOS;
  x_rsc_10_0_i_AWREGION <= x_rsc_10_0_AWREGION;
  x_rsc_10_0_i_AWUSER(0) <= x_rsc_10_0_AWUSER;
  x_rsc_10_0_i_WDATA <= x_rsc_10_0_WDATA;
  x_rsc_10_0_i_WSTRB <= x_rsc_10_0_WSTRB;
  x_rsc_10_0_i_WUSER(0) <= x_rsc_10_0_WUSER;
  x_rsc_10_0_BID <= x_rsc_10_0_i_BID(0);
  x_rsc_10_0_BRESP <= x_rsc_10_0_i_BRESP;
  x_rsc_10_0_BUSER <= x_rsc_10_0_i_BUSER(0);
  x_rsc_10_0_i_ARID(0) <= x_rsc_10_0_ARID;
  x_rsc_10_0_i_ARADDR <= x_rsc_10_0_ARADDR;
  x_rsc_10_0_i_ARLEN <= x_rsc_10_0_ARLEN;
  x_rsc_10_0_i_ARSIZE <= x_rsc_10_0_ARSIZE;
  x_rsc_10_0_i_ARBURST <= x_rsc_10_0_ARBURST;
  x_rsc_10_0_i_ARCACHE <= x_rsc_10_0_ARCACHE;
  x_rsc_10_0_i_ARPROT <= x_rsc_10_0_ARPROT;
  x_rsc_10_0_i_ARQOS <= x_rsc_10_0_ARQOS;
  x_rsc_10_0_i_ARREGION <= x_rsc_10_0_ARREGION;
  x_rsc_10_0_i_ARUSER(0) <= x_rsc_10_0_ARUSER;
  x_rsc_10_0_RID <= x_rsc_10_0_i_RID(0);
  x_rsc_10_0_RDATA <= x_rsc_10_0_i_RDATA;
  x_rsc_10_0_RRESP <= x_rsc_10_0_i_RRESP;
  x_rsc_10_0_RUSER <= x_rsc_10_0_i_RUSER(0);
  x_rsc_10_0_i_s_raddr_1 <= x_rsc_10_0_i_s_raddr;
  x_rsc_10_0_i_s_waddr_1 <= x_rsc_10_0_i_s_waddr;
  x_rsc_10_0_i_s_din <= x_rsc_10_0_i_s_din_1;
  x_rsc_10_0_i_s_dout_1 <= x_rsc_10_0_i_s_dout;

  hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl_inst : hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_10_0_i_oswt => x_rsc_10_0_i_oswt,
      x_rsc_10_0_i_oswt_1 => x_rsc_10_0_i_oswt_1,
      x_rsc_10_0_i_biwt => x_rsc_10_0_i_biwt,
      x_rsc_10_0_i_bdwt => x_rsc_10_0_i_bdwt,
      x_rsc_10_0_i_bcwt => x_rsc_10_0_i_bcwt,
      x_rsc_10_0_i_s_re_core_sct => x_rsc_10_0_i_s_re_core_sct,
      x_rsc_10_0_i_biwt_1 => x_rsc_10_0_i_biwt_1,
      x_rsc_10_0_i_bdwt_2 => x_rsc_10_0_i_bdwt_2,
      x_rsc_10_0_i_bcwt_1 => x_rsc_10_0_i_bcwt_1,
      x_rsc_10_0_i_s_we_core_sct => x_rsc_10_0_i_s_we_core_sct,
      x_rsc_10_0_i_s_rrdy => x_rsc_10_0_i_s_rrdy,
      x_rsc_10_0_i_s_wrdy => x_rsc_10_0_i_s_wrdy
    );
  hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst : hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_10_0_i_oswt => x_rsc_10_0_i_oswt,
      x_rsc_10_0_i_wen_comp => x_rsc_10_0_i_wen_comp,
      x_rsc_10_0_i_oswt_1 => x_rsc_10_0_i_oswt_1,
      x_rsc_10_0_i_wen_comp_1 => x_rsc_10_0_i_wen_comp_1,
      x_rsc_10_0_i_s_raddr_core => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_raddr_core,
      x_rsc_10_0_i_s_waddr_core => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_waddr_core,
      x_rsc_10_0_i_s_din_mxwt => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_din_mxwt,
      x_rsc_10_0_i_s_dout_core => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_dout_core,
      x_rsc_10_0_i_biwt => x_rsc_10_0_i_biwt,
      x_rsc_10_0_i_bdwt => x_rsc_10_0_i_bdwt,
      x_rsc_10_0_i_bcwt => x_rsc_10_0_i_bcwt,
      x_rsc_10_0_i_biwt_1 => x_rsc_10_0_i_biwt_1,
      x_rsc_10_0_i_bdwt_2 => x_rsc_10_0_i_bdwt_2,
      x_rsc_10_0_i_bcwt_1 => x_rsc_10_0_i_bcwt_1,
      x_rsc_10_0_i_s_raddr => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_raddr,
      x_rsc_10_0_i_s_raddr_core_sct => x_rsc_10_0_i_s_re_core_sct,
      x_rsc_10_0_i_s_waddr => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_waddr,
      x_rsc_10_0_i_s_waddr_core_sct => x_rsc_10_0_i_s_we_core_sct,
      x_rsc_10_0_i_s_din => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_din,
      x_rsc_10_0_i_s_dout => hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_dout
    );
  hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_raddr_core <= x_rsc_10_0_i_s_raddr_core;
  hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_waddr_core <= x_rsc_10_0_i_s_waddr_core;
  x_rsc_10_0_i_s_din_mxwt <= hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_din_mxwt;
  hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_dout_core <= x_rsc_10_0_i_s_dout_core;
  x_rsc_10_0_i_s_raddr <= hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_raddr;
  x_rsc_10_0_i_s_waddr <= hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_waddr;
  hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_din <= x_rsc_10_0_i_s_din;
  x_rsc_10_0_i_s_dout <= hybrid_core_x_rsc_10_0_i_x_rsc_10_0_wait_dp_inst_x_rsc_10_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_9_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_9_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_9_0_s_tdone : IN STD_LOGIC;
    x_rsc_9_0_tr_write_done : IN STD_LOGIC;
    x_rsc_9_0_RREADY : IN STD_LOGIC;
    x_rsc_9_0_RVALID : OUT STD_LOGIC;
    x_rsc_9_0_RUSER : OUT STD_LOGIC;
    x_rsc_9_0_RLAST : OUT STD_LOGIC;
    x_rsc_9_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_RID : OUT STD_LOGIC;
    x_rsc_9_0_ARREADY : OUT STD_LOGIC;
    x_rsc_9_0_ARVALID : IN STD_LOGIC;
    x_rsc_9_0_ARUSER : IN STD_LOGIC;
    x_rsc_9_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARLOCK : IN STD_LOGIC;
    x_rsc_9_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_9_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_9_0_ARID : IN STD_LOGIC;
    x_rsc_9_0_BREADY : IN STD_LOGIC;
    x_rsc_9_0_BVALID : OUT STD_LOGIC;
    x_rsc_9_0_BUSER : OUT STD_LOGIC;
    x_rsc_9_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_BID : OUT STD_LOGIC;
    x_rsc_9_0_WREADY : OUT STD_LOGIC;
    x_rsc_9_0_WVALID : IN STD_LOGIC;
    x_rsc_9_0_WUSER : IN STD_LOGIC;
    x_rsc_9_0_WLAST : IN STD_LOGIC;
    x_rsc_9_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_AWREADY : OUT STD_LOGIC;
    x_rsc_9_0_AWVALID : IN STD_LOGIC;
    x_rsc_9_0_AWUSER : IN STD_LOGIC;
    x_rsc_9_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWLOCK : IN STD_LOGIC;
    x_rsc_9_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_9_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_9_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_9_0_i_oswt : IN STD_LOGIC;
    x_rsc_9_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_9_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_9_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_9_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_9_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_9_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_9_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_9_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_9_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_9_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_9_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_9_0_i_oswt : IN STD_LOGIC;
      x_rsc_9_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_9_0_i_biwt : OUT STD_LOGIC;
      x_rsc_9_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_9_0_i_bcwt : IN STD_LOGIC;
      x_rsc_9_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_9_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_9_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_9_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_9_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_9_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_9_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_9_0_i_oswt : IN STD_LOGIC;
      x_rsc_9_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_9_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_9_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_9_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_9_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_9_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_i_biwt : IN STD_LOGIC;
      x_rsc_9_0_i_bdwt : IN STD_LOGIC;
      x_rsc_9_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_9_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_9_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_9_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_9_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_9_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_9_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_9_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_9_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_9_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_9_0_i_AWID,
      AWADDR => x_rsc_9_0_i_AWADDR,
      AWLEN => x_rsc_9_0_i_AWLEN,
      AWSIZE => x_rsc_9_0_i_AWSIZE,
      AWBURST => x_rsc_9_0_i_AWBURST,
      AWLOCK => x_rsc_9_0_AWLOCK,
      AWCACHE => x_rsc_9_0_i_AWCACHE,
      AWPROT => x_rsc_9_0_i_AWPROT,
      AWQOS => x_rsc_9_0_i_AWQOS,
      AWREGION => x_rsc_9_0_i_AWREGION,
      AWUSER => x_rsc_9_0_i_AWUSER,
      AWVALID => x_rsc_9_0_AWVALID,
      AWREADY => x_rsc_9_0_AWREADY,
      WDATA => x_rsc_9_0_i_WDATA,
      WSTRB => x_rsc_9_0_i_WSTRB,
      WLAST => x_rsc_9_0_WLAST,
      WUSER => x_rsc_9_0_i_WUSER,
      WVALID => x_rsc_9_0_WVALID,
      WREADY => x_rsc_9_0_WREADY,
      BID => x_rsc_9_0_i_BID,
      BRESP => x_rsc_9_0_i_BRESP,
      BUSER => x_rsc_9_0_i_BUSER,
      BVALID => x_rsc_9_0_BVALID,
      BREADY => x_rsc_9_0_BREADY,
      ARID => x_rsc_9_0_i_ARID,
      ARADDR => x_rsc_9_0_i_ARADDR,
      ARLEN => x_rsc_9_0_i_ARLEN,
      ARSIZE => x_rsc_9_0_i_ARSIZE,
      ARBURST => x_rsc_9_0_i_ARBURST,
      ARLOCK => x_rsc_9_0_ARLOCK,
      ARCACHE => x_rsc_9_0_i_ARCACHE,
      ARPROT => x_rsc_9_0_i_ARPROT,
      ARQOS => x_rsc_9_0_i_ARQOS,
      ARREGION => x_rsc_9_0_i_ARREGION,
      ARUSER => x_rsc_9_0_i_ARUSER,
      ARVALID => x_rsc_9_0_ARVALID,
      ARREADY => x_rsc_9_0_ARREADY,
      RID => x_rsc_9_0_i_RID,
      RDATA => x_rsc_9_0_i_RDATA,
      RRESP => x_rsc_9_0_i_RRESP,
      RLAST => x_rsc_9_0_RLAST,
      RUSER => x_rsc_9_0_i_RUSER,
      RVALID => x_rsc_9_0_RVALID,
      RREADY => x_rsc_9_0_RREADY,
      s_re => x_rsc_9_0_i_s_re_core_sct,
      s_we => x_rsc_9_0_i_s_we_core_sct,
      s_raddr => x_rsc_9_0_i_s_raddr_1,
      s_waddr => x_rsc_9_0_i_s_waddr_1,
      s_din => x_rsc_9_0_i_s_din_1,
      s_dout => x_rsc_9_0_i_s_dout_1,
      s_rrdy => x_rsc_9_0_i_s_rrdy,
      s_wrdy => x_rsc_9_0_i_s_wrdy,
      is_idle => x_rsc_9_0_is_idle_1,
      tr_write_done => x_rsc_9_0_tr_write_done,
      s_tdone => x_rsc_9_0_s_tdone
    );
  x_rsc_9_0_i_AWID(0) <= x_rsc_9_0_AWID;
  x_rsc_9_0_i_AWADDR <= x_rsc_9_0_AWADDR;
  x_rsc_9_0_i_AWLEN <= x_rsc_9_0_AWLEN;
  x_rsc_9_0_i_AWSIZE <= x_rsc_9_0_AWSIZE;
  x_rsc_9_0_i_AWBURST <= x_rsc_9_0_AWBURST;
  x_rsc_9_0_i_AWCACHE <= x_rsc_9_0_AWCACHE;
  x_rsc_9_0_i_AWPROT <= x_rsc_9_0_AWPROT;
  x_rsc_9_0_i_AWQOS <= x_rsc_9_0_AWQOS;
  x_rsc_9_0_i_AWREGION <= x_rsc_9_0_AWREGION;
  x_rsc_9_0_i_AWUSER(0) <= x_rsc_9_0_AWUSER;
  x_rsc_9_0_i_WDATA <= x_rsc_9_0_WDATA;
  x_rsc_9_0_i_WSTRB <= x_rsc_9_0_WSTRB;
  x_rsc_9_0_i_WUSER(0) <= x_rsc_9_0_WUSER;
  x_rsc_9_0_BID <= x_rsc_9_0_i_BID(0);
  x_rsc_9_0_BRESP <= x_rsc_9_0_i_BRESP;
  x_rsc_9_0_BUSER <= x_rsc_9_0_i_BUSER(0);
  x_rsc_9_0_i_ARID(0) <= x_rsc_9_0_ARID;
  x_rsc_9_0_i_ARADDR <= x_rsc_9_0_ARADDR;
  x_rsc_9_0_i_ARLEN <= x_rsc_9_0_ARLEN;
  x_rsc_9_0_i_ARSIZE <= x_rsc_9_0_ARSIZE;
  x_rsc_9_0_i_ARBURST <= x_rsc_9_0_ARBURST;
  x_rsc_9_0_i_ARCACHE <= x_rsc_9_0_ARCACHE;
  x_rsc_9_0_i_ARPROT <= x_rsc_9_0_ARPROT;
  x_rsc_9_0_i_ARQOS <= x_rsc_9_0_ARQOS;
  x_rsc_9_0_i_ARREGION <= x_rsc_9_0_ARREGION;
  x_rsc_9_0_i_ARUSER(0) <= x_rsc_9_0_ARUSER;
  x_rsc_9_0_RID <= x_rsc_9_0_i_RID(0);
  x_rsc_9_0_RDATA <= x_rsc_9_0_i_RDATA;
  x_rsc_9_0_RRESP <= x_rsc_9_0_i_RRESP;
  x_rsc_9_0_RUSER <= x_rsc_9_0_i_RUSER(0);
  x_rsc_9_0_i_s_raddr_1 <= x_rsc_9_0_i_s_raddr;
  x_rsc_9_0_i_s_waddr_1 <= x_rsc_9_0_i_s_waddr;
  x_rsc_9_0_i_s_din <= x_rsc_9_0_i_s_din_1;
  x_rsc_9_0_i_s_dout_1 <= x_rsc_9_0_i_s_dout;

  hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl_inst : hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_9_0_i_oswt => x_rsc_9_0_i_oswt,
      x_rsc_9_0_i_oswt_1 => x_rsc_9_0_i_oswt_1,
      x_rsc_9_0_i_biwt => x_rsc_9_0_i_biwt,
      x_rsc_9_0_i_bdwt => x_rsc_9_0_i_bdwt,
      x_rsc_9_0_i_bcwt => x_rsc_9_0_i_bcwt,
      x_rsc_9_0_i_s_re_core_sct => x_rsc_9_0_i_s_re_core_sct,
      x_rsc_9_0_i_biwt_1 => x_rsc_9_0_i_biwt_1,
      x_rsc_9_0_i_bdwt_2 => x_rsc_9_0_i_bdwt_2,
      x_rsc_9_0_i_bcwt_1 => x_rsc_9_0_i_bcwt_1,
      x_rsc_9_0_i_s_we_core_sct => x_rsc_9_0_i_s_we_core_sct,
      x_rsc_9_0_i_s_rrdy => x_rsc_9_0_i_s_rrdy,
      x_rsc_9_0_i_s_wrdy => x_rsc_9_0_i_s_wrdy
    );
  hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst : hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_9_0_i_oswt => x_rsc_9_0_i_oswt,
      x_rsc_9_0_i_wen_comp => x_rsc_9_0_i_wen_comp,
      x_rsc_9_0_i_oswt_1 => x_rsc_9_0_i_oswt_1,
      x_rsc_9_0_i_wen_comp_1 => x_rsc_9_0_i_wen_comp_1,
      x_rsc_9_0_i_s_raddr_core => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_raddr_core,
      x_rsc_9_0_i_s_waddr_core => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_waddr_core,
      x_rsc_9_0_i_s_din_mxwt => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_din_mxwt,
      x_rsc_9_0_i_s_dout_core => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_dout_core,
      x_rsc_9_0_i_biwt => x_rsc_9_0_i_biwt,
      x_rsc_9_0_i_bdwt => x_rsc_9_0_i_bdwt,
      x_rsc_9_0_i_bcwt => x_rsc_9_0_i_bcwt,
      x_rsc_9_0_i_biwt_1 => x_rsc_9_0_i_biwt_1,
      x_rsc_9_0_i_bdwt_2 => x_rsc_9_0_i_bdwt_2,
      x_rsc_9_0_i_bcwt_1 => x_rsc_9_0_i_bcwt_1,
      x_rsc_9_0_i_s_raddr => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_raddr,
      x_rsc_9_0_i_s_raddr_core_sct => x_rsc_9_0_i_s_re_core_sct,
      x_rsc_9_0_i_s_waddr => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_waddr,
      x_rsc_9_0_i_s_waddr_core_sct => x_rsc_9_0_i_s_we_core_sct,
      x_rsc_9_0_i_s_din => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_din,
      x_rsc_9_0_i_s_dout => hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_dout
    );
  hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_raddr_core <= x_rsc_9_0_i_s_raddr_core;
  hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_waddr_core <= x_rsc_9_0_i_s_waddr_core;
  x_rsc_9_0_i_s_din_mxwt <= hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_din_mxwt;
  hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_dout_core <= x_rsc_9_0_i_s_dout_core;
  x_rsc_9_0_i_s_raddr <= hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_raddr;
  x_rsc_9_0_i_s_waddr <= hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_waddr;
  hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_din <= x_rsc_9_0_i_s_din;
  x_rsc_9_0_i_s_dout <= hybrid_core_x_rsc_9_0_i_x_rsc_9_0_wait_dp_inst_x_rsc_9_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_8_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_8_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_8_0_s_tdone : IN STD_LOGIC;
    x_rsc_8_0_tr_write_done : IN STD_LOGIC;
    x_rsc_8_0_RREADY : IN STD_LOGIC;
    x_rsc_8_0_RVALID : OUT STD_LOGIC;
    x_rsc_8_0_RUSER : OUT STD_LOGIC;
    x_rsc_8_0_RLAST : OUT STD_LOGIC;
    x_rsc_8_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_RID : OUT STD_LOGIC;
    x_rsc_8_0_ARREADY : OUT STD_LOGIC;
    x_rsc_8_0_ARVALID : IN STD_LOGIC;
    x_rsc_8_0_ARUSER : IN STD_LOGIC;
    x_rsc_8_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARLOCK : IN STD_LOGIC;
    x_rsc_8_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_8_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_8_0_ARID : IN STD_LOGIC;
    x_rsc_8_0_BREADY : IN STD_LOGIC;
    x_rsc_8_0_BVALID : OUT STD_LOGIC;
    x_rsc_8_0_BUSER : OUT STD_LOGIC;
    x_rsc_8_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_BID : OUT STD_LOGIC;
    x_rsc_8_0_WREADY : OUT STD_LOGIC;
    x_rsc_8_0_WVALID : IN STD_LOGIC;
    x_rsc_8_0_WUSER : IN STD_LOGIC;
    x_rsc_8_0_WLAST : IN STD_LOGIC;
    x_rsc_8_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_AWREADY : OUT STD_LOGIC;
    x_rsc_8_0_AWVALID : IN STD_LOGIC;
    x_rsc_8_0_AWUSER : IN STD_LOGIC;
    x_rsc_8_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWLOCK : IN STD_LOGIC;
    x_rsc_8_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_8_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_8_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_8_0_i_oswt : IN STD_LOGIC;
    x_rsc_8_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_8_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_8_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_8_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_8_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_8_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_8_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_8_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_8_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_8_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_8_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_8_0_i_oswt : IN STD_LOGIC;
      x_rsc_8_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_8_0_i_biwt : OUT STD_LOGIC;
      x_rsc_8_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_8_0_i_bcwt : IN STD_LOGIC;
      x_rsc_8_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_8_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_8_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_8_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_8_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_8_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_8_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_8_0_i_oswt : IN STD_LOGIC;
      x_rsc_8_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_8_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_8_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_8_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_8_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_8_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_i_biwt : IN STD_LOGIC;
      x_rsc_8_0_i_bdwt : IN STD_LOGIC;
      x_rsc_8_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_8_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_8_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_8_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_8_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_8_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_8_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_8_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_8_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_8_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_8_0_i_AWID,
      AWADDR => x_rsc_8_0_i_AWADDR,
      AWLEN => x_rsc_8_0_i_AWLEN,
      AWSIZE => x_rsc_8_0_i_AWSIZE,
      AWBURST => x_rsc_8_0_i_AWBURST,
      AWLOCK => x_rsc_8_0_AWLOCK,
      AWCACHE => x_rsc_8_0_i_AWCACHE,
      AWPROT => x_rsc_8_0_i_AWPROT,
      AWQOS => x_rsc_8_0_i_AWQOS,
      AWREGION => x_rsc_8_0_i_AWREGION,
      AWUSER => x_rsc_8_0_i_AWUSER,
      AWVALID => x_rsc_8_0_AWVALID,
      AWREADY => x_rsc_8_0_AWREADY,
      WDATA => x_rsc_8_0_i_WDATA,
      WSTRB => x_rsc_8_0_i_WSTRB,
      WLAST => x_rsc_8_0_WLAST,
      WUSER => x_rsc_8_0_i_WUSER,
      WVALID => x_rsc_8_0_WVALID,
      WREADY => x_rsc_8_0_WREADY,
      BID => x_rsc_8_0_i_BID,
      BRESP => x_rsc_8_0_i_BRESP,
      BUSER => x_rsc_8_0_i_BUSER,
      BVALID => x_rsc_8_0_BVALID,
      BREADY => x_rsc_8_0_BREADY,
      ARID => x_rsc_8_0_i_ARID,
      ARADDR => x_rsc_8_0_i_ARADDR,
      ARLEN => x_rsc_8_0_i_ARLEN,
      ARSIZE => x_rsc_8_0_i_ARSIZE,
      ARBURST => x_rsc_8_0_i_ARBURST,
      ARLOCK => x_rsc_8_0_ARLOCK,
      ARCACHE => x_rsc_8_0_i_ARCACHE,
      ARPROT => x_rsc_8_0_i_ARPROT,
      ARQOS => x_rsc_8_0_i_ARQOS,
      ARREGION => x_rsc_8_0_i_ARREGION,
      ARUSER => x_rsc_8_0_i_ARUSER,
      ARVALID => x_rsc_8_0_ARVALID,
      ARREADY => x_rsc_8_0_ARREADY,
      RID => x_rsc_8_0_i_RID,
      RDATA => x_rsc_8_0_i_RDATA,
      RRESP => x_rsc_8_0_i_RRESP,
      RLAST => x_rsc_8_0_RLAST,
      RUSER => x_rsc_8_0_i_RUSER,
      RVALID => x_rsc_8_0_RVALID,
      RREADY => x_rsc_8_0_RREADY,
      s_re => x_rsc_8_0_i_s_re_core_sct,
      s_we => x_rsc_8_0_i_s_we_core_sct,
      s_raddr => x_rsc_8_0_i_s_raddr_1,
      s_waddr => x_rsc_8_0_i_s_waddr_1,
      s_din => x_rsc_8_0_i_s_din_1,
      s_dout => x_rsc_8_0_i_s_dout_1,
      s_rrdy => x_rsc_8_0_i_s_rrdy,
      s_wrdy => x_rsc_8_0_i_s_wrdy,
      is_idle => x_rsc_8_0_is_idle_1,
      tr_write_done => x_rsc_8_0_tr_write_done,
      s_tdone => x_rsc_8_0_s_tdone
    );
  x_rsc_8_0_i_AWID(0) <= x_rsc_8_0_AWID;
  x_rsc_8_0_i_AWADDR <= x_rsc_8_0_AWADDR;
  x_rsc_8_0_i_AWLEN <= x_rsc_8_0_AWLEN;
  x_rsc_8_0_i_AWSIZE <= x_rsc_8_0_AWSIZE;
  x_rsc_8_0_i_AWBURST <= x_rsc_8_0_AWBURST;
  x_rsc_8_0_i_AWCACHE <= x_rsc_8_0_AWCACHE;
  x_rsc_8_0_i_AWPROT <= x_rsc_8_0_AWPROT;
  x_rsc_8_0_i_AWQOS <= x_rsc_8_0_AWQOS;
  x_rsc_8_0_i_AWREGION <= x_rsc_8_0_AWREGION;
  x_rsc_8_0_i_AWUSER(0) <= x_rsc_8_0_AWUSER;
  x_rsc_8_0_i_WDATA <= x_rsc_8_0_WDATA;
  x_rsc_8_0_i_WSTRB <= x_rsc_8_0_WSTRB;
  x_rsc_8_0_i_WUSER(0) <= x_rsc_8_0_WUSER;
  x_rsc_8_0_BID <= x_rsc_8_0_i_BID(0);
  x_rsc_8_0_BRESP <= x_rsc_8_0_i_BRESP;
  x_rsc_8_0_BUSER <= x_rsc_8_0_i_BUSER(0);
  x_rsc_8_0_i_ARID(0) <= x_rsc_8_0_ARID;
  x_rsc_8_0_i_ARADDR <= x_rsc_8_0_ARADDR;
  x_rsc_8_0_i_ARLEN <= x_rsc_8_0_ARLEN;
  x_rsc_8_0_i_ARSIZE <= x_rsc_8_0_ARSIZE;
  x_rsc_8_0_i_ARBURST <= x_rsc_8_0_ARBURST;
  x_rsc_8_0_i_ARCACHE <= x_rsc_8_0_ARCACHE;
  x_rsc_8_0_i_ARPROT <= x_rsc_8_0_ARPROT;
  x_rsc_8_0_i_ARQOS <= x_rsc_8_0_ARQOS;
  x_rsc_8_0_i_ARREGION <= x_rsc_8_0_ARREGION;
  x_rsc_8_0_i_ARUSER(0) <= x_rsc_8_0_ARUSER;
  x_rsc_8_0_RID <= x_rsc_8_0_i_RID(0);
  x_rsc_8_0_RDATA <= x_rsc_8_0_i_RDATA;
  x_rsc_8_0_RRESP <= x_rsc_8_0_i_RRESP;
  x_rsc_8_0_RUSER <= x_rsc_8_0_i_RUSER(0);
  x_rsc_8_0_i_s_raddr_1 <= x_rsc_8_0_i_s_raddr;
  x_rsc_8_0_i_s_waddr_1 <= x_rsc_8_0_i_s_waddr;
  x_rsc_8_0_i_s_din <= x_rsc_8_0_i_s_din_1;
  x_rsc_8_0_i_s_dout_1 <= x_rsc_8_0_i_s_dout;

  hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl_inst : hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_8_0_i_oswt => x_rsc_8_0_i_oswt,
      x_rsc_8_0_i_oswt_1 => x_rsc_8_0_i_oswt_1,
      x_rsc_8_0_i_biwt => x_rsc_8_0_i_biwt,
      x_rsc_8_0_i_bdwt => x_rsc_8_0_i_bdwt,
      x_rsc_8_0_i_bcwt => x_rsc_8_0_i_bcwt,
      x_rsc_8_0_i_s_re_core_sct => x_rsc_8_0_i_s_re_core_sct,
      x_rsc_8_0_i_biwt_1 => x_rsc_8_0_i_biwt_1,
      x_rsc_8_0_i_bdwt_2 => x_rsc_8_0_i_bdwt_2,
      x_rsc_8_0_i_bcwt_1 => x_rsc_8_0_i_bcwt_1,
      x_rsc_8_0_i_s_we_core_sct => x_rsc_8_0_i_s_we_core_sct,
      x_rsc_8_0_i_s_rrdy => x_rsc_8_0_i_s_rrdy,
      x_rsc_8_0_i_s_wrdy => x_rsc_8_0_i_s_wrdy
    );
  hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst : hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_8_0_i_oswt => x_rsc_8_0_i_oswt,
      x_rsc_8_0_i_wen_comp => x_rsc_8_0_i_wen_comp,
      x_rsc_8_0_i_oswt_1 => x_rsc_8_0_i_oswt_1,
      x_rsc_8_0_i_wen_comp_1 => x_rsc_8_0_i_wen_comp_1,
      x_rsc_8_0_i_s_raddr_core => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_raddr_core,
      x_rsc_8_0_i_s_waddr_core => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_waddr_core,
      x_rsc_8_0_i_s_din_mxwt => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_din_mxwt,
      x_rsc_8_0_i_s_dout_core => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_dout_core,
      x_rsc_8_0_i_biwt => x_rsc_8_0_i_biwt,
      x_rsc_8_0_i_bdwt => x_rsc_8_0_i_bdwt,
      x_rsc_8_0_i_bcwt => x_rsc_8_0_i_bcwt,
      x_rsc_8_0_i_biwt_1 => x_rsc_8_0_i_biwt_1,
      x_rsc_8_0_i_bdwt_2 => x_rsc_8_0_i_bdwt_2,
      x_rsc_8_0_i_bcwt_1 => x_rsc_8_0_i_bcwt_1,
      x_rsc_8_0_i_s_raddr => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_raddr,
      x_rsc_8_0_i_s_raddr_core_sct => x_rsc_8_0_i_s_re_core_sct,
      x_rsc_8_0_i_s_waddr => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_waddr,
      x_rsc_8_0_i_s_waddr_core_sct => x_rsc_8_0_i_s_we_core_sct,
      x_rsc_8_0_i_s_din => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_din,
      x_rsc_8_0_i_s_dout => hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_dout
    );
  hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_raddr_core <= x_rsc_8_0_i_s_raddr_core;
  hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_waddr_core <= x_rsc_8_0_i_s_waddr_core;
  x_rsc_8_0_i_s_din_mxwt <= hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_din_mxwt;
  hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_dout_core <= x_rsc_8_0_i_s_dout_core;
  x_rsc_8_0_i_s_raddr <= hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_raddr;
  x_rsc_8_0_i_s_waddr <= hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_waddr;
  hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_din <= x_rsc_8_0_i_s_din;
  x_rsc_8_0_i_s_dout <= hybrid_core_x_rsc_8_0_i_x_rsc_8_0_wait_dp_inst_x_rsc_8_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_7_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_7_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_7_0_s_tdone : IN STD_LOGIC;
    x_rsc_7_0_tr_write_done : IN STD_LOGIC;
    x_rsc_7_0_RREADY : IN STD_LOGIC;
    x_rsc_7_0_RVALID : OUT STD_LOGIC;
    x_rsc_7_0_RUSER : OUT STD_LOGIC;
    x_rsc_7_0_RLAST : OUT STD_LOGIC;
    x_rsc_7_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_RID : OUT STD_LOGIC;
    x_rsc_7_0_ARREADY : OUT STD_LOGIC;
    x_rsc_7_0_ARVALID : IN STD_LOGIC;
    x_rsc_7_0_ARUSER : IN STD_LOGIC;
    x_rsc_7_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARLOCK : IN STD_LOGIC;
    x_rsc_7_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_7_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_7_0_ARID : IN STD_LOGIC;
    x_rsc_7_0_BREADY : IN STD_LOGIC;
    x_rsc_7_0_BVALID : OUT STD_LOGIC;
    x_rsc_7_0_BUSER : OUT STD_LOGIC;
    x_rsc_7_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_BID : OUT STD_LOGIC;
    x_rsc_7_0_WREADY : OUT STD_LOGIC;
    x_rsc_7_0_WVALID : IN STD_LOGIC;
    x_rsc_7_0_WUSER : IN STD_LOGIC;
    x_rsc_7_0_WLAST : IN STD_LOGIC;
    x_rsc_7_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_AWREADY : OUT STD_LOGIC;
    x_rsc_7_0_AWVALID : IN STD_LOGIC;
    x_rsc_7_0_AWUSER : IN STD_LOGIC;
    x_rsc_7_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWLOCK : IN STD_LOGIC;
    x_rsc_7_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_7_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_7_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_7_0_i_oswt : IN STD_LOGIC;
    x_rsc_7_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_7_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_7_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_7_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_7_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_7_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_7_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_7_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_7_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_7_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_7_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_7_0_i_oswt : IN STD_LOGIC;
      x_rsc_7_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_7_0_i_biwt : OUT STD_LOGIC;
      x_rsc_7_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_7_0_i_bcwt : IN STD_LOGIC;
      x_rsc_7_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_7_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_7_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_7_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_7_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_7_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_7_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_7_0_i_oswt : IN STD_LOGIC;
      x_rsc_7_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_7_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_7_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_7_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_7_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_7_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_i_biwt : IN STD_LOGIC;
      x_rsc_7_0_i_bdwt : IN STD_LOGIC;
      x_rsc_7_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_7_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_7_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_7_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_7_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_7_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_7_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_7_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_7_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_7_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_7_0_i_AWID,
      AWADDR => x_rsc_7_0_i_AWADDR,
      AWLEN => x_rsc_7_0_i_AWLEN,
      AWSIZE => x_rsc_7_0_i_AWSIZE,
      AWBURST => x_rsc_7_0_i_AWBURST,
      AWLOCK => x_rsc_7_0_AWLOCK,
      AWCACHE => x_rsc_7_0_i_AWCACHE,
      AWPROT => x_rsc_7_0_i_AWPROT,
      AWQOS => x_rsc_7_0_i_AWQOS,
      AWREGION => x_rsc_7_0_i_AWREGION,
      AWUSER => x_rsc_7_0_i_AWUSER,
      AWVALID => x_rsc_7_0_AWVALID,
      AWREADY => x_rsc_7_0_AWREADY,
      WDATA => x_rsc_7_0_i_WDATA,
      WSTRB => x_rsc_7_0_i_WSTRB,
      WLAST => x_rsc_7_0_WLAST,
      WUSER => x_rsc_7_0_i_WUSER,
      WVALID => x_rsc_7_0_WVALID,
      WREADY => x_rsc_7_0_WREADY,
      BID => x_rsc_7_0_i_BID,
      BRESP => x_rsc_7_0_i_BRESP,
      BUSER => x_rsc_7_0_i_BUSER,
      BVALID => x_rsc_7_0_BVALID,
      BREADY => x_rsc_7_0_BREADY,
      ARID => x_rsc_7_0_i_ARID,
      ARADDR => x_rsc_7_0_i_ARADDR,
      ARLEN => x_rsc_7_0_i_ARLEN,
      ARSIZE => x_rsc_7_0_i_ARSIZE,
      ARBURST => x_rsc_7_0_i_ARBURST,
      ARLOCK => x_rsc_7_0_ARLOCK,
      ARCACHE => x_rsc_7_0_i_ARCACHE,
      ARPROT => x_rsc_7_0_i_ARPROT,
      ARQOS => x_rsc_7_0_i_ARQOS,
      ARREGION => x_rsc_7_0_i_ARREGION,
      ARUSER => x_rsc_7_0_i_ARUSER,
      ARVALID => x_rsc_7_0_ARVALID,
      ARREADY => x_rsc_7_0_ARREADY,
      RID => x_rsc_7_0_i_RID,
      RDATA => x_rsc_7_0_i_RDATA,
      RRESP => x_rsc_7_0_i_RRESP,
      RLAST => x_rsc_7_0_RLAST,
      RUSER => x_rsc_7_0_i_RUSER,
      RVALID => x_rsc_7_0_RVALID,
      RREADY => x_rsc_7_0_RREADY,
      s_re => x_rsc_7_0_i_s_re_core_sct,
      s_we => x_rsc_7_0_i_s_we_core_sct,
      s_raddr => x_rsc_7_0_i_s_raddr_1,
      s_waddr => x_rsc_7_0_i_s_waddr_1,
      s_din => x_rsc_7_0_i_s_din_1,
      s_dout => x_rsc_7_0_i_s_dout_1,
      s_rrdy => x_rsc_7_0_i_s_rrdy,
      s_wrdy => x_rsc_7_0_i_s_wrdy,
      is_idle => x_rsc_7_0_is_idle_1,
      tr_write_done => x_rsc_7_0_tr_write_done,
      s_tdone => x_rsc_7_0_s_tdone
    );
  x_rsc_7_0_i_AWID(0) <= x_rsc_7_0_AWID;
  x_rsc_7_0_i_AWADDR <= x_rsc_7_0_AWADDR;
  x_rsc_7_0_i_AWLEN <= x_rsc_7_0_AWLEN;
  x_rsc_7_0_i_AWSIZE <= x_rsc_7_0_AWSIZE;
  x_rsc_7_0_i_AWBURST <= x_rsc_7_0_AWBURST;
  x_rsc_7_0_i_AWCACHE <= x_rsc_7_0_AWCACHE;
  x_rsc_7_0_i_AWPROT <= x_rsc_7_0_AWPROT;
  x_rsc_7_0_i_AWQOS <= x_rsc_7_0_AWQOS;
  x_rsc_7_0_i_AWREGION <= x_rsc_7_0_AWREGION;
  x_rsc_7_0_i_AWUSER(0) <= x_rsc_7_0_AWUSER;
  x_rsc_7_0_i_WDATA <= x_rsc_7_0_WDATA;
  x_rsc_7_0_i_WSTRB <= x_rsc_7_0_WSTRB;
  x_rsc_7_0_i_WUSER(0) <= x_rsc_7_0_WUSER;
  x_rsc_7_0_BID <= x_rsc_7_0_i_BID(0);
  x_rsc_7_0_BRESP <= x_rsc_7_0_i_BRESP;
  x_rsc_7_0_BUSER <= x_rsc_7_0_i_BUSER(0);
  x_rsc_7_0_i_ARID(0) <= x_rsc_7_0_ARID;
  x_rsc_7_0_i_ARADDR <= x_rsc_7_0_ARADDR;
  x_rsc_7_0_i_ARLEN <= x_rsc_7_0_ARLEN;
  x_rsc_7_0_i_ARSIZE <= x_rsc_7_0_ARSIZE;
  x_rsc_7_0_i_ARBURST <= x_rsc_7_0_ARBURST;
  x_rsc_7_0_i_ARCACHE <= x_rsc_7_0_ARCACHE;
  x_rsc_7_0_i_ARPROT <= x_rsc_7_0_ARPROT;
  x_rsc_7_0_i_ARQOS <= x_rsc_7_0_ARQOS;
  x_rsc_7_0_i_ARREGION <= x_rsc_7_0_ARREGION;
  x_rsc_7_0_i_ARUSER(0) <= x_rsc_7_0_ARUSER;
  x_rsc_7_0_RID <= x_rsc_7_0_i_RID(0);
  x_rsc_7_0_RDATA <= x_rsc_7_0_i_RDATA;
  x_rsc_7_0_RRESP <= x_rsc_7_0_i_RRESP;
  x_rsc_7_0_RUSER <= x_rsc_7_0_i_RUSER(0);
  x_rsc_7_0_i_s_raddr_1 <= x_rsc_7_0_i_s_raddr;
  x_rsc_7_0_i_s_waddr_1 <= x_rsc_7_0_i_s_waddr;
  x_rsc_7_0_i_s_din <= x_rsc_7_0_i_s_din_1;
  x_rsc_7_0_i_s_dout_1 <= x_rsc_7_0_i_s_dout;

  hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl_inst : hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_7_0_i_oswt => x_rsc_7_0_i_oswt,
      x_rsc_7_0_i_oswt_1 => x_rsc_7_0_i_oswt_1,
      x_rsc_7_0_i_biwt => x_rsc_7_0_i_biwt,
      x_rsc_7_0_i_bdwt => x_rsc_7_0_i_bdwt,
      x_rsc_7_0_i_bcwt => x_rsc_7_0_i_bcwt,
      x_rsc_7_0_i_s_re_core_sct => x_rsc_7_0_i_s_re_core_sct,
      x_rsc_7_0_i_biwt_1 => x_rsc_7_0_i_biwt_1,
      x_rsc_7_0_i_bdwt_2 => x_rsc_7_0_i_bdwt_2,
      x_rsc_7_0_i_bcwt_1 => x_rsc_7_0_i_bcwt_1,
      x_rsc_7_0_i_s_we_core_sct => x_rsc_7_0_i_s_we_core_sct,
      x_rsc_7_0_i_s_rrdy => x_rsc_7_0_i_s_rrdy,
      x_rsc_7_0_i_s_wrdy => x_rsc_7_0_i_s_wrdy
    );
  hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst : hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_7_0_i_oswt => x_rsc_7_0_i_oswt,
      x_rsc_7_0_i_wen_comp => x_rsc_7_0_i_wen_comp,
      x_rsc_7_0_i_oswt_1 => x_rsc_7_0_i_oswt_1,
      x_rsc_7_0_i_wen_comp_1 => x_rsc_7_0_i_wen_comp_1,
      x_rsc_7_0_i_s_raddr_core => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_raddr_core,
      x_rsc_7_0_i_s_waddr_core => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_waddr_core,
      x_rsc_7_0_i_s_din_mxwt => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_din_mxwt,
      x_rsc_7_0_i_s_dout_core => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_dout_core,
      x_rsc_7_0_i_biwt => x_rsc_7_0_i_biwt,
      x_rsc_7_0_i_bdwt => x_rsc_7_0_i_bdwt,
      x_rsc_7_0_i_bcwt => x_rsc_7_0_i_bcwt,
      x_rsc_7_0_i_biwt_1 => x_rsc_7_0_i_biwt_1,
      x_rsc_7_0_i_bdwt_2 => x_rsc_7_0_i_bdwt_2,
      x_rsc_7_0_i_bcwt_1 => x_rsc_7_0_i_bcwt_1,
      x_rsc_7_0_i_s_raddr => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_raddr,
      x_rsc_7_0_i_s_raddr_core_sct => x_rsc_7_0_i_s_re_core_sct,
      x_rsc_7_0_i_s_waddr => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_waddr,
      x_rsc_7_0_i_s_waddr_core_sct => x_rsc_7_0_i_s_we_core_sct,
      x_rsc_7_0_i_s_din => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_din,
      x_rsc_7_0_i_s_dout => hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_dout
    );
  hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_raddr_core <= x_rsc_7_0_i_s_raddr_core;
  hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_waddr_core <= x_rsc_7_0_i_s_waddr_core;
  x_rsc_7_0_i_s_din_mxwt <= hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_din_mxwt;
  hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_dout_core <= x_rsc_7_0_i_s_dout_core;
  x_rsc_7_0_i_s_raddr <= hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_raddr;
  x_rsc_7_0_i_s_waddr <= hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_waddr;
  hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_din <= x_rsc_7_0_i_s_din;
  x_rsc_7_0_i_s_dout <= hybrid_core_x_rsc_7_0_i_x_rsc_7_0_wait_dp_inst_x_rsc_7_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_6_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_6_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_6_0_s_tdone : IN STD_LOGIC;
    x_rsc_6_0_tr_write_done : IN STD_LOGIC;
    x_rsc_6_0_RREADY : IN STD_LOGIC;
    x_rsc_6_0_RVALID : OUT STD_LOGIC;
    x_rsc_6_0_RUSER : OUT STD_LOGIC;
    x_rsc_6_0_RLAST : OUT STD_LOGIC;
    x_rsc_6_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_RID : OUT STD_LOGIC;
    x_rsc_6_0_ARREADY : OUT STD_LOGIC;
    x_rsc_6_0_ARVALID : IN STD_LOGIC;
    x_rsc_6_0_ARUSER : IN STD_LOGIC;
    x_rsc_6_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARLOCK : IN STD_LOGIC;
    x_rsc_6_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_6_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_6_0_ARID : IN STD_LOGIC;
    x_rsc_6_0_BREADY : IN STD_LOGIC;
    x_rsc_6_0_BVALID : OUT STD_LOGIC;
    x_rsc_6_0_BUSER : OUT STD_LOGIC;
    x_rsc_6_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_BID : OUT STD_LOGIC;
    x_rsc_6_0_WREADY : OUT STD_LOGIC;
    x_rsc_6_0_WVALID : IN STD_LOGIC;
    x_rsc_6_0_WUSER : IN STD_LOGIC;
    x_rsc_6_0_WLAST : IN STD_LOGIC;
    x_rsc_6_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_AWREADY : OUT STD_LOGIC;
    x_rsc_6_0_AWVALID : IN STD_LOGIC;
    x_rsc_6_0_AWUSER : IN STD_LOGIC;
    x_rsc_6_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWLOCK : IN STD_LOGIC;
    x_rsc_6_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_6_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_6_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_6_0_i_oswt : IN STD_LOGIC;
    x_rsc_6_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_6_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_6_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_6_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_6_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_6_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_6_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_6_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_6_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_6_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_6_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_6_0_i_oswt : IN STD_LOGIC;
      x_rsc_6_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_6_0_i_biwt : OUT STD_LOGIC;
      x_rsc_6_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_6_0_i_bcwt : IN STD_LOGIC;
      x_rsc_6_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_6_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_6_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_6_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_6_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_6_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_6_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_6_0_i_oswt : IN STD_LOGIC;
      x_rsc_6_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_6_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_6_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_6_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_6_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_6_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_i_biwt : IN STD_LOGIC;
      x_rsc_6_0_i_bdwt : IN STD_LOGIC;
      x_rsc_6_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_6_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_6_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_6_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_6_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_6_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_6_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_6_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_6_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_6_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_6_0_i_AWID,
      AWADDR => x_rsc_6_0_i_AWADDR,
      AWLEN => x_rsc_6_0_i_AWLEN,
      AWSIZE => x_rsc_6_0_i_AWSIZE,
      AWBURST => x_rsc_6_0_i_AWBURST,
      AWLOCK => x_rsc_6_0_AWLOCK,
      AWCACHE => x_rsc_6_0_i_AWCACHE,
      AWPROT => x_rsc_6_0_i_AWPROT,
      AWQOS => x_rsc_6_0_i_AWQOS,
      AWREGION => x_rsc_6_0_i_AWREGION,
      AWUSER => x_rsc_6_0_i_AWUSER,
      AWVALID => x_rsc_6_0_AWVALID,
      AWREADY => x_rsc_6_0_AWREADY,
      WDATA => x_rsc_6_0_i_WDATA,
      WSTRB => x_rsc_6_0_i_WSTRB,
      WLAST => x_rsc_6_0_WLAST,
      WUSER => x_rsc_6_0_i_WUSER,
      WVALID => x_rsc_6_0_WVALID,
      WREADY => x_rsc_6_0_WREADY,
      BID => x_rsc_6_0_i_BID,
      BRESP => x_rsc_6_0_i_BRESP,
      BUSER => x_rsc_6_0_i_BUSER,
      BVALID => x_rsc_6_0_BVALID,
      BREADY => x_rsc_6_0_BREADY,
      ARID => x_rsc_6_0_i_ARID,
      ARADDR => x_rsc_6_0_i_ARADDR,
      ARLEN => x_rsc_6_0_i_ARLEN,
      ARSIZE => x_rsc_6_0_i_ARSIZE,
      ARBURST => x_rsc_6_0_i_ARBURST,
      ARLOCK => x_rsc_6_0_ARLOCK,
      ARCACHE => x_rsc_6_0_i_ARCACHE,
      ARPROT => x_rsc_6_0_i_ARPROT,
      ARQOS => x_rsc_6_0_i_ARQOS,
      ARREGION => x_rsc_6_0_i_ARREGION,
      ARUSER => x_rsc_6_0_i_ARUSER,
      ARVALID => x_rsc_6_0_ARVALID,
      ARREADY => x_rsc_6_0_ARREADY,
      RID => x_rsc_6_0_i_RID,
      RDATA => x_rsc_6_0_i_RDATA,
      RRESP => x_rsc_6_0_i_RRESP,
      RLAST => x_rsc_6_0_RLAST,
      RUSER => x_rsc_6_0_i_RUSER,
      RVALID => x_rsc_6_0_RVALID,
      RREADY => x_rsc_6_0_RREADY,
      s_re => x_rsc_6_0_i_s_re_core_sct,
      s_we => x_rsc_6_0_i_s_we_core_sct,
      s_raddr => x_rsc_6_0_i_s_raddr_1,
      s_waddr => x_rsc_6_0_i_s_waddr_1,
      s_din => x_rsc_6_0_i_s_din_1,
      s_dout => x_rsc_6_0_i_s_dout_1,
      s_rrdy => x_rsc_6_0_i_s_rrdy,
      s_wrdy => x_rsc_6_0_i_s_wrdy,
      is_idle => x_rsc_6_0_is_idle_1,
      tr_write_done => x_rsc_6_0_tr_write_done,
      s_tdone => x_rsc_6_0_s_tdone
    );
  x_rsc_6_0_i_AWID(0) <= x_rsc_6_0_AWID;
  x_rsc_6_0_i_AWADDR <= x_rsc_6_0_AWADDR;
  x_rsc_6_0_i_AWLEN <= x_rsc_6_0_AWLEN;
  x_rsc_6_0_i_AWSIZE <= x_rsc_6_0_AWSIZE;
  x_rsc_6_0_i_AWBURST <= x_rsc_6_0_AWBURST;
  x_rsc_6_0_i_AWCACHE <= x_rsc_6_0_AWCACHE;
  x_rsc_6_0_i_AWPROT <= x_rsc_6_0_AWPROT;
  x_rsc_6_0_i_AWQOS <= x_rsc_6_0_AWQOS;
  x_rsc_6_0_i_AWREGION <= x_rsc_6_0_AWREGION;
  x_rsc_6_0_i_AWUSER(0) <= x_rsc_6_0_AWUSER;
  x_rsc_6_0_i_WDATA <= x_rsc_6_0_WDATA;
  x_rsc_6_0_i_WSTRB <= x_rsc_6_0_WSTRB;
  x_rsc_6_0_i_WUSER(0) <= x_rsc_6_0_WUSER;
  x_rsc_6_0_BID <= x_rsc_6_0_i_BID(0);
  x_rsc_6_0_BRESP <= x_rsc_6_0_i_BRESP;
  x_rsc_6_0_BUSER <= x_rsc_6_0_i_BUSER(0);
  x_rsc_6_0_i_ARID(0) <= x_rsc_6_0_ARID;
  x_rsc_6_0_i_ARADDR <= x_rsc_6_0_ARADDR;
  x_rsc_6_0_i_ARLEN <= x_rsc_6_0_ARLEN;
  x_rsc_6_0_i_ARSIZE <= x_rsc_6_0_ARSIZE;
  x_rsc_6_0_i_ARBURST <= x_rsc_6_0_ARBURST;
  x_rsc_6_0_i_ARCACHE <= x_rsc_6_0_ARCACHE;
  x_rsc_6_0_i_ARPROT <= x_rsc_6_0_ARPROT;
  x_rsc_6_0_i_ARQOS <= x_rsc_6_0_ARQOS;
  x_rsc_6_0_i_ARREGION <= x_rsc_6_0_ARREGION;
  x_rsc_6_0_i_ARUSER(0) <= x_rsc_6_0_ARUSER;
  x_rsc_6_0_RID <= x_rsc_6_0_i_RID(0);
  x_rsc_6_0_RDATA <= x_rsc_6_0_i_RDATA;
  x_rsc_6_0_RRESP <= x_rsc_6_0_i_RRESP;
  x_rsc_6_0_RUSER <= x_rsc_6_0_i_RUSER(0);
  x_rsc_6_0_i_s_raddr_1 <= x_rsc_6_0_i_s_raddr;
  x_rsc_6_0_i_s_waddr_1 <= x_rsc_6_0_i_s_waddr;
  x_rsc_6_0_i_s_din <= x_rsc_6_0_i_s_din_1;
  x_rsc_6_0_i_s_dout_1 <= x_rsc_6_0_i_s_dout;

  hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl_inst : hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_6_0_i_oswt => x_rsc_6_0_i_oswt,
      x_rsc_6_0_i_oswt_1 => x_rsc_6_0_i_oswt_1,
      x_rsc_6_0_i_biwt => x_rsc_6_0_i_biwt,
      x_rsc_6_0_i_bdwt => x_rsc_6_0_i_bdwt,
      x_rsc_6_0_i_bcwt => x_rsc_6_0_i_bcwt,
      x_rsc_6_0_i_s_re_core_sct => x_rsc_6_0_i_s_re_core_sct,
      x_rsc_6_0_i_biwt_1 => x_rsc_6_0_i_biwt_1,
      x_rsc_6_0_i_bdwt_2 => x_rsc_6_0_i_bdwt_2,
      x_rsc_6_0_i_bcwt_1 => x_rsc_6_0_i_bcwt_1,
      x_rsc_6_0_i_s_we_core_sct => x_rsc_6_0_i_s_we_core_sct,
      x_rsc_6_0_i_s_rrdy => x_rsc_6_0_i_s_rrdy,
      x_rsc_6_0_i_s_wrdy => x_rsc_6_0_i_s_wrdy
    );
  hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst : hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_6_0_i_oswt => x_rsc_6_0_i_oswt,
      x_rsc_6_0_i_wen_comp => x_rsc_6_0_i_wen_comp,
      x_rsc_6_0_i_oswt_1 => x_rsc_6_0_i_oswt_1,
      x_rsc_6_0_i_wen_comp_1 => x_rsc_6_0_i_wen_comp_1,
      x_rsc_6_0_i_s_raddr_core => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_raddr_core,
      x_rsc_6_0_i_s_waddr_core => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_waddr_core,
      x_rsc_6_0_i_s_din_mxwt => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_din_mxwt,
      x_rsc_6_0_i_s_dout_core => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_dout_core,
      x_rsc_6_0_i_biwt => x_rsc_6_0_i_biwt,
      x_rsc_6_0_i_bdwt => x_rsc_6_0_i_bdwt,
      x_rsc_6_0_i_bcwt => x_rsc_6_0_i_bcwt,
      x_rsc_6_0_i_biwt_1 => x_rsc_6_0_i_biwt_1,
      x_rsc_6_0_i_bdwt_2 => x_rsc_6_0_i_bdwt_2,
      x_rsc_6_0_i_bcwt_1 => x_rsc_6_0_i_bcwt_1,
      x_rsc_6_0_i_s_raddr => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_raddr,
      x_rsc_6_0_i_s_raddr_core_sct => x_rsc_6_0_i_s_re_core_sct,
      x_rsc_6_0_i_s_waddr => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_waddr,
      x_rsc_6_0_i_s_waddr_core_sct => x_rsc_6_0_i_s_we_core_sct,
      x_rsc_6_0_i_s_din => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_din,
      x_rsc_6_0_i_s_dout => hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_dout
    );
  hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_raddr_core <= x_rsc_6_0_i_s_raddr_core;
  hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_waddr_core <= x_rsc_6_0_i_s_waddr_core;
  x_rsc_6_0_i_s_din_mxwt <= hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_din_mxwt;
  hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_dout_core <= x_rsc_6_0_i_s_dout_core;
  x_rsc_6_0_i_s_raddr <= hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_raddr;
  x_rsc_6_0_i_s_waddr <= hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_waddr;
  hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_din <= x_rsc_6_0_i_s_din;
  x_rsc_6_0_i_s_dout <= hybrid_core_x_rsc_6_0_i_x_rsc_6_0_wait_dp_inst_x_rsc_6_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_5_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_5_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_5_0_s_tdone : IN STD_LOGIC;
    x_rsc_5_0_tr_write_done : IN STD_LOGIC;
    x_rsc_5_0_RREADY : IN STD_LOGIC;
    x_rsc_5_0_RVALID : OUT STD_LOGIC;
    x_rsc_5_0_RUSER : OUT STD_LOGIC;
    x_rsc_5_0_RLAST : OUT STD_LOGIC;
    x_rsc_5_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_RID : OUT STD_LOGIC;
    x_rsc_5_0_ARREADY : OUT STD_LOGIC;
    x_rsc_5_0_ARVALID : IN STD_LOGIC;
    x_rsc_5_0_ARUSER : IN STD_LOGIC;
    x_rsc_5_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARLOCK : IN STD_LOGIC;
    x_rsc_5_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_5_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_5_0_ARID : IN STD_LOGIC;
    x_rsc_5_0_BREADY : IN STD_LOGIC;
    x_rsc_5_0_BVALID : OUT STD_LOGIC;
    x_rsc_5_0_BUSER : OUT STD_LOGIC;
    x_rsc_5_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_BID : OUT STD_LOGIC;
    x_rsc_5_0_WREADY : OUT STD_LOGIC;
    x_rsc_5_0_WVALID : IN STD_LOGIC;
    x_rsc_5_0_WUSER : IN STD_LOGIC;
    x_rsc_5_0_WLAST : IN STD_LOGIC;
    x_rsc_5_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_AWREADY : OUT STD_LOGIC;
    x_rsc_5_0_AWVALID : IN STD_LOGIC;
    x_rsc_5_0_AWUSER : IN STD_LOGIC;
    x_rsc_5_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWLOCK : IN STD_LOGIC;
    x_rsc_5_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_5_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_5_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_5_0_i_oswt : IN STD_LOGIC;
    x_rsc_5_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_5_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_5_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_5_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_5_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_5_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_5_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_5_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_5_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_5_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_5_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_5_0_i_oswt : IN STD_LOGIC;
      x_rsc_5_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_5_0_i_biwt : OUT STD_LOGIC;
      x_rsc_5_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_5_0_i_bcwt : IN STD_LOGIC;
      x_rsc_5_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_5_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_5_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_5_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_5_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_5_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_5_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_5_0_i_oswt : IN STD_LOGIC;
      x_rsc_5_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_5_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_5_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_5_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_5_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_5_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_i_biwt : IN STD_LOGIC;
      x_rsc_5_0_i_bdwt : IN STD_LOGIC;
      x_rsc_5_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_5_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_5_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_5_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_5_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_5_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_5_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_5_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_5_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_5_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_5_0_i_AWID,
      AWADDR => x_rsc_5_0_i_AWADDR,
      AWLEN => x_rsc_5_0_i_AWLEN,
      AWSIZE => x_rsc_5_0_i_AWSIZE,
      AWBURST => x_rsc_5_0_i_AWBURST,
      AWLOCK => x_rsc_5_0_AWLOCK,
      AWCACHE => x_rsc_5_0_i_AWCACHE,
      AWPROT => x_rsc_5_0_i_AWPROT,
      AWQOS => x_rsc_5_0_i_AWQOS,
      AWREGION => x_rsc_5_0_i_AWREGION,
      AWUSER => x_rsc_5_0_i_AWUSER,
      AWVALID => x_rsc_5_0_AWVALID,
      AWREADY => x_rsc_5_0_AWREADY,
      WDATA => x_rsc_5_0_i_WDATA,
      WSTRB => x_rsc_5_0_i_WSTRB,
      WLAST => x_rsc_5_0_WLAST,
      WUSER => x_rsc_5_0_i_WUSER,
      WVALID => x_rsc_5_0_WVALID,
      WREADY => x_rsc_5_0_WREADY,
      BID => x_rsc_5_0_i_BID,
      BRESP => x_rsc_5_0_i_BRESP,
      BUSER => x_rsc_5_0_i_BUSER,
      BVALID => x_rsc_5_0_BVALID,
      BREADY => x_rsc_5_0_BREADY,
      ARID => x_rsc_5_0_i_ARID,
      ARADDR => x_rsc_5_0_i_ARADDR,
      ARLEN => x_rsc_5_0_i_ARLEN,
      ARSIZE => x_rsc_5_0_i_ARSIZE,
      ARBURST => x_rsc_5_0_i_ARBURST,
      ARLOCK => x_rsc_5_0_ARLOCK,
      ARCACHE => x_rsc_5_0_i_ARCACHE,
      ARPROT => x_rsc_5_0_i_ARPROT,
      ARQOS => x_rsc_5_0_i_ARQOS,
      ARREGION => x_rsc_5_0_i_ARREGION,
      ARUSER => x_rsc_5_0_i_ARUSER,
      ARVALID => x_rsc_5_0_ARVALID,
      ARREADY => x_rsc_5_0_ARREADY,
      RID => x_rsc_5_0_i_RID,
      RDATA => x_rsc_5_0_i_RDATA,
      RRESP => x_rsc_5_0_i_RRESP,
      RLAST => x_rsc_5_0_RLAST,
      RUSER => x_rsc_5_0_i_RUSER,
      RVALID => x_rsc_5_0_RVALID,
      RREADY => x_rsc_5_0_RREADY,
      s_re => x_rsc_5_0_i_s_re_core_sct,
      s_we => x_rsc_5_0_i_s_we_core_sct,
      s_raddr => x_rsc_5_0_i_s_raddr_1,
      s_waddr => x_rsc_5_0_i_s_waddr_1,
      s_din => x_rsc_5_0_i_s_din_1,
      s_dout => x_rsc_5_0_i_s_dout_1,
      s_rrdy => x_rsc_5_0_i_s_rrdy,
      s_wrdy => x_rsc_5_0_i_s_wrdy,
      is_idle => x_rsc_5_0_is_idle_1,
      tr_write_done => x_rsc_5_0_tr_write_done,
      s_tdone => x_rsc_5_0_s_tdone
    );
  x_rsc_5_0_i_AWID(0) <= x_rsc_5_0_AWID;
  x_rsc_5_0_i_AWADDR <= x_rsc_5_0_AWADDR;
  x_rsc_5_0_i_AWLEN <= x_rsc_5_0_AWLEN;
  x_rsc_5_0_i_AWSIZE <= x_rsc_5_0_AWSIZE;
  x_rsc_5_0_i_AWBURST <= x_rsc_5_0_AWBURST;
  x_rsc_5_0_i_AWCACHE <= x_rsc_5_0_AWCACHE;
  x_rsc_5_0_i_AWPROT <= x_rsc_5_0_AWPROT;
  x_rsc_5_0_i_AWQOS <= x_rsc_5_0_AWQOS;
  x_rsc_5_0_i_AWREGION <= x_rsc_5_0_AWREGION;
  x_rsc_5_0_i_AWUSER(0) <= x_rsc_5_0_AWUSER;
  x_rsc_5_0_i_WDATA <= x_rsc_5_0_WDATA;
  x_rsc_5_0_i_WSTRB <= x_rsc_5_0_WSTRB;
  x_rsc_5_0_i_WUSER(0) <= x_rsc_5_0_WUSER;
  x_rsc_5_0_BID <= x_rsc_5_0_i_BID(0);
  x_rsc_5_0_BRESP <= x_rsc_5_0_i_BRESP;
  x_rsc_5_0_BUSER <= x_rsc_5_0_i_BUSER(0);
  x_rsc_5_0_i_ARID(0) <= x_rsc_5_0_ARID;
  x_rsc_5_0_i_ARADDR <= x_rsc_5_0_ARADDR;
  x_rsc_5_0_i_ARLEN <= x_rsc_5_0_ARLEN;
  x_rsc_5_0_i_ARSIZE <= x_rsc_5_0_ARSIZE;
  x_rsc_5_0_i_ARBURST <= x_rsc_5_0_ARBURST;
  x_rsc_5_0_i_ARCACHE <= x_rsc_5_0_ARCACHE;
  x_rsc_5_0_i_ARPROT <= x_rsc_5_0_ARPROT;
  x_rsc_5_0_i_ARQOS <= x_rsc_5_0_ARQOS;
  x_rsc_5_0_i_ARREGION <= x_rsc_5_0_ARREGION;
  x_rsc_5_0_i_ARUSER(0) <= x_rsc_5_0_ARUSER;
  x_rsc_5_0_RID <= x_rsc_5_0_i_RID(0);
  x_rsc_5_0_RDATA <= x_rsc_5_0_i_RDATA;
  x_rsc_5_0_RRESP <= x_rsc_5_0_i_RRESP;
  x_rsc_5_0_RUSER <= x_rsc_5_0_i_RUSER(0);
  x_rsc_5_0_i_s_raddr_1 <= x_rsc_5_0_i_s_raddr;
  x_rsc_5_0_i_s_waddr_1 <= x_rsc_5_0_i_s_waddr;
  x_rsc_5_0_i_s_din <= x_rsc_5_0_i_s_din_1;
  x_rsc_5_0_i_s_dout_1 <= x_rsc_5_0_i_s_dout;

  hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl_inst : hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_5_0_i_oswt => x_rsc_5_0_i_oswt,
      x_rsc_5_0_i_oswt_1 => x_rsc_5_0_i_oswt_1,
      x_rsc_5_0_i_biwt => x_rsc_5_0_i_biwt,
      x_rsc_5_0_i_bdwt => x_rsc_5_0_i_bdwt,
      x_rsc_5_0_i_bcwt => x_rsc_5_0_i_bcwt,
      x_rsc_5_0_i_s_re_core_sct => x_rsc_5_0_i_s_re_core_sct,
      x_rsc_5_0_i_biwt_1 => x_rsc_5_0_i_biwt_1,
      x_rsc_5_0_i_bdwt_2 => x_rsc_5_0_i_bdwt_2,
      x_rsc_5_0_i_bcwt_1 => x_rsc_5_0_i_bcwt_1,
      x_rsc_5_0_i_s_we_core_sct => x_rsc_5_0_i_s_we_core_sct,
      x_rsc_5_0_i_s_rrdy => x_rsc_5_0_i_s_rrdy,
      x_rsc_5_0_i_s_wrdy => x_rsc_5_0_i_s_wrdy
    );
  hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst : hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_5_0_i_oswt => x_rsc_5_0_i_oswt,
      x_rsc_5_0_i_wen_comp => x_rsc_5_0_i_wen_comp,
      x_rsc_5_0_i_oswt_1 => x_rsc_5_0_i_oswt_1,
      x_rsc_5_0_i_wen_comp_1 => x_rsc_5_0_i_wen_comp_1,
      x_rsc_5_0_i_s_raddr_core => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_raddr_core,
      x_rsc_5_0_i_s_waddr_core => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_waddr_core,
      x_rsc_5_0_i_s_din_mxwt => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_din_mxwt,
      x_rsc_5_0_i_s_dout_core => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_dout_core,
      x_rsc_5_0_i_biwt => x_rsc_5_0_i_biwt,
      x_rsc_5_0_i_bdwt => x_rsc_5_0_i_bdwt,
      x_rsc_5_0_i_bcwt => x_rsc_5_0_i_bcwt,
      x_rsc_5_0_i_biwt_1 => x_rsc_5_0_i_biwt_1,
      x_rsc_5_0_i_bdwt_2 => x_rsc_5_0_i_bdwt_2,
      x_rsc_5_0_i_bcwt_1 => x_rsc_5_0_i_bcwt_1,
      x_rsc_5_0_i_s_raddr => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_raddr,
      x_rsc_5_0_i_s_raddr_core_sct => x_rsc_5_0_i_s_re_core_sct,
      x_rsc_5_0_i_s_waddr => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_waddr,
      x_rsc_5_0_i_s_waddr_core_sct => x_rsc_5_0_i_s_we_core_sct,
      x_rsc_5_0_i_s_din => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_din,
      x_rsc_5_0_i_s_dout => hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_dout
    );
  hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_raddr_core <= x_rsc_5_0_i_s_raddr_core;
  hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_waddr_core <= x_rsc_5_0_i_s_waddr_core;
  x_rsc_5_0_i_s_din_mxwt <= hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_din_mxwt;
  hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_dout_core <= x_rsc_5_0_i_s_dout_core;
  x_rsc_5_0_i_s_raddr <= hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_raddr;
  x_rsc_5_0_i_s_waddr <= hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_waddr;
  hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_din <= x_rsc_5_0_i_s_din;
  x_rsc_5_0_i_s_dout <= hybrid_core_x_rsc_5_0_i_x_rsc_5_0_wait_dp_inst_x_rsc_5_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_4_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_4_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_4_0_s_tdone : IN STD_LOGIC;
    x_rsc_4_0_tr_write_done : IN STD_LOGIC;
    x_rsc_4_0_RREADY : IN STD_LOGIC;
    x_rsc_4_0_RVALID : OUT STD_LOGIC;
    x_rsc_4_0_RUSER : OUT STD_LOGIC;
    x_rsc_4_0_RLAST : OUT STD_LOGIC;
    x_rsc_4_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_RID : OUT STD_LOGIC;
    x_rsc_4_0_ARREADY : OUT STD_LOGIC;
    x_rsc_4_0_ARVALID : IN STD_LOGIC;
    x_rsc_4_0_ARUSER : IN STD_LOGIC;
    x_rsc_4_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARLOCK : IN STD_LOGIC;
    x_rsc_4_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_4_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_4_0_ARID : IN STD_LOGIC;
    x_rsc_4_0_BREADY : IN STD_LOGIC;
    x_rsc_4_0_BVALID : OUT STD_LOGIC;
    x_rsc_4_0_BUSER : OUT STD_LOGIC;
    x_rsc_4_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_BID : OUT STD_LOGIC;
    x_rsc_4_0_WREADY : OUT STD_LOGIC;
    x_rsc_4_0_WVALID : IN STD_LOGIC;
    x_rsc_4_0_WUSER : IN STD_LOGIC;
    x_rsc_4_0_WLAST : IN STD_LOGIC;
    x_rsc_4_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_AWREADY : OUT STD_LOGIC;
    x_rsc_4_0_AWVALID : IN STD_LOGIC;
    x_rsc_4_0_AWUSER : IN STD_LOGIC;
    x_rsc_4_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWLOCK : IN STD_LOGIC;
    x_rsc_4_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_4_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_4_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_4_0_i_oswt : IN STD_LOGIC;
    x_rsc_4_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_4_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_4_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_4_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_4_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_4_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_4_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_4_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_4_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_4_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_4_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_4_0_i_oswt : IN STD_LOGIC;
      x_rsc_4_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_4_0_i_biwt : OUT STD_LOGIC;
      x_rsc_4_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_4_0_i_bcwt : IN STD_LOGIC;
      x_rsc_4_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_4_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_4_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_4_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_4_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_4_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_4_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_4_0_i_oswt : IN STD_LOGIC;
      x_rsc_4_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_4_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_4_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_4_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_4_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_4_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_i_biwt : IN STD_LOGIC;
      x_rsc_4_0_i_bdwt : IN STD_LOGIC;
      x_rsc_4_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_4_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_4_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_4_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_4_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_4_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_4_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_4_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_4_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_4_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_4_0_i_AWID,
      AWADDR => x_rsc_4_0_i_AWADDR,
      AWLEN => x_rsc_4_0_i_AWLEN,
      AWSIZE => x_rsc_4_0_i_AWSIZE,
      AWBURST => x_rsc_4_0_i_AWBURST,
      AWLOCK => x_rsc_4_0_AWLOCK,
      AWCACHE => x_rsc_4_0_i_AWCACHE,
      AWPROT => x_rsc_4_0_i_AWPROT,
      AWQOS => x_rsc_4_0_i_AWQOS,
      AWREGION => x_rsc_4_0_i_AWREGION,
      AWUSER => x_rsc_4_0_i_AWUSER,
      AWVALID => x_rsc_4_0_AWVALID,
      AWREADY => x_rsc_4_0_AWREADY,
      WDATA => x_rsc_4_0_i_WDATA,
      WSTRB => x_rsc_4_0_i_WSTRB,
      WLAST => x_rsc_4_0_WLAST,
      WUSER => x_rsc_4_0_i_WUSER,
      WVALID => x_rsc_4_0_WVALID,
      WREADY => x_rsc_4_0_WREADY,
      BID => x_rsc_4_0_i_BID,
      BRESP => x_rsc_4_0_i_BRESP,
      BUSER => x_rsc_4_0_i_BUSER,
      BVALID => x_rsc_4_0_BVALID,
      BREADY => x_rsc_4_0_BREADY,
      ARID => x_rsc_4_0_i_ARID,
      ARADDR => x_rsc_4_0_i_ARADDR,
      ARLEN => x_rsc_4_0_i_ARLEN,
      ARSIZE => x_rsc_4_0_i_ARSIZE,
      ARBURST => x_rsc_4_0_i_ARBURST,
      ARLOCK => x_rsc_4_0_ARLOCK,
      ARCACHE => x_rsc_4_0_i_ARCACHE,
      ARPROT => x_rsc_4_0_i_ARPROT,
      ARQOS => x_rsc_4_0_i_ARQOS,
      ARREGION => x_rsc_4_0_i_ARREGION,
      ARUSER => x_rsc_4_0_i_ARUSER,
      ARVALID => x_rsc_4_0_ARVALID,
      ARREADY => x_rsc_4_0_ARREADY,
      RID => x_rsc_4_0_i_RID,
      RDATA => x_rsc_4_0_i_RDATA,
      RRESP => x_rsc_4_0_i_RRESP,
      RLAST => x_rsc_4_0_RLAST,
      RUSER => x_rsc_4_0_i_RUSER,
      RVALID => x_rsc_4_0_RVALID,
      RREADY => x_rsc_4_0_RREADY,
      s_re => x_rsc_4_0_i_s_re_core_sct,
      s_we => x_rsc_4_0_i_s_we_core_sct,
      s_raddr => x_rsc_4_0_i_s_raddr_1,
      s_waddr => x_rsc_4_0_i_s_waddr_1,
      s_din => x_rsc_4_0_i_s_din_1,
      s_dout => x_rsc_4_0_i_s_dout_1,
      s_rrdy => x_rsc_4_0_i_s_rrdy,
      s_wrdy => x_rsc_4_0_i_s_wrdy,
      is_idle => x_rsc_4_0_is_idle_1,
      tr_write_done => x_rsc_4_0_tr_write_done,
      s_tdone => x_rsc_4_0_s_tdone
    );
  x_rsc_4_0_i_AWID(0) <= x_rsc_4_0_AWID;
  x_rsc_4_0_i_AWADDR <= x_rsc_4_0_AWADDR;
  x_rsc_4_0_i_AWLEN <= x_rsc_4_0_AWLEN;
  x_rsc_4_0_i_AWSIZE <= x_rsc_4_0_AWSIZE;
  x_rsc_4_0_i_AWBURST <= x_rsc_4_0_AWBURST;
  x_rsc_4_0_i_AWCACHE <= x_rsc_4_0_AWCACHE;
  x_rsc_4_0_i_AWPROT <= x_rsc_4_0_AWPROT;
  x_rsc_4_0_i_AWQOS <= x_rsc_4_0_AWQOS;
  x_rsc_4_0_i_AWREGION <= x_rsc_4_0_AWREGION;
  x_rsc_4_0_i_AWUSER(0) <= x_rsc_4_0_AWUSER;
  x_rsc_4_0_i_WDATA <= x_rsc_4_0_WDATA;
  x_rsc_4_0_i_WSTRB <= x_rsc_4_0_WSTRB;
  x_rsc_4_0_i_WUSER(0) <= x_rsc_4_0_WUSER;
  x_rsc_4_0_BID <= x_rsc_4_0_i_BID(0);
  x_rsc_4_0_BRESP <= x_rsc_4_0_i_BRESP;
  x_rsc_4_0_BUSER <= x_rsc_4_0_i_BUSER(0);
  x_rsc_4_0_i_ARID(0) <= x_rsc_4_0_ARID;
  x_rsc_4_0_i_ARADDR <= x_rsc_4_0_ARADDR;
  x_rsc_4_0_i_ARLEN <= x_rsc_4_0_ARLEN;
  x_rsc_4_0_i_ARSIZE <= x_rsc_4_0_ARSIZE;
  x_rsc_4_0_i_ARBURST <= x_rsc_4_0_ARBURST;
  x_rsc_4_0_i_ARCACHE <= x_rsc_4_0_ARCACHE;
  x_rsc_4_0_i_ARPROT <= x_rsc_4_0_ARPROT;
  x_rsc_4_0_i_ARQOS <= x_rsc_4_0_ARQOS;
  x_rsc_4_0_i_ARREGION <= x_rsc_4_0_ARREGION;
  x_rsc_4_0_i_ARUSER(0) <= x_rsc_4_0_ARUSER;
  x_rsc_4_0_RID <= x_rsc_4_0_i_RID(0);
  x_rsc_4_0_RDATA <= x_rsc_4_0_i_RDATA;
  x_rsc_4_0_RRESP <= x_rsc_4_0_i_RRESP;
  x_rsc_4_0_RUSER <= x_rsc_4_0_i_RUSER(0);
  x_rsc_4_0_i_s_raddr_1 <= x_rsc_4_0_i_s_raddr;
  x_rsc_4_0_i_s_waddr_1 <= x_rsc_4_0_i_s_waddr;
  x_rsc_4_0_i_s_din <= x_rsc_4_0_i_s_din_1;
  x_rsc_4_0_i_s_dout_1 <= x_rsc_4_0_i_s_dout;

  hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl_inst : hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_4_0_i_oswt => x_rsc_4_0_i_oswt,
      x_rsc_4_0_i_oswt_1 => x_rsc_4_0_i_oswt_1,
      x_rsc_4_0_i_biwt => x_rsc_4_0_i_biwt,
      x_rsc_4_0_i_bdwt => x_rsc_4_0_i_bdwt,
      x_rsc_4_0_i_bcwt => x_rsc_4_0_i_bcwt,
      x_rsc_4_0_i_s_re_core_sct => x_rsc_4_0_i_s_re_core_sct,
      x_rsc_4_0_i_biwt_1 => x_rsc_4_0_i_biwt_1,
      x_rsc_4_0_i_bdwt_2 => x_rsc_4_0_i_bdwt_2,
      x_rsc_4_0_i_bcwt_1 => x_rsc_4_0_i_bcwt_1,
      x_rsc_4_0_i_s_we_core_sct => x_rsc_4_0_i_s_we_core_sct,
      x_rsc_4_0_i_s_rrdy => x_rsc_4_0_i_s_rrdy,
      x_rsc_4_0_i_s_wrdy => x_rsc_4_0_i_s_wrdy
    );
  hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst : hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_4_0_i_oswt => x_rsc_4_0_i_oswt,
      x_rsc_4_0_i_wen_comp => x_rsc_4_0_i_wen_comp,
      x_rsc_4_0_i_oswt_1 => x_rsc_4_0_i_oswt_1,
      x_rsc_4_0_i_wen_comp_1 => x_rsc_4_0_i_wen_comp_1,
      x_rsc_4_0_i_s_raddr_core => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_raddr_core,
      x_rsc_4_0_i_s_waddr_core => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_waddr_core,
      x_rsc_4_0_i_s_din_mxwt => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_din_mxwt,
      x_rsc_4_0_i_s_dout_core => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_dout_core,
      x_rsc_4_0_i_biwt => x_rsc_4_0_i_biwt,
      x_rsc_4_0_i_bdwt => x_rsc_4_0_i_bdwt,
      x_rsc_4_0_i_bcwt => x_rsc_4_0_i_bcwt,
      x_rsc_4_0_i_biwt_1 => x_rsc_4_0_i_biwt_1,
      x_rsc_4_0_i_bdwt_2 => x_rsc_4_0_i_bdwt_2,
      x_rsc_4_0_i_bcwt_1 => x_rsc_4_0_i_bcwt_1,
      x_rsc_4_0_i_s_raddr => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_raddr,
      x_rsc_4_0_i_s_raddr_core_sct => x_rsc_4_0_i_s_re_core_sct,
      x_rsc_4_0_i_s_waddr => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_waddr,
      x_rsc_4_0_i_s_waddr_core_sct => x_rsc_4_0_i_s_we_core_sct,
      x_rsc_4_0_i_s_din => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_din,
      x_rsc_4_0_i_s_dout => hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_dout
    );
  hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_raddr_core <= x_rsc_4_0_i_s_raddr_core;
  hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_waddr_core <= x_rsc_4_0_i_s_waddr_core;
  x_rsc_4_0_i_s_din_mxwt <= hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_din_mxwt;
  hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_dout_core <= x_rsc_4_0_i_s_dout_core;
  x_rsc_4_0_i_s_raddr <= hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_raddr;
  x_rsc_4_0_i_s_waddr <= hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_waddr;
  hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_din <= x_rsc_4_0_i_s_din;
  x_rsc_4_0_i_s_dout <= hybrid_core_x_rsc_4_0_i_x_rsc_4_0_wait_dp_inst_x_rsc_4_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_3_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_3_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_3_0_s_tdone : IN STD_LOGIC;
    x_rsc_3_0_tr_write_done : IN STD_LOGIC;
    x_rsc_3_0_RREADY : IN STD_LOGIC;
    x_rsc_3_0_RVALID : OUT STD_LOGIC;
    x_rsc_3_0_RUSER : OUT STD_LOGIC;
    x_rsc_3_0_RLAST : OUT STD_LOGIC;
    x_rsc_3_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_RID : OUT STD_LOGIC;
    x_rsc_3_0_ARREADY : OUT STD_LOGIC;
    x_rsc_3_0_ARVALID : IN STD_LOGIC;
    x_rsc_3_0_ARUSER : IN STD_LOGIC;
    x_rsc_3_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARLOCK : IN STD_LOGIC;
    x_rsc_3_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_3_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_3_0_ARID : IN STD_LOGIC;
    x_rsc_3_0_BREADY : IN STD_LOGIC;
    x_rsc_3_0_BVALID : OUT STD_LOGIC;
    x_rsc_3_0_BUSER : OUT STD_LOGIC;
    x_rsc_3_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_BID : OUT STD_LOGIC;
    x_rsc_3_0_WREADY : OUT STD_LOGIC;
    x_rsc_3_0_WVALID : IN STD_LOGIC;
    x_rsc_3_0_WUSER : IN STD_LOGIC;
    x_rsc_3_0_WLAST : IN STD_LOGIC;
    x_rsc_3_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_AWREADY : OUT STD_LOGIC;
    x_rsc_3_0_AWVALID : IN STD_LOGIC;
    x_rsc_3_0_AWUSER : IN STD_LOGIC;
    x_rsc_3_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWLOCK : IN STD_LOGIC;
    x_rsc_3_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_3_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_3_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_3_0_i_oswt : IN STD_LOGIC;
    x_rsc_3_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_3_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_3_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_3_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_3_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_3_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_3_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_3_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_3_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_3_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_3_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_3_0_i_oswt : IN STD_LOGIC;
      x_rsc_3_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_3_0_i_biwt : OUT STD_LOGIC;
      x_rsc_3_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_3_0_i_bcwt : IN STD_LOGIC;
      x_rsc_3_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_3_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_3_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_3_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_3_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_3_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_3_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_3_0_i_oswt : IN STD_LOGIC;
      x_rsc_3_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_3_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_3_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_3_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_3_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_3_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_i_biwt : IN STD_LOGIC;
      x_rsc_3_0_i_bdwt : IN STD_LOGIC;
      x_rsc_3_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_3_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_3_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_3_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_3_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_3_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_3_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_3_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_3_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_3_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_3_0_i_AWID,
      AWADDR => x_rsc_3_0_i_AWADDR,
      AWLEN => x_rsc_3_0_i_AWLEN,
      AWSIZE => x_rsc_3_0_i_AWSIZE,
      AWBURST => x_rsc_3_0_i_AWBURST,
      AWLOCK => x_rsc_3_0_AWLOCK,
      AWCACHE => x_rsc_3_0_i_AWCACHE,
      AWPROT => x_rsc_3_0_i_AWPROT,
      AWQOS => x_rsc_3_0_i_AWQOS,
      AWREGION => x_rsc_3_0_i_AWREGION,
      AWUSER => x_rsc_3_0_i_AWUSER,
      AWVALID => x_rsc_3_0_AWVALID,
      AWREADY => x_rsc_3_0_AWREADY,
      WDATA => x_rsc_3_0_i_WDATA,
      WSTRB => x_rsc_3_0_i_WSTRB,
      WLAST => x_rsc_3_0_WLAST,
      WUSER => x_rsc_3_0_i_WUSER,
      WVALID => x_rsc_3_0_WVALID,
      WREADY => x_rsc_3_0_WREADY,
      BID => x_rsc_3_0_i_BID,
      BRESP => x_rsc_3_0_i_BRESP,
      BUSER => x_rsc_3_0_i_BUSER,
      BVALID => x_rsc_3_0_BVALID,
      BREADY => x_rsc_3_0_BREADY,
      ARID => x_rsc_3_0_i_ARID,
      ARADDR => x_rsc_3_0_i_ARADDR,
      ARLEN => x_rsc_3_0_i_ARLEN,
      ARSIZE => x_rsc_3_0_i_ARSIZE,
      ARBURST => x_rsc_3_0_i_ARBURST,
      ARLOCK => x_rsc_3_0_ARLOCK,
      ARCACHE => x_rsc_3_0_i_ARCACHE,
      ARPROT => x_rsc_3_0_i_ARPROT,
      ARQOS => x_rsc_3_0_i_ARQOS,
      ARREGION => x_rsc_3_0_i_ARREGION,
      ARUSER => x_rsc_3_0_i_ARUSER,
      ARVALID => x_rsc_3_0_ARVALID,
      ARREADY => x_rsc_3_0_ARREADY,
      RID => x_rsc_3_0_i_RID,
      RDATA => x_rsc_3_0_i_RDATA,
      RRESP => x_rsc_3_0_i_RRESP,
      RLAST => x_rsc_3_0_RLAST,
      RUSER => x_rsc_3_0_i_RUSER,
      RVALID => x_rsc_3_0_RVALID,
      RREADY => x_rsc_3_0_RREADY,
      s_re => x_rsc_3_0_i_s_re_core_sct,
      s_we => x_rsc_3_0_i_s_we_core_sct,
      s_raddr => x_rsc_3_0_i_s_raddr_1,
      s_waddr => x_rsc_3_0_i_s_waddr_1,
      s_din => x_rsc_3_0_i_s_din_1,
      s_dout => x_rsc_3_0_i_s_dout_1,
      s_rrdy => x_rsc_3_0_i_s_rrdy,
      s_wrdy => x_rsc_3_0_i_s_wrdy,
      is_idle => x_rsc_3_0_is_idle_1,
      tr_write_done => x_rsc_3_0_tr_write_done,
      s_tdone => x_rsc_3_0_s_tdone
    );
  x_rsc_3_0_i_AWID(0) <= x_rsc_3_0_AWID;
  x_rsc_3_0_i_AWADDR <= x_rsc_3_0_AWADDR;
  x_rsc_3_0_i_AWLEN <= x_rsc_3_0_AWLEN;
  x_rsc_3_0_i_AWSIZE <= x_rsc_3_0_AWSIZE;
  x_rsc_3_0_i_AWBURST <= x_rsc_3_0_AWBURST;
  x_rsc_3_0_i_AWCACHE <= x_rsc_3_0_AWCACHE;
  x_rsc_3_0_i_AWPROT <= x_rsc_3_0_AWPROT;
  x_rsc_3_0_i_AWQOS <= x_rsc_3_0_AWQOS;
  x_rsc_3_0_i_AWREGION <= x_rsc_3_0_AWREGION;
  x_rsc_3_0_i_AWUSER(0) <= x_rsc_3_0_AWUSER;
  x_rsc_3_0_i_WDATA <= x_rsc_3_0_WDATA;
  x_rsc_3_0_i_WSTRB <= x_rsc_3_0_WSTRB;
  x_rsc_3_0_i_WUSER(0) <= x_rsc_3_0_WUSER;
  x_rsc_3_0_BID <= x_rsc_3_0_i_BID(0);
  x_rsc_3_0_BRESP <= x_rsc_3_0_i_BRESP;
  x_rsc_3_0_BUSER <= x_rsc_3_0_i_BUSER(0);
  x_rsc_3_0_i_ARID(0) <= x_rsc_3_0_ARID;
  x_rsc_3_0_i_ARADDR <= x_rsc_3_0_ARADDR;
  x_rsc_3_0_i_ARLEN <= x_rsc_3_0_ARLEN;
  x_rsc_3_0_i_ARSIZE <= x_rsc_3_0_ARSIZE;
  x_rsc_3_0_i_ARBURST <= x_rsc_3_0_ARBURST;
  x_rsc_3_0_i_ARCACHE <= x_rsc_3_0_ARCACHE;
  x_rsc_3_0_i_ARPROT <= x_rsc_3_0_ARPROT;
  x_rsc_3_0_i_ARQOS <= x_rsc_3_0_ARQOS;
  x_rsc_3_0_i_ARREGION <= x_rsc_3_0_ARREGION;
  x_rsc_3_0_i_ARUSER(0) <= x_rsc_3_0_ARUSER;
  x_rsc_3_0_RID <= x_rsc_3_0_i_RID(0);
  x_rsc_3_0_RDATA <= x_rsc_3_0_i_RDATA;
  x_rsc_3_0_RRESP <= x_rsc_3_0_i_RRESP;
  x_rsc_3_0_RUSER <= x_rsc_3_0_i_RUSER(0);
  x_rsc_3_0_i_s_raddr_1 <= x_rsc_3_0_i_s_raddr;
  x_rsc_3_0_i_s_waddr_1 <= x_rsc_3_0_i_s_waddr;
  x_rsc_3_0_i_s_din <= x_rsc_3_0_i_s_din_1;
  x_rsc_3_0_i_s_dout_1 <= x_rsc_3_0_i_s_dout;

  hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl_inst : hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_3_0_i_oswt => x_rsc_3_0_i_oswt,
      x_rsc_3_0_i_oswt_1 => x_rsc_3_0_i_oswt_1,
      x_rsc_3_0_i_biwt => x_rsc_3_0_i_biwt,
      x_rsc_3_0_i_bdwt => x_rsc_3_0_i_bdwt,
      x_rsc_3_0_i_bcwt => x_rsc_3_0_i_bcwt,
      x_rsc_3_0_i_s_re_core_sct => x_rsc_3_0_i_s_re_core_sct,
      x_rsc_3_0_i_biwt_1 => x_rsc_3_0_i_biwt_1,
      x_rsc_3_0_i_bdwt_2 => x_rsc_3_0_i_bdwt_2,
      x_rsc_3_0_i_bcwt_1 => x_rsc_3_0_i_bcwt_1,
      x_rsc_3_0_i_s_we_core_sct => x_rsc_3_0_i_s_we_core_sct,
      x_rsc_3_0_i_s_rrdy => x_rsc_3_0_i_s_rrdy,
      x_rsc_3_0_i_s_wrdy => x_rsc_3_0_i_s_wrdy
    );
  hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst : hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_3_0_i_oswt => x_rsc_3_0_i_oswt,
      x_rsc_3_0_i_wen_comp => x_rsc_3_0_i_wen_comp,
      x_rsc_3_0_i_oswt_1 => x_rsc_3_0_i_oswt_1,
      x_rsc_3_0_i_wen_comp_1 => x_rsc_3_0_i_wen_comp_1,
      x_rsc_3_0_i_s_raddr_core => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_raddr_core,
      x_rsc_3_0_i_s_waddr_core => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_waddr_core,
      x_rsc_3_0_i_s_din_mxwt => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_din_mxwt,
      x_rsc_3_0_i_s_dout_core => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_dout_core,
      x_rsc_3_0_i_biwt => x_rsc_3_0_i_biwt,
      x_rsc_3_0_i_bdwt => x_rsc_3_0_i_bdwt,
      x_rsc_3_0_i_bcwt => x_rsc_3_0_i_bcwt,
      x_rsc_3_0_i_biwt_1 => x_rsc_3_0_i_biwt_1,
      x_rsc_3_0_i_bdwt_2 => x_rsc_3_0_i_bdwt_2,
      x_rsc_3_0_i_bcwt_1 => x_rsc_3_0_i_bcwt_1,
      x_rsc_3_0_i_s_raddr => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_raddr,
      x_rsc_3_0_i_s_raddr_core_sct => x_rsc_3_0_i_s_re_core_sct,
      x_rsc_3_0_i_s_waddr => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_waddr,
      x_rsc_3_0_i_s_waddr_core_sct => x_rsc_3_0_i_s_we_core_sct,
      x_rsc_3_0_i_s_din => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_din,
      x_rsc_3_0_i_s_dout => hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_dout
    );
  hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_raddr_core <= x_rsc_3_0_i_s_raddr_core;
  hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_waddr_core <= x_rsc_3_0_i_s_waddr_core;
  x_rsc_3_0_i_s_din_mxwt <= hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_din_mxwt;
  hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_dout_core <= x_rsc_3_0_i_s_dout_core;
  x_rsc_3_0_i_s_raddr <= hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_raddr;
  x_rsc_3_0_i_s_waddr <= hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_waddr;
  hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_din <= x_rsc_3_0_i_s_din;
  x_rsc_3_0_i_s_dout <= hybrid_core_x_rsc_3_0_i_x_rsc_3_0_wait_dp_inst_x_rsc_3_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_2_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_2_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_2_0_s_tdone : IN STD_LOGIC;
    x_rsc_2_0_tr_write_done : IN STD_LOGIC;
    x_rsc_2_0_RREADY : IN STD_LOGIC;
    x_rsc_2_0_RVALID : OUT STD_LOGIC;
    x_rsc_2_0_RUSER : OUT STD_LOGIC;
    x_rsc_2_0_RLAST : OUT STD_LOGIC;
    x_rsc_2_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_RID : OUT STD_LOGIC;
    x_rsc_2_0_ARREADY : OUT STD_LOGIC;
    x_rsc_2_0_ARVALID : IN STD_LOGIC;
    x_rsc_2_0_ARUSER : IN STD_LOGIC;
    x_rsc_2_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARLOCK : IN STD_LOGIC;
    x_rsc_2_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_2_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_2_0_ARID : IN STD_LOGIC;
    x_rsc_2_0_BREADY : IN STD_LOGIC;
    x_rsc_2_0_BVALID : OUT STD_LOGIC;
    x_rsc_2_0_BUSER : OUT STD_LOGIC;
    x_rsc_2_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_BID : OUT STD_LOGIC;
    x_rsc_2_0_WREADY : OUT STD_LOGIC;
    x_rsc_2_0_WVALID : IN STD_LOGIC;
    x_rsc_2_0_WUSER : IN STD_LOGIC;
    x_rsc_2_0_WLAST : IN STD_LOGIC;
    x_rsc_2_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_AWREADY : OUT STD_LOGIC;
    x_rsc_2_0_AWVALID : IN STD_LOGIC;
    x_rsc_2_0_AWUSER : IN STD_LOGIC;
    x_rsc_2_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWLOCK : IN STD_LOGIC;
    x_rsc_2_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_2_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_2_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_2_0_i_oswt : IN STD_LOGIC;
    x_rsc_2_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_2_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_2_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_2_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_2_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_2_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_2_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_2_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_2_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_2_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_2_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_2_0_i_oswt : IN STD_LOGIC;
      x_rsc_2_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_2_0_i_biwt : OUT STD_LOGIC;
      x_rsc_2_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_2_0_i_bcwt : IN STD_LOGIC;
      x_rsc_2_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_2_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_2_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_2_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_2_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_2_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_2_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_2_0_i_oswt : IN STD_LOGIC;
      x_rsc_2_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_2_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_2_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_2_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_2_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_2_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_i_biwt : IN STD_LOGIC;
      x_rsc_2_0_i_bdwt : IN STD_LOGIC;
      x_rsc_2_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_2_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_2_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_2_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_2_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_2_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_2_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_2_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_2_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_2_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_2_0_i_AWID,
      AWADDR => x_rsc_2_0_i_AWADDR,
      AWLEN => x_rsc_2_0_i_AWLEN,
      AWSIZE => x_rsc_2_0_i_AWSIZE,
      AWBURST => x_rsc_2_0_i_AWBURST,
      AWLOCK => x_rsc_2_0_AWLOCK,
      AWCACHE => x_rsc_2_0_i_AWCACHE,
      AWPROT => x_rsc_2_0_i_AWPROT,
      AWQOS => x_rsc_2_0_i_AWQOS,
      AWREGION => x_rsc_2_0_i_AWREGION,
      AWUSER => x_rsc_2_0_i_AWUSER,
      AWVALID => x_rsc_2_0_AWVALID,
      AWREADY => x_rsc_2_0_AWREADY,
      WDATA => x_rsc_2_0_i_WDATA,
      WSTRB => x_rsc_2_0_i_WSTRB,
      WLAST => x_rsc_2_0_WLAST,
      WUSER => x_rsc_2_0_i_WUSER,
      WVALID => x_rsc_2_0_WVALID,
      WREADY => x_rsc_2_0_WREADY,
      BID => x_rsc_2_0_i_BID,
      BRESP => x_rsc_2_0_i_BRESP,
      BUSER => x_rsc_2_0_i_BUSER,
      BVALID => x_rsc_2_0_BVALID,
      BREADY => x_rsc_2_0_BREADY,
      ARID => x_rsc_2_0_i_ARID,
      ARADDR => x_rsc_2_0_i_ARADDR,
      ARLEN => x_rsc_2_0_i_ARLEN,
      ARSIZE => x_rsc_2_0_i_ARSIZE,
      ARBURST => x_rsc_2_0_i_ARBURST,
      ARLOCK => x_rsc_2_0_ARLOCK,
      ARCACHE => x_rsc_2_0_i_ARCACHE,
      ARPROT => x_rsc_2_0_i_ARPROT,
      ARQOS => x_rsc_2_0_i_ARQOS,
      ARREGION => x_rsc_2_0_i_ARREGION,
      ARUSER => x_rsc_2_0_i_ARUSER,
      ARVALID => x_rsc_2_0_ARVALID,
      ARREADY => x_rsc_2_0_ARREADY,
      RID => x_rsc_2_0_i_RID,
      RDATA => x_rsc_2_0_i_RDATA,
      RRESP => x_rsc_2_0_i_RRESP,
      RLAST => x_rsc_2_0_RLAST,
      RUSER => x_rsc_2_0_i_RUSER,
      RVALID => x_rsc_2_0_RVALID,
      RREADY => x_rsc_2_0_RREADY,
      s_re => x_rsc_2_0_i_s_re_core_sct,
      s_we => x_rsc_2_0_i_s_we_core_sct,
      s_raddr => x_rsc_2_0_i_s_raddr_1,
      s_waddr => x_rsc_2_0_i_s_waddr_1,
      s_din => x_rsc_2_0_i_s_din_1,
      s_dout => x_rsc_2_0_i_s_dout_1,
      s_rrdy => x_rsc_2_0_i_s_rrdy,
      s_wrdy => x_rsc_2_0_i_s_wrdy,
      is_idle => x_rsc_2_0_is_idle_1,
      tr_write_done => x_rsc_2_0_tr_write_done,
      s_tdone => x_rsc_2_0_s_tdone
    );
  x_rsc_2_0_i_AWID(0) <= x_rsc_2_0_AWID;
  x_rsc_2_0_i_AWADDR <= x_rsc_2_0_AWADDR;
  x_rsc_2_0_i_AWLEN <= x_rsc_2_0_AWLEN;
  x_rsc_2_0_i_AWSIZE <= x_rsc_2_0_AWSIZE;
  x_rsc_2_0_i_AWBURST <= x_rsc_2_0_AWBURST;
  x_rsc_2_0_i_AWCACHE <= x_rsc_2_0_AWCACHE;
  x_rsc_2_0_i_AWPROT <= x_rsc_2_0_AWPROT;
  x_rsc_2_0_i_AWQOS <= x_rsc_2_0_AWQOS;
  x_rsc_2_0_i_AWREGION <= x_rsc_2_0_AWREGION;
  x_rsc_2_0_i_AWUSER(0) <= x_rsc_2_0_AWUSER;
  x_rsc_2_0_i_WDATA <= x_rsc_2_0_WDATA;
  x_rsc_2_0_i_WSTRB <= x_rsc_2_0_WSTRB;
  x_rsc_2_0_i_WUSER(0) <= x_rsc_2_0_WUSER;
  x_rsc_2_0_BID <= x_rsc_2_0_i_BID(0);
  x_rsc_2_0_BRESP <= x_rsc_2_0_i_BRESP;
  x_rsc_2_0_BUSER <= x_rsc_2_0_i_BUSER(0);
  x_rsc_2_0_i_ARID(0) <= x_rsc_2_0_ARID;
  x_rsc_2_0_i_ARADDR <= x_rsc_2_0_ARADDR;
  x_rsc_2_0_i_ARLEN <= x_rsc_2_0_ARLEN;
  x_rsc_2_0_i_ARSIZE <= x_rsc_2_0_ARSIZE;
  x_rsc_2_0_i_ARBURST <= x_rsc_2_0_ARBURST;
  x_rsc_2_0_i_ARCACHE <= x_rsc_2_0_ARCACHE;
  x_rsc_2_0_i_ARPROT <= x_rsc_2_0_ARPROT;
  x_rsc_2_0_i_ARQOS <= x_rsc_2_0_ARQOS;
  x_rsc_2_0_i_ARREGION <= x_rsc_2_0_ARREGION;
  x_rsc_2_0_i_ARUSER(0) <= x_rsc_2_0_ARUSER;
  x_rsc_2_0_RID <= x_rsc_2_0_i_RID(0);
  x_rsc_2_0_RDATA <= x_rsc_2_0_i_RDATA;
  x_rsc_2_0_RRESP <= x_rsc_2_0_i_RRESP;
  x_rsc_2_0_RUSER <= x_rsc_2_0_i_RUSER(0);
  x_rsc_2_0_i_s_raddr_1 <= x_rsc_2_0_i_s_raddr;
  x_rsc_2_0_i_s_waddr_1 <= x_rsc_2_0_i_s_waddr;
  x_rsc_2_0_i_s_din <= x_rsc_2_0_i_s_din_1;
  x_rsc_2_0_i_s_dout_1 <= x_rsc_2_0_i_s_dout;

  hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl_inst : hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_2_0_i_oswt => x_rsc_2_0_i_oswt,
      x_rsc_2_0_i_oswt_1 => x_rsc_2_0_i_oswt_1,
      x_rsc_2_0_i_biwt => x_rsc_2_0_i_biwt,
      x_rsc_2_0_i_bdwt => x_rsc_2_0_i_bdwt,
      x_rsc_2_0_i_bcwt => x_rsc_2_0_i_bcwt,
      x_rsc_2_0_i_s_re_core_sct => x_rsc_2_0_i_s_re_core_sct,
      x_rsc_2_0_i_biwt_1 => x_rsc_2_0_i_biwt_1,
      x_rsc_2_0_i_bdwt_2 => x_rsc_2_0_i_bdwt_2,
      x_rsc_2_0_i_bcwt_1 => x_rsc_2_0_i_bcwt_1,
      x_rsc_2_0_i_s_we_core_sct => x_rsc_2_0_i_s_we_core_sct,
      x_rsc_2_0_i_s_rrdy => x_rsc_2_0_i_s_rrdy,
      x_rsc_2_0_i_s_wrdy => x_rsc_2_0_i_s_wrdy
    );
  hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst : hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_2_0_i_oswt => x_rsc_2_0_i_oswt,
      x_rsc_2_0_i_wen_comp => x_rsc_2_0_i_wen_comp,
      x_rsc_2_0_i_oswt_1 => x_rsc_2_0_i_oswt_1,
      x_rsc_2_0_i_wen_comp_1 => x_rsc_2_0_i_wen_comp_1,
      x_rsc_2_0_i_s_raddr_core => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_raddr_core,
      x_rsc_2_0_i_s_waddr_core => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_waddr_core,
      x_rsc_2_0_i_s_din_mxwt => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_din_mxwt,
      x_rsc_2_0_i_s_dout_core => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_dout_core,
      x_rsc_2_0_i_biwt => x_rsc_2_0_i_biwt,
      x_rsc_2_0_i_bdwt => x_rsc_2_0_i_bdwt,
      x_rsc_2_0_i_bcwt => x_rsc_2_0_i_bcwt,
      x_rsc_2_0_i_biwt_1 => x_rsc_2_0_i_biwt_1,
      x_rsc_2_0_i_bdwt_2 => x_rsc_2_0_i_bdwt_2,
      x_rsc_2_0_i_bcwt_1 => x_rsc_2_0_i_bcwt_1,
      x_rsc_2_0_i_s_raddr => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_raddr,
      x_rsc_2_0_i_s_raddr_core_sct => x_rsc_2_0_i_s_re_core_sct,
      x_rsc_2_0_i_s_waddr => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_waddr,
      x_rsc_2_0_i_s_waddr_core_sct => x_rsc_2_0_i_s_we_core_sct,
      x_rsc_2_0_i_s_din => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_din,
      x_rsc_2_0_i_s_dout => hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_dout
    );
  hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_raddr_core <= x_rsc_2_0_i_s_raddr_core;
  hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_waddr_core <= x_rsc_2_0_i_s_waddr_core;
  x_rsc_2_0_i_s_din_mxwt <= hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_din_mxwt;
  hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_dout_core <= x_rsc_2_0_i_s_dout_core;
  x_rsc_2_0_i_s_raddr <= hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_raddr;
  x_rsc_2_0_i_s_waddr <= hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_waddr;
  hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_din <= x_rsc_2_0_i_s_din;
  x_rsc_2_0_i_s_dout <= hybrid_core_x_rsc_2_0_i_x_rsc_2_0_wait_dp_inst_x_rsc_2_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_1_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_1_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_1_0_s_tdone : IN STD_LOGIC;
    x_rsc_1_0_tr_write_done : IN STD_LOGIC;
    x_rsc_1_0_RREADY : IN STD_LOGIC;
    x_rsc_1_0_RVALID : OUT STD_LOGIC;
    x_rsc_1_0_RUSER : OUT STD_LOGIC;
    x_rsc_1_0_RLAST : OUT STD_LOGIC;
    x_rsc_1_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_RID : OUT STD_LOGIC;
    x_rsc_1_0_ARREADY : OUT STD_LOGIC;
    x_rsc_1_0_ARVALID : IN STD_LOGIC;
    x_rsc_1_0_ARUSER : IN STD_LOGIC;
    x_rsc_1_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARLOCK : IN STD_LOGIC;
    x_rsc_1_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_1_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_1_0_ARID : IN STD_LOGIC;
    x_rsc_1_0_BREADY : IN STD_LOGIC;
    x_rsc_1_0_BVALID : OUT STD_LOGIC;
    x_rsc_1_0_BUSER : OUT STD_LOGIC;
    x_rsc_1_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_BID : OUT STD_LOGIC;
    x_rsc_1_0_WREADY : OUT STD_LOGIC;
    x_rsc_1_0_WVALID : IN STD_LOGIC;
    x_rsc_1_0_WUSER : IN STD_LOGIC;
    x_rsc_1_0_WLAST : IN STD_LOGIC;
    x_rsc_1_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_AWREADY : OUT STD_LOGIC;
    x_rsc_1_0_AWVALID : IN STD_LOGIC;
    x_rsc_1_0_AWUSER : IN STD_LOGIC;
    x_rsc_1_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWLOCK : IN STD_LOGIC;
    x_rsc_1_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_1_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_1_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_1_0_i_oswt : IN STD_LOGIC;
    x_rsc_1_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_1_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_1_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_1_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_1_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_1_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_1_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_1_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_1_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_1_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_1_0_i_oswt : IN STD_LOGIC;
      x_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_1_0_i_biwt : OUT STD_LOGIC;
      x_rsc_1_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_1_0_i_bcwt : IN STD_LOGIC;
      x_rsc_1_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_1_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_1_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_1_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_1_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_1_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_1_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_1_0_i_oswt : IN STD_LOGIC;
      x_rsc_1_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_1_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_1_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_1_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_1_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_i_biwt : IN STD_LOGIC;
      x_rsc_1_0_i_bdwt : IN STD_LOGIC;
      x_rsc_1_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_1_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_1_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_1_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_1_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_1_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_1_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_1_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_1_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_1_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_1_0_i_AWID,
      AWADDR => x_rsc_1_0_i_AWADDR,
      AWLEN => x_rsc_1_0_i_AWLEN,
      AWSIZE => x_rsc_1_0_i_AWSIZE,
      AWBURST => x_rsc_1_0_i_AWBURST,
      AWLOCK => x_rsc_1_0_AWLOCK,
      AWCACHE => x_rsc_1_0_i_AWCACHE,
      AWPROT => x_rsc_1_0_i_AWPROT,
      AWQOS => x_rsc_1_0_i_AWQOS,
      AWREGION => x_rsc_1_0_i_AWREGION,
      AWUSER => x_rsc_1_0_i_AWUSER,
      AWVALID => x_rsc_1_0_AWVALID,
      AWREADY => x_rsc_1_0_AWREADY,
      WDATA => x_rsc_1_0_i_WDATA,
      WSTRB => x_rsc_1_0_i_WSTRB,
      WLAST => x_rsc_1_0_WLAST,
      WUSER => x_rsc_1_0_i_WUSER,
      WVALID => x_rsc_1_0_WVALID,
      WREADY => x_rsc_1_0_WREADY,
      BID => x_rsc_1_0_i_BID,
      BRESP => x_rsc_1_0_i_BRESP,
      BUSER => x_rsc_1_0_i_BUSER,
      BVALID => x_rsc_1_0_BVALID,
      BREADY => x_rsc_1_0_BREADY,
      ARID => x_rsc_1_0_i_ARID,
      ARADDR => x_rsc_1_0_i_ARADDR,
      ARLEN => x_rsc_1_0_i_ARLEN,
      ARSIZE => x_rsc_1_0_i_ARSIZE,
      ARBURST => x_rsc_1_0_i_ARBURST,
      ARLOCK => x_rsc_1_0_ARLOCK,
      ARCACHE => x_rsc_1_0_i_ARCACHE,
      ARPROT => x_rsc_1_0_i_ARPROT,
      ARQOS => x_rsc_1_0_i_ARQOS,
      ARREGION => x_rsc_1_0_i_ARREGION,
      ARUSER => x_rsc_1_0_i_ARUSER,
      ARVALID => x_rsc_1_0_ARVALID,
      ARREADY => x_rsc_1_0_ARREADY,
      RID => x_rsc_1_0_i_RID,
      RDATA => x_rsc_1_0_i_RDATA,
      RRESP => x_rsc_1_0_i_RRESP,
      RLAST => x_rsc_1_0_RLAST,
      RUSER => x_rsc_1_0_i_RUSER,
      RVALID => x_rsc_1_0_RVALID,
      RREADY => x_rsc_1_0_RREADY,
      s_re => x_rsc_1_0_i_s_re_core_sct,
      s_we => x_rsc_1_0_i_s_we_core_sct,
      s_raddr => x_rsc_1_0_i_s_raddr_1,
      s_waddr => x_rsc_1_0_i_s_waddr_1,
      s_din => x_rsc_1_0_i_s_din_1,
      s_dout => x_rsc_1_0_i_s_dout_1,
      s_rrdy => x_rsc_1_0_i_s_rrdy,
      s_wrdy => x_rsc_1_0_i_s_wrdy,
      is_idle => x_rsc_1_0_is_idle_1,
      tr_write_done => x_rsc_1_0_tr_write_done,
      s_tdone => x_rsc_1_0_s_tdone
    );
  x_rsc_1_0_i_AWID(0) <= x_rsc_1_0_AWID;
  x_rsc_1_0_i_AWADDR <= x_rsc_1_0_AWADDR;
  x_rsc_1_0_i_AWLEN <= x_rsc_1_0_AWLEN;
  x_rsc_1_0_i_AWSIZE <= x_rsc_1_0_AWSIZE;
  x_rsc_1_0_i_AWBURST <= x_rsc_1_0_AWBURST;
  x_rsc_1_0_i_AWCACHE <= x_rsc_1_0_AWCACHE;
  x_rsc_1_0_i_AWPROT <= x_rsc_1_0_AWPROT;
  x_rsc_1_0_i_AWQOS <= x_rsc_1_0_AWQOS;
  x_rsc_1_0_i_AWREGION <= x_rsc_1_0_AWREGION;
  x_rsc_1_0_i_AWUSER(0) <= x_rsc_1_0_AWUSER;
  x_rsc_1_0_i_WDATA <= x_rsc_1_0_WDATA;
  x_rsc_1_0_i_WSTRB <= x_rsc_1_0_WSTRB;
  x_rsc_1_0_i_WUSER(0) <= x_rsc_1_0_WUSER;
  x_rsc_1_0_BID <= x_rsc_1_0_i_BID(0);
  x_rsc_1_0_BRESP <= x_rsc_1_0_i_BRESP;
  x_rsc_1_0_BUSER <= x_rsc_1_0_i_BUSER(0);
  x_rsc_1_0_i_ARID(0) <= x_rsc_1_0_ARID;
  x_rsc_1_0_i_ARADDR <= x_rsc_1_0_ARADDR;
  x_rsc_1_0_i_ARLEN <= x_rsc_1_0_ARLEN;
  x_rsc_1_0_i_ARSIZE <= x_rsc_1_0_ARSIZE;
  x_rsc_1_0_i_ARBURST <= x_rsc_1_0_ARBURST;
  x_rsc_1_0_i_ARCACHE <= x_rsc_1_0_ARCACHE;
  x_rsc_1_0_i_ARPROT <= x_rsc_1_0_ARPROT;
  x_rsc_1_0_i_ARQOS <= x_rsc_1_0_ARQOS;
  x_rsc_1_0_i_ARREGION <= x_rsc_1_0_ARREGION;
  x_rsc_1_0_i_ARUSER(0) <= x_rsc_1_0_ARUSER;
  x_rsc_1_0_RID <= x_rsc_1_0_i_RID(0);
  x_rsc_1_0_RDATA <= x_rsc_1_0_i_RDATA;
  x_rsc_1_0_RRESP <= x_rsc_1_0_i_RRESP;
  x_rsc_1_0_RUSER <= x_rsc_1_0_i_RUSER(0);
  x_rsc_1_0_i_s_raddr_1 <= x_rsc_1_0_i_s_raddr;
  x_rsc_1_0_i_s_waddr_1 <= x_rsc_1_0_i_s_waddr;
  x_rsc_1_0_i_s_din <= x_rsc_1_0_i_s_din_1;
  x_rsc_1_0_i_s_dout_1 <= x_rsc_1_0_i_s_dout;

  hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl_inst : hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_1_0_i_oswt => x_rsc_1_0_i_oswt,
      x_rsc_1_0_i_oswt_1 => x_rsc_1_0_i_oswt_1,
      x_rsc_1_0_i_biwt => x_rsc_1_0_i_biwt,
      x_rsc_1_0_i_bdwt => x_rsc_1_0_i_bdwt,
      x_rsc_1_0_i_bcwt => x_rsc_1_0_i_bcwt,
      x_rsc_1_0_i_s_re_core_sct => x_rsc_1_0_i_s_re_core_sct,
      x_rsc_1_0_i_biwt_1 => x_rsc_1_0_i_biwt_1,
      x_rsc_1_0_i_bdwt_2 => x_rsc_1_0_i_bdwt_2,
      x_rsc_1_0_i_bcwt_1 => x_rsc_1_0_i_bcwt_1,
      x_rsc_1_0_i_s_we_core_sct => x_rsc_1_0_i_s_we_core_sct,
      x_rsc_1_0_i_s_rrdy => x_rsc_1_0_i_s_rrdy,
      x_rsc_1_0_i_s_wrdy => x_rsc_1_0_i_s_wrdy
    );
  hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst : hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_1_0_i_oswt => x_rsc_1_0_i_oswt,
      x_rsc_1_0_i_wen_comp => x_rsc_1_0_i_wen_comp,
      x_rsc_1_0_i_oswt_1 => x_rsc_1_0_i_oswt_1,
      x_rsc_1_0_i_wen_comp_1 => x_rsc_1_0_i_wen_comp_1,
      x_rsc_1_0_i_s_raddr_core => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_raddr_core,
      x_rsc_1_0_i_s_waddr_core => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_waddr_core,
      x_rsc_1_0_i_s_din_mxwt => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_din_mxwt,
      x_rsc_1_0_i_s_dout_core => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_dout_core,
      x_rsc_1_0_i_biwt => x_rsc_1_0_i_biwt,
      x_rsc_1_0_i_bdwt => x_rsc_1_0_i_bdwt,
      x_rsc_1_0_i_bcwt => x_rsc_1_0_i_bcwt,
      x_rsc_1_0_i_biwt_1 => x_rsc_1_0_i_biwt_1,
      x_rsc_1_0_i_bdwt_2 => x_rsc_1_0_i_bdwt_2,
      x_rsc_1_0_i_bcwt_1 => x_rsc_1_0_i_bcwt_1,
      x_rsc_1_0_i_s_raddr => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_raddr,
      x_rsc_1_0_i_s_raddr_core_sct => x_rsc_1_0_i_s_re_core_sct,
      x_rsc_1_0_i_s_waddr => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_waddr,
      x_rsc_1_0_i_s_waddr_core_sct => x_rsc_1_0_i_s_we_core_sct,
      x_rsc_1_0_i_s_din => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_din,
      x_rsc_1_0_i_s_dout => hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_dout
    );
  hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_raddr_core <= x_rsc_1_0_i_s_raddr_core;
  hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_waddr_core <= x_rsc_1_0_i_s_waddr_core;
  x_rsc_1_0_i_s_din_mxwt <= hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_din_mxwt;
  hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_dout_core <= x_rsc_1_0_i_s_dout_core;
  x_rsc_1_0_i_s_raddr <= hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_raddr;
  x_rsc_1_0_i_s_waddr <= hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_waddr;
  hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_din <= x_rsc_1_0_i_s_din;
  x_rsc_1_0_i_s_dout <= hybrid_core_x_rsc_1_0_i_x_rsc_1_0_wait_dp_inst_x_rsc_1_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_x_rsc_0_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_x_rsc_0_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_0_0_s_tdone : IN STD_LOGIC;
    x_rsc_0_0_tr_write_done : IN STD_LOGIC;
    x_rsc_0_0_RREADY : IN STD_LOGIC;
    x_rsc_0_0_RVALID : OUT STD_LOGIC;
    x_rsc_0_0_RUSER : OUT STD_LOGIC;
    x_rsc_0_0_RLAST : OUT STD_LOGIC;
    x_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_RID : OUT STD_LOGIC;
    x_rsc_0_0_ARREADY : OUT STD_LOGIC;
    x_rsc_0_0_ARVALID : IN STD_LOGIC;
    x_rsc_0_0_ARUSER : IN STD_LOGIC;
    x_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARLOCK : IN STD_LOGIC;
    x_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_0_0_ARID : IN STD_LOGIC;
    x_rsc_0_0_BREADY : IN STD_LOGIC;
    x_rsc_0_0_BVALID : OUT STD_LOGIC;
    x_rsc_0_0_BUSER : OUT STD_LOGIC;
    x_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_BID : OUT STD_LOGIC;
    x_rsc_0_0_WREADY : OUT STD_LOGIC;
    x_rsc_0_0_WVALID : IN STD_LOGIC;
    x_rsc_0_0_WUSER : IN STD_LOGIC;
    x_rsc_0_0_WLAST : IN STD_LOGIC;
    x_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_AWREADY : OUT STD_LOGIC;
    x_rsc_0_0_AWVALID : IN STD_LOGIC;
    x_rsc_0_0_AWUSER : IN STD_LOGIC;
    x_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWLOCK : IN STD_LOGIC;
    x_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_0_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    x_rsc_0_0_i_oswt : IN STD_LOGIC;
    x_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
    x_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
    x_rsc_0_0_i_wen_comp_1 : OUT STD_LOGIC;
    x_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_0_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    x_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END hybrid_core_x_rsc_0_0_i;

ARCHITECTURE v14 OF hybrid_core_x_rsc_0_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL x_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_biwt_1 : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_bdwt_2 : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_bcwt_1 : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_s_we_core_sct : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_rrdy : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_s_wrdy : STD_LOGIC;
  SIGNAL x_rsc_0_0_is_idle_1 : STD_LOGIC;

  SIGNAL x_rsc_0_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_waddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_s_dout_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      x_rsc_0_0_i_oswt : IN STD_LOGIC;
      x_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_0_0_i_biwt : OUT STD_LOGIC;
      x_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      x_rsc_0_0_i_bcwt : IN STD_LOGIC;
      x_rsc_0_0_i_s_re_core_sct : OUT STD_LOGIC;
      x_rsc_0_0_i_biwt_1 : OUT STD_LOGIC;
      x_rsc_0_0_i_bdwt_2 : OUT STD_LOGIC;
      x_rsc_0_0_i_bcwt_1 : IN STD_LOGIC;
      x_rsc_0_0_i_s_we_core_sct : OUT STD_LOGIC;
      x_rsc_0_0_i_s_rrdy : IN STD_LOGIC;
      x_rsc_0_0_i_s_wrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_0_0_i_oswt : IN STD_LOGIC;
      x_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_0_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_0_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_i_biwt : IN STD_LOGIC;
      x_rsc_0_0_i_bdwt : IN STD_LOGIC;
      x_rsc_0_0_i_bcwt : OUT STD_LOGIC;
      x_rsc_0_0_i_biwt_1 : IN STD_LOGIC;
      x_rsc_0_0_i_bdwt_2 : IN STD_LOGIC;
      x_rsc_0_0_i_bcwt_1 : OUT STD_LOGIC;
      x_rsc_0_0_i_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_0_0_i_s_raddr_core_sct : IN STD_LOGIC;
      x_rsc_0_0_i_s_waddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_0_0_i_s_waddr_core_sct : IN STD_LOGIC;
      x_rsc_0_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_i_s_dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_waddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_dout_core :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_waddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_dout : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  x_rsc_0_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 32,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => x_rsc_0_0_i_AWID,
      AWADDR => x_rsc_0_0_i_AWADDR,
      AWLEN => x_rsc_0_0_i_AWLEN,
      AWSIZE => x_rsc_0_0_i_AWSIZE,
      AWBURST => x_rsc_0_0_i_AWBURST,
      AWLOCK => x_rsc_0_0_AWLOCK,
      AWCACHE => x_rsc_0_0_i_AWCACHE,
      AWPROT => x_rsc_0_0_i_AWPROT,
      AWQOS => x_rsc_0_0_i_AWQOS,
      AWREGION => x_rsc_0_0_i_AWREGION,
      AWUSER => x_rsc_0_0_i_AWUSER,
      AWVALID => x_rsc_0_0_AWVALID,
      AWREADY => x_rsc_0_0_AWREADY,
      WDATA => x_rsc_0_0_i_WDATA,
      WSTRB => x_rsc_0_0_i_WSTRB,
      WLAST => x_rsc_0_0_WLAST,
      WUSER => x_rsc_0_0_i_WUSER,
      WVALID => x_rsc_0_0_WVALID,
      WREADY => x_rsc_0_0_WREADY,
      BID => x_rsc_0_0_i_BID,
      BRESP => x_rsc_0_0_i_BRESP,
      BUSER => x_rsc_0_0_i_BUSER,
      BVALID => x_rsc_0_0_BVALID,
      BREADY => x_rsc_0_0_BREADY,
      ARID => x_rsc_0_0_i_ARID,
      ARADDR => x_rsc_0_0_i_ARADDR,
      ARLEN => x_rsc_0_0_i_ARLEN,
      ARSIZE => x_rsc_0_0_i_ARSIZE,
      ARBURST => x_rsc_0_0_i_ARBURST,
      ARLOCK => x_rsc_0_0_ARLOCK,
      ARCACHE => x_rsc_0_0_i_ARCACHE,
      ARPROT => x_rsc_0_0_i_ARPROT,
      ARQOS => x_rsc_0_0_i_ARQOS,
      ARREGION => x_rsc_0_0_i_ARREGION,
      ARUSER => x_rsc_0_0_i_ARUSER,
      ARVALID => x_rsc_0_0_ARVALID,
      ARREADY => x_rsc_0_0_ARREADY,
      RID => x_rsc_0_0_i_RID,
      RDATA => x_rsc_0_0_i_RDATA,
      RRESP => x_rsc_0_0_i_RRESP,
      RLAST => x_rsc_0_0_RLAST,
      RUSER => x_rsc_0_0_i_RUSER,
      RVALID => x_rsc_0_0_RVALID,
      RREADY => x_rsc_0_0_RREADY,
      s_re => x_rsc_0_0_i_s_re_core_sct,
      s_we => x_rsc_0_0_i_s_we_core_sct,
      s_raddr => x_rsc_0_0_i_s_raddr_1,
      s_waddr => x_rsc_0_0_i_s_waddr_1,
      s_din => x_rsc_0_0_i_s_din_1,
      s_dout => x_rsc_0_0_i_s_dout_1,
      s_rrdy => x_rsc_0_0_i_s_rrdy,
      s_wrdy => x_rsc_0_0_i_s_wrdy,
      is_idle => x_rsc_0_0_is_idle_1,
      tr_write_done => x_rsc_0_0_tr_write_done,
      s_tdone => x_rsc_0_0_s_tdone
    );
  x_rsc_0_0_i_AWID(0) <= x_rsc_0_0_AWID;
  x_rsc_0_0_i_AWADDR <= x_rsc_0_0_AWADDR;
  x_rsc_0_0_i_AWLEN <= x_rsc_0_0_AWLEN;
  x_rsc_0_0_i_AWSIZE <= x_rsc_0_0_AWSIZE;
  x_rsc_0_0_i_AWBURST <= x_rsc_0_0_AWBURST;
  x_rsc_0_0_i_AWCACHE <= x_rsc_0_0_AWCACHE;
  x_rsc_0_0_i_AWPROT <= x_rsc_0_0_AWPROT;
  x_rsc_0_0_i_AWQOS <= x_rsc_0_0_AWQOS;
  x_rsc_0_0_i_AWREGION <= x_rsc_0_0_AWREGION;
  x_rsc_0_0_i_AWUSER(0) <= x_rsc_0_0_AWUSER;
  x_rsc_0_0_i_WDATA <= x_rsc_0_0_WDATA;
  x_rsc_0_0_i_WSTRB <= x_rsc_0_0_WSTRB;
  x_rsc_0_0_i_WUSER(0) <= x_rsc_0_0_WUSER;
  x_rsc_0_0_BID <= x_rsc_0_0_i_BID(0);
  x_rsc_0_0_BRESP <= x_rsc_0_0_i_BRESP;
  x_rsc_0_0_BUSER <= x_rsc_0_0_i_BUSER(0);
  x_rsc_0_0_i_ARID(0) <= x_rsc_0_0_ARID;
  x_rsc_0_0_i_ARADDR <= x_rsc_0_0_ARADDR;
  x_rsc_0_0_i_ARLEN <= x_rsc_0_0_ARLEN;
  x_rsc_0_0_i_ARSIZE <= x_rsc_0_0_ARSIZE;
  x_rsc_0_0_i_ARBURST <= x_rsc_0_0_ARBURST;
  x_rsc_0_0_i_ARCACHE <= x_rsc_0_0_ARCACHE;
  x_rsc_0_0_i_ARPROT <= x_rsc_0_0_ARPROT;
  x_rsc_0_0_i_ARQOS <= x_rsc_0_0_ARQOS;
  x_rsc_0_0_i_ARREGION <= x_rsc_0_0_ARREGION;
  x_rsc_0_0_i_ARUSER(0) <= x_rsc_0_0_ARUSER;
  x_rsc_0_0_RID <= x_rsc_0_0_i_RID(0);
  x_rsc_0_0_RDATA <= x_rsc_0_0_i_RDATA;
  x_rsc_0_0_RRESP <= x_rsc_0_0_i_RRESP;
  x_rsc_0_0_RUSER <= x_rsc_0_0_i_RUSER(0);
  x_rsc_0_0_i_s_raddr_1 <= x_rsc_0_0_i_s_raddr;
  x_rsc_0_0_i_s_waddr_1 <= x_rsc_0_0_i_s_waddr;
  x_rsc_0_0_i_s_din <= x_rsc_0_0_i_s_din_1;
  x_rsc_0_0_i_s_dout_1 <= x_rsc_0_0_i_s_dout;

  hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl_inst : hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      x_rsc_0_0_i_oswt => x_rsc_0_0_i_oswt,
      x_rsc_0_0_i_oswt_1 => x_rsc_0_0_i_oswt_1,
      x_rsc_0_0_i_biwt => x_rsc_0_0_i_biwt,
      x_rsc_0_0_i_bdwt => x_rsc_0_0_i_bdwt,
      x_rsc_0_0_i_bcwt => x_rsc_0_0_i_bcwt,
      x_rsc_0_0_i_s_re_core_sct => x_rsc_0_0_i_s_re_core_sct,
      x_rsc_0_0_i_biwt_1 => x_rsc_0_0_i_biwt_1,
      x_rsc_0_0_i_bdwt_2 => x_rsc_0_0_i_bdwt_2,
      x_rsc_0_0_i_bcwt_1 => x_rsc_0_0_i_bcwt_1,
      x_rsc_0_0_i_s_we_core_sct => x_rsc_0_0_i_s_we_core_sct,
      x_rsc_0_0_i_s_rrdy => x_rsc_0_0_i_s_rrdy,
      x_rsc_0_0_i_s_wrdy => x_rsc_0_0_i_s_wrdy
    );
  hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst : hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_0_0_i_oswt => x_rsc_0_0_i_oswt,
      x_rsc_0_0_i_wen_comp => x_rsc_0_0_i_wen_comp,
      x_rsc_0_0_i_oswt_1 => x_rsc_0_0_i_oswt_1,
      x_rsc_0_0_i_wen_comp_1 => x_rsc_0_0_i_wen_comp_1,
      x_rsc_0_0_i_s_raddr_core => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_raddr_core,
      x_rsc_0_0_i_s_waddr_core => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_waddr_core,
      x_rsc_0_0_i_s_din_mxwt => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_din_mxwt,
      x_rsc_0_0_i_s_dout_core => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_dout_core,
      x_rsc_0_0_i_biwt => x_rsc_0_0_i_biwt,
      x_rsc_0_0_i_bdwt => x_rsc_0_0_i_bdwt,
      x_rsc_0_0_i_bcwt => x_rsc_0_0_i_bcwt,
      x_rsc_0_0_i_biwt_1 => x_rsc_0_0_i_biwt_1,
      x_rsc_0_0_i_bdwt_2 => x_rsc_0_0_i_bdwt_2,
      x_rsc_0_0_i_bcwt_1 => x_rsc_0_0_i_bcwt_1,
      x_rsc_0_0_i_s_raddr => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_raddr,
      x_rsc_0_0_i_s_raddr_core_sct => x_rsc_0_0_i_s_re_core_sct,
      x_rsc_0_0_i_s_waddr => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_waddr,
      x_rsc_0_0_i_s_waddr_core_sct => x_rsc_0_0_i_s_we_core_sct,
      x_rsc_0_0_i_s_din => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_din,
      x_rsc_0_0_i_s_dout => hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_dout
    );
  hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_raddr_core <= x_rsc_0_0_i_s_raddr_core;
  hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_waddr_core <= x_rsc_0_0_i_s_waddr_core;
  x_rsc_0_0_i_s_din_mxwt <= hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_din_mxwt;
  hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_dout_core <= x_rsc_0_0_i_s_dout_core;
  x_rsc_0_0_i_s_raddr <= hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_raddr;
  x_rsc_0_0_i_s_waddr <= hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_waddr;
  hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_din <= x_rsc_0_0_i_s_din;
  x_rsc_0_0_i_s_dout <= hybrid_core_x_rsc_0_0_i_x_rsc_0_0_wait_dp_inst_x_rsc_0_0_i_s_dout;

END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_h_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_h_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    tw_h_rsc_s_tdone : IN STD_LOGIC;
    tw_h_rsc_tr_write_done : IN STD_LOGIC;
    tw_h_rsc_RREADY : IN STD_LOGIC;
    tw_h_rsc_RVALID : OUT STD_LOGIC;
    tw_h_rsc_RUSER : OUT STD_LOGIC;
    tw_h_rsc_RLAST : OUT STD_LOGIC;
    tw_h_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_h_rsc_RID : OUT STD_LOGIC;
    tw_h_rsc_ARREADY : OUT STD_LOGIC;
    tw_h_rsc_ARVALID : IN STD_LOGIC;
    tw_h_rsc_ARUSER : IN STD_LOGIC;
    tw_h_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARLOCK : IN STD_LOGIC;
    tw_h_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_h_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_h_rsc_ARID : IN STD_LOGIC;
    tw_h_rsc_BREADY : IN STD_LOGIC;
    tw_h_rsc_BVALID : OUT STD_LOGIC;
    tw_h_rsc_BUSER : OUT STD_LOGIC;
    tw_h_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_BID : OUT STD_LOGIC;
    tw_h_rsc_WREADY : OUT STD_LOGIC;
    tw_h_rsc_WVALID : IN STD_LOGIC;
    tw_h_rsc_WUSER : IN STD_LOGIC;
    tw_h_rsc_WLAST : IN STD_LOGIC;
    tw_h_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_h_rsc_AWREADY : OUT STD_LOGIC;
    tw_h_rsc_AWVALID : IN STD_LOGIC;
    tw_h_rsc_AWUSER : IN STD_LOGIC;
    tw_h_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWLOCK : IN STD_LOGIC;
    tw_h_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_h_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_h_rsc_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    tw_h_rsci_oswt : IN STD_LOGIC;
    tw_h_rsci_wen_comp : OUT STD_LOGIC;
    tw_h_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    tw_h_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0)
  );
END hybrid_core_tw_h_rsci;

ARCHITECTURE v14 OF hybrid_core_tw_h_rsci IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL tw_h_rsci_biwt : STD_LOGIC;
  SIGNAL tw_h_rsci_bdwt : STD_LOGIC;
  SIGNAL tw_h_rsci_bcwt : STD_LOGIC;
  SIGNAL tw_h_rsci_s_re_core_sct : STD_LOGIC;
  SIGNAL tw_h_rsci_s_raddr : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_h_rsci_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_h_rsci_s_rrdy : STD_LOGIC;
  SIGNAL tw_h_rsci_s_wrdy : STD_LOGIC;
  SIGNAL tw_h_rsc_is_idle : STD_LOGIC;
  SIGNAL tw_h_rsci_s_din_mxwt_pconst : STD_LOGIC_VECTOR (19 DOWNTO 0);

  SIGNAL tw_h_rsci_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL tw_h_rsci_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL tw_h_rsci_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_h_rsci_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_h_rsci_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_h_rsci_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_h_rsci_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_h_rsci_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL tw_h_rsci_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL tw_h_rsci_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_h_rsci_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_h_rsci_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_h_rsci_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_h_rsci_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_h_rsci_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_h_rsci_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_h_rsci_s_raddr_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_h_rsci_s_waddr : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_h_rsci_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_h_rsci_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      tw_h_rsci_oswt : IN STD_LOGIC;
      tw_h_rsci_biwt : OUT STD_LOGIC;
      tw_h_rsci_bdwt : OUT STD_LOGIC;
      tw_h_rsci_bcwt : IN STD_LOGIC;
      tw_h_rsci_s_re_core_sct : OUT STD_LOGIC;
      tw_h_rsci_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      tw_h_rsci_oswt : IN STD_LOGIC;
      tw_h_rsci_wen_comp : OUT STD_LOGIC;
      tw_h_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      tw_h_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
      tw_h_rsci_biwt : IN STD_LOGIC;
      tw_h_rsci_bdwt : IN STD_LOGIC;
      tw_h_rsci_bcwt : OUT STD_LOGIC;
      tw_h_rsci_s_raddr : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      tw_h_rsci_s_raddr_core_sct : IN STD_LOGIC;
      tw_h_rsci_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_raddr_core : STD_LOGIC_VECTOR
      (9 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_din_mxwt : STD_LOGIC_VECTOR
      (19 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_raddr : STD_LOGIC_VECTOR
      (9 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  tw_h_rsci : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 1024,
      op_width => 32,
      cwidth => 32,
      addr_w => 10,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => tw_h_rsci_AWID,
      AWADDR => tw_h_rsci_AWADDR,
      AWLEN => tw_h_rsci_AWLEN,
      AWSIZE => tw_h_rsci_AWSIZE,
      AWBURST => tw_h_rsci_AWBURST,
      AWLOCK => tw_h_rsc_AWLOCK,
      AWCACHE => tw_h_rsci_AWCACHE,
      AWPROT => tw_h_rsci_AWPROT,
      AWQOS => tw_h_rsci_AWQOS,
      AWREGION => tw_h_rsci_AWREGION,
      AWUSER => tw_h_rsci_AWUSER,
      AWVALID => tw_h_rsc_AWVALID,
      AWREADY => tw_h_rsc_AWREADY,
      WDATA => tw_h_rsci_WDATA,
      WSTRB => tw_h_rsci_WSTRB,
      WLAST => tw_h_rsc_WLAST,
      WUSER => tw_h_rsci_WUSER,
      WVALID => tw_h_rsc_WVALID,
      WREADY => tw_h_rsc_WREADY,
      BID => tw_h_rsci_BID,
      BRESP => tw_h_rsci_BRESP,
      BUSER => tw_h_rsci_BUSER,
      BVALID => tw_h_rsc_BVALID,
      BREADY => tw_h_rsc_BREADY,
      ARID => tw_h_rsci_ARID,
      ARADDR => tw_h_rsci_ARADDR,
      ARLEN => tw_h_rsci_ARLEN,
      ARSIZE => tw_h_rsci_ARSIZE,
      ARBURST => tw_h_rsci_ARBURST,
      ARLOCK => tw_h_rsc_ARLOCK,
      ARCACHE => tw_h_rsci_ARCACHE,
      ARPROT => tw_h_rsci_ARPROT,
      ARQOS => tw_h_rsci_ARQOS,
      ARREGION => tw_h_rsci_ARREGION,
      ARUSER => tw_h_rsci_ARUSER,
      ARVALID => tw_h_rsc_ARVALID,
      ARREADY => tw_h_rsc_ARREADY,
      RID => tw_h_rsci_RID,
      RDATA => tw_h_rsci_RDATA,
      RRESP => tw_h_rsci_RRESP,
      RLAST => tw_h_rsc_RLAST,
      RUSER => tw_h_rsci_RUSER,
      RVALID => tw_h_rsc_RVALID,
      RREADY => tw_h_rsc_RREADY,
      s_re => tw_h_rsci_s_re_core_sct,
      s_we => '0',
      s_raddr => tw_h_rsci_s_raddr_1,
      s_waddr => tw_h_rsci_s_waddr,
      s_din => tw_h_rsci_s_din_1,
      s_dout => tw_h_rsci_s_dout,
      s_rrdy => tw_h_rsci_s_rrdy,
      s_wrdy => tw_h_rsci_s_wrdy,
      is_idle => tw_h_rsc_is_idle,
      tr_write_done => tw_h_rsc_tr_write_done,
      s_tdone => tw_h_rsc_s_tdone
    );
  tw_h_rsci_AWID(0) <= tw_h_rsc_AWID;
  tw_h_rsci_AWADDR <= tw_h_rsc_AWADDR;
  tw_h_rsci_AWLEN <= tw_h_rsc_AWLEN;
  tw_h_rsci_AWSIZE <= tw_h_rsc_AWSIZE;
  tw_h_rsci_AWBURST <= tw_h_rsc_AWBURST;
  tw_h_rsci_AWCACHE <= tw_h_rsc_AWCACHE;
  tw_h_rsci_AWPROT <= tw_h_rsc_AWPROT;
  tw_h_rsci_AWQOS <= tw_h_rsc_AWQOS;
  tw_h_rsci_AWREGION <= tw_h_rsc_AWREGION;
  tw_h_rsci_AWUSER(0) <= tw_h_rsc_AWUSER;
  tw_h_rsci_WDATA <= tw_h_rsc_WDATA;
  tw_h_rsci_WSTRB <= tw_h_rsc_WSTRB;
  tw_h_rsci_WUSER(0) <= tw_h_rsc_WUSER;
  tw_h_rsc_BID <= tw_h_rsci_BID(0);
  tw_h_rsc_BRESP <= tw_h_rsci_BRESP;
  tw_h_rsc_BUSER <= tw_h_rsci_BUSER(0);
  tw_h_rsci_ARID(0) <= tw_h_rsc_ARID;
  tw_h_rsci_ARADDR <= tw_h_rsc_ARADDR;
  tw_h_rsci_ARLEN <= tw_h_rsc_ARLEN;
  tw_h_rsci_ARSIZE <= tw_h_rsc_ARSIZE;
  tw_h_rsci_ARBURST <= tw_h_rsc_ARBURST;
  tw_h_rsci_ARCACHE <= tw_h_rsc_ARCACHE;
  tw_h_rsci_ARPROT <= tw_h_rsc_ARPROT;
  tw_h_rsci_ARQOS <= tw_h_rsc_ARQOS;
  tw_h_rsci_ARREGION <= tw_h_rsc_ARREGION;
  tw_h_rsci_ARUSER(0) <= tw_h_rsc_ARUSER;
  tw_h_rsc_RID <= tw_h_rsci_RID(0);
  tw_h_rsc_RDATA <= tw_h_rsci_RDATA;
  tw_h_rsc_RRESP <= tw_h_rsci_RRESP;
  tw_h_rsc_RUSER <= tw_h_rsci_RUSER(0);
  tw_h_rsci_s_raddr_1 <= tw_h_rsci_s_raddr;
  tw_h_rsci_s_waddr <= STD_LOGIC_VECTOR'( "0000000000");
  tw_h_rsci_s_din <= tw_h_rsci_s_din_1;
  tw_h_rsci_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl_inst : hybrid_core_tw_h_rsci_tw_h_rsc_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      tw_h_rsci_oswt => tw_h_rsci_oswt,
      tw_h_rsci_biwt => tw_h_rsci_biwt,
      tw_h_rsci_bdwt => tw_h_rsci_bdwt,
      tw_h_rsci_bcwt => tw_h_rsci_bcwt,
      tw_h_rsci_s_re_core_sct => tw_h_rsci_s_re_core_sct,
      tw_h_rsci_s_rrdy => tw_h_rsci_s_rrdy
    );
  hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst : hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      tw_h_rsci_oswt => tw_h_rsci_oswt,
      tw_h_rsci_wen_comp => tw_h_rsci_wen_comp,
      tw_h_rsci_s_raddr_core => hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_raddr_core,
      tw_h_rsci_s_din_mxwt => hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_din_mxwt,
      tw_h_rsci_biwt => tw_h_rsci_biwt,
      tw_h_rsci_bdwt => tw_h_rsci_bdwt,
      tw_h_rsci_bcwt => tw_h_rsci_bcwt,
      tw_h_rsci_s_raddr => hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_raddr,
      tw_h_rsci_s_raddr_core_sct => tw_h_rsci_s_re_core_sct,
      tw_h_rsci_s_din => hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_din
    );
  hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_raddr_core <= tw_h_rsci_s_raddr_core;
  tw_h_rsci_s_din_mxwt_pconst <= hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_din_mxwt;
  tw_h_rsci_s_raddr <= hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_raddr;
  hybrid_core_tw_h_rsci_tw_h_rsc_wait_dp_inst_tw_h_rsci_s_din <= tw_h_rsci_s_din;

  tw_h_rsci_s_din_mxwt <= tw_h_rsci_s_din_mxwt_pconst;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_tw_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_tw_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    tw_rsc_s_tdone : IN STD_LOGIC;
    tw_rsc_tr_write_done : IN STD_LOGIC;
    tw_rsc_RREADY : IN STD_LOGIC;
    tw_rsc_RVALID : OUT STD_LOGIC;
    tw_rsc_RUSER : OUT STD_LOGIC;
    tw_rsc_RLAST : OUT STD_LOGIC;
    tw_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_rsc_RID : OUT STD_LOGIC;
    tw_rsc_ARREADY : OUT STD_LOGIC;
    tw_rsc_ARVALID : IN STD_LOGIC;
    tw_rsc_ARUSER : IN STD_LOGIC;
    tw_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARLOCK : IN STD_LOGIC;
    tw_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_rsc_ARID : IN STD_LOGIC;
    tw_rsc_BREADY : IN STD_LOGIC;
    tw_rsc_BVALID : OUT STD_LOGIC;
    tw_rsc_BUSER : OUT STD_LOGIC;
    tw_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_BID : OUT STD_LOGIC;
    tw_rsc_WREADY : OUT STD_LOGIC;
    tw_rsc_WVALID : IN STD_LOGIC;
    tw_rsc_WUSER : IN STD_LOGIC;
    tw_rsc_WLAST : IN STD_LOGIC;
    tw_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_rsc_AWREADY : OUT STD_LOGIC;
    tw_rsc_AWVALID : IN STD_LOGIC;
    tw_rsc_AWUSER : IN STD_LOGIC;
    tw_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWLOCK : IN STD_LOGIC;
    tw_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_rsc_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    tw_rsci_oswt : IN STD_LOGIC;
    tw_rsci_wen_comp : OUT STD_LOGIC;
    tw_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    tw_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0)
  );
END hybrid_core_tw_rsci;

ARCHITECTURE v14 OF hybrid_core_tw_rsci IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL tw_rsci_biwt : STD_LOGIC;
  SIGNAL tw_rsci_bdwt : STD_LOGIC;
  SIGNAL tw_rsci_bcwt : STD_LOGIC;
  SIGNAL tw_rsci_s_re_core_sct : STD_LOGIC;
  SIGNAL tw_rsci_s_raddr : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_rsci_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_rsci_s_rrdy : STD_LOGIC;
  SIGNAL tw_rsci_s_wrdy : STD_LOGIC;
  SIGNAL tw_rsc_is_idle : STD_LOGIC;
  SIGNAL tw_rsci_s_din_mxwt_pconst : STD_LOGIC_VECTOR (19 DOWNTO 0);

  SIGNAL tw_rsci_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL tw_rsci_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL tw_rsci_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_rsci_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_rsci_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_rsci_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_rsci_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_rsci_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL tw_rsci_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL tw_rsci_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_rsci_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_rsci_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL tw_rsci_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tw_rsci_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_rsci_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL tw_rsci_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL tw_rsci_s_raddr_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_rsci_s_waddr : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_rsci_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tw_rsci_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_tw_rsci_tw_rsc_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      tw_rsci_oswt : IN STD_LOGIC;
      tw_rsci_biwt : OUT STD_LOGIC;
      tw_rsci_bdwt : OUT STD_LOGIC;
      tw_rsci_bcwt : IN STD_LOGIC;
      tw_rsci_s_re_core_sct : OUT STD_LOGIC;
      tw_rsci_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_tw_rsci_tw_rsc_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      tw_rsci_oswt : IN STD_LOGIC;
      tw_rsci_wen_comp : OUT STD_LOGIC;
      tw_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      tw_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0);
      tw_rsci_biwt : IN STD_LOGIC;
      tw_rsci_bdwt : IN STD_LOGIC;
      tw_rsci_bcwt : OUT STD_LOGIC;
      tw_rsci_s_raddr : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      tw_rsci_s_raddr_core_sct : IN STD_LOGIC;
      tw_rsci_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_raddr_core : STD_LOGIC_VECTOR
      (9 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_din_mxwt : STD_LOGIC_VECTOR
      (19 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_raddr : STD_LOGIC_VECTOR
      (9 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  tw_rsci : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 1024,
      op_width => 32,
      cwidth => 32,
      addr_w => 10,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => tw_rsci_AWID,
      AWADDR => tw_rsci_AWADDR,
      AWLEN => tw_rsci_AWLEN,
      AWSIZE => tw_rsci_AWSIZE,
      AWBURST => tw_rsci_AWBURST,
      AWLOCK => tw_rsc_AWLOCK,
      AWCACHE => tw_rsci_AWCACHE,
      AWPROT => tw_rsci_AWPROT,
      AWQOS => tw_rsci_AWQOS,
      AWREGION => tw_rsci_AWREGION,
      AWUSER => tw_rsci_AWUSER,
      AWVALID => tw_rsc_AWVALID,
      AWREADY => tw_rsc_AWREADY,
      WDATA => tw_rsci_WDATA,
      WSTRB => tw_rsci_WSTRB,
      WLAST => tw_rsc_WLAST,
      WUSER => tw_rsci_WUSER,
      WVALID => tw_rsc_WVALID,
      WREADY => tw_rsc_WREADY,
      BID => tw_rsci_BID,
      BRESP => tw_rsci_BRESP,
      BUSER => tw_rsci_BUSER,
      BVALID => tw_rsc_BVALID,
      BREADY => tw_rsc_BREADY,
      ARID => tw_rsci_ARID,
      ARADDR => tw_rsci_ARADDR,
      ARLEN => tw_rsci_ARLEN,
      ARSIZE => tw_rsci_ARSIZE,
      ARBURST => tw_rsci_ARBURST,
      ARLOCK => tw_rsc_ARLOCK,
      ARCACHE => tw_rsci_ARCACHE,
      ARPROT => tw_rsci_ARPROT,
      ARQOS => tw_rsci_ARQOS,
      ARREGION => tw_rsci_ARREGION,
      ARUSER => tw_rsci_ARUSER,
      ARVALID => tw_rsc_ARVALID,
      ARREADY => tw_rsc_ARREADY,
      RID => tw_rsci_RID,
      RDATA => tw_rsci_RDATA,
      RRESP => tw_rsci_RRESP,
      RLAST => tw_rsc_RLAST,
      RUSER => tw_rsci_RUSER,
      RVALID => tw_rsc_RVALID,
      RREADY => tw_rsc_RREADY,
      s_re => tw_rsci_s_re_core_sct,
      s_we => '0',
      s_raddr => tw_rsci_s_raddr_1,
      s_waddr => tw_rsci_s_waddr,
      s_din => tw_rsci_s_din_1,
      s_dout => tw_rsci_s_dout,
      s_rrdy => tw_rsci_s_rrdy,
      s_wrdy => tw_rsci_s_wrdy,
      is_idle => tw_rsc_is_idle,
      tr_write_done => tw_rsc_tr_write_done,
      s_tdone => tw_rsc_s_tdone
    );
  tw_rsci_AWID(0) <= tw_rsc_AWID;
  tw_rsci_AWADDR <= tw_rsc_AWADDR;
  tw_rsci_AWLEN <= tw_rsc_AWLEN;
  tw_rsci_AWSIZE <= tw_rsc_AWSIZE;
  tw_rsci_AWBURST <= tw_rsc_AWBURST;
  tw_rsci_AWCACHE <= tw_rsc_AWCACHE;
  tw_rsci_AWPROT <= tw_rsc_AWPROT;
  tw_rsci_AWQOS <= tw_rsc_AWQOS;
  tw_rsci_AWREGION <= tw_rsc_AWREGION;
  tw_rsci_AWUSER(0) <= tw_rsc_AWUSER;
  tw_rsci_WDATA <= tw_rsc_WDATA;
  tw_rsci_WSTRB <= tw_rsc_WSTRB;
  tw_rsci_WUSER(0) <= tw_rsc_WUSER;
  tw_rsc_BID <= tw_rsci_BID(0);
  tw_rsc_BRESP <= tw_rsci_BRESP;
  tw_rsc_BUSER <= tw_rsci_BUSER(0);
  tw_rsci_ARID(0) <= tw_rsc_ARID;
  tw_rsci_ARADDR <= tw_rsc_ARADDR;
  tw_rsci_ARLEN <= tw_rsc_ARLEN;
  tw_rsci_ARSIZE <= tw_rsc_ARSIZE;
  tw_rsci_ARBURST <= tw_rsc_ARBURST;
  tw_rsci_ARCACHE <= tw_rsc_ARCACHE;
  tw_rsci_ARPROT <= tw_rsc_ARPROT;
  tw_rsci_ARQOS <= tw_rsc_ARQOS;
  tw_rsci_ARREGION <= tw_rsc_ARREGION;
  tw_rsci_ARUSER(0) <= tw_rsc_ARUSER;
  tw_rsc_RID <= tw_rsci_RID(0);
  tw_rsc_RDATA <= tw_rsci_RDATA;
  tw_rsc_RRESP <= tw_rsci_RRESP;
  tw_rsc_RUSER <= tw_rsci_RUSER(0);
  tw_rsci_s_raddr_1 <= tw_rsci_s_raddr;
  tw_rsci_s_waddr <= STD_LOGIC_VECTOR'( "0000000000");
  tw_rsci_s_din <= tw_rsci_s_din_1;
  tw_rsci_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  hybrid_core_tw_rsci_tw_rsc_wait_ctrl_inst : hybrid_core_tw_rsci_tw_rsc_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      tw_rsci_oswt => tw_rsci_oswt,
      tw_rsci_biwt => tw_rsci_biwt,
      tw_rsci_bdwt => tw_rsci_bdwt,
      tw_rsci_bcwt => tw_rsci_bcwt,
      tw_rsci_s_re_core_sct => tw_rsci_s_re_core_sct,
      tw_rsci_s_rrdy => tw_rsci_s_rrdy
    );
  hybrid_core_tw_rsci_tw_rsc_wait_dp_inst : hybrid_core_tw_rsci_tw_rsc_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      tw_rsci_oswt => tw_rsci_oswt,
      tw_rsci_wen_comp => tw_rsci_wen_comp,
      tw_rsci_s_raddr_core => hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_raddr_core,
      tw_rsci_s_din_mxwt => hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_din_mxwt,
      tw_rsci_biwt => tw_rsci_biwt,
      tw_rsci_bdwt => tw_rsci_bdwt,
      tw_rsci_bcwt => tw_rsci_bcwt,
      tw_rsci_s_raddr => hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_raddr,
      tw_rsci_s_raddr_core_sct => tw_rsci_s_re_core_sct,
      tw_rsci_s_din => hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_din
    );
  hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_raddr_core <= tw_rsci_s_raddr_core;
  tw_rsci_s_din_mxwt_pconst <= hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_din_mxwt;
  tw_rsci_s_raddr <= hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_raddr;
  hybrid_core_tw_rsci_tw_rsc_wait_dp_inst_tw_rsci_s_din <= tw_rsci_s_din;

  tw_rsci_s_din_mxwt <= tw_rsci_s_din_mxwt_pconst;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_revArr_rsci
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_revArr_rsci IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    revArr_rsc_s_tdone : IN STD_LOGIC;
    revArr_rsc_tr_write_done : IN STD_LOGIC;
    revArr_rsc_RREADY : IN STD_LOGIC;
    revArr_rsc_RVALID : OUT STD_LOGIC;
    revArr_rsc_RUSER : OUT STD_LOGIC;
    revArr_rsc_RLAST : OUT STD_LOGIC;
    revArr_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    revArr_rsc_RID : OUT STD_LOGIC;
    revArr_rsc_ARREADY : OUT STD_LOGIC;
    revArr_rsc_ARVALID : IN STD_LOGIC;
    revArr_rsc_ARUSER : IN STD_LOGIC;
    revArr_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARLOCK : IN STD_LOGIC;
    revArr_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    revArr_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    revArr_rsc_ARID : IN STD_LOGIC;
    revArr_rsc_BREADY : IN STD_LOGIC;
    revArr_rsc_BVALID : OUT STD_LOGIC;
    revArr_rsc_BUSER : OUT STD_LOGIC;
    revArr_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_BID : OUT STD_LOGIC;
    revArr_rsc_WREADY : OUT STD_LOGIC;
    revArr_rsc_WVALID : IN STD_LOGIC;
    revArr_rsc_WUSER : IN STD_LOGIC;
    revArr_rsc_WLAST : IN STD_LOGIC;
    revArr_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    revArr_rsc_AWREADY : OUT STD_LOGIC;
    revArr_rsc_AWVALID : IN STD_LOGIC;
    revArr_rsc_AWUSER : IN STD_LOGIC;
    revArr_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWLOCK : IN STD_LOGIC;
    revArr_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    revArr_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    revArr_rsc_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    revArr_rsci_oswt : IN STD_LOGIC;
    revArr_rsci_wen_comp : OUT STD_LOGIC;
    revArr_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    revArr_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
  );
END hybrid_core_revArr_rsci;

ARCHITECTURE v14 OF hybrid_core_revArr_rsci IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL revArr_rsci_biwt : STD_LOGIC;
  SIGNAL revArr_rsci_bdwt : STD_LOGIC;
  SIGNAL revArr_rsci_bcwt : STD_LOGIC;
  SIGNAL revArr_rsci_s_re_core_sct : STD_LOGIC;
  SIGNAL revArr_rsci_s_raddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL revArr_rsci_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL revArr_rsci_s_rrdy : STD_LOGIC;
  SIGNAL revArr_rsci_s_wrdy : STD_LOGIC;
  SIGNAL revArr_rsc_is_idle : STD_LOGIC;
  SIGNAL revArr_rsci_s_din_mxwt_pconst : STD_LOGIC_VECTOR (9 DOWNTO 0);

  SIGNAL revArr_rsci_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL revArr_rsci_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL revArr_rsci_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL revArr_rsci_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL revArr_rsci_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL revArr_rsci_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL revArr_rsci_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL revArr_rsci_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL revArr_rsci_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL revArr_rsci_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL revArr_rsci_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL revArr_rsci_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL revArr_rsci_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL revArr_rsci_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL revArr_rsci_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL revArr_rsci_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL revArr_rsci_s_raddr_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL revArr_rsci_s_waddr : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL revArr_rsci_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL revArr_rsci_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      revArr_rsci_oswt : IN STD_LOGIC;
      revArr_rsci_biwt : OUT STD_LOGIC;
      revArr_rsci_bdwt : OUT STD_LOGIC;
      revArr_rsci_bcwt : IN STD_LOGIC;
      revArr_rsci_s_re_core_sct : OUT STD_LOGIC;
      revArr_rsci_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_revArr_rsci_revArr_rsc_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      revArr_rsci_oswt : IN STD_LOGIC;
      revArr_rsci_wen_comp : OUT STD_LOGIC;
      revArr_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      revArr_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      revArr_rsci_biwt : IN STD_LOGIC;
      revArr_rsci_bdwt : IN STD_LOGIC;
      revArr_rsci_bcwt : OUT STD_LOGIC;
      revArr_rsci_s_raddr : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      revArr_rsci_s_raddr_core_sct : IN STD_LOGIC;
      revArr_rsci_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_raddr_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_din_mxwt :
      STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_raddr : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_din : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

BEGIN
  revArr_rsci : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 32,
      op_width => 20,
      cwidth => 32,
      addr_w => 5,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => revArr_rsci_AWID,
      AWADDR => revArr_rsci_AWADDR,
      AWLEN => revArr_rsci_AWLEN,
      AWSIZE => revArr_rsci_AWSIZE,
      AWBURST => revArr_rsci_AWBURST,
      AWLOCK => revArr_rsc_AWLOCK,
      AWCACHE => revArr_rsci_AWCACHE,
      AWPROT => revArr_rsci_AWPROT,
      AWQOS => revArr_rsci_AWQOS,
      AWREGION => revArr_rsci_AWREGION,
      AWUSER => revArr_rsci_AWUSER,
      AWVALID => revArr_rsc_AWVALID,
      AWREADY => revArr_rsc_AWREADY,
      WDATA => revArr_rsci_WDATA,
      WSTRB => revArr_rsci_WSTRB,
      WLAST => revArr_rsc_WLAST,
      WUSER => revArr_rsci_WUSER,
      WVALID => revArr_rsc_WVALID,
      WREADY => revArr_rsc_WREADY,
      BID => revArr_rsci_BID,
      BRESP => revArr_rsci_BRESP,
      BUSER => revArr_rsci_BUSER,
      BVALID => revArr_rsc_BVALID,
      BREADY => revArr_rsc_BREADY,
      ARID => revArr_rsci_ARID,
      ARADDR => revArr_rsci_ARADDR,
      ARLEN => revArr_rsci_ARLEN,
      ARSIZE => revArr_rsci_ARSIZE,
      ARBURST => revArr_rsci_ARBURST,
      ARLOCK => revArr_rsc_ARLOCK,
      ARCACHE => revArr_rsci_ARCACHE,
      ARPROT => revArr_rsci_ARPROT,
      ARQOS => revArr_rsci_ARQOS,
      ARREGION => revArr_rsci_ARREGION,
      ARUSER => revArr_rsci_ARUSER,
      ARVALID => revArr_rsc_ARVALID,
      ARREADY => revArr_rsc_ARREADY,
      RID => revArr_rsci_RID,
      RDATA => revArr_rsci_RDATA,
      RRESP => revArr_rsci_RRESP,
      RLAST => revArr_rsc_RLAST,
      RUSER => revArr_rsci_RUSER,
      RVALID => revArr_rsc_RVALID,
      RREADY => revArr_rsc_RREADY,
      s_re => revArr_rsci_s_re_core_sct,
      s_we => '0',
      s_raddr => revArr_rsci_s_raddr_1,
      s_waddr => revArr_rsci_s_waddr,
      s_din => revArr_rsci_s_din_1,
      s_dout => revArr_rsci_s_dout,
      s_rrdy => revArr_rsci_s_rrdy,
      s_wrdy => revArr_rsci_s_wrdy,
      is_idle => revArr_rsc_is_idle,
      tr_write_done => revArr_rsc_tr_write_done,
      s_tdone => revArr_rsc_s_tdone
    );
  revArr_rsci_AWID(0) <= revArr_rsc_AWID;
  revArr_rsci_AWADDR <= revArr_rsc_AWADDR;
  revArr_rsci_AWLEN <= revArr_rsc_AWLEN;
  revArr_rsci_AWSIZE <= revArr_rsc_AWSIZE;
  revArr_rsci_AWBURST <= revArr_rsc_AWBURST;
  revArr_rsci_AWCACHE <= revArr_rsc_AWCACHE;
  revArr_rsci_AWPROT <= revArr_rsc_AWPROT;
  revArr_rsci_AWQOS <= revArr_rsc_AWQOS;
  revArr_rsci_AWREGION <= revArr_rsc_AWREGION;
  revArr_rsci_AWUSER(0) <= revArr_rsc_AWUSER;
  revArr_rsci_WDATA <= revArr_rsc_WDATA;
  revArr_rsci_WSTRB <= revArr_rsc_WSTRB;
  revArr_rsci_WUSER(0) <= revArr_rsc_WUSER;
  revArr_rsc_BID <= revArr_rsci_BID(0);
  revArr_rsc_BRESP <= revArr_rsci_BRESP;
  revArr_rsc_BUSER <= revArr_rsci_BUSER(0);
  revArr_rsci_ARID(0) <= revArr_rsc_ARID;
  revArr_rsci_ARADDR <= revArr_rsc_ARADDR;
  revArr_rsci_ARLEN <= revArr_rsc_ARLEN;
  revArr_rsci_ARSIZE <= revArr_rsc_ARSIZE;
  revArr_rsci_ARBURST <= revArr_rsc_ARBURST;
  revArr_rsci_ARCACHE <= revArr_rsc_ARCACHE;
  revArr_rsci_ARPROT <= revArr_rsc_ARPROT;
  revArr_rsci_ARQOS <= revArr_rsc_ARQOS;
  revArr_rsci_ARREGION <= revArr_rsc_ARREGION;
  revArr_rsci_ARUSER(0) <= revArr_rsc_ARUSER;
  revArr_rsc_RID <= revArr_rsci_RID(0);
  revArr_rsc_RDATA <= revArr_rsci_RDATA;
  revArr_rsc_RRESP <= revArr_rsci_RRESP;
  revArr_rsc_RUSER <= revArr_rsci_RUSER(0);
  revArr_rsci_s_raddr_1 <= revArr_rsci_s_raddr;
  revArr_rsci_s_waddr <= STD_LOGIC_VECTOR'( "00000");
  revArr_rsci_s_din <= revArr_rsci_s_din_1;
  revArr_rsci_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl_inst : hybrid_core_revArr_rsci_revArr_rsc_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      revArr_rsci_oswt => revArr_rsci_oswt,
      revArr_rsci_biwt => revArr_rsci_biwt,
      revArr_rsci_bdwt => revArr_rsci_bdwt,
      revArr_rsci_bcwt => revArr_rsci_bcwt,
      revArr_rsci_s_re_core_sct => revArr_rsci_s_re_core_sct,
      revArr_rsci_s_rrdy => revArr_rsci_s_rrdy
    );
  hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst : hybrid_core_revArr_rsci_revArr_rsc_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      revArr_rsci_oswt => revArr_rsci_oswt,
      revArr_rsci_wen_comp => revArr_rsci_wen_comp,
      revArr_rsci_s_raddr_core => hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_raddr_core,
      revArr_rsci_s_din_mxwt => hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_din_mxwt,
      revArr_rsci_biwt => revArr_rsci_biwt,
      revArr_rsci_bdwt => revArr_rsci_bdwt,
      revArr_rsci_bcwt => revArr_rsci_bcwt,
      revArr_rsci_s_raddr => hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_raddr,
      revArr_rsci_s_raddr_core_sct => revArr_rsci_s_re_core_sct,
      revArr_rsci_s_din => hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_din
    );
  hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_raddr_core <= revArr_rsci_s_raddr_core;
  revArr_rsci_s_din_mxwt_pconst <= hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_din_mxwt;
  revArr_rsci_s_raddr <= hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_raddr;
  hybrid_core_revArr_rsci_revArr_rsc_wait_dp_inst_revArr_rsci_s_din <= revArr_rsci_s_din;

  revArr_rsci_s_din_mxwt <= revArr_rsci_s_din_mxwt_pconst;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_h_rsci_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_h_rsci_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_h_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsci_oswt : IN STD_LOGIC;
    twiddle_h_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_h_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsci_oswt_pff : IN STD_LOGIC
  );
END hybrid_core_twiddle_h_rsci_1;

ARCHITECTURE v14 OF hybrid_core_twiddle_h_rsci_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsci_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsci_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsci_adrb_d_reg : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_h_rsci_adrb_d_core_sct_iff : STD_LOGIC;

  COMPONENT hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsci_oswt : IN STD_LOGIC;
      twiddle_h_rsci_biwt : OUT STD_LOGIC;
      twiddle_h_rsci_bdwt : OUT STD_LOGIC;
      twiddle_h_rsci_adrb_d_core_sct_pff : OUT STD_LOGIC;
      twiddle_h_rsci_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_h_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_h_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsci_biwt : IN STD_LOGIC;
      twiddle_h_rsci_bdwt : IN STD_LOGIC;
      twiddle_h_rsci_adrb_d_core_sct : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_adrb_d
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_qb_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_adrb_d_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl_inst : hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsci_oswt => twiddle_h_rsci_oswt,
      twiddle_h_rsci_biwt => twiddle_h_rsci_biwt,
      twiddle_h_rsci_bdwt => twiddle_h_rsci_bdwt,
      twiddle_h_rsci_adrb_d_core_sct_pff => twiddle_h_rsci_adrb_d_core_sct_iff,
      twiddle_h_rsci_oswt_pff => twiddle_h_rsci_oswt_pff
    );
  hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst : hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsci_adrb_d => hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_adrb_d,
      twiddle_h_rsci_qb_d => hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_qb_d,
      twiddle_h_rsci_adrb_d_core => hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_adrb_d_core,
      twiddle_h_rsci_qb_d_mxwt => hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_qb_d_mxwt,
      twiddle_h_rsci_biwt => twiddle_h_rsci_biwt,
      twiddle_h_rsci_bdwt => twiddle_h_rsci_bdwt,
      twiddle_h_rsci_adrb_d_core_sct => twiddle_h_rsci_adrb_d_core_sct_iff
    );
  twiddle_h_rsci_adrb_d_reg <= hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_adrb_d;
  hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_qb_d <=
      twiddle_h_rsci_qb_d;
  hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_adrb_d_core
      <= '0' & (twiddle_h_rsci_adrb_d_core(3 DOWNTO 0));
  twiddle_h_rsci_qb_d_mxwt <= hybrid_core_twiddle_h_rsci_1_twiddle_h_rsc_wait_dp_inst_twiddle_h_rsci_qb_d_mxwt;

  twiddle_h_rsci_adrb_d <= twiddle_h_rsci_adrb_d_reg;
  twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsci_adrb_d_core_sct_iff;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core_twiddle_rsci_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core_twiddle_rsci_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsci_oswt : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsci_oswt_pff : IN STD_LOGIC
  );
END hybrid_core_twiddle_rsci_1;

ARCHITECTURE v14 OF hybrid_core_twiddle_rsci_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsci_biwt : STD_LOGIC;
  SIGNAL twiddle_rsci_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsci_adrb_d_reg : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsci_adrb_d_core_sct_iff : STD_LOGIC;

  COMPONENT hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsci_oswt : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsci_biwt : OUT STD_LOGIC;
      twiddle_rsci_bdwt : OUT STD_LOGIC;
      twiddle_rsci_adrb_d_core_sct_pff : OUT STD_LOGIC;
      twiddle_rsci_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsci_biwt : IN STD_LOGIC;
      twiddle_rsci_bdwt : IN STD_LOGIC;
      twiddle_rsci_adrb_d_core_sct : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_adrb_d
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_qb_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_adrb_d_core
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_qb_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl_inst : hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsci_oswt => twiddle_rsci_oswt,
      core_wten => core_wten,
      twiddle_rsci_biwt => twiddle_rsci_biwt,
      twiddle_rsci_bdwt => twiddle_rsci_bdwt,
      twiddle_rsci_adrb_d_core_sct_pff => twiddle_rsci_adrb_d_core_sct_iff,
      twiddle_rsci_oswt_pff => twiddle_rsci_oswt_pff
    );
  hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst : hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsci_adrb_d => hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_adrb_d,
      twiddle_rsci_qb_d => hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_qb_d,
      twiddle_rsci_adrb_d_core => hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_adrb_d_core,
      twiddle_rsci_qb_d_mxwt => hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_qb_d_mxwt,
      twiddle_rsci_biwt => twiddle_rsci_biwt,
      twiddle_rsci_bdwt => twiddle_rsci_bdwt,
      twiddle_rsci_adrb_d_core_sct => twiddle_rsci_adrb_d_core_sct_iff
    );
  twiddle_rsci_adrb_d_reg <= hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_adrb_d;
  hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_qb_d <= twiddle_rsci_qb_d;
  hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_adrb_d_core <=
      '0' & (twiddle_rsci_adrb_d_core(3 DOWNTO 0));
  twiddle_rsci_qb_d_mxwt <= hybrid_core_twiddle_rsci_1_twiddle_rsc_wait_dp_inst_twiddle_rsci_qb_d_mxwt;

  twiddle_rsci_adrb_d <= twiddle_rsci_adrb_d_reg;
  twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsci_adrb_d_core_sct_iff;
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_0_0_s_tdone : IN STD_LOGIC;
    x_rsc_0_0_tr_write_done : IN STD_LOGIC;
    x_rsc_0_0_RREADY : IN STD_LOGIC;
    x_rsc_0_0_RVALID : OUT STD_LOGIC;
    x_rsc_0_0_RUSER : OUT STD_LOGIC;
    x_rsc_0_0_RLAST : OUT STD_LOGIC;
    x_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_RID : OUT STD_LOGIC;
    x_rsc_0_0_ARREADY : OUT STD_LOGIC;
    x_rsc_0_0_ARVALID : IN STD_LOGIC;
    x_rsc_0_0_ARUSER : IN STD_LOGIC;
    x_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARLOCK : IN STD_LOGIC;
    x_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_0_0_ARID : IN STD_LOGIC;
    x_rsc_0_0_BREADY : IN STD_LOGIC;
    x_rsc_0_0_BVALID : OUT STD_LOGIC;
    x_rsc_0_0_BUSER : OUT STD_LOGIC;
    x_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_BID : OUT STD_LOGIC;
    x_rsc_0_0_WREADY : OUT STD_LOGIC;
    x_rsc_0_0_WVALID : IN STD_LOGIC;
    x_rsc_0_0_WUSER : IN STD_LOGIC;
    x_rsc_0_0_WLAST : IN STD_LOGIC;
    x_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_AWREADY : OUT STD_LOGIC;
    x_rsc_0_0_AWVALID : IN STD_LOGIC;
    x_rsc_0_0_AWUSER : IN STD_LOGIC;
    x_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWLOCK : IN STD_LOGIC;
    x_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_0_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    x_rsc_1_0_s_tdone : IN STD_LOGIC;
    x_rsc_1_0_tr_write_done : IN STD_LOGIC;
    x_rsc_1_0_RREADY : IN STD_LOGIC;
    x_rsc_1_0_RVALID : OUT STD_LOGIC;
    x_rsc_1_0_RUSER : OUT STD_LOGIC;
    x_rsc_1_0_RLAST : OUT STD_LOGIC;
    x_rsc_1_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_RID : OUT STD_LOGIC;
    x_rsc_1_0_ARREADY : OUT STD_LOGIC;
    x_rsc_1_0_ARVALID : IN STD_LOGIC;
    x_rsc_1_0_ARUSER : IN STD_LOGIC;
    x_rsc_1_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARLOCK : IN STD_LOGIC;
    x_rsc_1_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_1_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_1_0_ARID : IN STD_LOGIC;
    x_rsc_1_0_BREADY : IN STD_LOGIC;
    x_rsc_1_0_BVALID : OUT STD_LOGIC;
    x_rsc_1_0_BUSER : OUT STD_LOGIC;
    x_rsc_1_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_BID : OUT STD_LOGIC;
    x_rsc_1_0_WREADY : OUT STD_LOGIC;
    x_rsc_1_0_WVALID : IN STD_LOGIC;
    x_rsc_1_0_WUSER : IN STD_LOGIC;
    x_rsc_1_0_WLAST : IN STD_LOGIC;
    x_rsc_1_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_AWREADY : OUT STD_LOGIC;
    x_rsc_1_0_AWVALID : IN STD_LOGIC;
    x_rsc_1_0_AWUSER : IN STD_LOGIC;
    x_rsc_1_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWLOCK : IN STD_LOGIC;
    x_rsc_1_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_1_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_1_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    x_rsc_2_0_s_tdone : IN STD_LOGIC;
    x_rsc_2_0_tr_write_done : IN STD_LOGIC;
    x_rsc_2_0_RREADY : IN STD_LOGIC;
    x_rsc_2_0_RVALID : OUT STD_LOGIC;
    x_rsc_2_0_RUSER : OUT STD_LOGIC;
    x_rsc_2_0_RLAST : OUT STD_LOGIC;
    x_rsc_2_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_RID : OUT STD_LOGIC;
    x_rsc_2_0_ARREADY : OUT STD_LOGIC;
    x_rsc_2_0_ARVALID : IN STD_LOGIC;
    x_rsc_2_0_ARUSER : IN STD_LOGIC;
    x_rsc_2_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARLOCK : IN STD_LOGIC;
    x_rsc_2_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_2_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_2_0_ARID : IN STD_LOGIC;
    x_rsc_2_0_BREADY : IN STD_LOGIC;
    x_rsc_2_0_BVALID : OUT STD_LOGIC;
    x_rsc_2_0_BUSER : OUT STD_LOGIC;
    x_rsc_2_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_BID : OUT STD_LOGIC;
    x_rsc_2_0_WREADY : OUT STD_LOGIC;
    x_rsc_2_0_WVALID : IN STD_LOGIC;
    x_rsc_2_0_WUSER : IN STD_LOGIC;
    x_rsc_2_0_WLAST : IN STD_LOGIC;
    x_rsc_2_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_AWREADY : OUT STD_LOGIC;
    x_rsc_2_0_AWVALID : IN STD_LOGIC;
    x_rsc_2_0_AWUSER : IN STD_LOGIC;
    x_rsc_2_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWLOCK : IN STD_LOGIC;
    x_rsc_2_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_2_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_2_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_2_0_lz : OUT STD_LOGIC;
    x_rsc_3_0_s_tdone : IN STD_LOGIC;
    x_rsc_3_0_tr_write_done : IN STD_LOGIC;
    x_rsc_3_0_RREADY : IN STD_LOGIC;
    x_rsc_3_0_RVALID : OUT STD_LOGIC;
    x_rsc_3_0_RUSER : OUT STD_LOGIC;
    x_rsc_3_0_RLAST : OUT STD_LOGIC;
    x_rsc_3_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_RID : OUT STD_LOGIC;
    x_rsc_3_0_ARREADY : OUT STD_LOGIC;
    x_rsc_3_0_ARVALID : IN STD_LOGIC;
    x_rsc_3_0_ARUSER : IN STD_LOGIC;
    x_rsc_3_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARLOCK : IN STD_LOGIC;
    x_rsc_3_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_3_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_3_0_ARID : IN STD_LOGIC;
    x_rsc_3_0_BREADY : IN STD_LOGIC;
    x_rsc_3_0_BVALID : OUT STD_LOGIC;
    x_rsc_3_0_BUSER : OUT STD_LOGIC;
    x_rsc_3_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_BID : OUT STD_LOGIC;
    x_rsc_3_0_WREADY : OUT STD_LOGIC;
    x_rsc_3_0_WVALID : IN STD_LOGIC;
    x_rsc_3_0_WUSER : IN STD_LOGIC;
    x_rsc_3_0_WLAST : IN STD_LOGIC;
    x_rsc_3_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_AWREADY : OUT STD_LOGIC;
    x_rsc_3_0_AWVALID : IN STD_LOGIC;
    x_rsc_3_0_AWUSER : IN STD_LOGIC;
    x_rsc_3_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWLOCK : IN STD_LOGIC;
    x_rsc_3_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_3_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_3_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_3_0_lz : OUT STD_LOGIC;
    x_rsc_4_0_s_tdone : IN STD_LOGIC;
    x_rsc_4_0_tr_write_done : IN STD_LOGIC;
    x_rsc_4_0_RREADY : IN STD_LOGIC;
    x_rsc_4_0_RVALID : OUT STD_LOGIC;
    x_rsc_4_0_RUSER : OUT STD_LOGIC;
    x_rsc_4_0_RLAST : OUT STD_LOGIC;
    x_rsc_4_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_RID : OUT STD_LOGIC;
    x_rsc_4_0_ARREADY : OUT STD_LOGIC;
    x_rsc_4_0_ARVALID : IN STD_LOGIC;
    x_rsc_4_0_ARUSER : IN STD_LOGIC;
    x_rsc_4_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARLOCK : IN STD_LOGIC;
    x_rsc_4_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_4_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_4_0_ARID : IN STD_LOGIC;
    x_rsc_4_0_BREADY : IN STD_LOGIC;
    x_rsc_4_0_BVALID : OUT STD_LOGIC;
    x_rsc_4_0_BUSER : OUT STD_LOGIC;
    x_rsc_4_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_BID : OUT STD_LOGIC;
    x_rsc_4_0_WREADY : OUT STD_LOGIC;
    x_rsc_4_0_WVALID : IN STD_LOGIC;
    x_rsc_4_0_WUSER : IN STD_LOGIC;
    x_rsc_4_0_WLAST : IN STD_LOGIC;
    x_rsc_4_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_AWREADY : OUT STD_LOGIC;
    x_rsc_4_0_AWVALID : IN STD_LOGIC;
    x_rsc_4_0_AWUSER : IN STD_LOGIC;
    x_rsc_4_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWLOCK : IN STD_LOGIC;
    x_rsc_4_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_4_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_4_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_4_0_lz : OUT STD_LOGIC;
    x_rsc_5_0_s_tdone : IN STD_LOGIC;
    x_rsc_5_0_tr_write_done : IN STD_LOGIC;
    x_rsc_5_0_RREADY : IN STD_LOGIC;
    x_rsc_5_0_RVALID : OUT STD_LOGIC;
    x_rsc_5_0_RUSER : OUT STD_LOGIC;
    x_rsc_5_0_RLAST : OUT STD_LOGIC;
    x_rsc_5_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_RID : OUT STD_LOGIC;
    x_rsc_5_0_ARREADY : OUT STD_LOGIC;
    x_rsc_5_0_ARVALID : IN STD_LOGIC;
    x_rsc_5_0_ARUSER : IN STD_LOGIC;
    x_rsc_5_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARLOCK : IN STD_LOGIC;
    x_rsc_5_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_5_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_5_0_ARID : IN STD_LOGIC;
    x_rsc_5_0_BREADY : IN STD_LOGIC;
    x_rsc_5_0_BVALID : OUT STD_LOGIC;
    x_rsc_5_0_BUSER : OUT STD_LOGIC;
    x_rsc_5_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_BID : OUT STD_LOGIC;
    x_rsc_5_0_WREADY : OUT STD_LOGIC;
    x_rsc_5_0_WVALID : IN STD_LOGIC;
    x_rsc_5_0_WUSER : IN STD_LOGIC;
    x_rsc_5_0_WLAST : IN STD_LOGIC;
    x_rsc_5_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_AWREADY : OUT STD_LOGIC;
    x_rsc_5_0_AWVALID : IN STD_LOGIC;
    x_rsc_5_0_AWUSER : IN STD_LOGIC;
    x_rsc_5_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWLOCK : IN STD_LOGIC;
    x_rsc_5_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_5_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_5_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_5_0_lz : OUT STD_LOGIC;
    x_rsc_6_0_s_tdone : IN STD_LOGIC;
    x_rsc_6_0_tr_write_done : IN STD_LOGIC;
    x_rsc_6_0_RREADY : IN STD_LOGIC;
    x_rsc_6_0_RVALID : OUT STD_LOGIC;
    x_rsc_6_0_RUSER : OUT STD_LOGIC;
    x_rsc_6_0_RLAST : OUT STD_LOGIC;
    x_rsc_6_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_RID : OUT STD_LOGIC;
    x_rsc_6_0_ARREADY : OUT STD_LOGIC;
    x_rsc_6_0_ARVALID : IN STD_LOGIC;
    x_rsc_6_0_ARUSER : IN STD_LOGIC;
    x_rsc_6_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARLOCK : IN STD_LOGIC;
    x_rsc_6_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_6_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_6_0_ARID : IN STD_LOGIC;
    x_rsc_6_0_BREADY : IN STD_LOGIC;
    x_rsc_6_0_BVALID : OUT STD_LOGIC;
    x_rsc_6_0_BUSER : OUT STD_LOGIC;
    x_rsc_6_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_BID : OUT STD_LOGIC;
    x_rsc_6_0_WREADY : OUT STD_LOGIC;
    x_rsc_6_0_WVALID : IN STD_LOGIC;
    x_rsc_6_0_WUSER : IN STD_LOGIC;
    x_rsc_6_0_WLAST : IN STD_LOGIC;
    x_rsc_6_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_AWREADY : OUT STD_LOGIC;
    x_rsc_6_0_AWVALID : IN STD_LOGIC;
    x_rsc_6_0_AWUSER : IN STD_LOGIC;
    x_rsc_6_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWLOCK : IN STD_LOGIC;
    x_rsc_6_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_6_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_6_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_6_0_lz : OUT STD_LOGIC;
    x_rsc_7_0_s_tdone : IN STD_LOGIC;
    x_rsc_7_0_tr_write_done : IN STD_LOGIC;
    x_rsc_7_0_RREADY : IN STD_LOGIC;
    x_rsc_7_0_RVALID : OUT STD_LOGIC;
    x_rsc_7_0_RUSER : OUT STD_LOGIC;
    x_rsc_7_0_RLAST : OUT STD_LOGIC;
    x_rsc_7_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_RID : OUT STD_LOGIC;
    x_rsc_7_0_ARREADY : OUT STD_LOGIC;
    x_rsc_7_0_ARVALID : IN STD_LOGIC;
    x_rsc_7_0_ARUSER : IN STD_LOGIC;
    x_rsc_7_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARLOCK : IN STD_LOGIC;
    x_rsc_7_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_7_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_7_0_ARID : IN STD_LOGIC;
    x_rsc_7_0_BREADY : IN STD_LOGIC;
    x_rsc_7_0_BVALID : OUT STD_LOGIC;
    x_rsc_7_0_BUSER : OUT STD_LOGIC;
    x_rsc_7_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_BID : OUT STD_LOGIC;
    x_rsc_7_0_WREADY : OUT STD_LOGIC;
    x_rsc_7_0_WVALID : IN STD_LOGIC;
    x_rsc_7_0_WUSER : IN STD_LOGIC;
    x_rsc_7_0_WLAST : IN STD_LOGIC;
    x_rsc_7_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_AWREADY : OUT STD_LOGIC;
    x_rsc_7_0_AWVALID : IN STD_LOGIC;
    x_rsc_7_0_AWUSER : IN STD_LOGIC;
    x_rsc_7_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWLOCK : IN STD_LOGIC;
    x_rsc_7_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_7_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_7_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_7_0_lz : OUT STD_LOGIC;
    x_rsc_8_0_s_tdone : IN STD_LOGIC;
    x_rsc_8_0_tr_write_done : IN STD_LOGIC;
    x_rsc_8_0_RREADY : IN STD_LOGIC;
    x_rsc_8_0_RVALID : OUT STD_LOGIC;
    x_rsc_8_0_RUSER : OUT STD_LOGIC;
    x_rsc_8_0_RLAST : OUT STD_LOGIC;
    x_rsc_8_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_RID : OUT STD_LOGIC;
    x_rsc_8_0_ARREADY : OUT STD_LOGIC;
    x_rsc_8_0_ARVALID : IN STD_LOGIC;
    x_rsc_8_0_ARUSER : IN STD_LOGIC;
    x_rsc_8_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARLOCK : IN STD_LOGIC;
    x_rsc_8_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_8_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_8_0_ARID : IN STD_LOGIC;
    x_rsc_8_0_BREADY : IN STD_LOGIC;
    x_rsc_8_0_BVALID : OUT STD_LOGIC;
    x_rsc_8_0_BUSER : OUT STD_LOGIC;
    x_rsc_8_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_BID : OUT STD_LOGIC;
    x_rsc_8_0_WREADY : OUT STD_LOGIC;
    x_rsc_8_0_WVALID : IN STD_LOGIC;
    x_rsc_8_0_WUSER : IN STD_LOGIC;
    x_rsc_8_0_WLAST : IN STD_LOGIC;
    x_rsc_8_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_AWREADY : OUT STD_LOGIC;
    x_rsc_8_0_AWVALID : IN STD_LOGIC;
    x_rsc_8_0_AWUSER : IN STD_LOGIC;
    x_rsc_8_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWLOCK : IN STD_LOGIC;
    x_rsc_8_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_8_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_8_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_8_0_lz : OUT STD_LOGIC;
    x_rsc_9_0_s_tdone : IN STD_LOGIC;
    x_rsc_9_0_tr_write_done : IN STD_LOGIC;
    x_rsc_9_0_RREADY : IN STD_LOGIC;
    x_rsc_9_0_RVALID : OUT STD_LOGIC;
    x_rsc_9_0_RUSER : OUT STD_LOGIC;
    x_rsc_9_0_RLAST : OUT STD_LOGIC;
    x_rsc_9_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_RID : OUT STD_LOGIC;
    x_rsc_9_0_ARREADY : OUT STD_LOGIC;
    x_rsc_9_0_ARVALID : IN STD_LOGIC;
    x_rsc_9_0_ARUSER : IN STD_LOGIC;
    x_rsc_9_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARLOCK : IN STD_LOGIC;
    x_rsc_9_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_9_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_9_0_ARID : IN STD_LOGIC;
    x_rsc_9_0_BREADY : IN STD_LOGIC;
    x_rsc_9_0_BVALID : OUT STD_LOGIC;
    x_rsc_9_0_BUSER : OUT STD_LOGIC;
    x_rsc_9_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_BID : OUT STD_LOGIC;
    x_rsc_9_0_WREADY : OUT STD_LOGIC;
    x_rsc_9_0_WVALID : IN STD_LOGIC;
    x_rsc_9_0_WUSER : IN STD_LOGIC;
    x_rsc_9_0_WLAST : IN STD_LOGIC;
    x_rsc_9_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_AWREADY : OUT STD_LOGIC;
    x_rsc_9_0_AWVALID : IN STD_LOGIC;
    x_rsc_9_0_AWUSER : IN STD_LOGIC;
    x_rsc_9_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWLOCK : IN STD_LOGIC;
    x_rsc_9_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_9_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_9_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_9_0_lz : OUT STD_LOGIC;
    x_rsc_10_0_s_tdone : IN STD_LOGIC;
    x_rsc_10_0_tr_write_done : IN STD_LOGIC;
    x_rsc_10_0_RREADY : IN STD_LOGIC;
    x_rsc_10_0_RVALID : OUT STD_LOGIC;
    x_rsc_10_0_RUSER : OUT STD_LOGIC;
    x_rsc_10_0_RLAST : OUT STD_LOGIC;
    x_rsc_10_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_RID : OUT STD_LOGIC;
    x_rsc_10_0_ARREADY : OUT STD_LOGIC;
    x_rsc_10_0_ARVALID : IN STD_LOGIC;
    x_rsc_10_0_ARUSER : IN STD_LOGIC;
    x_rsc_10_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARLOCK : IN STD_LOGIC;
    x_rsc_10_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_10_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_10_0_ARID : IN STD_LOGIC;
    x_rsc_10_0_BREADY : IN STD_LOGIC;
    x_rsc_10_0_BVALID : OUT STD_LOGIC;
    x_rsc_10_0_BUSER : OUT STD_LOGIC;
    x_rsc_10_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_BID : OUT STD_LOGIC;
    x_rsc_10_0_WREADY : OUT STD_LOGIC;
    x_rsc_10_0_WVALID : IN STD_LOGIC;
    x_rsc_10_0_WUSER : IN STD_LOGIC;
    x_rsc_10_0_WLAST : IN STD_LOGIC;
    x_rsc_10_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_AWREADY : OUT STD_LOGIC;
    x_rsc_10_0_AWVALID : IN STD_LOGIC;
    x_rsc_10_0_AWUSER : IN STD_LOGIC;
    x_rsc_10_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWLOCK : IN STD_LOGIC;
    x_rsc_10_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_10_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_10_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_10_0_lz : OUT STD_LOGIC;
    x_rsc_11_0_s_tdone : IN STD_LOGIC;
    x_rsc_11_0_tr_write_done : IN STD_LOGIC;
    x_rsc_11_0_RREADY : IN STD_LOGIC;
    x_rsc_11_0_RVALID : OUT STD_LOGIC;
    x_rsc_11_0_RUSER : OUT STD_LOGIC;
    x_rsc_11_0_RLAST : OUT STD_LOGIC;
    x_rsc_11_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_RID : OUT STD_LOGIC;
    x_rsc_11_0_ARREADY : OUT STD_LOGIC;
    x_rsc_11_0_ARVALID : IN STD_LOGIC;
    x_rsc_11_0_ARUSER : IN STD_LOGIC;
    x_rsc_11_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARLOCK : IN STD_LOGIC;
    x_rsc_11_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_11_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_11_0_ARID : IN STD_LOGIC;
    x_rsc_11_0_BREADY : IN STD_LOGIC;
    x_rsc_11_0_BVALID : OUT STD_LOGIC;
    x_rsc_11_0_BUSER : OUT STD_LOGIC;
    x_rsc_11_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_BID : OUT STD_LOGIC;
    x_rsc_11_0_WREADY : OUT STD_LOGIC;
    x_rsc_11_0_WVALID : IN STD_LOGIC;
    x_rsc_11_0_WUSER : IN STD_LOGIC;
    x_rsc_11_0_WLAST : IN STD_LOGIC;
    x_rsc_11_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_AWREADY : OUT STD_LOGIC;
    x_rsc_11_0_AWVALID : IN STD_LOGIC;
    x_rsc_11_0_AWUSER : IN STD_LOGIC;
    x_rsc_11_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWLOCK : IN STD_LOGIC;
    x_rsc_11_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_11_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_11_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_11_0_lz : OUT STD_LOGIC;
    x_rsc_12_0_s_tdone : IN STD_LOGIC;
    x_rsc_12_0_tr_write_done : IN STD_LOGIC;
    x_rsc_12_0_RREADY : IN STD_LOGIC;
    x_rsc_12_0_RVALID : OUT STD_LOGIC;
    x_rsc_12_0_RUSER : OUT STD_LOGIC;
    x_rsc_12_0_RLAST : OUT STD_LOGIC;
    x_rsc_12_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_RID : OUT STD_LOGIC;
    x_rsc_12_0_ARREADY : OUT STD_LOGIC;
    x_rsc_12_0_ARVALID : IN STD_LOGIC;
    x_rsc_12_0_ARUSER : IN STD_LOGIC;
    x_rsc_12_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARLOCK : IN STD_LOGIC;
    x_rsc_12_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_12_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_12_0_ARID : IN STD_LOGIC;
    x_rsc_12_0_BREADY : IN STD_LOGIC;
    x_rsc_12_0_BVALID : OUT STD_LOGIC;
    x_rsc_12_0_BUSER : OUT STD_LOGIC;
    x_rsc_12_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_BID : OUT STD_LOGIC;
    x_rsc_12_0_WREADY : OUT STD_LOGIC;
    x_rsc_12_0_WVALID : IN STD_LOGIC;
    x_rsc_12_0_WUSER : IN STD_LOGIC;
    x_rsc_12_0_WLAST : IN STD_LOGIC;
    x_rsc_12_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_AWREADY : OUT STD_LOGIC;
    x_rsc_12_0_AWVALID : IN STD_LOGIC;
    x_rsc_12_0_AWUSER : IN STD_LOGIC;
    x_rsc_12_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWLOCK : IN STD_LOGIC;
    x_rsc_12_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_12_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_12_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_12_0_lz : OUT STD_LOGIC;
    x_rsc_13_0_s_tdone : IN STD_LOGIC;
    x_rsc_13_0_tr_write_done : IN STD_LOGIC;
    x_rsc_13_0_RREADY : IN STD_LOGIC;
    x_rsc_13_0_RVALID : OUT STD_LOGIC;
    x_rsc_13_0_RUSER : OUT STD_LOGIC;
    x_rsc_13_0_RLAST : OUT STD_LOGIC;
    x_rsc_13_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_RID : OUT STD_LOGIC;
    x_rsc_13_0_ARREADY : OUT STD_LOGIC;
    x_rsc_13_0_ARVALID : IN STD_LOGIC;
    x_rsc_13_0_ARUSER : IN STD_LOGIC;
    x_rsc_13_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARLOCK : IN STD_LOGIC;
    x_rsc_13_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_13_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_13_0_ARID : IN STD_LOGIC;
    x_rsc_13_0_BREADY : IN STD_LOGIC;
    x_rsc_13_0_BVALID : OUT STD_LOGIC;
    x_rsc_13_0_BUSER : OUT STD_LOGIC;
    x_rsc_13_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_BID : OUT STD_LOGIC;
    x_rsc_13_0_WREADY : OUT STD_LOGIC;
    x_rsc_13_0_WVALID : IN STD_LOGIC;
    x_rsc_13_0_WUSER : IN STD_LOGIC;
    x_rsc_13_0_WLAST : IN STD_LOGIC;
    x_rsc_13_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_AWREADY : OUT STD_LOGIC;
    x_rsc_13_0_AWVALID : IN STD_LOGIC;
    x_rsc_13_0_AWUSER : IN STD_LOGIC;
    x_rsc_13_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWLOCK : IN STD_LOGIC;
    x_rsc_13_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_13_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_13_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_13_0_lz : OUT STD_LOGIC;
    x_rsc_14_0_s_tdone : IN STD_LOGIC;
    x_rsc_14_0_tr_write_done : IN STD_LOGIC;
    x_rsc_14_0_RREADY : IN STD_LOGIC;
    x_rsc_14_0_RVALID : OUT STD_LOGIC;
    x_rsc_14_0_RUSER : OUT STD_LOGIC;
    x_rsc_14_0_RLAST : OUT STD_LOGIC;
    x_rsc_14_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_RID : OUT STD_LOGIC;
    x_rsc_14_0_ARREADY : OUT STD_LOGIC;
    x_rsc_14_0_ARVALID : IN STD_LOGIC;
    x_rsc_14_0_ARUSER : IN STD_LOGIC;
    x_rsc_14_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARLOCK : IN STD_LOGIC;
    x_rsc_14_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_14_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_14_0_ARID : IN STD_LOGIC;
    x_rsc_14_0_BREADY : IN STD_LOGIC;
    x_rsc_14_0_BVALID : OUT STD_LOGIC;
    x_rsc_14_0_BUSER : OUT STD_LOGIC;
    x_rsc_14_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_BID : OUT STD_LOGIC;
    x_rsc_14_0_WREADY : OUT STD_LOGIC;
    x_rsc_14_0_WVALID : IN STD_LOGIC;
    x_rsc_14_0_WUSER : IN STD_LOGIC;
    x_rsc_14_0_WLAST : IN STD_LOGIC;
    x_rsc_14_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_AWREADY : OUT STD_LOGIC;
    x_rsc_14_0_AWVALID : IN STD_LOGIC;
    x_rsc_14_0_AWUSER : IN STD_LOGIC;
    x_rsc_14_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWLOCK : IN STD_LOGIC;
    x_rsc_14_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_14_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_14_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_14_0_lz : OUT STD_LOGIC;
    x_rsc_15_0_s_tdone : IN STD_LOGIC;
    x_rsc_15_0_tr_write_done : IN STD_LOGIC;
    x_rsc_15_0_RREADY : IN STD_LOGIC;
    x_rsc_15_0_RVALID : OUT STD_LOGIC;
    x_rsc_15_0_RUSER : OUT STD_LOGIC;
    x_rsc_15_0_RLAST : OUT STD_LOGIC;
    x_rsc_15_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_RID : OUT STD_LOGIC;
    x_rsc_15_0_ARREADY : OUT STD_LOGIC;
    x_rsc_15_0_ARVALID : IN STD_LOGIC;
    x_rsc_15_0_ARUSER : IN STD_LOGIC;
    x_rsc_15_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARLOCK : IN STD_LOGIC;
    x_rsc_15_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_15_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_15_0_ARID : IN STD_LOGIC;
    x_rsc_15_0_BREADY : IN STD_LOGIC;
    x_rsc_15_0_BVALID : OUT STD_LOGIC;
    x_rsc_15_0_BUSER : OUT STD_LOGIC;
    x_rsc_15_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_BID : OUT STD_LOGIC;
    x_rsc_15_0_WREADY : OUT STD_LOGIC;
    x_rsc_15_0_WVALID : IN STD_LOGIC;
    x_rsc_15_0_WUSER : IN STD_LOGIC;
    x_rsc_15_0_WLAST : IN STD_LOGIC;
    x_rsc_15_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_AWREADY : OUT STD_LOGIC;
    x_rsc_15_0_AWVALID : IN STD_LOGIC;
    x_rsc_15_0_AWUSER : IN STD_LOGIC;
    x_rsc_15_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWLOCK : IN STD_LOGIC;
    x_rsc_15_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_15_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_15_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_15_0_lz : OUT STD_LOGIC;
    x_rsc_16_0_s_tdone : IN STD_LOGIC;
    x_rsc_16_0_tr_write_done : IN STD_LOGIC;
    x_rsc_16_0_RREADY : IN STD_LOGIC;
    x_rsc_16_0_RVALID : OUT STD_LOGIC;
    x_rsc_16_0_RUSER : OUT STD_LOGIC;
    x_rsc_16_0_RLAST : OUT STD_LOGIC;
    x_rsc_16_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_RID : OUT STD_LOGIC;
    x_rsc_16_0_ARREADY : OUT STD_LOGIC;
    x_rsc_16_0_ARVALID : IN STD_LOGIC;
    x_rsc_16_0_ARUSER : IN STD_LOGIC;
    x_rsc_16_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARLOCK : IN STD_LOGIC;
    x_rsc_16_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_16_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_16_0_ARID : IN STD_LOGIC;
    x_rsc_16_0_BREADY : IN STD_LOGIC;
    x_rsc_16_0_BVALID : OUT STD_LOGIC;
    x_rsc_16_0_BUSER : OUT STD_LOGIC;
    x_rsc_16_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_BID : OUT STD_LOGIC;
    x_rsc_16_0_WREADY : OUT STD_LOGIC;
    x_rsc_16_0_WVALID : IN STD_LOGIC;
    x_rsc_16_0_WUSER : IN STD_LOGIC;
    x_rsc_16_0_WLAST : IN STD_LOGIC;
    x_rsc_16_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_AWREADY : OUT STD_LOGIC;
    x_rsc_16_0_AWVALID : IN STD_LOGIC;
    x_rsc_16_0_AWUSER : IN STD_LOGIC;
    x_rsc_16_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWLOCK : IN STD_LOGIC;
    x_rsc_16_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_16_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_16_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_16_0_lz : OUT STD_LOGIC;
    x_rsc_17_0_s_tdone : IN STD_LOGIC;
    x_rsc_17_0_tr_write_done : IN STD_LOGIC;
    x_rsc_17_0_RREADY : IN STD_LOGIC;
    x_rsc_17_0_RVALID : OUT STD_LOGIC;
    x_rsc_17_0_RUSER : OUT STD_LOGIC;
    x_rsc_17_0_RLAST : OUT STD_LOGIC;
    x_rsc_17_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_RID : OUT STD_LOGIC;
    x_rsc_17_0_ARREADY : OUT STD_LOGIC;
    x_rsc_17_0_ARVALID : IN STD_LOGIC;
    x_rsc_17_0_ARUSER : IN STD_LOGIC;
    x_rsc_17_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARLOCK : IN STD_LOGIC;
    x_rsc_17_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_17_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_17_0_ARID : IN STD_LOGIC;
    x_rsc_17_0_BREADY : IN STD_LOGIC;
    x_rsc_17_0_BVALID : OUT STD_LOGIC;
    x_rsc_17_0_BUSER : OUT STD_LOGIC;
    x_rsc_17_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_BID : OUT STD_LOGIC;
    x_rsc_17_0_WREADY : OUT STD_LOGIC;
    x_rsc_17_0_WVALID : IN STD_LOGIC;
    x_rsc_17_0_WUSER : IN STD_LOGIC;
    x_rsc_17_0_WLAST : IN STD_LOGIC;
    x_rsc_17_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_AWREADY : OUT STD_LOGIC;
    x_rsc_17_0_AWVALID : IN STD_LOGIC;
    x_rsc_17_0_AWUSER : IN STD_LOGIC;
    x_rsc_17_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWLOCK : IN STD_LOGIC;
    x_rsc_17_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_17_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_17_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_17_0_lz : OUT STD_LOGIC;
    x_rsc_18_0_s_tdone : IN STD_LOGIC;
    x_rsc_18_0_tr_write_done : IN STD_LOGIC;
    x_rsc_18_0_RREADY : IN STD_LOGIC;
    x_rsc_18_0_RVALID : OUT STD_LOGIC;
    x_rsc_18_0_RUSER : OUT STD_LOGIC;
    x_rsc_18_0_RLAST : OUT STD_LOGIC;
    x_rsc_18_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_RID : OUT STD_LOGIC;
    x_rsc_18_0_ARREADY : OUT STD_LOGIC;
    x_rsc_18_0_ARVALID : IN STD_LOGIC;
    x_rsc_18_0_ARUSER : IN STD_LOGIC;
    x_rsc_18_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARLOCK : IN STD_LOGIC;
    x_rsc_18_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_18_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_18_0_ARID : IN STD_LOGIC;
    x_rsc_18_0_BREADY : IN STD_LOGIC;
    x_rsc_18_0_BVALID : OUT STD_LOGIC;
    x_rsc_18_0_BUSER : OUT STD_LOGIC;
    x_rsc_18_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_BID : OUT STD_LOGIC;
    x_rsc_18_0_WREADY : OUT STD_LOGIC;
    x_rsc_18_0_WVALID : IN STD_LOGIC;
    x_rsc_18_0_WUSER : IN STD_LOGIC;
    x_rsc_18_0_WLAST : IN STD_LOGIC;
    x_rsc_18_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_AWREADY : OUT STD_LOGIC;
    x_rsc_18_0_AWVALID : IN STD_LOGIC;
    x_rsc_18_0_AWUSER : IN STD_LOGIC;
    x_rsc_18_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWLOCK : IN STD_LOGIC;
    x_rsc_18_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_18_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_18_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_18_0_lz : OUT STD_LOGIC;
    x_rsc_19_0_s_tdone : IN STD_LOGIC;
    x_rsc_19_0_tr_write_done : IN STD_LOGIC;
    x_rsc_19_0_RREADY : IN STD_LOGIC;
    x_rsc_19_0_RVALID : OUT STD_LOGIC;
    x_rsc_19_0_RUSER : OUT STD_LOGIC;
    x_rsc_19_0_RLAST : OUT STD_LOGIC;
    x_rsc_19_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_RID : OUT STD_LOGIC;
    x_rsc_19_0_ARREADY : OUT STD_LOGIC;
    x_rsc_19_0_ARVALID : IN STD_LOGIC;
    x_rsc_19_0_ARUSER : IN STD_LOGIC;
    x_rsc_19_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARLOCK : IN STD_LOGIC;
    x_rsc_19_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_19_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_19_0_ARID : IN STD_LOGIC;
    x_rsc_19_0_BREADY : IN STD_LOGIC;
    x_rsc_19_0_BVALID : OUT STD_LOGIC;
    x_rsc_19_0_BUSER : OUT STD_LOGIC;
    x_rsc_19_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_BID : OUT STD_LOGIC;
    x_rsc_19_0_WREADY : OUT STD_LOGIC;
    x_rsc_19_0_WVALID : IN STD_LOGIC;
    x_rsc_19_0_WUSER : IN STD_LOGIC;
    x_rsc_19_0_WLAST : IN STD_LOGIC;
    x_rsc_19_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_AWREADY : OUT STD_LOGIC;
    x_rsc_19_0_AWVALID : IN STD_LOGIC;
    x_rsc_19_0_AWUSER : IN STD_LOGIC;
    x_rsc_19_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWLOCK : IN STD_LOGIC;
    x_rsc_19_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_19_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_19_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_19_0_lz : OUT STD_LOGIC;
    x_rsc_20_0_s_tdone : IN STD_LOGIC;
    x_rsc_20_0_tr_write_done : IN STD_LOGIC;
    x_rsc_20_0_RREADY : IN STD_LOGIC;
    x_rsc_20_0_RVALID : OUT STD_LOGIC;
    x_rsc_20_0_RUSER : OUT STD_LOGIC;
    x_rsc_20_0_RLAST : OUT STD_LOGIC;
    x_rsc_20_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_RID : OUT STD_LOGIC;
    x_rsc_20_0_ARREADY : OUT STD_LOGIC;
    x_rsc_20_0_ARVALID : IN STD_LOGIC;
    x_rsc_20_0_ARUSER : IN STD_LOGIC;
    x_rsc_20_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARLOCK : IN STD_LOGIC;
    x_rsc_20_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_20_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_20_0_ARID : IN STD_LOGIC;
    x_rsc_20_0_BREADY : IN STD_LOGIC;
    x_rsc_20_0_BVALID : OUT STD_LOGIC;
    x_rsc_20_0_BUSER : OUT STD_LOGIC;
    x_rsc_20_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_BID : OUT STD_LOGIC;
    x_rsc_20_0_WREADY : OUT STD_LOGIC;
    x_rsc_20_0_WVALID : IN STD_LOGIC;
    x_rsc_20_0_WUSER : IN STD_LOGIC;
    x_rsc_20_0_WLAST : IN STD_LOGIC;
    x_rsc_20_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_AWREADY : OUT STD_LOGIC;
    x_rsc_20_0_AWVALID : IN STD_LOGIC;
    x_rsc_20_0_AWUSER : IN STD_LOGIC;
    x_rsc_20_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWLOCK : IN STD_LOGIC;
    x_rsc_20_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_20_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_20_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_20_0_lz : OUT STD_LOGIC;
    x_rsc_21_0_s_tdone : IN STD_LOGIC;
    x_rsc_21_0_tr_write_done : IN STD_LOGIC;
    x_rsc_21_0_RREADY : IN STD_LOGIC;
    x_rsc_21_0_RVALID : OUT STD_LOGIC;
    x_rsc_21_0_RUSER : OUT STD_LOGIC;
    x_rsc_21_0_RLAST : OUT STD_LOGIC;
    x_rsc_21_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_RID : OUT STD_LOGIC;
    x_rsc_21_0_ARREADY : OUT STD_LOGIC;
    x_rsc_21_0_ARVALID : IN STD_LOGIC;
    x_rsc_21_0_ARUSER : IN STD_LOGIC;
    x_rsc_21_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARLOCK : IN STD_LOGIC;
    x_rsc_21_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_21_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_21_0_ARID : IN STD_LOGIC;
    x_rsc_21_0_BREADY : IN STD_LOGIC;
    x_rsc_21_0_BVALID : OUT STD_LOGIC;
    x_rsc_21_0_BUSER : OUT STD_LOGIC;
    x_rsc_21_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_BID : OUT STD_LOGIC;
    x_rsc_21_0_WREADY : OUT STD_LOGIC;
    x_rsc_21_0_WVALID : IN STD_LOGIC;
    x_rsc_21_0_WUSER : IN STD_LOGIC;
    x_rsc_21_0_WLAST : IN STD_LOGIC;
    x_rsc_21_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_AWREADY : OUT STD_LOGIC;
    x_rsc_21_0_AWVALID : IN STD_LOGIC;
    x_rsc_21_0_AWUSER : IN STD_LOGIC;
    x_rsc_21_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWLOCK : IN STD_LOGIC;
    x_rsc_21_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_21_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_21_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_21_0_lz : OUT STD_LOGIC;
    x_rsc_22_0_s_tdone : IN STD_LOGIC;
    x_rsc_22_0_tr_write_done : IN STD_LOGIC;
    x_rsc_22_0_RREADY : IN STD_LOGIC;
    x_rsc_22_0_RVALID : OUT STD_LOGIC;
    x_rsc_22_0_RUSER : OUT STD_LOGIC;
    x_rsc_22_0_RLAST : OUT STD_LOGIC;
    x_rsc_22_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_RID : OUT STD_LOGIC;
    x_rsc_22_0_ARREADY : OUT STD_LOGIC;
    x_rsc_22_0_ARVALID : IN STD_LOGIC;
    x_rsc_22_0_ARUSER : IN STD_LOGIC;
    x_rsc_22_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARLOCK : IN STD_LOGIC;
    x_rsc_22_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_22_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_22_0_ARID : IN STD_LOGIC;
    x_rsc_22_0_BREADY : IN STD_LOGIC;
    x_rsc_22_0_BVALID : OUT STD_LOGIC;
    x_rsc_22_0_BUSER : OUT STD_LOGIC;
    x_rsc_22_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_BID : OUT STD_LOGIC;
    x_rsc_22_0_WREADY : OUT STD_LOGIC;
    x_rsc_22_0_WVALID : IN STD_LOGIC;
    x_rsc_22_0_WUSER : IN STD_LOGIC;
    x_rsc_22_0_WLAST : IN STD_LOGIC;
    x_rsc_22_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_AWREADY : OUT STD_LOGIC;
    x_rsc_22_0_AWVALID : IN STD_LOGIC;
    x_rsc_22_0_AWUSER : IN STD_LOGIC;
    x_rsc_22_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWLOCK : IN STD_LOGIC;
    x_rsc_22_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_22_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_22_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_22_0_lz : OUT STD_LOGIC;
    x_rsc_23_0_s_tdone : IN STD_LOGIC;
    x_rsc_23_0_tr_write_done : IN STD_LOGIC;
    x_rsc_23_0_RREADY : IN STD_LOGIC;
    x_rsc_23_0_RVALID : OUT STD_LOGIC;
    x_rsc_23_0_RUSER : OUT STD_LOGIC;
    x_rsc_23_0_RLAST : OUT STD_LOGIC;
    x_rsc_23_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_RID : OUT STD_LOGIC;
    x_rsc_23_0_ARREADY : OUT STD_LOGIC;
    x_rsc_23_0_ARVALID : IN STD_LOGIC;
    x_rsc_23_0_ARUSER : IN STD_LOGIC;
    x_rsc_23_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARLOCK : IN STD_LOGIC;
    x_rsc_23_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_23_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_23_0_ARID : IN STD_LOGIC;
    x_rsc_23_0_BREADY : IN STD_LOGIC;
    x_rsc_23_0_BVALID : OUT STD_LOGIC;
    x_rsc_23_0_BUSER : OUT STD_LOGIC;
    x_rsc_23_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_BID : OUT STD_LOGIC;
    x_rsc_23_0_WREADY : OUT STD_LOGIC;
    x_rsc_23_0_WVALID : IN STD_LOGIC;
    x_rsc_23_0_WUSER : IN STD_LOGIC;
    x_rsc_23_0_WLAST : IN STD_LOGIC;
    x_rsc_23_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_AWREADY : OUT STD_LOGIC;
    x_rsc_23_0_AWVALID : IN STD_LOGIC;
    x_rsc_23_0_AWUSER : IN STD_LOGIC;
    x_rsc_23_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWLOCK : IN STD_LOGIC;
    x_rsc_23_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_23_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_23_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_23_0_lz : OUT STD_LOGIC;
    x_rsc_24_0_s_tdone : IN STD_LOGIC;
    x_rsc_24_0_tr_write_done : IN STD_LOGIC;
    x_rsc_24_0_RREADY : IN STD_LOGIC;
    x_rsc_24_0_RVALID : OUT STD_LOGIC;
    x_rsc_24_0_RUSER : OUT STD_LOGIC;
    x_rsc_24_0_RLAST : OUT STD_LOGIC;
    x_rsc_24_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_RID : OUT STD_LOGIC;
    x_rsc_24_0_ARREADY : OUT STD_LOGIC;
    x_rsc_24_0_ARVALID : IN STD_LOGIC;
    x_rsc_24_0_ARUSER : IN STD_LOGIC;
    x_rsc_24_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARLOCK : IN STD_LOGIC;
    x_rsc_24_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_24_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_24_0_ARID : IN STD_LOGIC;
    x_rsc_24_0_BREADY : IN STD_LOGIC;
    x_rsc_24_0_BVALID : OUT STD_LOGIC;
    x_rsc_24_0_BUSER : OUT STD_LOGIC;
    x_rsc_24_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_BID : OUT STD_LOGIC;
    x_rsc_24_0_WREADY : OUT STD_LOGIC;
    x_rsc_24_0_WVALID : IN STD_LOGIC;
    x_rsc_24_0_WUSER : IN STD_LOGIC;
    x_rsc_24_0_WLAST : IN STD_LOGIC;
    x_rsc_24_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_AWREADY : OUT STD_LOGIC;
    x_rsc_24_0_AWVALID : IN STD_LOGIC;
    x_rsc_24_0_AWUSER : IN STD_LOGIC;
    x_rsc_24_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWLOCK : IN STD_LOGIC;
    x_rsc_24_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_24_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_24_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_24_0_lz : OUT STD_LOGIC;
    x_rsc_25_0_s_tdone : IN STD_LOGIC;
    x_rsc_25_0_tr_write_done : IN STD_LOGIC;
    x_rsc_25_0_RREADY : IN STD_LOGIC;
    x_rsc_25_0_RVALID : OUT STD_LOGIC;
    x_rsc_25_0_RUSER : OUT STD_LOGIC;
    x_rsc_25_0_RLAST : OUT STD_LOGIC;
    x_rsc_25_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_RID : OUT STD_LOGIC;
    x_rsc_25_0_ARREADY : OUT STD_LOGIC;
    x_rsc_25_0_ARVALID : IN STD_LOGIC;
    x_rsc_25_0_ARUSER : IN STD_LOGIC;
    x_rsc_25_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARLOCK : IN STD_LOGIC;
    x_rsc_25_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_25_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_25_0_ARID : IN STD_LOGIC;
    x_rsc_25_0_BREADY : IN STD_LOGIC;
    x_rsc_25_0_BVALID : OUT STD_LOGIC;
    x_rsc_25_0_BUSER : OUT STD_LOGIC;
    x_rsc_25_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_BID : OUT STD_LOGIC;
    x_rsc_25_0_WREADY : OUT STD_LOGIC;
    x_rsc_25_0_WVALID : IN STD_LOGIC;
    x_rsc_25_0_WUSER : IN STD_LOGIC;
    x_rsc_25_0_WLAST : IN STD_LOGIC;
    x_rsc_25_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_AWREADY : OUT STD_LOGIC;
    x_rsc_25_0_AWVALID : IN STD_LOGIC;
    x_rsc_25_0_AWUSER : IN STD_LOGIC;
    x_rsc_25_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWLOCK : IN STD_LOGIC;
    x_rsc_25_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_25_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_25_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_25_0_lz : OUT STD_LOGIC;
    x_rsc_26_0_s_tdone : IN STD_LOGIC;
    x_rsc_26_0_tr_write_done : IN STD_LOGIC;
    x_rsc_26_0_RREADY : IN STD_LOGIC;
    x_rsc_26_0_RVALID : OUT STD_LOGIC;
    x_rsc_26_0_RUSER : OUT STD_LOGIC;
    x_rsc_26_0_RLAST : OUT STD_LOGIC;
    x_rsc_26_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_RID : OUT STD_LOGIC;
    x_rsc_26_0_ARREADY : OUT STD_LOGIC;
    x_rsc_26_0_ARVALID : IN STD_LOGIC;
    x_rsc_26_0_ARUSER : IN STD_LOGIC;
    x_rsc_26_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARLOCK : IN STD_LOGIC;
    x_rsc_26_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_26_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_26_0_ARID : IN STD_LOGIC;
    x_rsc_26_0_BREADY : IN STD_LOGIC;
    x_rsc_26_0_BVALID : OUT STD_LOGIC;
    x_rsc_26_0_BUSER : OUT STD_LOGIC;
    x_rsc_26_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_BID : OUT STD_LOGIC;
    x_rsc_26_0_WREADY : OUT STD_LOGIC;
    x_rsc_26_0_WVALID : IN STD_LOGIC;
    x_rsc_26_0_WUSER : IN STD_LOGIC;
    x_rsc_26_0_WLAST : IN STD_LOGIC;
    x_rsc_26_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_AWREADY : OUT STD_LOGIC;
    x_rsc_26_0_AWVALID : IN STD_LOGIC;
    x_rsc_26_0_AWUSER : IN STD_LOGIC;
    x_rsc_26_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWLOCK : IN STD_LOGIC;
    x_rsc_26_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_26_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_26_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_26_0_lz : OUT STD_LOGIC;
    x_rsc_27_0_s_tdone : IN STD_LOGIC;
    x_rsc_27_0_tr_write_done : IN STD_LOGIC;
    x_rsc_27_0_RREADY : IN STD_LOGIC;
    x_rsc_27_0_RVALID : OUT STD_LOGIC;
    x_rsc_27_0_RUSER : OUT STD_LOGIC;
    x_rsc_27_0_RLAST : OUT STD_LOGIC;
    x_rsc_27_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_RID : OUT STD_LOGIC;
    x_rsc_27_0_ARREADY : OUT STD_LOGIC;
    x_rsc_27_0_ARVALID : IN STD_LOGIC;
    x_rsc_27_0_ARUSER : IN STD_LOGIC;
    x_rsc_27_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARLOCK : IN STD_LOGIC;
    x_rsc_27_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_27_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_27_0_ARID : IN STD_LOGIC;
    x_rsc_27_0_BREADY : IN STD_LOGIC;
    x_rsc_27_0_BVALID : OUT STD_LOGIC;
    x_rsc_27_0_BUSER : OUT STD_LOGIC;
    x_rsc_27_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_BID : OUT STD_LOGIC;
    x_rsc_27_0_WREADY : OUT STD_LOGIC;
    x_rsc_27_0_WVALID : IN STD_LOGIC;
    x_rsc_27_0_WUSER : IN STD_LOGIC;
    x_rsc_27_0_WLAST : IN STD_LOGIC;
    x_rsc_27_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_AWREADY : OUT STD_LOGIC;
    x_rsc_27_0_AWVALID : IN STD_LOGIC;
    x_rsc_27_0_AWUSER : IN STD_LOGIC;
    x_rsc_27_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWLOCK : IN STD_LOGIC;
    x_rsc_27_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_27_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_27_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_27_0_lz : OUT STD_LOGIC;
    x_rsc_28_0_s_tdone : IN STD_LOGIC;
    x_rsc_28_0_tr_write_done : IN STD_LOGIC;
    x_rsc_28_0_RREADY : IN STD_LOGIC;
    x_rsc_28_0_RVALID : OUT STD_LOGIC;
    x_rsc_28_0_RUSER : OUT STD_LOGIC;
    x_rsc_28_0_RLAST : OUT STD_LOGIC;
    x_rsc_28_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_RID : OUT STD_LOGIC;
    x_rsc_28_0_ARREADY : OUT STD_LOGIC;
    x_rsc_28_0_ARVALID : IN STD_LOGIC;
    x_rsc_28_0_ARUSER : IN STD_LOGIC;
    x_rsc_28_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARLOCK : IN STD_LOGIC;
    x_rsc_28_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_28_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_28_0_ARID : IN STD_LOGIC;
    x_rsc_28_0_BREADY : IN STD_LOGIC;
    x_rsc_28_0_BVALID : OUT STD_LOGIC;
    x_rsc_28_0_BUSER : OUT STD_LOGIC;
    x_rsc_28_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_BID : OUT STD_LOGIC;
    x_rsc_28_0_WREADY : OUT STD_LOGIC;
    x_rsc_28_0_WVALID : IN STD_LOGIC;
    x_rsc_28_0_WUSER : IN STD_LOGIC;
    x_rsc_28_0_WLAST : IN STD_LOGIC;
    x_rsc_28_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_AWREADY : OUT STD_LOGIC;
    x_rsc_28_0_AWVALID : IN STD_LOGIC;
    x_rsc_28_0_AWUSER : IN STD_LOGIC;
    x_rsc_28_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWLOCK : IN STD_LOGIC;
    x_rsc_28_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_28_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_28_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_28_0_lz : OUT STD_LOGIC;
    x_rsc_29_0_s_tdone : IN STD_LOGIC;
    x_rsc_29_0_tr_write_done : IN STD_LOGIC;
    x_rsc_29_0_RREADY : IN STD_LOGIC;
    x_rsc_29_0_RVALID : OUT STD_LOGIC;
    x_rsc_29_0_RUSER : OUT STD_LOGIC;
    x_rsc_29_0_RLAST : OUT STD_LOGIC;
    x_rsc_29_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_RID : OUT STD_LOGIC;
    x_rsc_29_0_ARREADY : OUT STD_LOGIC;
    x_rsc_29_0_ARVALID : IN STD_LOGIC;
    x_rsc_29_0_ARUSER : IN STD_LOGIC;
    x_rsc_29_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARLOCK : IN STD_LOGIC;
    x_rsc_29_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_29_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_29_0_ARID : IN STD_LOGIC;
    x_rsc_29_0_BREADY : IN STD_LOGIC;
    x_rsc_29_0_BVALID : OUT STD_LOGIC;
    x_rsc_29_0_BUSER : OUT STD_LOGIC;
    x_rsc_29_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_BID : OUT STD_LOGIC;
    x_rsc_29_0_WREADY : OUT STD_LOGIC;
    x_rsc_29_0_WVALID : IN STD_LOGIC;
    x_rsc_29_0_WUSER : IN STD_LOGIC;
    x_rsc_29_0_WLAST : IN STD_LOGIC;
    x_rsc_29_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_AWREADY : OUT STD_LOGIC;
    x_rsc_29_0_AWVALID : IN STD_LOGIC;
    x_rsc_29_0_AWUSER : IN STD_LOGIC;
    x_rsc_29_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWLOCK : IN STD_LOGIC;
    x_rsc_29_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_29_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_29_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_29_0_lz : OUT STD_LOGIC;
    x_rsc_30_0_s_tdone : IN STD_LOGIC;
    x_rsc_30_0_tr_write_done : IN STD_LOGIC;
    x_rsc_30_0_RREADY : IN STD_LOGIC;
    x_rsc_30_0_RVALID : OUT STD_LOGIC;
    x_rsc_30_0_RUSER : OUT STD_LOGIC;
    x_rsc_30_0_RLAST : OUT STD_LOGIC;
    x_rsc_30_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_RID : OUT STD_LOGIC;
    x_rsc_30_0_ARREADY : OUT STD_LOGIC;
    x_rsc_30_0_ARVALID : IN STD_LOGIC;
    x_rsc_30_0_ARUSER : IN STD_LOGIC;
    x_rsc_30_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARLOCK : IN STD_LOGIC;
    x_rsc_30_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_30_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_30_0_ARID : IN STD_LOGIC;
    x_rsc_30_0_BREADY : IN STD_LOGIC;
    x_rsc_30_0_BVALID : OUT STD_LOGIC;
    x_rsc_30_0_BUSER : OUT STD_LOGIC;
    x_rsc_30_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_BID : OUT STD_LOGIC;
    x_rsc_30_0_WREADY : OUT STD_LOGIC;
    x_rsc_30_0_WVALID : IN STD_LOGIC;
    x_rsc_30_0_WUSER : IN STD_LOGIC;
    x_rsc_30_0_WLAST : IN STD_LOGIC;
    x_rsc_30_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_AWREADY : OUT STD_LOGIC;
    x_rsc_30_0_AWVALID : IN STD_LOGIC;
    x_rsc_30_0_AWUSER : IN STD_LOGIC;
    x_rsc_30_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWLOCK : IN STD_LOGIC;
    x_rsc_30_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_30_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_30_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_30_0_lz : OUT STD_LOGIC;
    x_rsc_31_0_s_tdone : IN STD_LOGIC;
    x_rsc_31_0_tr_write_done : IN STD_LOGIC;
    x_rsc_31_0_RREADY : IN STD_LOGIC;
    x_rsc_31_0_RVALID : OUT STD_LOGIC;
    x_rsc_31_0_RUSER : OUT STD_LOGIC;
    x_rsc_31_0_RLAST : OUT STD_LOGIC;
    x_rsc_31_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_RID : OUT STD_LOGIC;
    x_rsc_31_0_ARREADY : OUT STD_LOGIC;
    x_rsc_31_0_ARVALID : IN STD_LOGIC;
    x_rsc_31_0_ARUSER : IN STD_LOGIC;
    x_rsc_31_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARLOCK : IN STD_LOGIC;
    x_rsc_31_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_31_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_31_0_ARID : IN STD_LOGIC;
    x_rsc_31_0_BREADY : IN STD_LOGIC;
    x_rsc_31_0_BVALID : OUT STD_LOGIC;
    x_rsc_31_0_BUSER : OUT STD_LOGIC;
    x_rsc_31_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_BID : OUT STD_LOGIC;
    x_rsc_31_0_WREADY : OUT STD_LOGIC;
    x_rsc_31_0_WVALID : IN STD_LOGIC;
    x_rsc_31_0_WUSER : IN STD_LOGIC;
    x_rsc_31_0_WLAST : IN STD_LOGIC;
    x_rsc_31_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_AWREADY : OUT STD_LOGIC;
    x_rsc_31_0_AWVALID : IN STD_LOGIC;
    x_rsc_31_0_AWUSER : IN STD_LOGIC;
    x_rsc_31_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWLOCK : IN STD_LOGIC;
    x_rsc_31_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_31_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_31_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_31_0_lz : OUT STD_LOGIC;
    m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    m_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_h_rsc_triosy_lz : OUT STD_LOGIC;
    revArr_rsc_s_tdone : IN STD_LOGIC;
    revArr_rsc_tr_write_done : IN STD_LOGIC;
    revArr_rsc_RREADY : IN STD_LOGIC;
    revArr_rsc_RVALID : OUT STD_LOGIC;
    revArr_rsc_RUSER : OUT STD_LOGIC;
    revArr_rsc_RLAST : OUT STD_LOGIC;
    revArr_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    revArr_rsc_RID : OUT STD_LOGIC;
    revArr_rsc_ARREADY : OUT STD_LOGIC;
    revArr_rsc_ARVALID : IN STD_LOGIC;
    revArr_rsc_ARUSER : IN STD_LOGIC;
    revArr_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARLOCK : IN STD_LOGIC;
    revArr_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    revArr_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    revArr_rsc_ARID : IN STD_LOGIC;
    revArr_rsc_BREADY : IN STD_LOGIC;
    revArr_rsc_BVALID : OUT STD_LOGIC;
    revArr_rsc_BUSER : OUT STD_LOGIC;
    revArr_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_BID : OUT STD_LOGIC;
    revArr_rsc_WREADY : OUT STD_LOGIC;
    revArr_rsc_WVALID : IN STD_LOGIC;
    revArr_rsc_WUSER : IN STD_LOGIC;
    revArr_rsc_WLAST : IN STD_LOGIC;
    revArr_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    revArr_rsc_AWREADY : OUT STD_LOGIC;
    revArr_rsc_AWVALID : IN STD_LOGIC;
    revArr_rsc_AWUSER : IN STD_LOGIC;
    revArr_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWLOCK : IN STD_LOGIC;
    revArr_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    revArr_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    revArr_rsc_AWID : IN STD_LOGIC;
    revArr_rsc_triosy_lz : OUT STD_LOGIC;
    tw_rsc_s_tdone : IN STD_LOGIC;
    tw_rsc_tr_write_done : IN STD_LOGIC;
    tw_rsc_RREADY : IN STD_LOGIC;
    tw_rsc_RVALID : OUT STD_LOGIC;
    tw_rsc_RUSER : OUT STD_LOGIC;
    tw_rsc_RLAST : OUT STD_LOGIC;
    tw_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_rsc_RID : OUT STD_LOGIC;
    tw_rsc_ARREADY : OUT STD_LOGIC;
    tw_rsc_ARVALID : IN STD_LOGIC;
    tw_rsc_ARUSER : IN STD_LOGIC;
    tw_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARLOCK : IN STD_LOGIC;
    tw_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_rsc_ARID : IN STD_LOGIC;
    tw_rsc_BREADY : IN STD_LOGIC;
    tw_rsc_BVALID : OUT STD_LOGIC;
    tw_rsc_BUSER : OUT STD_LOGIC;
    tw_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_BID : OUT STD_LOGIC;
    tw_rsc_WREADY : OUT STD_LOGIC;
    tw_rsc_WVALID : IN STD_LOGIC;
    tw_rsc_WUSER : IN STD_LOGIC;
    tw_rsc_WLAST : IN STD_LOGIC;
    tw_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_rsc_AWREADY : OUT STD_LOGIC;
    tw_rsc_AWVALID : IN STD_LOGIC;
    tw_rsc_AWUSER : IN STD_LOGIC;
    tw_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWLOCK : IN STD_LOGIC;
    tw_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_rsc_AWID : IN STD_LOGIC;
    tw_rsc_triosy_lz : OUT STD_LOGIC;
    tw_h_rsc_s_tdone : IN STD_LOGIC;
    tw_h_rsc_tr_write_done : IN STD_LOGIC;
    tw_h_rsc_RREADY : IN STD_LOGIC;
    tw_h_rsc_RVALID : OUT STD_LOGIC;
    tw_h_rsc_RUSER : OUT STD_LOGIC;
    tw_h_rsc_RLAST : OUT STD_LOGIC;
    tw_h_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_h_rsc_RID : OUT STD_LOGIC;
    tw_h_rsc_ARREADY : OUT STD_LOGIC;
    tw_h_rsc_ARVALID : IN STD_LOGIC;
    tw_h_rsc_ARUSER : IN STD_LOGIC;
    tw_h_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARLOCK : IN STD_LOGIC;
    tw_h_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_h_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_h_rsc_ARID : IN STD_LOGIC;
    tw_h_rsc_BREADY : IN STD_LOGIC;
    tw_h_rsc_BVALID : OUT STD_LOGIC;
    tw_h_rsc_BUSER : OUT STD_LOGIC;
    tw_h_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_BID : OUT STD_LOGIC;
    tw_h_rsc_WREADY : OUT STD_LOGIC;
    tw_h_rsc_WVALID : IN STD_LOGIC;
    tw_h_rsc_WUSER : IN STD_LOGIC;
    tw_h_rsc_WLAST : IN STD_LOGIC;
    tw_h_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_h_rsc_AWREADY : OUT STD_LOGIC;
    tw_h_rsc_AWVALID : IN STD_LOGIC;
    tw_h_rsc_AWUSER : IN STD_LOGIC;
    tw_h_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWLOCK : IN STD_LOGIC;
    tw_h_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_h_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_h_rsc_AWID : IN STD_LOGIC;
    tw_h_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    twiddle_h_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_h_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xx_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_1_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_2_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_2_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_2_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_3_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_3_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_3_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_4_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_4_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_4_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_5_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_5_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_5_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_6_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_6_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_6_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_7_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_7_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_7_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_8_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_8_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_8_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_9_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_9_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_9_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_10_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_10_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_10_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_11_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_11_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_11_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_12_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_12_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_12_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_13_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_13_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_13_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_14_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_14_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_14_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_15_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_15_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_15_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_16_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_16_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_16_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_17_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_17_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_17_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_18_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_18_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_18_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_19_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_19_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_19_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_20_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_20_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_20_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_21_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_21_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_21_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_22_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_22_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_22_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_23_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_23_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_23_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_24_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_24_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_24_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_25_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_25_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_25_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_26_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_26_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_26_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_27_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_27_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_27_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_28_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_28_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_28_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_29_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_29_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_29_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_30_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_30_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_30_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_31_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
    xx_rsc_31_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_31_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_1_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_2_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_2_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_2_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_3_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_3_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_3_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_4_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_4_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_4_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_5_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_5_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_5_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_6_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_6_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_6_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_7_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_7_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_7_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_8_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_8_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_8_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_9_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_9_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_9_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_10_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_10_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_10_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_11_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_11_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_11_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_12_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_12_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_12_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_13_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_13_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_13_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_14_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_14_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_14_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_15_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_15_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_15_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_16_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_16_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_16_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_17_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_17_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_17_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_18_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_18_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_18_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_19_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_19_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_19_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_20_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_20_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_20_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_21_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_21_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_21_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_22_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_22_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_22_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_23_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_23_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_23_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_24_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_24_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_24_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_25_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_25_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_25_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_26_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_26_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_26_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_27_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_27_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_27_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_28_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_28_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_28_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_29_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_29_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_29_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_30_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_30_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_30_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_31_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    yy_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
    yy_rsc_31_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_31_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
        0);
    S34_OUTER_LOOP_for_tf_mul_cmp_a : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    S34_OUTER_LOOP_for_tf_mul_cmp_b : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    S34_OUTER_LOOP_for_tf_mul_cmp_z : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
    xx_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_1_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_2_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    xx_rsc_3_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_1_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_2_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
    yy_rsc_3_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
  );
END hybrid_core;

ARCHITECTURE v14 OF hybrid_core IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL core_wen : STD_LOGIC;
  SIGNAL m_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL core_wten : STD_LOGIC;
  SIGNAL twiddle_rsci_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsci_qb_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL revArr_rsci_wen_comp : STD_LOGIC;
  SIGNAL revArr_rsci_s_din_mxwt : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL tw_rsci_wen_comp : STD_LOGIC;
  SIGNAL tw_rsci_s_din_mxwt : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL tw_h_rsci_wen_comp : STD_LOGIC;
  SIGNAL tw_h_rsci_s_din_mxwt : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL x_rsc_0_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_0_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_1_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_1_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_2_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_2_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_3_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_3_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_4_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_4_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_5_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_5_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_6_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_6_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_7_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_7_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_8_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_8_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_9_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_9_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_10_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_10_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_11_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_11_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_12_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_12_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_13_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_13_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_14_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_14_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_15_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_15_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_16_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_16_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_17_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_17_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_18_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_18_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_19_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_19_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_20_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_20_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_21_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_21_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_22_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_22_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_23_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_23_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_24_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_24_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_25_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_25_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_26_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_26_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_27_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_27_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_28_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_28_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_29_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_29_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_30_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_30_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL x_rsc_31_0_i_wen_comp : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_wen_comp_1 : STD_LOGIC;
  SIGNAL x_rsc_31_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_mul_cmp_en : STD_LOGIC;
  SIGNAL mult_12_z_mul_cmp_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_en : STD_LOGIC;
  SIGNAL mult_z_mul_cmp_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL S34_OUTER_LOOP_for_k_slc_S34_OUTER_LOOP_for_k_sva_19_5_4_0_1 : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL S34_OUTER_LOOP_for_k_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL fsm_output : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL S6_OUTER_LOOP_for_acc_tmp : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL S34_OUTER_LOOP_for_a_acc_2_tmp : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL operator_20_true_28_acc_tmp : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL and_dcpl_42 : STD_LOGIC;
  SIGNAL not_tmp_28 : STD_LOGIC;
  SIGNAL nor_tmp_3 : STD_LOGIC;
  SIGNAL nor_tmp_4 : STD_LOGIC;
  SIGNAL or_tmp_35 : STD_LOGIC;
  SIGNAL nor_tmp_8 : STD_LOGIC;
  SIGNAL or_tmp_48 : STD_LOGIC;
  SIGNAL or_tmp_59 : STD_LOGIC;
  SIGNAL or_tmp_77 : STD_LOGIC;
  SIGNAL and_dcpl_53 : STD_LOGIC;
  SIGNAL and_dcpl_54 : STD_LOGIC;
  SIGNAL and_dcpl_57 : STD_LOGIC;
  SIGNAL and_dcpl_60 : STD_LOGIC;
  SIGNAL and_dcpl_61 : STD_LOGIC;
  SIGNAL and_dcpl_64 : STD_LOGIC;
  SIGNAL and_dcpl_66 : STD_LOGIC;
  SIGNAL and_dcpl_67 : STD_LOGIC;
  SIGNAL and_dcpl_69 : STD_LOGIC;
  SIGNAL and_dcpl_70 : STD_LOGIC;
  SIGNAL and_dcpl_71 : STD_LOGIC;
  SIGNAL and_dcpl_72 : STD_LOGIC;
  SIGNAL and_dcpl_74 : STD_LOGIC;
  SIGNAL and_dcpl_75 : STD_LOGIC;
  SIGNAL and_dcpl_76 : STD_LOGIC;
  SIGNAL and_dcpl_77 : STD_LOGIC;
  SIGNAL and_dcpl_79 : STD_LOGIC;
  SIGNAL and_dcpl_82 : STD_LOGIC;
  SIGNAL and_dcpl_84 : STD_LOGIC;
  SIGNAL and_dcpl_86 : STD_LOGIC;
  SIGNAL not_tmp_116 : STD_LOGIC;
  SIGNAL and_dcpl_88 : STD_LOGIC;
  SIGNAL and_dcpl_89 : STD_LOGIC;
  SIGNAL and_dcpl_90 : STD_LOGIC;
  SIGNAL and_dcpl_91 : STD_LOGIC;
  SIGNAL and_dcpl_92 : STD_LOGIC;
  SIGNAL and_dcpl_93 : STD_LOGIC;
  SIGNAL or_tmp_131 : STD_LOGIC;
  SIGNAL or_tmp_134 : STD_LOGIC;
  SIGNAL mux_tmp_121 : STD_LOGIC;
  SIGNAL mux_tmp_128 : STD_LOGIC;
  SIGNAL or_tmp_156 : STD_LOGIC;
  SIGNAL and_dcpl_94 : STD_LOGIC;
  SIGNAL and_dcpl_95 : STD_LOGIC;
  SIGNAL and_dcpl_96 : STD_LOGIC;
  SIGNAL and_dcpl_97 : STD_LOGIC;
  SIGNAL and_dcpl_98 : STD_LOGIC;
  SIGNAL and_dcpl_99 : STD_LOGIC;
  SIGNAL or_tmp_166 : STD_LOGIC;
  SIGNAL mux_tmp_139 : STD_LOGIC;
  SIGNAL and_dcpl_100 : STD_LOGIC;
  SIGNAL and_dcpl_101 : STD_LOGIC;
  SIGNAL and_dcpl_102 : STD_LOGIC;
  SIGNAL and_dcpl_103 : STD_LOGIC;
  SIGNAL and_dcpl_105 : STD_LOGIC;
  SIGNAL or_tmp_169 : STD_LOGIC;
  SIGNAL and_dcpl_107 : STD_LOGIC;
  SIGNAL and_dcpl_108 : STD_LOGIC;
  SIGNAL and_dcpl_109 : STD_LOGIC;
  SIGNAL and_dcpl_110 : STD_LOGIC;
  SIGNAL and_dcpl_111 : STD_LOGIC;
  SIGNAL and_dcpl_112 : STD_LOGIC;
  SIGNAL and_dcpl_113 : STD_LOGIC;
  SIGNAL or_tmp_170 : STD_LOGIC;
  SIGNAL and_dcpl_114 : STD_LOGIC;
  SIGNAL and_dcpl_115 : STD_LOGIC;
  SIGNAL and_dcpl_116 : STD_LOGIC;
  SIGNAL and_dcpl_117 : STD_LOGIC;
  SIGNAL and_dcpl_119 : STD_LOGIC;
  SIGNAL and_dcpl_121 : STD_LOGIC;
  SIGNAL and_dcpl_123 : STD_LOGIC;
  SIGNAL and_dcpl_125 : STD_LOGIC;
  SIGNAL and_dcpl_126 : STD_LOGIC;
  SIGNAL and_dcpl_127 : STD_LOGIC;
  SIGNAL and_dcpl_128 : STD_LOGIC;
  SIGNAL and_dcpl_129 : STD_LOGIC;
  SIGNAL and_dcpl_130 : STD_LOGIC;
  SIGNAL and_dcpl_131 : STD_LOGIC;
  SIGNAL nor_tmp_31 : STD_LOGIC;
  SIGNAL and_dcpl_135 : STD_LOGIC;
  SIGNAL and_dcpl_136 : STD_LOGIC;
  SIGNAL and_dcpl_137 : STD_LOGIC;
  SIGNAL nor_tmp_35 : STD_LOGIC;
  SIGNAL nor_tmp_36 : STD_LOGIC;
  SIGNAL and_dcpl_140 : STD_LOGIC;
  SIGNAL and_dcpl_141 : STD_LOGIC;
  SIGNAL and_dcpl_142 : STD_LOGIC;
  SIGNAL not_tmp_149 : STD_LOGIC;
  SIGNAL or_dcpl_177 : STD_LOGIC;
  SIGNAL or_dcpl_178 : STD_LOGIC;
  SIGNAL or_dcpl_179 : STD_LOGIC;
  SIGNAL or_dcpl_180 : STD_LOGIC;
  SIGNAL or_tmp_207 : STD_LOGIC;
  SIGNAL mux_tmp_186 : STD_LOGIC;
  SIGNAL and_dcpl_148 : STD_LOGIC;
  SIGNAL and_dcpl_149 : STD_LOGIC;
  SIGNAL and_dcpl_151 : STD_LOGIC;
  SIGNAL and_dcpl_152 : STD_LOGIC;
  SIGNAL mux_tmp_193 : STD_LOGIC;
  SIGNAL and_dcpl_154 : STD_LOGIC;
  SIGNAL and_dcpl_155 : STD_LOGIC;
  SIGNAL and_dcpl_157 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_162 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL or_tmp_245 : STD_LOGIC;
  SIGNAL or_tmp_246 : STD_LOGIC;
  SIGNAL not_tmp_169 : STD_LOGIC;
  SIGNAL and_dcpl_168 : STD_LOGIC;
  SIGNAL or_dcpl_181 : STD_LOGIC;
  SIGNAL or_dcpl_182 : STD_LOGIC;
  SIGNAL or_tmp_263 : STD_LOGIC;
  SIGNAL mux_tmp_231 : STD_LOGIC;
  SIGNAL and_dcpl_170 : STD_LOGIC;
  SIGNAL and_dcpl_171 : STD_LOGIC;
  SIGNAL and_dcpl_173 : STD_LOGIC;
  SIGNAL and_dcpl_174 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_177 : STD_LOGIC;
  SIGNAL and_dcpl_178 : STD_LOGIC;
  SIGNAL and_dcpl_179 : STD_LOGIC;
  SIGNAL and_dcpl_180 : STD_LOGIC;
  SIGNAL or_tmp_301 : STD_LOGIC;
  SIGNAL not_tmp_188 : STD_LOGIC;
  SIGNAL or_dcpl_183 : STD_LOGIC;
  SIGNAL or_dcpl_184 : STD_LOGIC;
  SIGNAL or_tmp_317 : STD_LOGIC;
  SIGNAL and_dcpl_184 : STD_LOGIC;
  SIGNAL and_dcpl_187 : STD_LOGIC;
  SIGNAL and_dcpl_188 : STD_LOGIC;
  SIGNAL and_dcpl_190 : STD_LOGIC;
  SIGNAL and_dcpl_191 : STD_LOGIC;
  SIGNAL and_dcpl_192 : STD_LOGIC;
  SIGNAL mux_tmp_302 : STD_LOGIC;
  SIGNAL not_tmp_209 : STD_LOGIC;
  SIGNAL or_dcpl_185 : STD_LOGIC;
  SIGNAL or_tmp_362 : STD_LOGIC;
  SIGNAL or_tmp_365 : STD_LOGIC;
  SIGNAL mux_tmp_340 : STD_LOGIC;
  SIGNAL mux_tmp_347 : STD_LOGIC;
  SIGNAL or_tmp_386 : STD_LOGIC;
  SIGNAL and_dcpl_199 : STD_LOGIC;
  SIGNAL and_dcpl_201 : STD_LOGIC;
  SIGNAL and_dcpl_203 : STD_LOGIC;
  SIGNAL nor_tmp_96 : STD_LOGIC;
  SIGNAL and_dcpl_206 : STD_LOGIC;
  SIGNAL and_dcpl_207 : STD_LOGIC;
  SIGNAL or_dcpl_186 : STD_LOGIC;
  SIGNAL or_dcpl_187 : STD_LOGIC;
  SIGNAL or_dcpl_188 : STD_LOGIC;
  SIGNAL mux_tmp_391 : STD_LOGIC;
  SIGNAL mux_tmp_403 : STD_LOGIC;
  SIGNAL and_dcpl_213 : STD_LOGIC;
  SIGNAL and_dcpl_215 : STD_LOGIC;
  SIGNAL and_dcpl_216 : STD_LOGIC;
  SIGNAL and_dcpl_220 : STD_LOGIC;
  SIGNAL or_dcpl_189 : STD_LOGIC;
  SIGNAL or_tmp_493 : STD_LOGIC;
  SIGNAL mux_tmp_445 : STD_LOGIC;
  SIGNAL and_dcpl_224 : STD_LOGIC;
  SIGNAL or_dcpl_190 : STD_LOGIC;
  SIGNAL or_dcpl_191 : STD_LOGIC;
  SIGNAL or_tmp_545 : STD_LOGIC;
  SIGNAL and_dcpl_230 : STD_LOGIC;
  SIGNAL mux_tmp_516 : STD_LOGIC;
  SIGNAL or_dcpl_192 : STD_LOGIC;
  SIGNAL or_tmp_595 : STD_LOGIC;
  SIGNAL or_tmp_598 : STD_LOGIC;
  SIGNAL mux_tmp_549 : STD_LOGIC;
  SIGNAL mux_tmp_556 : STD_LOGIC;
  SIGNAL or_tmp_620 : STD_LOGIC;
  SIGNAL and_dcpl_236 : STD_LOGIC;
  SIGNAL and_dcpl_237 : STD_LOGIC;
  SIGNAL and_dcpl_239 : STD_LOGIC;
  SIGNAL and_dcpl_241 : STD_LOGIC;
  SIGNAL and_dcpl_242 : STD_LOGIC;
  SIGNAL nor_tmp_165 : STD_LOGIC;
  SIGNAL and_dcpl_245 : STD_LOGIC;
  SIGNAL or_dcpl_193 : STD_LOGIC;
  SIGNAL or_dcpl_194 : STD_LOGIC;
  SIGNAL mux_tmp_609 : STD_LOGIC;
  SIGNAL and_dcpl_250 : STD_LOGIC;
  SIGNAL and_dcpl_252 : STD_LOGIC;
  SIGNAL and_dcpl_254 : STD_LOGIC;
  SIGNAL and_dcpl_255 : STD_LOGIC;
  SIGNAL and_dcpl_257 : STD_LOGIC;
  SIGNAL and_dcpl_259 : STD_LOGIC;
  SIGNAL or_dcpl_195 : STD_LOGIC;
  SIGNAL or_dcpl_196 : STD_LOGIC;
  SIGNAL mux_tmp_651 : STD_LOGIC;
  SIGNAL and_dcpl_262 : STD_LOGIC;
  SIGNAL and_dcpl_263 : STD_LOGIC;
  SIGNAL and_dcpl_265 : STD_LOGIC;
  SIGNAL or_dcpl_197 : STD_LOGIC;
  SIGNAL or_tmp_759 : STD_LOGIC;
  SIGNAL and_dcpl_270 : STD_LOGIC;
  SIGNAL and_dcpl_272 : STD_LOGIC;
  SIGNAL mux_tmp_719 : STD_LOGIC;
  SIGNAL or_dcpl_198 : STD_LOGIC;
  SIGNAL or_tmp_806 : STD_LOGIC;
  SIGNAL or_tmp_809 : STD_LOGIC;
  SIGNAL mux_tmp_755 : STD_LOGIC;
  SIGNAL mux_tmp_762 : STD_LOGIC;
  SIGNAL or_tmp_830 : STD_LOGIC;
  SIGNAL and_dcpl_279 : STD_LOGIC;
  SIGNAL and_dcpl_281 : STD_LOGIC;
  SIGNAL nor_tmp_225 : STD_LOGIC;
  SIGNAL or_dcpl_199 : STD_LOGIC;
  SIGNAL or_tmp_875 : STD_LOGIC;
  SIGNAL not_tmp_389 : STD_LOGIC;
  SIGNAL mux_tmp_815 : STD_LOGIC;
  SIGNAL and_dcpl_289 : STD_LOGIC;
  SIGNAL and_dcpl_291 : STD_LOGIC;
  SIGNAL and_dcpl_293 : STD_LOGIC;
  SIGNAL and_dcpl_295 : STD_LOGIC;
  SIGNAL or_dcpl_200 : STD_LOGIC;
  SIGNAL or_tmp_931 : STD_LOGIC;
  SIGNAL mux_tmp_857 : STD_LOGIC;
  SIGNAL and_dcpl_299 : STD_LOGIC;
  SIGNAL or_dcpl_201 : STD_LOGIC;
  SIGNAL or_tmp_982 : STD_LOGIC;
  SIGNAL and_dcpl_305 : STD_LOGIC;
  SIGNAL mux_tmp_928 : STD_LOGIC;
  SIGNAL or_dcpl_202 : STD_LOGIC;
  SIGNAL or_tmp_1030 : STD_LOGIC;
  SIGNAL or_tmp_1033 : STD_LOGIC;
  SIGNAL mux_tmp_962 : STD_LOGIC;
  SIGNAL mux_tmp_969 : STD_LOGIC;
  SIGNAL or_tmp_1054 : STD_LOGIC;
  SIGNAL not_tmp_451 : STD_LOGIC;
  SIGNAL and_dcpl_312 : STD_LOGIC;
  SIGNAL and_dcpl_314 : STD_LOGIC;
  SIGNAL or_tmp_1079 : STD_LOGIC;
  SIGNAL and_dcpl_316 : STD_LOGIC;
  SIGNAL nor_tmp_299 : STD_LOGIC;
  SIGNAL and_dcpl_319 : STD_LOGIC;
  SIGNAL or_dcpl_203 : STD_LOGIC;
  SIGNAL or_dcpl_204 : STD_LOGIC;
  SIGNAL or_dcpl_205 : STD_LOGIC;
  SIGNAL or_tmp_1110 : STD_LOGIC;
  SIGNAL mux_tmp_1025 : STD_LOGIC;
  SIGNAL and_dcpl_325 : STD_LOGIC;
  SIGNAL or_tmp_1133 : STD_LOGIC;
  SIGNAL and_dcpl_327 : STD_LOGIC;
  SIGNAL and_dcpl_328 : STD_LOGIC;
  SIGNAL and_dcpl_330 : STD_LOGIC;
  SIGNAL and_dcpl_332 : STD_LOGIC;
  SIGNAL or_dcpl_206 : STD_LOGIC;
  SIGNAL mux_tmp_1069 : STD_LOGIC;
  SIGNAL or_tmp_1162 : STD_LOGIC;
  SIGNAL and_dcpl_336 : STD_LOGIC;
  SIGNAL or_tmp_1185 : STD_LOGIC;
  SIGNAL or_dcpl_207 : STD_LOGIC;
  SIGNAL or_dcpl_208 : STD_LOGIC;
  SIGNAL or_tmp_1200 : STD_LOGIC;
  SIGNAL or_tmp_1212 : STD_LOGIC;
  SIGNAL and_dcpl_342 : STD_LOGIC;
  SIGNAL mux_tmp_1142 : STD_LOGIC;
  SIGNAL or_tmp_1235 : STD_LOGIC;
  SIGNAL or_dcpl_209 : STD_LOGIC;
  SIGNAL or_tmp_1248 : STD_LOGIC;
  SIGNAL or_tmp_1251 : STD_LOGIC;
  SIGNAL mux_tmp_1179 : STD_LOGIC;
  SIGNAL mux_tmp_1186 : STD_LOGIC;
  SIGNAL or_tmp_1271 : STD_LOGIC;
  SIGNAL not_tmp_542 : STD_LOGIC;
  SIGNAL and_dcpl_349 : STD_LOGIC;
  SIGNAL and_dcpl_351 : STD_LOGIC;
  SIGNAL not_tmp_551 : STD_LOGIC;
  SIGNAL or_tmp_1298 : STD_LOGIC;
  SIGNAL nor_tmp_366 : STD_LOGIC;
  SIGNAL and_dcpl_355 : STD_LOGIC;
  SIGNAL or_dcpl_210 : STD_LOGIC;
  SIGNAL or_dcpl_211 : STD_LOGIC;
  SIGNAL or_dcpl_212 : STD_LOGIC;
  SIGNAL or_tmp_1316 : STD_LOGIC;
  SIGNAL or_tmp_1319 : STD_LOGIC;
  SIGNAL or_tmp_1324 : STD_LOGIC;
  SIGNAL or_tmp_1340 : STD_LOGIC;
  SIGNAL mux_tmp_1243 : STD_LOGIC;
  SIGNAL and_dcpl_361 : STD_LOGIC;
  SIGNAL or_tmp_1363 : STD_LOGIC;
  SIGNAL and_dcpl_363 : STD_LOGIC;
  SIGNAL and_dcpl_365 : STD_LOGIC;
  SIGNAL and_dcpl_367 : STD_LOGIC;
  SIGNAL or_dcpl_213 : STD_LOGIC;
  SIGNAL or_tmp_1379 : STD_LOGIC;
  SIGNAL not_tmp_590 : STD_LOGIC;
  SIGNAL mux_tmp_1287 : STD_LOGIC;
  SIGNAL or_tmp_1397 : STD_LOGIC;
  SIGNAL not_tmp_598 : STD_LOGIC;
  SIGNAL and_dcpl_371 : STD_LOGIC;
  SIGNAL or_tmp_1422 : STD_LOGIC;
  SIGNAL or_dcpl_214 : STD_LOGIC;
  SIGNAL or_dcpl_215 : STD_LOGIC;
  SIGNAL or_tmp_1437 : STD_LOGIC;
  SIGNAL or_tmp_1452 : STD_LOGIC;
  SIGNAL and_dcpl_377 : STD_LOGIC;
  SIGNAL mux_tmp_1363 : STD_LOGIC;
  SIGNAL or_tmp_1479 : STD_LOGIC;
  SIGNAL or_dcpl_216 : STD_LOGIC;
  SIGNAL or_tmp_1492 : STD_LOGIC;
  SIGNAL or_tmp_1495 : STD_LOGIC;
  SIGNAL mux_tmp_1397 : STD_LOGIC;
  SIGNAL mux_tmp_1404 : STD_LOGIC;
  SIGNAL or_tmp_1516 : STD_LOGIC;
  SIGNAL and_dcpl_384 : STD_LOGIC;
  SIGNAL or_tmp_1540 : STD_LOGIC;
  SIGNAL nor_tmp_445 : STD_LOGIC;
  SIGNAL or_dcpl_217 : STD_LOGIC;
  SIGNAL or_tmp_1558 : STD_LOGIC;
  SIGNAL or_tmp_1572 : STD_LOGIC;
  SIGNAL mux_tmp_1460 : STD_LOGIC;
  SIGNAL and_dcpl_393 : STD_LOGIC;
  SIGNAL or_tmp_1595 : STD_LOGIC;
  SIGNAL and_dcpl_395 : STD_LOGIC;
  SIGNAL and_dcpl_396 : STD_LOGIC;
  SIGNAL and_dcpl_398 : STD_LOGIC;
  SIGNAL and_dcpl_400 : STD_LOGIC;
  SIGNAL or_dcpl_218 : STD_LOGIC;
  SIGNAL or_tmp_1610 : STD_LOGIC;
  SIGNAL mux_tmp_1504 : STD_LOGIC;
  SIGNAL or_tmp_1624 : STD_LOGIC;
  SIGNAL and_dcpl_404 : STD_LOGIC;
  SIGNAL or_tmp_1647 : STD_LOGIC;
  SIGNAL or_dcpl_219 : STD_LOGIC;
  SIGNAL or_tmp_1662 : STD_LOGIC;
  SIGNAL or_tmp_1677 : STD_LOGIC;
  SIGNAL and_dcpl_410 : STD_LOGIC;
  SIGNAL mux_tmp_1577 : STD_LOGIC;
  SIGNAL or_tmp_1703 : STD_LOGIC;
  SIGNAL or_dcpl_220 : STD_LOGIC;
  SIGNAL or_tmp_1716 : STD_LOGIC;
  SIGNAL or_tmp_1719 : STD_LOGIC;
  SIGNAL mux_tmp_1614 : STD_LOGIC;
  SIGNAL mux_tmp_1621 : STD_LOGIC;
  SIGNAL or_tmp_1739 : STD_LOGIC;
  SIGNAL and_dcpl_417 : STD_LOGIC;
  SIGNAL not_tmp_741 : STD_LOGIC;
  SIGNAL or_tmp_1765 : STD_LOGIC;
  SIGNAL nor_tmp_525 : STD_LOGIC;
  SIGNAL or_dcpl_221 : STD_LOGIC;
  SIGNAL or_tmp_1783 : STD_LOGIC;
  SIGNAL or_tmp_1796 : STD_LOGIC;
  SIGNAL mux_tmp_1677 : STD_LOGIC;
  SIGNAL and_dcpl_426 : STD_LOGIC;
  SIGNAL or_tmp_1818 : STD_LOGIC;
  SIGNAL and_dcpl_428 : STD_LOGIC;
  SIGNAL and_dcpl_430 : STD_LOGIC;
  SIGNAL and_dcpl_432 : STD_LOGIC;
  SIGNAL or_dcpl_222 : STD_LOGIC;
  SIGNAL or_tmp_1833 : STD_LOGIC;
  SIGNAL mux_tmp_1721 : STD_LOGIC;
  SIGNAL or_tmp_1845 : STD_LOGIC;
  SIGNAL and_dcpl_436 : STD_LOGIC;
  SIGNAL or_tmp_1867 : STD_LOGIC;
  SIGNAL or_dcpl_223 : STD_LOGIC;
  SIGNAL and_dcpl_442 : STD_LOGIC;
  SIGNAL mux_tmp_1793 : STD_LOGIC;
  SIGNAL mux_tmp_1820 : STD_LOGIC;
  SIGNAL mux_tmp_1821 : STD_LOGIC;
  SIGNAL or_tmp_1918 : STD_LOGIC;
  SIGNAL or_tmp_1924 : STD_LOGIC;
  SIGNAL mux_tmp_1832 : STD_LOGIC;
  SIGNAL or_tmp_1928 : STD_LOGIC;
  SIGNAL and_dcpl_447 : STD_LOGIC;
  SIGNAL and_dcpl_448 : STD_LOGIC;
  SIGNAL and_dcpl_449 : STD_LOGIC;
  SIGNAL and_dcpl_450 : STD_LOGIC;
  SIGNAL and_dcpl_451 : STD_LOGIC;
  SIGNAL not_tmp_833 : STD_LOGIC;
  SIGNAL and_dcpl_454 : STD_LOGIC;
  SIGNAL and_dcpl_456 : STD_LOGIC;
  SIGNAL and_dcpl_457 : STD_LOGIC;
  SIGNAL and_dcpl_458 : STD_LOGIC;
  SIGNAL and_dcpl_459 : STD_LOGIC;
  SIGNAL and_dcpl_460 : STD_LOGIC;
  SIGNAL and_dcpl_461 : STD_LOGIC;
  SIGNAL and_dcpl_462 : STD_LOGIC;
  SIGNAL and_dcpl_464 : STD_LOGIC;
  SIGNAL and_dcpl_466 : STD_LOGIC;
  SIGNAL and_dcpl_467 : STD_LOGIC;
  SIGNAL and_dcpl_468 : STD_LOGIC;
  SIGNAL and_dcpl_469 : STD_LOGIC;
  SIGNAL and_dcpl_470 : STD_LOGIC;
  SIGNAL and_dcpl_472 : STD_LOGIC;
  SIGNAL and_dcpl_475 : STD_LOGIC;
  SIGNAL and_dcpl_476 : STD_LOGIC;
  SIGNAL and_dcpl_477 : STD_LOGIC;
  SIGNAL and_dcpl_478 : STD_LOGIC;
  SIGNAL and_dcpl_479 : STD_LOGIC;
  SIGNAL and_dcpl_480 : STD_LOGIC;
  SIGNAL and_dcpl_483 : STD_LOGIC;
  SIGNAL and_dcpl_484 : STD_LOGIC;
  SIGNAL not_tmp_843 : STD_LOGIC;
  SIGNAL and_dcpl_488 : STD_LOGIC;
  SIGNAL and_dcpl_489 : STD_LOGIC;
  SIGNAL and_dcpl_490 : STD_LOGIC;
  SIGNAL and_dcpl_492 : STD_LOGIC;
  SIGNAL and_dcpl_493 : STD_LOGIC;
  SIGNAL and_dcpl_494 : STD_LOGIC;
  SIGNAL and_dcpl_497 : STD_LOGIC;
  SIGNAL and_dcpl_499 : STD_LOGIC;
  SIGNAL and_dcpl_501 : STD_LOGIC;
  SIGNAL and_dcpl_503 : STD_LOGIC;
  SIGNAL or_dcpl_225 : STD_LOGIC;
  SIGNAL or_dcpl_226 : STD_LOGIC;
  SIGNAL or_dcpl_227 : STD_LOGIC;
  SIGNAL or_tmp_1976 : STD_LOGIC;
  SIGNAL mux_tmp_1887 : STD_LOGIC;
  SIGNAL or_tmp_1981 : STD_LOGIC;
  SIGNAL or_tmp_1983 : STD_LOGIC;
  SIGNAL and_dcpl_506 : STD_LOGIC;
  SIGNAL and_dcpl_507 : STD_LOGIC;
  SIGNAL and_dcpl_508 : STD_LOGIC;
  SIGNAL and_dcpl_510 : STD_LOGIC;
  SIGNAL and_dcpl_511 : STD_LOGIC;
  SIGNAL not_tmp_865 : STD_LOGIC;
  SIGNAL and_dcpl_519 : STD_LOGIC;
  SIGNAL and_dcpl_521 : STD_LOGIC;
  SIGNAL and_dcpl_522 : STD_LOGIC;
  SIGNAL and_dcpl_523 : STD_LOGIC;
  SIGNAL and_dcpl_525 : STD_LOGIC;
  SIGNAL and_dcpl_526 : STD_LOGIC;
  SIGNAL and_dcpl_528 : STD_LOGIC;
  SIGNAL or_dcpl_229 : STD_LOGIC;
  SIGNAL mux_tmp_1938 : STD_LOGIC;
  SIGNAL or_tmp_2035 : STD_LOGIC;
  SIGNAL and_dcpl_533 : STD_LOGIC;
  SIGNAL and_dcpl_534 : STD_LOGIC;
  SIGNAL and_dcpl_535 : STD_LOGIC;
  SIGNAL and_dcpl_536 : STD_LOGIC;
  SIGNAL and_dcpl_537 : STD_LOGIC;
  SIGNAL and_dcpl_540 : STD_LOGIC;
  SIGNAL and_dcpl_541 : STD_LOGIC;
  SIGNAL mux_tmp_1958 : STD_LOGIC;
  SIGNAL not_tmp_874 : STD_LOGIC;
  SIGNAL and_dcpl_544 : STD_LOGIC;
  SIGNAL and_dcpl_546 : STD_LOGIC;
  SIGNAL and_dcpl_548 : STD_LOGIC;
  SIGNAL or_dcpl_231 : STD_LOGIC;
  SIGNAL or_tmp_2071 : STD_LOGIC;
  SIGNAL or_tmp_2075 : STD_LOGIC;
  SIGNAL or_tmp_2076 : STD_LOGIC;
  SIGNAL mux_tmp_1996 : STD_LOGIC;
  SIGNAL mux_tmp_1999 : STD_LOGIC;
  SIGNAL and_dcpl_551 : STD_LOGIC;
  SIGNAL and_dcpl_552 : STD_LOGIC;
  SIGNAL and_dcpl_553 : STD_LOGIC;
  SIGNAL and_dcpl_556 : STD_LOGIC;
  SIGNAL and_dcpl_557 : STD_LOGIC;
  SIGNAL mux_tmp_2019 : STD_LOGIC;
  SIGNAL and_dcpl_559 : STD_LOGIC;
  SIGNAL nor_tmp_674 : STD_LOGIC;
  SIGNAL not_tmp_890 : STD_LOGIC;
  SIGNAL and_dcpl_564 : STD_LOGIC;
  SIGNAL or_dcpl_233 : STD_LOGIC;
  SIGNAL mux_tmp_2052 : STD_LOGIC;
  SIGNAL mux_tmp_2053 : STD_LOGIC;
  SIGNAL or_tmp_2119 : STD_LOGIC;
  SIGNAL or_tmp_2122 : STD_LOGIC;
  SIGNAL mux_tmp_2064 : STD_LOGIC;
  SIGNAL or_tmp_2126 : STD_LOGIC;
  SIGNAL and_dcpl_567 : STD_LOGIC;
  SIGNAL and_dcpl_568 : STD_LOGIC;
  SIGNAL and_dcpl_569 : STD_LOGIC;
  SIGNAL and_dcpl_570 : STD_LOGIC;
  SIGNAL and_dcpl_574 : STD_LOGIC;
  SIGNAL and_dcpl_577 : STD_LOGIC;
  SIGNAL and_dcpl_578 : STD_LOGIC;
  SIGNAL and_dcpl_580 : STD_LOGIC;
  SIGNAL and_dcpl_581 : STD_LOGIC;
  SIGNAL and_dcpl_585 : STD_LOGIC;
  SIGNAL or_dcpl_235 : STD_LOGIC;
  SIGNAL or_dcpl_236 : STD_LOGIC;
  SIGNAL or_tmp_2168 : STD_LOGIC;
  SIGNAL mux_tmp_2115 : STD_LOGIC;
  SIGNAL or_tmp_2176 : STD_LOGIC;
  SIGNAL or_tmp_2179 : STD_LOGIC;
  SIGNAL and_dcpl_588 : STD_LOGIC;
  SIGNAL and_dcpl_594 : STD_LOGIC;
  SIGNAL and_dcpl_596 : STD_LOGIC;
  SIGNAL mux_tmp_2163 : STD_LOGIC;
  SIGNAL or_tmp_2228 : STD_LOGIC;
  SIGNAL and_dcpl_599 : STD_LOGIC;
  SIGNAL and_dcpl_600 : STD_LOGIC;
  SIGNAL mux_tmp_2187 : STD_LOGIC;
  SIGNAL and_dcpl_605 : STD_LOGIC;
  SIGNAL or_tmp_2259 : STD_LOGIC;
  SIGNAL or_tmp_2265 : STD_LOGIC;
  SIGNAL or_tmp_2266 : STD_LOGIC;
  SIGNAL mux_tmp_2219 : STD_LOGIC;
  SIGNAL mux_tmp_2222 : STD_LOGIC;
  SIGNAL and_dcpl_609 : STD_LOGIC;
  SIGNAL mux_tmp_2245 : STD_LOGIC;
  SIGNAL and_dcpl_613 : STD_LOGIC;
  SIGNAL mux_tmp_2272 : STD_LOGIC;
  SIGNAL mux_tmp_2273 : STD_LOGIC;
  SIGNAL or_tmp_2300 : STD_LOGIC;
  SIGNAL or_tmp_2306 : STD_LOGIC;
  SIGNAL mux_tmp_2284 : STD_LOGIC;
  SIGNAL or_tmp_2310 : STD_LOGIC;
  SIGNAL and_dcpl_619 : STD_LOGIC;
  SIGNAL and_dcpl_620 : STD_LOGIC;
  SIGNAL and_dcpl_621 : STD_LOGIC;
  SIGNAL and_dcpl_622 : STD_LOGIC;
  SIGNAL and_dcpl_626 : STD_LOGIC;
  SIGNAL and_dcpl_629 : STD_LOGIC;
  SIGNAL and_dcpl_631 : STD_LOGIC;
  SIGNAL and_dcpl_634 : STD_LOGIC;
  SIGNAL and_dcpl_635 : STD_LOGIC;
  SIGNAL and_dcpl_637 : STD_LOGIC;
  SIGNAL or_dcpl_241 : STD_LOGIC;
  SIGNAL or_tmp_2348 : STD_LOGIC;
  SIGNAL mux_tmp_2335 : STD_LOGIC;
  SIGNAL or_tmp_2353 : STD_LOGIC;
  SIGNAL or_tmp_2355 : STD_LOGIC;
  SIGNAL and_dcpl_640 : STD_LOGIC;
  SIGNAL and_dcpl_646 : STD_LOGIC;
  SIGNAL and_dcpl_648 : STD_LOGIC;
  SIGNAL and_dcpl_650 : STD_LOGIC;
  SIGNAL mux_tmp_2383 : STD_LOGIC;
  SIGNAL or_tmp_2398 : STD_LOGIC;
  SIGNAL and_dcpl_653 : STD_LOGIC;
  SIGNAL and_dcpl_654 : STD_LOGIC;
  SIGNAL and_dcpl_655 : STD_LOGIC;
  SIGNAL mux_tmp_2403 : STD_LOGIC;
  SIGNAL and_dcpl_660 : STD_LOGIC;
  SIGNAL and_dcpl_662 : STD_LOGIC;
  SIGNAL and_dcpl_664 : STD_LOGIC;
  SIGNAL or_tmp_2428 : STD_LOGIC;
  SIGNAL or_tmp_2432 : STD_LOGIC;
  SIGNAL or_tmp_2433 : STD_LOGIC;
  SIGNAL mux_tmp_2439 : STD_LOGIC;
  SIGNAL mux_tmp_2442 : STD_LOGIC;
  SIGNAL and_dcpl_667 : STD_LOGIC;
  SIGNAL mux_tmp_2461 : STD_LOGIC;
  SIGNAL and_dcpl_675 : STD_LOGIC;
  SIGNAL mux_tmp_2492 : STD_LOGIC;
  SIGNAL mux_tmp_2493 : STD_LOGIC;
  SIGNAL or_tmp_2469 : STD_LOGIC;
  SIGNAL or_tmp_2472 : STD_LOGIC;
  SIGNAL mux_tmp_2504 : STD_LOGIC;
  SIGNAL or_tmp_2476 : STD_LOGIC;
  SIGNAL and_dcpl_678 : STD_LOGIC;
  SIGNAL and_dcpl_679 : STD_LOGIC;
  SIGNAL and_dcpl_683 : STD_LOGIC;
  SIGNAL and_dcpl_686 : STD_LOGIC;
  SIGNAL or_dcpl_246 : STD_LOGIC;
  SIGNAL or_tmp_2518 : STD_LOGIC;
  SIGNAL mux_tmp_2555 : STD_LOGIC;
  SIGNAL or_tmp_2526 : STD_LOGIC;
  SIGNAL or_tmp_2529 : STD_LOGIC;
  SIGNAL and_dcpl_692 : STD_LOGIC;
  SIGNAL and_dcpl_699 : STD_LOGIC;
  SIGNAL mux_tmp_2603 : STD_LOGIC;
  SIGNAL or_tmp_2578 : STD_LOGIC;
  SIGNAL and_dcpl_702 : STD_LOGIC;
  SIGNAL and_dcpl_703 : STD_LOGIC;
  SIGNAL mux_tmp_2627 : STD_LOGIC;
  SIGNAL and_dcpl_708 : STD_LOGIC;
  SIGNAL or_tmp_2609 : STD_LOGIC;
  SIGNAL or_tmp_2615 : STD_LOGIC;
  SIGNAL or_tmp_2616 : STD_LOGIC;
  SIGNAL mux_tmp_2659 : STD_LOGIC;
  SIGNAL mux_tmp_2662 : STD_LOGIC;
  SIGNAL and_dcpl_712 : STD_LOGIC;
  SIGNAL mux_tmp_2685 : STD_LOGIC;
  SIGNAL mux_tmp_2712 : STD_LOGIC;
  SIGNAL mux_tmp_2713 : STD_LOGIC;
  SIGNAL or_tmp_2656 : STD_LOGIC;
  SIGNAL or_tmp_2663 : STD_LOGIC;
  SIGNAL mux_tmp_2723 : STD_LOGIC;
  SIGNAL or_tmp_2666 : STD_LOGIC;
  SIGNAL and_dcpl_721 : STD_LOGIC;
  SIGNAL and_dcpl_722 : STD_LOGIC;
  SIGNAL and_dcpl_723 : STD_LOGIC;
  SIGNAL and_dcpl_724 : STD_LOGIC;
  SIGNAL and_dcpl_728 : STD_LOGIC;
  SIGNAL and_dcpl_731 : STD_LOGIC;
  SIGNAL and_dcpl_733 : STD_LOGIC;
  SIGNAL and_dcpl_736 : STD_LOGIC;
  SIGNAL and_dcpl_737 : STD_LOGIC;
  SIGNAL and_dcpl_739 : STD_LOGIC;
  SIGNAL or_dcpl_251 : STD_LOGIC;
  SIGNAL or_dcpl_252 : STD_LOGIC;
  SIGNAL or_tmp_2710 : STD_LOGIC;
  SIGNAL mux_tmp_2775 : STD_LOGIC;
  SIGNAL or_tmp_2716 : STD_LOGIC;
  SIGNAL or_tmp_2717 : STD_LOGIC;
  SIGNAL and_dcpl_742 : STD_LOGIC;
  SIGNAL and_dcpl_748 : STD_LOGIC;
  SIGNAL and_dcpl_749 : STD_LOGIC;
  SIGNAL and_dcpl_751 : STD_LOGIC;
  SIGNAL and_dcpl_753 : STD_LOGIC;
  SIGNAL mux_tmp_2823 : STD_LOGIC;
  SIGNAL or_tmp_2765 : STD_LOGIC;
  SIGNAL and_dcpl_756 : STD_LOGIC;
  SIGNAL and_dcpl_757 : STD_LOGIC;
  SIGNAL and_dcpl_758 : STD_LOGIC;
  SIGNAL mux_tmp_2843 : STD_LOGIC;
  SIGNAL and_dcpl_763 : STD_LOGIC;
  SIGNAL and_dcpl_765 : STD_LOGIC;
  SIGNAL and_dcpl_767 : STD_LOGIC;
  SIGNAL or_tmp_2802 : STD_LOGIC;
  SIGNAL or_tmp_2806 : STD_LOGIC;
  SIGNAL or_tmp_2808 : STD_LOGIC;
  SIGNAL mux_tmp_2879 : STD_LOGIC;
  SIGNAL mux_tmp_2880 : STD_LOGIC;
  SIGNAL and_dcpl_770 : STD_LOGIC;
  SIGNAL mux_tmp_2901 : STD_LOGIC;
  SIGNAL and_dcpl_778 : STD_LOGIC;
  SIGNAL mux_tmp_2932 : STD_LOGIC;
  SIGNAL mux_tmp_2933 : STD_LOGIC;
  SIGNAL or_tmp_2855 : STD_LOGIC;
  SIGNAL or_tmp_2858 : STD_LOGIC;
  SIGNAL mux_tmp_2943 : STD_LOGIC;
  SIGNAL or_tmp_2861 : STD_LOGIC;
  SIGNAL and_dcpl_781 : STD_LOGIC;
  SIGNAL and_dcpl_782 : STD_LOGIC;
  SIGNAL and_dcpl_788 : STD_LOGIC;
  SIGNAL and_dcpl_790 : STD_LOGIC;
  SIGNAL or_dcpl_257 : STD_LOGIC;
  SIGNAL or_dcpl_258 : STD_LOGIC;
  SIGNAL or_tmp_2909 : STD_LOGIC;
  SIGNAL mux_tmp_2995 : STD_LOGIC;
  SIGNAL or_tmp_2918 : STD_LOGIC;
  SIGNAL or_tmp_2920 : STD_LOGIC;
  SIGNAL and_dcpl_795 : STD_LOGIC;
  SIGNAL and_dcpl_802 : STD_LOGIC;
  SIGNAL mux_tmp_3043 : STD_LOGIC;
  SIGNAL or_tmp_2974 : STD_LOGIC;
  SIGNAL and_dcpl_805 : STD_LOGIC;
  SIGNAL and_dcpl_806 : STD_LOGIC;
  SIGNAL mux_tmp_3067 : STD_LOGIC;
  SIGNAL and_dcpl_811 : STD_LOGIC;
  SIGNAL or_tmp_3012 : STD_LOGIC;
  SIGNAL or_tmp_3018 : STD_LOGIC;
  SIGNAL or_tmp_3020 : STD_LOGIC;
  SIGNAL mux_tmp_3099 : STD_LOGIC;
  SIGNAL mux_tmp_3100 : STD_LOGIC;
  SIGNAL and_dcpl_815 : STD_LOGIC;
  SIGNAL mux_tmp_3125 : STD_LOGIC;
  SIGNAL not_tmp_1143 : STD_LOGIC;
  SIGNAL mux_tmp_3152 : STD_LOGIC;
  SIGNAL mux_tmp_3153 : STD_LOGIC;
  SIGNAL or_tmp_3064 : STD_LOGIC;
  SIGNAL or_tmp_3071 : STD_LOGIC;
  SIGNAL mux_tmp_3163 : STD_LOGIC;
  SIGNAL or_tmp_3074 : STD_LOGIC;
  SIGNAL and_dcpl_825 : STD_LOGIC;
  SIGNAL and_dcpl_826 : STD_LOGIC;
  SIGNAL and_dcpl_827 : STD_LOGIC;
  SIGNAL and_dcpl_833 : STD_LOGIC;
  SIGNAL and_dcpl_837 : STD_LOGIC;
  SIGNAL and_dcpl_838 : STD_LOGIC;
  SIGNAL and_dcpl_840 : STD_LOGIC;
  SIGNAL or_dcpl_263 : STD_LOGIC;
  SIGNAL or_tmp_3118 : STD_LOGIC;
  SIGNAL mux_tmp_3215 : STD_LOGIC;
  SIGNAL or_tmp_3124 : STD_LOGIC;
  SIGNAL or_tmp_3125 : STD_LOGIC;
  SIGNAL and_dcpl_843 : STD_LOGIC;
  SIGNAL and_dcpl_849 : STD_LOGIC;
  SIGNAL and_dcpl_851 : STD_LOGIC;
  SIGNAL and_dcpl_853 : STD_LOGIC;
  SIGNAL mux_tmp_3263 : STD_LOGIC;
  SIGNAL or_tmp_3173 : STD_LOGIC;
  SIGNAL and_dcpl_856 : STD_LOGIC;
  SIGNAL and_dcpl_857 : STD_LOGIC;
  SIGNAL and_dcpl_858 : STD_LOGIC;
  SIGNAL mux_tmp_3283 : STD_LOGIC;
  SIGNAL and_dcpl_863 : STD_LOGIC;
  SIGNAL and_dcpl_865 : STD_LOGIC;
  SIGNAL and_dcpl_867 : STD_LOGIC;
  SIGNAL or_tmp_3210 : STD_LOGIC;
  SIGNAL or_tmp_3214 : STD_LOGIC;
  SIGNAL or_tmp_3216 : STD_LOGIC;
  SIGNAL mux_tmp_3319 : STD_LOGIC;
  SIGNAL mux_tmp_3320 : STD_LOGIC;
  SIGNAL and_dcpl_870 : STD_LOGIC;
  SIGNAL mux_tmp_3341 : STD_LOGIC;
  SIGNAL and_dcpl_878 : STD_LOGIC;
  SIGNAL not_tmp_1199 : STD_LOGIC;
  SIGNAL mux_tmp_3372 : STD_LOGIC;
  SIGNAL mux_tmp_3373 : STD_LOGIC;
  SIGNAL or_tmp_3261 : STD_LOGIC;
  SIGNAL or_tmp_3264 : STD_LOGIC;
  SIGNAL mux_tmp_3383 : STD_LOGIC;
  SIGNAL or_tmp_3266 : STD_LOGIC;
  SIGNAL and_dcpl_881 : STD_LOGIC;
  SIGNAL and_dcpl_882 : STD_LOGIC;
  SIGNAL and_dcpl_888 : STD_LOGIC;
  SIGNAL or_dcpl_268 : STD_LOGIC;
  SIGNAL nor_tmp_1094 : STD_LOGIC;
  SIGNAL or_tmp_3312 : STD_LOGIC;
  SIGNAL mux_tmp_3435 : STD_LOGIC;
  SIGNAL or_tmp_3320 : STD_LOGIC;
  SIGNAL not_tmp_1218 : STD_LOGIC;
  SIGNAL and_dcpl_894 : STD_LOGIC;
  SIGNAL and_dcpl_901 : STD_LOGIC;
  SIGNAL not_tmp_1235 : STD_LOGIC;
  SIGNAL mux_tmp_3483 : STD_LOGIC;
  SIGNAL not_tmp_1239 : STD_LOGIC;
  SIGNAL and_dcpl_904 : STD_LOGIC;
  SIGNAL and_dcpl_905 : STD_LOGIC;
  SIGNAL mux_tmp_3507 : STD_LOGIC;
  SIGNAL and_dcpl_910 : STD_LOGIC;
  SIGNAL or_tmp_3410 : STD_LOGIC;
  SIGNAL not_tmp_1250 : STD_LOGIC;
  SIGNAL or_tmp_3413 : STD_LOGIC;
  SIGNAL or_tmp_3415 : STD_LOGIC;
  SIGNAL mux_tmp_3539 : STD_LOGIC;
  SIGNAL mux_tmp_3540 : STD_LOGIC;
  SIGNAL nor_tmp_1140 : STD_LOGIC;
  SIGNAL and_dcpl_914 : STD_LOGIC;
  SIGNAL or_dcpl_273 : STD_LOGIC;
  SIGNAL mux_tmp_3565 : STD_LOGIC;
  SIGNAL and_dcpl_924 : STD_LOGIC;
  SIGNAL and_dcpl_925 : STD_LOGIC;
  SIGNAL and_dcpl_927 : STD_LOGIC;
  SIGNAL and_dcpl_932 : STD_LOGIC;
  SIGNAL and_dcpl_934 : STD_LOGIC;
  SIGNAL and_dcpl_935 : STD_LOGIC;
  SIGNAL not_tmp_1278 : STD_LOGIC;
  SIGNAL not_tmp_1311 : STD_LOGIC;
  SIGNAL not_tmp_1328 : STD_LOGIC;
  SIGNAL and_dcpl_1000 : STD_LOGIC;
  SIGNAL and_dcpl_1007 : STD_LOGIC;
  SIGNAL and_dcpl_1008 : STD_LOGIC;
  SIGNAL and_dcpl_1010 : STD_LOGIC;
  SIGNAL or_tmp_3536 : STD_LOGIC;
  SIGNAL or_tmp_3537 : STD_LOGIC;
  SIGNAL or_tmp_3538 : STD_LOGIC;
  SIGNAL or_tmp_3540 : STD_LOGIC;
  SIGNAL mux_tmp_3659 : STD_LOGIC;
  SIGNAL or_tmp_3550 : STD_LOGIC;
  SIGNAL and_dcpl_1011 : STD_LOGIC;
  SIGNAL and_dcpl_1012 : STD_LOGIC;
  SIGNAL and_dcpl_1013 : STD_LOGIC;
  SIGNAL xor_dcpl_1 : STD_LOGIC;
  SIGNAL and_dcpl_1014 : STD_LOGIC;
  SIGNAL not_tmp_1345 : STD_LOGIC;
  SIGNAL not_tmp_1349 : STD_LOGIC;
  SIGNAL and_dcpl_1022 : STD_LOGIC;
  SIGNAL and_dcpl_1023 : STD_LOGIC;
  SIGNAL and_dcpl_1024 : STD_LOGIC;
  SIGNAL and_dcpl_1027 : STD_LOGIC;
  SIGNAL and_dcpl_1031 : STD_LOGIC;
  SIGNAL and_dcpl_1032 : STD_LOGIC;
  SIGNAL and_dcpl_1033 : STD_LOGIC;
  SIGNAL and_dcpl_1035 : STD_LOGIC;
  SIGNAL and_dcpl_1037 : STD_LOGIC;
  SIGNAL and_dcpl_1041 : STD_LOGIC;
  SIGNAL and_dcpl_1044 : STD_LOGIC;
  SIGNAL and_dcpl_1052 : STD_LOGIC;
  SIGNAL and_dcpl_1054 : STD_LOGIC;
  SIGNAL mux_tmp_3698 : STD_LOGIC;
  SIGNAL mux_tmp_3714 : STD_LOGIC;
  SIGNAL and_dcpl_1070 : STD_LOGIC;
  SIGNAL mux_tmp_3730 : STD_LOGIC;
  SIGNAL or_tmp_3658 : STD_LOGIC;
  SIGNAL or_tmp_3661 : STD_LOGIC;
  SIGNAL or_tmp_3662 : STD_LOGIC;
  SIGNAL mux_tmp_3769 : STD_LOGIC;
  SIGNAL and_dcpl_1082 : STD_LOGIC;
  SIGNAL and_dcpl_1083 : STD_LOGIC;
  SIGNAL and_dcpl_1084 : STD_LOGIC;
  SIGNAL or_dcpl_276 : STD_LOGIC;
  SIGNAL or_dcpl_277 : STD_LOGIC;
  SIGNAL and_dcpl_1085 : STD_LOGIC;
  SIGNAL and_dcpl_1086 : STD_LOGIC;
  SIGNAL mux_tmp_3812 : STD_LOGIC;
  SIGNAL and_dcpl_1088 : STD_LOGIC;
  SIGNAL or_tmp_3706 : STD_LOGIC;
  SIGNAL mux_tmp_3819 : STD_LOGIC;
  SIGNAL nor_tmp_1200 : STD_LOGIC;
  SIGNAL and_dcpl_1091 : STD_LOGIC;
  SIGNAL and_dcpl_1092 : STD_LOGIC;
  SIGNAL or_tmp_3740 : STD_LOGIC;
  SIGNAL and_dcpl_1095 : STD_LOGIC;
  SIGNAL not_tmp_1436 : STD_LOGIC;
  SIGNAL and_dcpl_1096 : STD_LOGIC;
  SIGNAL or_tmp_3812 : STD_LOGIC;
  SIGNAL or_tmp_3814 : STD_LOGIC;
  SIGNAL and_dcpl_1097 : STD_LOGIC;
  SIGNAL and_dcpl_1101 : STD_LOGIC;
  SIGNAL and_dcpl_1103 : STD_LOGIC;
  SIGNAL and_dcpl_1105 : STD_LOGIC;
  SIGNAL and_dcpl_1108 : STD_LOGIC;
  SIGNAL and_dcpl_1109 : STD_LOGIC;
  SIGNAL and_dcpl_1110 : STD_LOGIC;
  SIGNAL and_dcpl_1112 : STD_LOGIC;
  SIGNAL and_dcpl_1113 : STD_LOGIC;
  SIGNAL and_dcpl_1114 : STD_LOGIC;
  SIGNAL and_dcpl_1115 : STD_LOGIC;
  SIGNAL and_dcpl_1116 : STD_LOGIC;
  SIGNAL or_tmp_3871 : STD_LOGIC;
  SIGNAL not_tmp_1520 : STD_LOGIC;
  SIGNAL or_tmp_4011 : STD_LOGIC;
  SIGNAL mux_tmp_4062 : STD_LOGIC;
  SIGNAL mux_tmp_4069 : STD_LOGIC;
  SIGNAL and_dcpl_1136 : STD_LOGIC;
  SIGNAL or_tmp_4014 : STD_LOGIC;
  SIGNAL mux_tmp_4075 : STD_LOGIC;
  SIGNAL mux_tmp_4094 : STD_LOGIC;
  SIGNAL or_dcpl_286 : STD_LOGIC;
  SIGNAL or_dcpl_302 : STD_LOGIC;
  SIGNAL operator_20_true_15_slc_operator_20_true_15_acc_14_itm : STD_LOGIC;
  SIGNAL modulo_sub_base_20_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_21_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_23_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_16_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_17_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_19_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_12_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_13_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_14_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_15_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S1_OUTER_LOOP_k_5_0_sva_2 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL operator_20_true_8_slc_operator_20_true_8_acc_14_itm : STD_LOGIC;
  SIGNAL modulo_sub_base_8_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_9_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_10_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_11_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S2_INNER_LOOP1_r_4_0_sva_2 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL modulo_sub_base_4_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_5_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_6_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_7_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_1_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_2_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_3_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_20_true_1_slc_operator_20_true_1_acc_14_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_21_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_53_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_22_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_25_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_61_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_30_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_40_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_35_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_36_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_20_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_51_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_24_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_55_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_57_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_26_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_27_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_59_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_28_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_29_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_60_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_6_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_37_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_42_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_47_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_33_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_39_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_41_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_43_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_44_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_18_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_49_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_1_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_4_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_36_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_44_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_33_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_37_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_45_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_48_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_52_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_56_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_41_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_54_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_58_itm : STD_LOGIC;
  SIGNAL S2_OUTER_LOOP_c_1_sva : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_39_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_25_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_8_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_26_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_3_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_7_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_14_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_2_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_49_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_1_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_43_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_51_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_55_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_35_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_40_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_42_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_47_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_50_itm : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_39_itm : STD_LOGIC;
  SIGNAL modulo_add_13_slc_32_svs_st : STD_LOGIC;
  SIGNAL modulo_add_base_20_sva_mx0w33 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_21_sva_mx0w32 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_22_sva_mx0w31 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_23_sva_mx0w30 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_16_sva_mx0w29 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_17_sva_mx0w28 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_18_sva_mx0w27 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_19_sva_mx0w26 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_12_sva_mx0w24 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_13_sva_mx0w23 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_14_sva_mx0w22 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_15_sva_mx0w21 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_8_sva_mx0w17 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_9_sva_mx0w16 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_10_sva_mx0w15 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_11_sva_mx0w14 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_4_sva_mx0w12 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_5_sva_mx0w11 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_6_sva_mx0w10 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_7_sva_mx0w9 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_sva_mx0w7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_1_sva_mx0w6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_2_sva_mx0w5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_3_sva_mx0w4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S1_OUTER_LOOP_for_p_sva_1 : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL m_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_615_ssc : STD_LOGIC;
  SIGNAL and_616_ssc : STD_LOGIC;
  SIGNAL and_173_ssc : STD_LOGIC;
  SIGNAL and_174_ssc : STD_LOGIC;
  SIGNAL and_540_ssc : STD_LOGIC;
  SIGNAL and_532_ssc : STD_LOGIC;
  SIGNAL and_518_ssc : STD_LOGIC;
  SIGNAL and_507_ssc : STD_LOGIC;
  SIGNAL and_498_ssc : STD_LOGIC;
  SIGNAL and_490_ssc : STD_LOGIC;
  SIGNAL and_475_ssc : STD_LOGIC;
  SIGNAL and_464_ssc : STD_LOGIC;
  SIGNAL and_455_ssc : STD_LOGIC;
  SIGNAL and_447_ssc : STD_LOGIC;
  SIGNAL and_433_ssc : STD_LOGIC;
  SIGNAL and_419_ssc : STD_LOGIC;
  SIGNAL and_410_ssc : STD_LOGIC;
  SIGNAL and_402_ssc : STD_LOGIC;
  SIGNAL and_387_ssc : STD_LOGIC;
  SIGNAL and_372_ssc : STD_LOGIC;
  SIGNAL and_363_ssc : STD_LOGIC;
  SIGNAL and_354_ssc : STD_LOGIC;
  SIGNAL and_339_ssc : STD_LOGIC;
  SIGNAL and_326_ssc : STD_LOGIC;
  SIGNAL and_316_ssc : STD_LOGIC;
  SIGNAL and_305_ssc : STD_LOGIC;
  SIGNAL and_288_ssc : STD_LOGIC;
  SIGNAL and_271_ssc : STD_LOGIC;
  SIGNAL and_262_ssc : STD_LOGIC;
  SIGNAL and_253_ssc : STD_LOGIC;
  SIGNAL and_237_ssc : STD_LOGIC;
  SIGNAL and_221_ssc : STD_LOGIC;
  SIGNAL and_207_ssc : STD_LOGIC;
  SIGNAL and_191_ssc : STD_LOGIC;
  SIGNAL and_164_ssc : STD_LOGIC;
  SIGNAL and_116_ssc : STD_LOGIC;
  SIGNAL butterFly_7_or_ssc_28 : STD_LOGIC;
  SIGNAL butterFly_7_or_ssc_29 : STD_LOGIC;
  SIGNAL butterFly_7_or_ssc_30 : STD_LOGIC;
  SIGNAL butterFly_7_or_ssc_31 : STD_LOGIC;
  SIGNAL and_151_seb : STD_LOGIC;
  SIGNAL and_179_seb : STD_LOGIC;
  SIGNAL and_201_seb : STD_LOGIC;
  SIGNAL and_217_seb : STD_LOGIC;
  SIGNAL and_230_seb : STD_LOGIC;
  SIGNAL and_243_seb : STD_LOGIC;
  SIGNAL and_257_seb : STD_LOGIC;
  SIGNAL and_267_seb : STD_LOGIC;
  SIGNAL and_281_seb : STD_LOGIC;
  SIGNAL and_295_seb : STD_LOGIC;
  SIGNAL and_311_seb : STD_LOGIC;
  SIGNAL and_322_seb : STD_LOGIC;
  SIGNAL and_333_seb : STD_LOGIC;
  SIGNAL and_344_seb : STD_LOGIC;
  SIGNAL and_358_seb : STD_LOGIC;
  SIGNAL and_368_seb : STD_LOGIC;
  SIGNAL and_381_seb : STD_LOGIC;
  SIGNAL and_393_seb : STD_LOGIC;
  SIGNAL and_406_seb : STD_LOGIC;
  SIGNAL and_415_seb : STD_LOGIC;
  SIGNAL and_427_seb : STD_LOGIC;
  SIGNAL and_438_seb : STD_LOGIC;
  SIGNAL and_451_seb : STD_LOGIC;
  SIGNAL and_460_seb : STD_LOGIC;
  SIGNAL and_470_seb : STD_LOGIC;
  SIGNAL and_481_seb : STD_LOGIC;
  SIGNAL and_494_seb : STD_LOGIC;
  SIGNAL and_503_seb : STD_LOGIC;
  SIGNAL and_513_seb : STD_LOGIC;
  SIGNAL and_523_seb : STD_LOGIC;
  SIGNAL and_536_seb : STD_LOGIC;
  SIGNAL and_546_seb : STD_LOGIC;
  SIGNAL and_587_seb : STD_LOGIC;
  SIGNAL and_618_seb : STD_LOGIC;
  SIGNAL and_644_seb : STD_LOGIC;
  SIGNAL and_662_seb : STD_LOGIC;
  SIGNAL and_677_seb : STD_LOGIC;
  SIGNAL and_693_seb : STD_LOGIC;
  SIGNAL and_705_seb : STD_LOGIC;
  SIGNAL and_716_seb : STD_LOGIC;
  SIGNAL and_729_seb : STD_LOGIC;
  SIGNAL and_745_seb : STD_LOGIC;
  SIGNAL and_760_seb : STD_LOGIC;
  SIGNAL and_773_seb : STD_LOGIC;
  SIGNAL and_786_seb : STD_LOGIC;
  SIGNAL and_797_seb : STD_LOGIC;
  SIGNAL and_808_seb : STD_LOGIC;
  SIGNAL and_818_seb : STD_LOGIC;
  SIGNAL and_831_seb : STD_LOGIC;
  SIGNAL and_847_seb : STD_LOGIC;
  SIGNAL and_863_seb : STD_LOGIC;
  SIGNAL and_876_seb : STD_LOGIC;
  SIGNAL and_888_seb : STD_LOGIC;
  SIGNAL and_900_seb : STD_LOGIC;
  SIGNAL and_911_seb : STD_LOGIC;
  SIGNAL and_921_seb : STD_LOGIC;
  SIGNAL and_933_seb : STD_LOGIC;
  SIGNAL and_948_seb : STD_LOGIC;
  SIGNAL and_963_seb : STD_LOGIC;
  SIGNAL and_976_seb : STD_LOGIC;
  SIGNAL and_988_seb : STD_LOGIC;
  SIGNAL and_1000_seb : STD_LOGIC;
  SIGNAL and_1011_seb : STD_LOGIC;
  SIGNAL and_1022_seb : STD_LOGIC;
  SIGNAL reg_twiddle_rsci_oswt_cse : STD_LOGIC;
  SIGNAL reg_revArr_rsci_oswt_cse : STD_LOGIC;
  SIGNAL reg_tw_rsci_oswt_cse : STD_LOGIC;
  SIGNAL reg_tw_rsci_s_raddr_core_cse : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL reg_xx_rsc_0_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_1_0_cgo_cse : STD_LOGIC;
  SIGNAL mux_167_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_2_0_cgo_cse : STD_LOGIC;
  SIGNAL or_435_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_3_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_4_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_5_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_6_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_7_0_cgo_cse : STD_LOGIC;
  SIGNAL or_673_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_8_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_9_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_10_0_cgo_cse : STD_LOGIC;
  SIGNAL or_898_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_11_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_12_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_13_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_14_0_cgo_cse : STD_LOGIC;
  SIGNAL nor_245_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_15_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_16_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_17_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_18_0_cgo_cse : STD_LOGIC;
  SIGNAL or_1344_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_19_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_20_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_21_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_22_0_cgo_cse : STD_LOGIC;
  SIGNAL nor_389_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_23_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_24_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_25_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_26_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_27_0_cgo_cse : STD_LOGIC;
  SIGNAL or_1818_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_28_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_29_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_30_0_cgo_cse : STD_LOGIC;
  SIGNAL and_1737_cse : STD_LOGIC;
  SIGNAL reg_xx_rsc_31_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_0_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_1_0_cgo_cse : STD_LOGIC;
  SIGNAL nor_636_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_2_0_cgo_cse : STD_LOGIC;
  SIGNAL or_2242_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_3_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_4_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_5_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_6_0_cgo_cse : STD_LOGIC;
  SIGNAL nor_701_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_7_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_8_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_9_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_10_0_cgo_cse : STD_LOGIC;
  SIGNAL or_2619_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_11_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_12_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_13_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_14_0_cgo_cse : STD_LOGIC;
  SIGNAL nor_817_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_15_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_16_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_17_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_18_0_cgo_cse : STD_LOGIC;
  SIGNAL or_2999_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_19_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_20_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_21_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_22_0_cgo_cse : STD_LOGIC;
  SIGNAL nor_947_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_23_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_24_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_25_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_26_0_cgo_cse : STD_LOGIC;
  SIGNAL or_3418_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_27_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_28_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_29_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_30_0_cgo_cse : STD_LOGIC;
  SIGNAL and_1369_cse : STD_LOGIC;
  SIGNAL reg_yy_rsc_31_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_0_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_0_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_1_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_1_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_0_0_i_s_raddr_core_cse : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL reg_x_rsc_0_0_i_s_waddr_core_cse : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL reg_x_rsc_0_0_i_s_dout_core_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_x_rsc_2_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_2_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_3_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_3_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_4_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_4_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_5_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_5_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_6_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_6_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_7_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_7_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_8_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_8_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_9_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_9_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_10_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_10_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_11_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_11_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_12_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_12_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_13_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_13_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_14_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_14_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_15_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_15_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_16_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_16_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_17_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_17_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_18_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_18_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_19_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_19_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_20_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_20_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_21_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_21_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_22_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_22_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_23_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_23_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_24_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_24_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_25_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_25_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_26_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_26_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_27_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_27_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_28_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_28_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_29_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_29_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_30_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_30_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_31_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_31_0_i_oswt_1_cse : STD_LOGIC;
  SIGNAL reg_x_rsc_triosy_31_0_obj_iswt0_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_1_cse : STD_LOGIC;
  SIGNAL and_1317_cse : STD_LOGIC;
  SIGNAL or_3894_cse : STD_LOGIC;
  SIGNAL and_2141_cse : STD_LOGIC;
  SIGNAL nor_1730_cse : STD_LOGIC;
  SIGNAL nor_2152_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_2_cse : STD_LOGIC;
  SIGNAL operator_20_true_1_and_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_5_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_16_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_1_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_34_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_39_cse : STD_LOGIC;
  SIGNAL and_1380_cse : STD_LOGIC;
  SIGNAL and_1919_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_44_cse : STD_LOGIC;
  SIGNAL and_1827_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_47_cse : STD_LOGIC;
  SIGNAL and_1773_cse : STD_LOGIC;
  SIGNAL and_1740_cse : STD_LOGIC;
  SIGNAL and_1721_cse : STD_LOGIC;
  SIGNAL and_1692_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_55_cse : STD_LOGIC;
  SIGNAL nor_1368_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_60_cse : STD_LOGIC;
  SIGNAL butterFly_4_f1_butterFly_4_f1_nor_cse : STD_LOGIC;
  SIGNAL nor_1375_cse : STD_LOGIC;
  SIGNAL butterFly_f1_and_cse : STD_LOGIC;
  SIGNAL butterFly_4_f1_and_cse : STD_LOGIC;
  SIGNAL butterFly_8_f1_and_cse : STD_LOGIC;
  SIGNAL operator_20_true_8_and_cse : STD_LOGIC;
  SIGNAL butterFly_12_f1_and_cse : STD_LOGIC;
  SIGNAL butterFly_16_f1_and_cse : STD_LOGIC;
  SIGNAL butterFly_20_f1_and_cse : STD_LOGIC;
  SIGNAL operator_20_true_15_and_cse : STD_LOGIC;
  SIGNAL or_2664_cse : STD_LOGIC;
  SIGNAL or_2186_cse : STD_LOGIC;
  SIGNAL or_2189_cse : STD_LOGIC;
  SIGNAL or_309_cse : STD_LOGIC;
  SIGNAL nor_1311_cse : STD_LOGIC;
  SIGNAL or_2245_cse : STD_LOGIC;
  SIGNAL or_324_cse : STD_LOGIC;
  SIGNAL nor_2142_cse : STD_LOGIC;
  SIGNAL nor_2186_cse : STD_LOGIC;
  SIGNAL or_2294_cse : STD_LOGIC;
  SIGNAL or_394_cse : STD_LOGIC;
  SIGNAL or_2338_cse : STD_LOGIC;
  SIGNAL and_2080_cse : STD_LOGIC;
  SIGNAL nor_44_cse : STD_LOGIC;
  SIGNAL or_338_cse : STD_LOGIC;
  SIGNAL or_337_cse : STD_LOGIC;
  SIGNAL or_336_cse : STD_LOGIC;
  SIGNAL nor_690_cse : STD_LOGIC;
  SIGNAL or_2386_cse : STD_LOGIC;
  SIGNAL nor_2156_cse : STD_LOGIC;
  SIGNAL nor_2157_cse : STD_LOGIC;
  SIGNAL or_549_cse : STD_LOGIC;
  SIGNAL or_401_cse : STD_LOGIC;
  SIGNAL or_2440_cse : STD_LOGIC;
  SIGNAL nor_132_cse : STD_LOGIC;
  SIGNAL nor_2081_cse : STD_LOGIC;
  SIGNAL or_2487_cse : STD_LOGIC;
  SIGNAL or_632_cse : STD_LOGIC;
  SIGNAL or_2528_cse : STD_LOGIC;
  SIGNAL or_2574_cse : STD_LOGIC;
  SIGNAL or_2577_cse : STD_LOGIC;
  SIGNAL or_789_cse : STD_LOGIC;
  SIGNAL or_2622_cse : STD_LOGIC;
  SIGNAL nor_2030_cse : STD_LOGIC;
  SIGNAL or_863_cse : STD_LOGIC;
  SIGNAL or_2700_cse : STD_LOGIC;
  SIGNAL nand_492_cse : STD_LOGIC;
  SIGNAL nor_805_cse : STD_LOGIC;
  SIGNAL or_2747_cse : STD_LOGIC;
  SIGNAL or_1006_cse : STD_LOGIC;
  SIGNAL or_2800_cse : STD_LOGIC;
  SIGNAL or_2847_cse : STD_LOGIC;
  SIGNAL nand_317_cse : STD_LOGIC;
  SIGNAL or_2947_cse : STD_LOGIC;
  SIGNAL nor_873_cse : STD_LOGIC;
  SIGNAL nor_885_cse : STD_LOGIC;
  SIGNAL nor_1928_cse : STD_LOGIC;
  SIGNAL or_1309_cse : STD_LOGIC;
  SIGNAL nor_934_cse : STD_LOGIC;
  SIGNAL nor_938_cse : STD_LOGIC;
  SIGNAL nor_951_cse : STD_LOGIC;
  SIGNAL nand_479_cse : STD_LOGIC;
  SIGNAL or_3367_cse : STD_LOGIC;
  SIGNAL nor_1010_cse : STD_LOGIC;
  SIGNAL nor_1025_cse : STD_LOGIC;
  SIGNAL nor_1822_cse : STD_LOGIC;
  SIGNAL and_1812_cse : STD_LOGIC;
  SIGNAL or_1783_cse : STD_LOGIC;
  SIGNAL nand_520_cse : STD_LOGIC;
  SIGNAL nor_1089_cse : STD_LOGIC;
  SIGNAL and_1366_cse : STD_LOGIC;
  SIGNAL and_1329_cse : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_61_cse : STD_LOGIC;
  SIGNAL or_348_cse : STD_LOGIC;
  SIGNAL nor_2197_cse : STD_LOGIC;
  SIGNAL or_3918_cse : STD_LOGIC;
  SIGNAL or_119_cse : STD_LOGIC;
  SIGNAL or_2199_cse : STD_LOGIC;
  SIGNAL and_1674_cse : STD_LOGIC;
  SIGNAL or_4378_cse : STD_LOGIC;
  SIGNAL and_1665_cse : STD_LOGIC;
  SIGNAL or_2161_cse : STD_LOGIC;
  SIGNAL or_2158_cse : STD_LOGIC;
  SIGNAL or_2157_cse : STD_LOGIC;
  SIGNAL or_2147_cse : STD_LOGIC;
  SIGNAL nand_331_cse : STD_LOGIC;
  SIGNAL or_582_cse : STD_LOGIC;
  SIGNAL or_2215_cse : STD_LOGIC;
  SIGNAL or_2273_cse : STD_LOGIC;
  SIGNAL or_2272_cse : STD_LOGIC;
  SIGNAL or_2271_cse : STD_LOGIC;
  SIGNAL or_2396_cse : STD_LOGIC;
  SIGNAL nor_673_cse : STD_LOGIC;
  SIGNAL or_823_cse : STD_LOGIC;
  SIGNAL nand_330_cse : STD_LOGIC;
  SIGNAL or_2585_cse : STD_LOGIC;
  SIGNAL or_1039_cse : STD_LOGIC;
  SIGNAL nor_291_cse : STD_LOGIC;
  SIGNAL nor_901_cse : STD_LOGIC;
  SIGNAL or_2958_cse : STD_LOGIC;
  SIGNAL nor_920_cse : STD_LOGIC;
  SIGNAL nor_356_cse : STD_LOGIC;
  SIGNAL nand_327_cse : STD_LOGIC;
  SIGNAL nor_969_cse : STD_LOGIC;
  SIGNAL or_3159_cse : STD_LOGIC;
  SIGNAL and_1435_cse : STD_LOGIC;
  SIGNAL nor_437_cse : STD_LOGIC;
  SIGNAL nor_1044_cse : STD_LOGIC;
  SIGNAL or_3377_cse : STD_LOGIC;
  SIGNAL and_1391_cse : STD_LOGIC;
  SIGNAL and_1765_cse : STD_LOGIC;
  SIGNAL and_1350_cse : STD_LOGIC;
  SIGNAL nor_2144_cse : STD_LOGIC;
  SIGNAL nor_2032_cse : STD_LOGIC;
  SIGNAL nor_1930_cse : STD_LOGIC;
  SIGNAL nor_2183_cse : STD_LOGIC;
  SIGNAL or_4342_cse : STD_LOGIC;
  SIGNAL and_1532_cse : STD_LOGIC;
  SIGNAL and_1447_cse : STD_LOGIC;
  SIGNAL and_1403_cse : STD_LOGIC;
  SIGNAL and_1373_cse : STD_LOGIC;
  SIGNAL and_1344_cse : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_22_cse : STD_LOGIC;
  SIGNAL or_4376_cse : STD_LOGIC;
  SIGNAL and_1306_cse : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_44_cse : STD_LOGIC;
  SIGNAL and_2120_cse : STD_LOGIC;
  SIGNAL or_448_cse : STD_LOGIC;
  SIGNAL or_387_cse : STD_LOGIC;
  SIGNAL or_445_cse : STD_LOGIC;
  SIGNAL or_501_cse : STD_LOGIC;
  SIGNAL or_686_cse : STD_LOGIC;
  SIGNAL or_618_cse : STD_LOGIC;
  SIGNAL or_682_cse : STD_LOGIC;
  SIGNAL or_735_cse : STD_LOGIC;
  SIGNAL or_233_cse : STD_LOGIC;
  SIGNAL or_911_cse : STD_LOGIC;
  SIGNAL or_856_cse : STD_LOGIC;
  SIGNAL or_261_cse : STD_LOGIC;
  SIGNAL or_908_cse : STD_LOGIC;
  SIGNAL or_955_cse : STD_LOGIC;
  SIGNAL or_1073_cse : STD_LOGIC;
  SIGNAL or_1130_cse : STD_LOGIC;
  SIGNAL nand_449_cse : STD_LOGIC;
  SIGNAL or_1358_cse : STD_LOGIC;
  SIGNAL nand_508_cse : STD_LOGIC;
  SIGNAL or_1527_cse : STD_LOGIC;
  SIGNAL nand_480_cse : STD_LOGIC;
  SIGNAL nand_393_cse : STD_LOGIC;
  SIGNAL nand_517_cse : STD_LOGIC;
  SIGNAL nand_336_cse : STD_LOGIC;
  SIGNAL nand_351_cse : STD_LOGIC;
  SIGNAL and_1713_cse : STD_LOGIC;
  SIGNAL or_4679_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_76_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_90_cse : STD_LOGIC;
  SIGNAL or_395_cse : STD_LOGIC;
  SIGNAL or_2204_cse : STD_LOGIC;
  SIGNAL or_4699_cse : STD_LOGIC;
  SIGNAL nor_1712_cse : STD_LOGIC;
  SIGNAL or_634_cse : STD_LOGIC;
  SIGNAL or_2405_cse : STD_LOGIC;
  SIGNAL or_864_cse : STD_LOGIC;
  SIGNAL or_2590_cse : STD_LOGIC;
  SIGNAL or_1310_cse : STD_LOGIC;
  SIGNAL or_2962_cse : STD_LOGIC;
  SIGNAL or_1547_cse : STD_LOGIC;
  SIGNAL nand_542_cse : STD_LOGIC;
  SIGNAL or_1784_cse : STD_LOGIC;
  SIGNAL nand_300_cse : STD_LOGIC;
  SIGNAL nor_1711_cse : STD_LOGIC;
  SIGNAL and_2112_cse : STD_LOGIC;
  SIGNAL nand_242_cse : STD_LOGIC;
  SIGNAL mux_45_cse : STD_LOGIC;
  SIGNAL or_129_cse : STD_LOGIC;
  SIGNAL nor_1303_cse : STD_LOGIC;
  SIGNAL or_4162_cse : STD_LOGIC;
  SIGNAL or_4165_cse : STD_LOGIC;
  SIGNAL mux_108_cse : STD_LOGIC;
  SIGNAL and_1274_cse : STD_LOGIC;
  SIGNAL and_1272_cse : STD_LOGIC;
  SIGNAL or_3852_cse : STD_LOGIC;
  SIGNAL nor_2247_cse : STD_LOGIC;
  SIGNAL or_315_cse : STD_LOGIC;
  SIGNAL or_447_cse : STD_LOGIC;
  SIGNAL or_555_cse : STD_LOGIC;
  SIGNAL or_684_cse : STD_LOGIC;
  SIGNAL or_795_cse : STD_LOGIC;
  SIGNAL or_910_cse : STD_LOGIC;
  SIGNAL or_1012_cse : STD_LOGIC;
  SIGNAL or_1133_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_201_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_204_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_207_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_210_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_213_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_216_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_219_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_222_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_225_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_228_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_231_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_234_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_237_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_240_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_243_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_246_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_249_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_252_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_255_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_258_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_261_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_264_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_267_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_270_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_273_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_276_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_279_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_282_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_285_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_288_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_291_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_294_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_264_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_201_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_296_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_203_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_301_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_205_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_306_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_207_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_311_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_209_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_211_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_213_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_215_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_217_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_219_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_221_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_223_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_225_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_227_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_229_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_231_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_233_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_235_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_237_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_239_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_241_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_243_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_245_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_247_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_249_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_251_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_253_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_255_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_257_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_259_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_261_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_263_cse : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_66 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48 : STD_LOGIC;
  SIGNAL mux_162_cse : STD_LOGIC;
  SIGNAL mux_226_cse : STD_LOGIC;
  SIGNAL mux_213_cse : STD_LOGIC;
  SIGNAL mux_223_cse : STD_LOGIC;
  SIGNAL mux_435_cse : STD_LOGIC;
  SIGNAL mux_641_cse : STD_LOGIC;
  SIGNAL nor_1978_cse : STD_LOGIC;
  SIGNAL or_1083_cse : STD_LOGIC;
  SIGNAL mux_847_cse : STD_LOGIC;
  SIGNAL nor_1862_cse : STD_LOGIC;
  SIGNAL mux_1493_cse : STD_LOGIC;
  SIGNAL nor_1771_cse : STD_LOGIC;
  SIGNAL or_2011_cse : STD_LOGIC;
  SIGNAL mux_1877_cse : STD_LOGIC;
  SIGNAL mux_1872_cse : STD_LOGIC;
  SIGNAL mux_1868_cse : STD_LOGIC;
  SIGNAL mux_1865_cse : STD_LOGIC;
  SIGNAL or_2756_cse : STD_LOGIC;
  SIGNAL or_3574_cse : STD_LOGIC;
  SIGNAL mux_297_cse : STD_LOGIC;
  SIGNAL or_1135_cse : STD_LOGIC;
  SIGNAL mux_295_cse : STD_LOGIC;
  SIGNAL or_1085_cse : STD_LOGIC;
  SIGNAL or_2765_cse : STD_LOGIC;
  SIGNAL mux_37_cse : STD_LOGIC;
  SIGNAL or_124_cse : STD_LOGIC;
  SIGNAL mux_3678_cse : STD_LOGIC;
  SIGNAL mux_3731_cse : STD_LOGIC;
  SIGNAL mux_146_cse : STD_LOGIC;
  SIGNAL and_142_cse : STD_LOGIC;
  SIGNAL mux_309_cse : STD_LOGIC;
  SIGNAL mux_296_cse : STD_LOGIC;
  SIGNAL mux_1953_cse : STD_LOGIC;
  SIGNAL mux_1857_cse : STD_LOGIC;
  SIGNAL mux_1854_cse : STD_LOGIC;
  SIGNAL mux_1847_cse : STD_LOGIC;
  SIGNAL or_2224_cse : STD_LOGIC;
  SIGNAL mux_1967_cse : STD_LOGIC;
  SIGNAL mux_2028_cse : STD_LOGIC;
  SIGNAL butterFly_3_f1_asn_17 : STD_LOGIC;
  SIGNAL nor_2124_cse : STD_LOGIC;
  SIGNAL mux_171_cse : STD_LOGIC;
  SIGNAL mux_163_cse : STD_LOGIC;
  SIGNAL nor_2066_cse : STD_LOGIC;
  SIGNAL mux_440_cse : STD_LOGIC;
  SIGNAL mux_646_cse : STD_LOGIC;
  SIGNAL nor_2014_cse : STD_LOGIC;
  SIGNAL mux_852_cse : STD_LOGIC;
  SIGNAL nor_1963_cse : STD_LOGIC;
  SIGNAL mux_1063_cse : STD_LOGIC;
  SIGNAL nor_1914_cse : STD_LOGIC;
  SIGNAL mux_1281_cse : STD_LOGIC;
  SIGNAL nor_1860_cse : STD_LOGIC;
  SIGNAL nor_1810_cse : STD_LOGIC;
  SIGNAL mux_1498_cse : STD_LOGIC;
  SIGNAL mux_1715_cse : STD_LOGIC;
  SIGNAL nor_1758_cse : STD_LOGIC;
  SIGNAL mux_1927_cse : STD_LOGIC;
  SIGNAL mux_2152_cse : STD_LOGIC;
  SIGNAL mux_2372_cse : STD_LOGIC;
  SIGNAL mux_2592_cse : STD_LOGIC;
  SIGNAL mux_2812_cse : STD_LOGIC;
  SIGNAL mux_3032_cse : STD_LOGIC;
  SIGNAL mux_3252_cse : STD_LOGIC;
  SIGNAL mux_3472_cse : STD_LOGIC;
  SIGNAL mux_298_cse : STD_LOGIC;
  SIGNAL mux_308_cse : STD_LOGIC;
  SIGNAL mux_1966_cse : STD_LOGIC;
  SIGNAL mux_2027_cse : STD_LOGIC;
  SIGNAL twiddle_rsci_adrb_d_reg : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL mux_111_rmff : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_tfh_S2_INNER_LOOP1_tfh_mux_rmff : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_tfh_mux1h_rmff : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL twiddle_h_rsci_adrb_d_reg : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_rmff : STD_LOGIC;
  SIGNAL mux_191_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_2_rmff : STD_LOGIC;
  SIGNAL mux_241_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_4_rmff : STD_LOGIC;
  SIGNAL mux_293_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_6_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_8_rmff : STD_LOGIC;
  SIGNAL mux_408_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_10_rmff : STD_LOGIC;
  SIGNAL mux_455_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_12_rmff : STD_LOGIC;
  SIGNAL mux_504_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_14_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_16_rmff : STD_LOGIC;
  SIGNAL mux_614_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_18_rmff : STD_LOGIC;
  SIGNAL mux_661_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_20_rmff : STD_LOGIC;
  SIGNAL mux_710_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_22_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_24_rmff : STD_LOGIC;
  SIGNAL mux_820_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_26_rmff : STD_LOGIC;
  SIGNAL mux_867_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_28_rmff : STD_LOGIC;
  SIGNAL mux_916_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_30_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_32_rmff : STD_LOGIC;
  SIGNAL mux_1030_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_34_rmff : STD_LOGIC;
  SIGNAL mux_1080_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_36_rmff : STD_LOGIC;
  SIGNAL mux_1132_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_38_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_40_rmff : STD_LOGIC;
  SIGNAL mux_1248_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_42_rmff : STD_LOGIC;
  SIGNAL mux_1298_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_44_rmff : STD_LOGIC;
  SIGNAL mux_1350_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_46_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_48_rmff : STD_LOGIC;
  SIGNAL mux_1465_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_50_rmff : STD_LOGIC;
  SIGNAL mux_1515_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_52_rmff : STD_LOGIC;
  SIGNAL mux_1567_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_54_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_56_rmff : STD_LOGIC;
  SIGNAL mux_1682_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_58_rmff : STD_LOGIC;
  SIGNAL mux_1732_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_60_rmff : STD_LOGIC;
  SIGNAL mux_1781_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_62_rmff : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_rmff : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_butterFly_3_or_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_64_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_65_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_66_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_67_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_68_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_69_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_70_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_71_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_72_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_73_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_74_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_75_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_76_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_77_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_78_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_79_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_80_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_81_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_82_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_83_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_84_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_85_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_86_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_87_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_88_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_89_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_90_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_91_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_92_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_93_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_94_rmff : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_95_rmff : STD_LOGIC;
  SIGNAL and_1109_rmff : STD_LOGIC;
  SIGNAL mux_1880_seb : STD_LOGIC;
  SIGNAL mux_1932_seb : STD_LOGIC;
  SIGNAL mux_1990_seb : STD_LOGIC;
  SIGNAL mux_2051_seb : STD_LOGIC;
  SIGNAL mux_2108_seb : STD_LOGIC;
  SIGNAL mux_2157_seb : STD_LOGIC;
  SIGNAL mux_2213_seb : STD_LOGIC;
  SIGNAL mux_2271_seb : STD_LOGIC;
  SIGNAL mux_2328_seb : STD_LOGIC;
  SIGNAL mux_2377_seb : STD_LOGIC;
  SIGNAL mux_2433_seb : STD_LOGIC;
  SIGNAL mux_2491_seb : STD_LOGIC;
  SIGNAL mux_2548_seb : STD_LOGIC;
  SIGNAL mux_2597_seb : STD_LOGIC;
  SIGNAL mux_2653_seb : STD_LOGIC;
  SIGNAL mux_2711_seb : STD_LOGIC;
  SIGNAL mux_2768_seb : STD_LOGIC;
  SIGNAL mux_2817_seb : STD_LOGIC;
  SIGNAL mux_2873_seb : STD_LOGIC;
  SIGNAL mux_2931_seb : STD_LOGIC;
  SIGNAL mux_2988_seb : STD_LOGIC;
  SIGNAL mux_3037_seb : STD_LOGIC;
  SIGNAL mux_3093_seb : STD_LOGIC;
  SIGNAL mux_3151_seb : STD_LOGIC;
  SIGNAL mux_3208_seb : STD_LOGIC;
  SIGNAL mux_3257_seb : STD_LOGIC;
  SIGNAL mux_3313_seb : STD_LOGIC;
  SIGNAL mux_3371_seb : STD_LOGIC;
  SIGNAL mux_3428_seb : STD_LOGIC;
  SIGNAL mux_3477_seb : STD_LOGIC;
  SIGNAL mux_3533_seb : STD_LOGIC;
  SIGNAL mux_3591_seb : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_tf_sva : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL tmp_37_lpi_3_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_7_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_5_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_3_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_1_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_7_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_33_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_31_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_29_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_35_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_13_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_11_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_9_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_43_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_41_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_39_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_45_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_51_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_49_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_47_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_53_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S2_INNER_LOOP1_tfh_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S2_INNER_LOOP1_tf_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S34_OUTER_LOOP_for_tf_h_sva : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL modulo_sub_7_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_1_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_3_qr_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_15_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_23_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_4_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_12_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_20_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_5_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_13_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_21_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_6_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_14_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_3_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_19_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_55_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_11_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_16_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_8_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_1_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_17_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_9_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_2_qr_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_10_qr_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mux_138_itm : STD_LOGIC;
  SIGNAL mux_357_itm : STD_LOGIC;
  SIGNAL mux_566_itm : STD_LOGIC;
  SIGNAL mux_772_itm : STD_LOGIC;
  SIGNAL mux_979_itm : STD_LOGIC;
  SIGNAL mux_1196_itm : STD_LOGIC;
  SIGNAL mux_1414_itm : STD_LOGIC;
  SIGNAL mux_1631_itm : STD_LOGIC;
  SIGNAL mux_1843_itm : STD_LOGIC;
  SIGNAL mux_1902_itm : STD_LOGIC;
  SIGNAL mux_1950_itm : STD_LOGIC;
  SIGNAL mux_2010_itm : STD_LOGIC;
  SIGNAL mux_2075_itm : STD_LOGIC;
  SIGNAL mux_2130_itm : STD_LOGIC;
  SIGNAL mux_2175_itm : STD_LOGIC;
  SIGNAL mux_2233_itm : STD_LOGIC;
  SIGNAL mux_2295_itm : STD_LOGIC;
  SIGNAL mux_2350_itm : STD_LOGIC;
  SIGNAL mux_2395_itm : STD_LOGIC;
  SIGNAL mux_2453_itm : STD_LOGIC;
  SIGNAL mux_2515_itm : STD_LOGIC;
  SIGNAL mux_2570_itm : STD_LOGIC;
  SIGNAL mux_2615_itm : STD_LOGIC;
  SIGNAL mux_2673_itm : STD_LOGIC;
  SIGNAL mux_2735_itm : STD_LOGIC;
  SIGNAL mux_2790_itm : STD_LOGIC;
  SIGNAL mux_2835_itm : STD_LOGIC;
  SIGNAL mux_2893_itm : STD_LOGIC;
  SIGNAL mux_2955_itm : STD_LOGIC;
  SIGNAL mux_3010_itm : STD_LOGIC;
  SIGNAL mux_3055_itm : STD_LOGIC;
  SIGNAL mux_3113_itm : STD_LOGIC;
  SIGNAL mux_3175_itm : STD_LOGIC;
  SIGNAL mux_3230_itm : STD_LOGIC;
  SIGNAL mux_3275_itm : STD_LOGIC;
  SIGNAL mux_3333_itm : STD_LOGIC;
  SIGNAL mux_3395_itm : STD_LOGIC;
  SIGNAL mux_3450_itm : STD_LOGIC;
  SIGNAL mux_3495_itm : STD_LOGIC;
  SIGNAL mux_3553_itm : STD_LOGIC;
  SIGNAL mux_3669_itm : STD_LOGIC;
  SIGNAL mux_156_itm : STD_LOGIC;
  SIGNAL mux_3695_itm : STD_LOGIC;
  SIGNAL z_out : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL and_dcpl_1165 : STD_LOGIC;
  SIGNAL and_dcpl_1178 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL or_tmp_4090 : STD_LOGIC;
  SIGNAL and_dcpl_1206 : STD_LOGIC;
  SIGNAL and_dcpl_1210 : STD_LOGIC;
  SIGNAL and_dcpl_1222 : STD_LOGIC;
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_dcpl_1241 : STD_LOGIC;
  SIGNAL and_dcpl_1246 : STD_LOGIC;
  SIGNAL and_dcpl_1257 : STD_LOGIC;
  SIGNAL z_out_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_dcpl_1324 : STD_LOGIC;
  SIGNAL z_out_9 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_10 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_11 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_12 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_13 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_14 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_dcpl_1455 : STD_LOGIC;
  SIGNAL and_dcpl_1566 : STD_LOGIC;
  SIGNAL and_dcpl_1573 : STD_LOGIC;
  SIGNAL and_dcpl_1596 : STD_LOGIC;
  SIGNAL and_dcpl_1633 : STD_LOGIC;
  SIGNAL z_out_26 : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL S2_OUTER_LOOP_c_2_sva : STD_LOGIC;
  SIGNAL tmp_1_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_13_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_13_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_13_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_13_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_13_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_15_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_sva_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_sva_22 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_sva_23 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_sva_26 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_sva_31 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_17_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_19_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_sva_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_sva_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_23_lpi_4_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_10 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_26 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_27 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_sva_29 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_9_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_19_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_23_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_28_itm : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nor_32_itm : STD_LOGIC;
  SIGNAL mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL S1_OUTER_LOOP_for_p_sva_1_mx0c1 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_nor_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_9_itm_mx0w1 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_nor_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_nor_1_itm_mx0w1 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_nor_14_itm_mx0w1 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_5_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_25_itm_mx0w2 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_8_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_27_itm_mx0w2 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm_mx0w0 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_nor_itm_mx0w1 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_29_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_4_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_6_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_10_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_12_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_13_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_14_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_18_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_20_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_21_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_16_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_24_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_19_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_2_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_23_itm_mx0w1 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_11_itm_mx0w0 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_17_itm_mx0w0 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c3 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c4 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c9 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c14 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c18 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c21 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c26 : STD_LOGIC;
  SIGNAL modulo_add_base_1_sva_mx0c30 : STD_LOGIC;
  SIGNAL mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 : STD_LOGIC;
  SIGNAL mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c7 : STD_LOGIC;
  SIGNAL mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 : STD_LOGIC;
  SIGNAL mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 : STD_LOGIC;
  SIGNAL operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm_mx0c3
      : STD_LOGIC;
  SIGNAL operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm_mx0c3
      : STD_LOGIC;
  SIGNAL operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm_mx0c3
      : STD_LOGIC;
  SIGNAL S2_OUTER_LOOP_c_1_sva_mx0c1 : STD_LOGIC;
  SIGNAL S2_OUTER_LOOP_c_1_sva_mx0c2 : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_tf_and_psp_sva_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL tmp_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_1_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_3_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_5_lpi_4_dfm_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2383_ssc : STD_LOGIC;
  SIGNAL reg_tmp_54_lpi_3_dfm_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_modulo_add_3_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL reg_mult_res_lpi_4_dfm_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_3_res_lpi_4_dfm_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_2_res_lpi_4_dfm_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_1_res_lpi_4_dfm_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_modulo_add_5_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL reg_modulo_add_1_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL reg_modulo_add_6_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL reg_modulo_add_7_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL reg_modulo_add_2_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL reg_modulo_add_11_slc_32_svs_st_cse : STD_LOGIC;
  SIGNAL butterFly_3_or_456_cse : STD_LOGIC;
  SIGNAL nor_2307_cse : STD_LOGIC;
  SIGNAL mux_100_cse : STD_LOGIC;
  SIGNAL nor_1346_cse : STD_LOGIC;
  SIGNAL and_2083_cse : STD_LOGIC;
  SIGNAL nor_1395_cse : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_tf_and_1_cse : STD_LOGIC;
  SIGNAL reg_modulo_sub_18_qr_lpi_4_dfm_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2399_cse : STD_LOGIC;
  SIGNAL mux_tmp_4267 : STD_LOGIC;
  SIGNAL mux_tmp_4268 : STD_LOGIC;
  SIGNAL or_tmp_4112 : STD_LOGIC;
  SIGNAL or_tmp_4115 : STD_LOGIC;
  SIGNAL or_tmp_4117 : STD_LOGIC;
  SIGNAL or_tmp_4118 : STD_LOGIC;
  SIGNAL or_tmp_4121 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_p_asn_S2_COPY_LOOP_p_5_0_sva_4_0_S1_OUTER_LOOP_k_and_rgt :
      STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL or_tmp_4152 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_i_mux1h_2_rgt : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL mux_tmp_4334 : STD_LOGIC;
  SIGNAL or_tmp_4164 : STD_LOGIC;
  SIGNAL or_tmp_4177 : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_and_rgt : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL mux_tmp_4373 : STD_LOGIC;
  SIGNAL mux_tmp_4374 : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_S2_COPY_LOOP_for_mux_6_rgt : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  SIGNAL or_tmp_4199 : STD_LOGIC;
  SIGNAL mux_tmp_4396 : STD_LOGIC;
  SIGNAL or_tmp_4208 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_acc_svs_4 : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_acc_svs_3_0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL S2_COPY_LOOP_for_i_5_0_sva_1_5 : STD_LOGIC;
  SIGNAL operator_33_true_return_2_3_0_sva_3 : STD_LOGIC;
  SIGNAL operator_33_true_return_2_3_0_sva_2_0 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL revArr_rsci_s_raddr_core_4 : STD_LOGIC;
  SIGNAL revArr_rsci_s_raddr_core_3_0 : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL reg_drf_revArr_ptr_1_smx_9_0_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reg_drf_revArr_ptr_1_smx_9_0_1_reg : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_S2_COPY_LOOP_for_i_5_0_1_reg : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL reg_S2_COPY_LOOP_for_i_5_0_2_reg : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg : STD_LOGIC;
  SIGNAL reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_2348_ssc : STD_LOGIC;
  SIGNAL or_2194_cse : STD_LOGIC;
  SIGNAL nand_531_cse : STD_LOGIC;
  SIGNAL nor_2178_cse_1 : STD_LOGIC;
  SIGNAL nand_570_cse : STD_LOGIC;
  SIGNAL nand_569_cse : STD_LOGIC;
  SIGNAL and_2893_cse : STD_LOGIC;
  SIGNAL nor_1308_cse : STD_LOGIC;
  SIGNAL or_4805_cse : STD_LOGIC;
  SIGNAL nor_2412_cse : STD_LOGIC;
  SIGNAL nor_2411_cse : STD_LOGIC;
  SIGNAL nand_568_cse : STD_LOGIC;
  SIGNAL or_4854_cse : STD_LOGIC;
  SIGNAL or_4818_cse : STD_LOGIC;
  SIGNAL or_4781_cse : STD_LOGIC;
  SIGNAL and_2881_cse : STD_LOGIC;
  SIGNAL or_4797_cse : STD_LOGIC;
  SIGNAL butterFly_7_or_360_cse : STD_LOGIC;
  SIGNAL nand_536_cse : STD_LOGIC;
  SIGNAL or_4769_cse : STD_LOGIC;
  SIGNAL z_out_16_14 : STD_LOGIC;
  SIGNAL z_out_17_32 : STD_LOGIC;
  SIGNAL z_out_19_32 : STD_LOGIC;
  SIGNAL and_2913_cse : STD_LOGIC;

  SIGNAL mux_104_nl : STD_LOGIC;
  SIGNAL nor_2174_nl : STD_LOGIC;
  SIGNAL mux_103_nl : STD_LOGIC;
  SIGNAL mux_102_nl : STD_LOGIC;
  SIGNAL or_285_nl : STD_LOGIC;
  SIGNAL mux_101_nl : STD_LOGIC;
  SIGNAL mux_110_nl : STD_LOGIC;
  SIGNAL nor_2167_nl : STD_LOGIC;
  SIGNAL mux_109_nl : STD_LOGIC;
  SIGNAL or_299_nl : STD_LOGIC;
  SIGNAL or_298_nl : STD_LOGIC;
  SIGNAL and_2097_nl : STD_LOGIC;
  SIGNAL and_2098_nl : STD_LOGIC;
  SIGNAL mux_107_nl : STD_LOGIC;
  SIGNAL nor_2170_nl : STD_LOGIC;
  SIGNAL nor_2171_nl : STD_LOGIC;
  SIGNAL S2_INNER_LOOP2_tf_and_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL and_90_nl : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_tfh_or_nl : STD_LOGIC;
  SIGNAL mux_137_nl : STD_LOGIC;
  SIGNAL mux_136_nl : STD_LOGIC;
  SIGNAL mux_135_nl : STD_LOGIC;
  SIGNAL mux_134_nl : STD_LOGIC;
  SIGNAL mux_133_nl : STD_LOGIC;
  SIGNAL mux_132_nl : STD_LOGIC;
  SIGNAL or_340_nl : STD_LOGIC;
  SIGNAL mux_131_nl : STD_LOGIC;
  SIGNAL mux_130_nl : STD_LOGIC;
  SIGNAL mux_129_nl : STD_LOGIC;
  SIGNAL or_335_nl : STD_LOGIC;
  SIGNAL or_332_nl : STD_LOGIC;
  SIGNAL or_327_nl : STD_LOGIC;
  SIGNAL mux_126_nl : STD_LOGIC;
  SIGNAL mux_125_nl : STD_LOGIC;
  SIGNAL mux_124_nl : STD_LOGIC;
  SIGNAL or_326_nl : STD_LOGIC;
  SIGNAL mux_123_nl : STD_LOGIC;
  SIGNAL or_325_nl : STD_LOGIC;
  SIGNAL mux_122_nl : STD_LOGIC;
  SIGNAL or_323_nl : STD_LOGIC;
  SIGNAL mux_120_nl : STD_LOGIC;
  SIGNAL mux_119_nl : STD_LOGIC;
  SIGNAL or_317_nl : STD_LOGIC;
  SIGNAL or_316_nl : STD_LOGIC;
  SIGNAL mux_118_nl : STD_LOGIC;
  SIGNAL mux_117_nl : STD_LOGIC;
  SIGNAL or_313_nl : STD_LOGIC;
  SIGNAL nand_8_nl : STD_LOGIC;
  SIGNAL mux_116_nl : STD_LOGIC;
  SIGNAL or_312_nl : STD_LOGIC;
  SIGNAL mux_115_nl : STD_LOGIC;
  SIGNAL mux_170_nl : STD_LOGIC;
  SIGNAL mux_169_nl : STD_LOGIC;
  SIGNAL and_2086_nl : STD_LOGIC;
  SIGNAL mux_168_nl : STD_LOGIC;
  SIGNAL or_374_nl : STD_LOGIC;
  SIGNAL mux_190_nl : STD_LOGIC;
  SIGNAL mux_189_nl : STD_LOGIC;
  SIGNAL mux_188_nl : STD_LOGIC;
  SIGNAL and_2084_nl : STD_LOGIC;
  SIGNAL mux_187_nl : STD_LOGIC;
  SIGNAL nor_2139_nl : STD_LOGIC;
  SIGNAL nor_2140_nl : STD_LOGIC;
  SIGNAL nor_2141_nl : STD_LOGIC;
  SIGNAL and_2085_nl : STD_LOGIC;
  SIGNAL mux_185_nl : STD_LOGIC;
  SIGNAL nor_2143_nl : STD_LOGIC;
  SIGNAL mux_184_nl : STD_LOGIC;
  SIGNAL mux_183_nl : STD_LOGIC;
  SIGNAL mux_182_nl : STD_LOGIC;
  SIGNAL or_400_nl : STD_LOGIC;
  SIGNAL nor_2145_nl : STD_LOGIC;
  SIGNAL mux_181_nl : STD_LOGIC;
  SIGNAL or_396_nl : STD_LOGIC;
  SIGNAL mux_180_nl : STD_LOGIC;
  SIGNAL or_393_nl : STD_LOGIC;
  SIGNAL mux_179_nl : STD_LOGIC;
  SIGNAL or_392_nl : STD_LOGIC;
  SIGNAL mux_178_nl : STD_LOGIC;
  SIGNAL mux_177_nl : STD_LOGIC;
  SIGNAL mux_176_nl : STD_LOGIC;
  SIGNAL nor_2146_nl : STD_LOGIC;
  SIGNAL or_389_nl : STD_LOGIC;
  SIGNAL nand_10_nl : STD_LOGIC;
  SIGNAL and_2074_nl : STD_LOGIC;
  SIGNAL mux_222_nl : STD_LOGIC;
  SIGNAL mux_225_nl : STD_LOGIC;
  SIGNAL mux_224_nl : STD_LOGIC;
  SIGNAL mux_221_nl : STD_LOGIC;
  SIGNAL or_434_nl : STD_LOGIC;
  SIGNAL mux_240_nl : STD_LOGIC;
  SIGNAL mux_239_nl : STD_LOGIC;
  SIGNAL mux_238_nl : STD_LOGIC;
  SIGNAL and_2073_nl : STD_LOGIC;
  SIGNAL mux_237_nl : STD_LOGIC;
  SIGNAL nor_2122_nl : STD_LOGIC;
  SIGNAL nor_2123_nl : STD_LOGIC;
  SIGNAL nor_2125_nl : STD_LOGIC;
  SIGNAL mux_236_nl : STD_LOGIC;
  SIGNAL nor_2127_nl : STD_LOGIC;
  SIGNAL mux_235_nl : STD_LOGIC;
  SIGNAL mux_234_nl : STD_LOGIC;
  SIGNAL nand_494_nl : STD_LOGIC;
  SIGNAL or_458_nl : STD_LOGIC;
  SIGNAL nor_2130_nl : STD_LOGIC;
  SIGNAL mux_233_nl : STD_LOGIC;
  SIGNAL or_454_nl : STD_LOGIC;
  SIGNAL mux_232_nl : STD_LOGIC;
  SIGNAL or_453_nl : STD_LOGIC;
  SIGNAL or_449_nl : STD_LOGIC;
  SIGNAL mux_230_nl : STD_LOGIC;
  SIGNAL nand_14_nl : STD_LOGIC;
  SIGNAL mux_229_nl : STD_LOGIC;
  SIGNAL nand_495_nl : STD_LOGIC;
  SIGNAL nand_496_nl : STD_LOGIC;
  SIGNAL mux_292_nl : STD_LOGIC;
  SIGNAL mux_291_nl : STD_LOGIC;
  SIGNAL mux_290_nl : STD_LOGIC;
  SIGNAL and_2062_nl : STD_LOGIC;
  SIGNAL mux_289_nl : STD_LOGIC;
  SIGNAL nor_2103_nl : STD_LOGIC;
  SIGNAL nor_2104_nl : STD_LOGIC;
  SIGNAL and_2063_nl : STD_LOGIC;
  SIGNAL mux_288_nl : STD_LOGIC;
  SIGNAL nor_2106_nl : STD_LOGIC;
  SIGNAL nor_2107_nl : STD_LOGIC;
  SIGNAL mux_287_nl : STD_LOGIC;
  SIGNAL nor_2109_nl : STD_LOGIC;
  SIGNAL mux_286_nl : STD_LOGIC;
  SIGNAL mux_285_nl : STD_LOGIC;
  SIGNAL nand_491_nl : STD_LOGIC;
  SIGNAL or_512_nl : STD_LOGIC;
  SIGNAL nor_2112_nl : STD_LOGIC;
  SIGNAL mux_284_nl : STD_LOGIC;
  SIGNAL or_508_nl : STD_LOGIC;
  SIGNAL or_507_nl : STD_LOGIC;
  SIGNAL mux_283_nl : STD_LOGIC;
  SIGNAL nand_17_nl : STD_LOGIC;
  SIGNAL mux_281_nl : STD_LOGIC;
  SIGNAL mux_280_nl : STD_LOGIC;
  SIGNAL and_2064_nl : STD_LOGIC;
  SIGNAL or_503_nl : STD_LOGIC;
  SIGNAL and_203_nl : STD_LOGIC;
  SIGNAL mux_356_nl : STD_LOGIC;
  SIGNAL mux_355_nl : STD_LOGIC;
  SIGNAL mux_354_nl : STD_LOGIC;
  SIGNAL mux_353_nl : STD_LOGIC;
  SIGNAL or_579_nl : STD_LOGIC;
  SIGNAL or_577_nl : STD_LOGIC;
  SIGNAL mux_352_nl : STD_LOGIC;
  SIGNAL mux_351_nl : STD_LOGIC;
  SIGNAL mux_350_nl : STD_LOGIC;
  SIGNAL mux_349_nl : STD_LOGIC;
  SIGNAL or_576_nl : STD_LOGIC;
  SIGNAL mux_348_nl : STD_LOGIC;
  SIGNAL or_567_nl : STD_LOGIC;
  SIGNAL mux_345_nl : STD_LOGIC;
  SIGNAL mux_344_nl : STD_LOGIC;
  SIGNAL mux_343_nl : STD_LOGIC;
  SIGNAL or_566_nl : STD_LOGIC;
  SIGNAL mux_342_nl : STD_LOGIC;
  SIGNAL or_565_nl : STD_LOGIC;
  SIGNAL mux_341_nl : STD_LOGIC;
  SIGNAL or_563_nl : STD_LOGIC;
  SIGNAL mux_339_nl : STD_LOGIC;
  SIGNAL mux_338_nl : STD_LOGIC;
  SIGNAL or_557_nl : STD_LOGIC;
  SIGNAL or_556_nl : STD_LOGIC;
  SIGNAL mux_337_nl : STD_LOGIC;
  SIGNAL mux_336_nl : STD_LOGIC;
  SIGNAL or_553_nl : STD_LOGIC;
  SIGNAL nand_21_nl : STD_LOGIC;
  SIGNAL mux_335_nl : STD_LOGIC;
  SIGNAL or_552_nl : STD_LOGIC;
  SIGNAL mux_334_nl : STD_LOGIC;
  SIGNAL mux_407_nl : STD_LOGIC;
  SIGNAL mux_406_nl : STD_LOGIC;
  SIGNAL mux_405_nl : STD_LOGIC;
  SIGNAL and_2041_nl : STD_LOGIC;
  SIGNAL mux_404_nl : STD_LOGIC;
  SIGNAL nor_2078_nl : STD_LOGIC;
  SIGNAL nor_2079_nl : STD_LOGIC;
  SIGNAL nor_2080_nl : STD_LOGIC;
  SIGNAL and_2042_nl : STD_LOGIC;
  SIGNAL mux_402_nl : STD_LOGIC;
  SIGNAL nor_2082_nl : STD_LOGIC;
  SIGNAL mux_401_nl : STD_LOGIC;
  SIGNAL mux_400_nl : STD_LOGIC;
  SIGNAL mux_399_nl : STD_LOGIC;
  SIGNAL nor_2083_nl : STD_LOGIC;
  SIGNAL or_640_nl : STD_LOGIC;
  SIGNAL nor_2084_nl : STD_LOGIC;
  SIGNAL mux_398_nl : STD_LOGIC;
  SIGNAL or_635_nl : STD_LOGIC;
  SIGNAL mux_397_nl : STD_LOGIC;
  SIGNAL or_630_nl : STD_LOGIC;
  SIGNAL mux_396_nl : STD_LOGIC;
  SIGNAL or_629_nl : STD_LOGIC;
  SIGNAL mux_395_nl : STD_LOGIC;
  SIGNAL mux_394_nl : STD_LOGIC;
  SIGNAL mux_393_nl : STD_LOGIC;
  SIGNAL mux_392_nl : STD_LOGIC;
  SIGNAL or_627_nl : STD_LOGIC;
  SIGNAL or_621_nl : STD_LOGIC;
  SIGNAL mux_390_nl : STD_LOGIC;
  SIGNAL or_620_nl : STD_LOGIC;
  SIGNAL or_672_nl : STD_LOGIC;
  SIGNAL mux_439_nl : STD_LOGIC;
  SIGNAL mux_438_nl : STD_LOGIC;
  SIGNAL mux_454_nl : STD_LOGIC;
  SIGNAL mux_453_nl : STD_LOGIC;
  SIGNAL mux_452_nl : STD_LOGIC;
  SIGNAL and_2031_nl : STD_LOGIC;
  SIGNAL mux_451_nl : STD_LOGIC;
  SIGNAL nor_2064_nl : STD_LOGIC;
  SIGNAL nor_2065_nl : STD_LOGIC;
  SIGNAL nor_2067_nl : STD_LOGIC;
  SIGNAL mux_450_nl : STD_LOGIC;
  SIGNAL nor_2069_nl : STD_LOGIC;
  SIGNAL mux_449_nl : STD_LOGIC;
  SIGNAL mux_448_nl : STD_LOGIC;
  SIGNAL nand_482_nl : STD_LOGIC;
  SIGNAL or_699_nl : STD_LOGIC;
  SIGNAL nor_2072_nl : STD_LOGIC;
  SIGNAL mux_447_nl : STD_LOGIC;
  SIGNAL or_695_nl : STD_LOGIC;
  SIGNAL mux_446_nl : STD_LOGIC;
  SIGNAL or_694_nl : STD_LOGIC;
  SIGNAL or_687_nl : STD_LOGIC;
  SIGNAL mux_444_nl : STD_LOGIC;
  SIGNAL nand_26_nl : STD_LOGIC;
  SIGNAL mux_443_nl : STD_LOGIC;
  SIGNAL nand_483_nl : STD_LOGIC;
  SIGNAL nand_484_nl : STD_LOGIC;
  SIGNAL mux_503_nl : STD_LOGIC;
  SIGNAL mux_502_nl : STD_LOGIC;
  SIGNAL mux_501_nl : STD_LOGIC;
  SIGNAL and_2019_nl : STD_LOGIC;
  SIGNAL mux_500_nl : STD_LOGIC;
  SIGNAL and_2020_nl : STD_LOGIC;
  SIGNAL nor_2050_nl : STD_LOGIC;
  SIGNAL and_2021_nl : STD_LOGIC;
  SIGNAL mux_499_nl : STD_LOGIC;
  SIGNAL nor_2052_nl : STD_LOGIC;
  SIGNAL nor_2053_nl : STD_LOGIC;
  SIGNAL mux_498_nl : STD_LOGIC;
  SIGNAL nor_2055_nl : STD_LOGIC;
  SIGNAL mux_497_nl : STD_LOGIC;
  SIGNAL mux_496_nl : STD_LOGIC;
  SIGNAL nand_478_nl : STD_LOGIC;
  SIGNAL or_750_nl : STD_LOGIC;
  SIGNAL nor_2058_nl : STD_LOGIC;
  SIGNAL mux_495_nl : STD_LOGIC;
  SIGNAL or_746_nl : STD_LOGIC;
  SIGNAL or_744_nl : STD_LOGIC;
  SIGNAL mux_494_nl : STD_LOGIC;
  SIGNAL nand_29_nl : STD_LOGIC;
  SIGNAL mux_492_nl : STD_LOGIC;
  SIGNAL mux_491_nl : STD_LOGIC;
  SIGNAL and_2022_nl : STD_LOGIC;
  SIGNAL or_738_nl : STD_LOGIC;
  SIGNAL and_259_nl : STD_LOGIC;
  SIGNAL mux_565_nl : STD_LOGIC;
  SIGNAL mux_564_nl : STD_LOGIC;
  SIGNAL mux_563_nl : STD_LOGIC;
  SIGNAL mux_562_nl : STD_LOGIC;
  SIGNAL mux_561_nl : STD_LOGIC;
  SIGNAL mux_560_nl : STD_LOGIC;
  SIGNAL or_820_nl : STD_LOGIC;
  SIGNAL mux_559_nl : STD_LOGIC;
  SIGNAL mux_558_nl : STD_LOGIC;
  SIGNAL mux_557_nl : STD_LOGIC;
  SIGNAL or_815_nl : STD_LOGIC;
  SIGNAL or_812_nl : STD_LOGIC;
  SIGNAL or_807_nl : STD_LOGIC;
  SIGNAL mux_554_nl : STD_LOGIC;
  SIGNAL mux_553_nl : STD_LOGIC;
  SIGNAL mux_552_nl : STD_LOGIC;
  SIGNAL or_806_nl : STD_LOGIC;
  SIGNAL mux_551_nl : STD_LOGIC;
  SIGNAL or_805_nl : STD_LOGIC;
  SIGNAL mux_550_nl : STD_LOGIC;
  SIGNAL or_803_nl : STD_LOGIC;
  SIGNAL mux_548_nl : STD_LOGIC;
  SIGNAL mux_547_nl : STD_LOGIC;
  SIGNAL or_797_nl : STD_LOGIC;
  SIGNAL or_796_nl : STD_LOGIC;
  SIGNAL mux_546_nl : STD_LOGIC;
  SIGNAL mux_545_nl : STD_LOGIC;
  SIGNAL or_793_nl : STD_LOGIC;
  SIGNAL nand_33_nl : STD_LOGIC;
  SIGNAL mux_544_nl : STD_LOGIC;
  SIGNAL or_792_nl : STD_LOGIC;
  SIGNAL mux_543_nl : STD_LOGIC;
  SIGNAL mux_613_nl : STD_LOGIC;
  SIGNAL mux_612_nl : STD_LOGIC;
  SIGNAL mux_611_nl : STD_LOGIC;
  SIGNAL and_1999_nl : STD_LOGIC;
  SIGNAL mux_610_nl : STD_LOGIC;
  SIGNAL nor_2027_nl : STD_LOGIC;
  SIGNAL nor_2028_nl : STD_LOGIC;
  SIGNAL nor_2029_nl : STD_LOGIC;
  SIGNAL and_2000_nl : STD_LOGIC;
  SIGNAL mux_608_nl : STD_LOGIC;
  SIGNAL nor_2031_nl : STD_LOGIC;
  SIGNAL mux_607_nl : STD_LOGIC;
  SIGNAL mux_606_nl : STD_LOGIC;
  SIGNAL mux_605_nl : STD_LOGIC;
  SIGNAL or_869_nl : STD_LOGIC;
  SIGNAL nor_2033_nl : STD_LOGIC;
  SIGNAL mux_604_nl : STD_LOGIC;
  SIGNAL or_865_nl : STD_LOGIC;
  SIGNAL mux_603_nl : STD_LOGIC;
  SIGNAL or_862_nl : STD_LOGIC;
  SIGNAL mux_602_nl : STD_LOGIC;
  SIGNAL or_861_nl : STD_LOGIC;
  SIGNAL mux_601_nl : STD_LOGIC;
  SIGNAL mux_600_nl : STD_LOGIC;
  SIGNAL mux_599_nl : STD_LOGIC;
  SIGNAL nor_2034_nl : STD_LOGIC;
  SIGNAL or_858_nl : STD_LOGIC;
  SIGNAL nand_35_nl : STD_LOGIC;
  SIGNAL or_897_nl : STD_LOGIC;
  SIGNAL mux_645_nl : STD_LOGIC;
  SIGNAL mux_644_nl : STD_LOGIC;
  SIGNAL mux_660_nl : STD_LOGIC;
  SIGNAL mux_659_nl : STD_LOGIC;
  SIGNAL mux_658_nl : STD_LOGIC;
  SIGNAL and_1989_nl : STD_LOGIC;
  SIGNAL mux_657_nl : STD_LOGIC;
  SIGNAL nor_2012_nl : STD_LOGIC;
  SIGNAL nor_2013_nl : STD_LOGIC;
  SIGNAL nor_2015_nl : STD_LOGIC;
  SIGNAL mux_656_nl : STD_LOGIC;
  SIGNAL nor_2017_nl : STD_LOGIC;
  SIGNAL mux_655_nl : STD_LOGIC;
  SIGNAL mux_654_nl : STD_LOGIC;
  SIGNAL nand_468_nl : STD_LOGIC;
  SIGNAL or_921_nl : STD_LOGIC;
  SIGNAL nor_2020_nl : STD_LOGIC;
  SIGNAL mux_653_nl : STD_LOGIC;
  SIGNAL or_917_nl : STD_LOGIC;
  SIGNAL mux_652_nl : STD_LOGIC;
  SIGNAL or_916_nl : STD_LOGIC;
  SIGNAL or_912_nl : STD_LOGIC;
  SIGNAL mux_650_nl : STD_LOGIC;
  SIGNAL nand_39_nl : STD_LOGIC;
  SIGNAL mux_649_nl : STD_LOGIC;
  SIGNAL nand_469_nl : STD_LOGIC;
  SIGNAL nand_470_nl : STD_LOGIC;
  SIGNAL mux_709_nl : STD_LOGIC;
  SIGNAL mux_708_nl : STD_LOGIC;
  SIGNAL mux_707_nl : STD_LOGIC;
  SIGNAL and_1977_nl : STD_LOGIC;
  SIGNAL mux_706_nl : STD_LOGIC;
  SIGNAL and_1978_nl : STD_LOGIC;
  SIGNAL nor_1998_nl : STD_LOGIC;
  SIGNAL and_1979_nl : STD_LOGIC;
  SIGNAL mux_705_nl : STD_LOGIC;
  SIGNAL nor_2000_nl : STD_LOGIC;
  SIGNAL nor_2001_nl : STD_LOGIC;
  SIGNAL mux_704_nl : STD_LOGIC;
  SIGNAL nor_2003_nl : STD_LOGIC;
  SIGNAL mux_703_nl : STD_LOGIC;
  SIGNAL mux_702_nl : STD_LOGIC;
  SIGNAL nand_465_nl : STD_LOGIC;
  SIGNAL or_970_nl : STD_LOGIC;
  SIGNAL nor_2006_nl : STD_LOGIC;
  SIGNAL mux_701_nl : STD_LOGIC;
  SIGNAL or_966_nl : STD_LOGIC;
  SIGNAL or_964_nl : STD_LOGIC;
  SIGNAL mux_700_nl : STD_LOGIC;
  SIGNAL nand_42_nl : STD_LOGIC;
  SIGNAL mux_698_nl : STD_LOGIC;
  SIGNAL mux_697_nl : STD_LOGIC;
  SIGNAL and_1980_nl : STD_LOGIC;
  SIGNAL or_958_nl : STD_LOGIC;
  SIGNAL and_313_nl : STD_LOGIC;
  SIGNAL mux_771_nl : STD_LOGIC;
  SIGNAL mux_770_nl : STD_LOGIC;
  SIGNAL mux_769_nl : STD_LOGIC;
  SIGNAL mux_768_nl : STD_LOGIC;
  SIGNAL or_1036_nl : STD_LOGIC;
  SIGNAL or_1034_nl : STD_LOGIC;
  SIGNAL mux_767_nl : STD_LOGIC;
  SIGNAL mux_766_nl : STD_LOGIC;
  SIGNAL mux_765_nl : STD_LOGIC;
  SIGNAL mux_764_nl : STD_LOGIC;
  SIGNAL or_1033_nl : STD_LOGIC;
  SIGNAL mux_763_nl : STD_LOGIC;
  SIGNAL or_1024_nl : STD_LOGIC;
  SIGNAL mux_760_nl : STD_LOGIC;
  SIGNAL mux_759_nl : STD_LOGIC;
  SIGNAL mux_758_nl : STD_LOGIC;
  SIGNAL or_1023_nl : STD_LOGIC;
  SIGNAL mux_757_nl : STD_LOGIC;
  SIGNAL or_1022_nl : STD_LOGIC;
  SIGNAL mux_756_nl : STD_LOGIC;
  SIGNAL or_1020_nl : STD_LOGIC;
  SIGNAL mux_754_nl : STD_LOGIC;
  SIGNAL mux_753_nl : STD_LOGIC;
  SIGNAL or_1014_nl : STD_LOGIC;
  SIGNAL or_1013_nl : STD_LOGIC;
  SIGNAL mux_752_nl : STD_LOGIC;
  SIGNAL mux_751_nl : STD_LOGIC;
  SIGNAL or_1010_nl : STD_LOGIC;
  SIGNAL nand_46_nl : STD_LOGIC;
  SIGNAL mux_750_nl : STD_LOGIC;
  SIGNAL or_1009_nl : STD_LOGIC;
  SIGNAL mux_749_nl : STD_LOGIC;
  SIGNAL mux_819_nl : STD_LOGIC;
  SIGNAL mux_818_nl : STD_LOGIC;
  SIGNAL mux_817_nl : STD_LOGIC;
  SIGNAL and_1956_nl : STD_LOGIC;
  SIGNAL mux_816_nl : STD_LOGIC;
  SIGNAL and_1957_nl : STD_LOGIC;
  SIGNAL nor_1976_nl : STD_LOGIC;
  SIGNAL nor_1977_nl : STD_LOGIC;
  SIGNAL and_1958_nl : STD_LOGIC;
  SIGNAL mux_814_nl : STD_LOGIC;
  SIGNAL nor_1979_nl : STD_LOGIC;
  SIGNAL mux_813_nl : STD_LOGIC;
  SIGNAL mux_812_nl : STD_LOGIC;
  SIGNAL mux_811_nl : STD_LOGIC;
  SIGNAL nor_1980_nl : STD_LOGIC;
  SIGNAL or_1090_nl : STD_LOGIC;
  SIGNAL nor_1981_nl : STD_LOGIC;
  SIGNAL mux_810_nl : STD_LOGIC;
  SIGNAL or_1086_nl : STD_LOGIC;
  SIGNAL mux_809_nl : STD_LOGIC;
  SIGNAL or_1081_nl : STD_LOGIC;
  SIGNAL mux_808_nl : STD_LOGIC;
  SIGNAL or_1080_nl : STD_LOGIC;
  SIGNAL mux_807_nl : STD_LOGIC;
  SIGNAL mux_806_nl : STD_LOGIC;
  SIGNAL or_1078_nl : STD_LOGIC;
  SIGNAL mux_805_nl : STD_LOGIC;
  SIGNAL nor_1982_nl : STD_LOGIC;
  SIGNAL or_1076_nl : STD_LOGIC;
  SIGNAL nand_48_nl : STD_LOGIC;
  SIGNAL or_1121_nl : STD_LOGIC;
  SIGNAL mux_851_nl : STD_LOGIC;
  SIGNAL mux_850_nl : STD_LOGIC;
  SIGNAL mux_866_nl : STD_LOGIC;
  SIGNAL mux_865_nl : STD_LOGIC;
  SIGNAL mux_864_nl : STD_LOGIC;
  SIGNAL and_1944_nl : STD_LOGIC;
  SIGNAL mux_863_nl : STD_LOGIC;
  SIGNAL and_1945_nl : STD_LOGIC;
  SIGNAL nor_1962_nl : STD_LOGIC;
  SIGNAL nor_1964_nl : STD_LOGIC;
  SIGNAL mux_862_nl : STD_LOGIC;
  SIGNAL nor_1966_nl : STD_LOGIC;
  SIGNAL mux_861_nl : STD_LOGIC;
  SIGNAL mux_860_nl : STD_LOGIC;
  SIGNAL nand_453_nl : STD_LOGIC;
  SIGNAL or_1148_nl : STD_LOGIC;
  SIGNAL nor_1969_nl : STD_LOGIC;
  SIGNAL mux_859_nl : STD_LOGIC;
  SIGNAL or_1144_nl : STD_LOGIC;
  SIGNAL mux_858_nl : STD_LOGIC;
  SIGNAL or_1143_nl : STD_LOGIC;
  SIGNAL or_1136_nl : STD_LOGIC;
  SIGNAL mux_856_nl : STD_LOGIC;
  SIGNAL nand_52_nl : STD_LOGIC;
  SIGNAL mux_855_nl : STD_LOGIC;
  SIGNAL nand_454_nl : STD_LOGIC;
  SIGNAL nand_455_nl : STD_LOGIC;
  SIGNAL mux_915_nl : STD_LOGIC;
  SIGNAL mux_914_nl : STD_LOGIC;
  SIGNAL mux_913_nl : STD_LOGIC;
  SIGNAL and_1930_nl : STD_LOGIC;
  SIGNAL mux_912_nl : STD_LOGIC;
  SIGNAL and_1931_nl : STD_LOGIC;
  SIGNAL nor_1949_nl : STD_LOGIC;
  SIGNAL and_1932_nl : STD_LOGIC;
  SIGNAL mux_911_nl : STD_LOGIC;
  SIGNAL nor_1951_nl : STD_LOGIC;
  SIGNAL nor_1952_nl : STD_LOGIC;
  SIGNAL mux_910_nl : STD_LOGIC;
  SIGNAL nor_1954_nl : STD_LOGIC;
  SIGNAL mux_909_nl : STD_LOGIC;
  SIGNAL mux_908_nl : STD_LOGIC;
  SIGNAL nand_445_nl : STD_LOGIC;
  SIGNAL nand_446_nl : STD_LOGIC;
  SIGNAL nor_1956_nl : STD_LOGIC;
  SIGNAL mux_907_nl : STD_LOGIC;
  SIGNAL or_1192_nl : STD_LOGIC;
  SIGNAL or_1190_nl : STD_LOGIC;
  SIGNAL mux_906_nl : STD_LOGIC;
  SIGNAL nand_55_nl : STD_LOGIC;
  SIGNAL mux_904_nl : STD_LOGIC;
  SIGNAL mux_903_nl : STD_LOGIC;
  SIGNAL and_1934_nl : STD_LOGIC;
  SIGNAL and_360_nl : STD_LOGIC;
  SIGNAL mux_978_nl : STD_LOGIC;
  SIGNAL mux_977_nl : STD_LOGIC;
  SIGNAL mux_976_nl : STD_LOGIC;
  SIGNAL mux_975_nl : STD_LOGIC;
  SIGNAL mux_974_nl : STD_LOGIC;
  SIGNAL mux_973_nl : STD_LOGIC;
  SIGNAL or_1264_nl : STD_LOGIC;
  SIGNAL mux_972_nl : STD_LOGIC;
  SIGNAL mux_971_nl : STD_LOGIC;
  SIGNAL mux_970_nl : STD_LOGIC;
  SIGNAL or_1259_nl : STD_LOGIC;
  SIGNAL or_1256_nl : STD_LOGIC;
  SIGNAL or_1251_nl : STD_LOGIC;
  SIGNAL mux_967_nl : STD_LOGIC;
  SIGNAL mux_966_nl : STD_LOGIC;
  SIGNAL mux_965_nl : STD_LOGIC;
  SIGNAL or_1250_nl : STD_LOGIC;
  SIGNAL mux_964_nl : STD_LOGIC;
  SIGNAL or_1249_nl : STD_LOGIC;
  SIGNAL mux_963_nl : STD_LOGIC;
  SIGNAL or_1248_nl : STD_LOGIC;
  SIGNAL mux_961_nl : STD_LOGIC;
  SIGNAL mux_960_nl : STD_LOGIC;
  SIGNAL or_1242_nl : STD_LOGIC;
  SIGNAL or_1241_nl : STD_LOGIC;
  SIGNAL mux_959_nl : STD_LOGIC;
  SIGNAL or_1240_nl : STD_LOGIC;
  SIGNAL mux_958_nl : STD_LOGIC;
  SIGNAL or_1238_nl : STD_LOGIC;
  SIGNAL nand_59_nl : STD_LOGIC;
  SIGNAL mux_957_nl : STD_LOGIC;
  SIGNAL or_1237_nl : STD_LOGIC;
  SIGNAL mux_956_nl : STD_LOGIC;
  SIGNAL mux_955_nl : STD_LOGIC;
  SIGNAL or_1234_nl : STD_LOGIC;
  SIGNAL mux_1029_nl : STD_LOGIC;
  SIGNAL mux_1028_nl : STD_LOGIC;
  SIGNAL mux_1027_nl : STD_LOGIC;
  SIGNAL and_1905_nl : STD_LOGIC;
  SIGNAL mux_1026_nl : STD_LOGIC;
  SIGNAL nor_1925_nl : STD_LOGIC;
  SIGNAL nor_1926_nl : STD_LOGIC;
  SIGNAL nor_1927_nl : STD_LOGIC;
  SIGNAL and_1906_nl : STD_LOGIC;
  SIGNAL mux_1024_nl : STD_LOGIC;
  SIGNAL nor_1929_nl : STD_LOGIC;
  SIGNAL mux_1023_nl : STD_LOGIC;
  SIGNAL mux_1022_nl : STD_LOGIC;
  SIGNAL mux_1021_nl : STD_LOGIC;
  SIGNAL mux_1020_nl : STD_LOGIC;
  SIGNAL or_1314_nl : STD_LOGIC;
  SIGNAL nor_1931_nl : STD_LOGIC;
  SIGNAL mux_1019_nl : STD_LOGIC;
  SIGNAL or_1311_nl : STD_LOGIC;
  SIGNAL mux_1018_nl : STD_LOGIC;
  SIGNAL or_1308_nl : STD_LOGIC;
  SIGNAL mux_1017_nl : STD_LOGIC;
  SIGNAL or_1307_nl : STD_LOGIC;
  SIGNAL mux_1016_nl : STD_LOGIC;
  SIGNAL mux_1015_nl : STD_LOGIC;
  SIGNAL mux_1014_nl : STD_LOGIC;
  SIGNAL nor_1932_nl : STD_LOGIC;
  SIGNAL or_1304_nl : STD_LOGIC;
  SIGNAL nand_61_nl : STD_LOGIC;
  SIGNAL mux_1013_nl : STD_LOGIC;
  SIGNAL nor_1933_nl : STD_LOGIC;
  SIGNAL or_1301_nl : STD_LOGIC;
  SIGNAL mux_1062_nl : STD_LOGIC;
  SIGNAL mux_1061_nl : STD_LOGIC;
  SIGNAL mux_1058_nl : STD_LOGIC;
  SIGNAL or_1343_nl : STD_LOGIC;
  SIGNAL mux_1079_nl : STD_LOGIC;
  SIGNAL mux_1078_nl : STD_LOGIC;
  SIGNAL mux_1077_nl : STD_LOGIC;
  SIGNAL and_1895_nl : STD_LOGIC;
  SIGNAL mux_1076_nl : STD_LOGIC;
  SIGNAL nor_1912_nl : STD_LOGIC;
  SIGNAL nor_1913_nl : STD_LOGIC;
  SIGNAL nor_1915_nl : STD_LOGIC;
  SIGNAL mux_1075_nl : STD_LOGIC;
  SIGNAL nor_1917_nl : STD_LOGIC;
  SIGNAL mux_1074_nl : STD_LOGIC;
  SIGNAL mux_1073_nl : STD_LOGIC;
  SIGNAL mux_1072_nl : STD_LOGIC;
  SIGNAL nand_434_nl : STD_LOGIC;
  SIGNAL or_1367_nl : STD_LOGIC;
  SIGNAL nor_1920_nl : STD_LOGIC;
  SIGNAL mux_1071_nl : STD_LOGIC;
  SIGNAL or_1364_nl : STD_LOGIC;
  SIGNAL mux_1070_nl : STD_LOGIC;
  SIGNAL or_1363_nl : STD_LOGIC;
  SIGNAL or_1359_nl : STD_LOGIC;
  SIGNAL mux_1068_nl : STD_LOGIC;
  SIGNAL nand_65_nl : STD_LOGIC;
  SIGNAL mux_1067_nl : STD_LOGIC;
  SIGNAL and_399_nl : STD_LOGIC;
  SIGNAL mux_1066_nl : STD_LOGIC;
  SIGNAL nor_1921_nl : STD_LOGIC;
  SIGNAL or_1354_nl : STD_LOGIC;
  SIGNAL mux_1131_nl : STD_LOGIC;
  SIGNAL mux_1130_nl : STD_LOGIC;
  SIGNAL mux_1129_nl : STD_LOGIC;
  SIGNAL and_1884_nl : STD_LOGIC;
  SIGNAL mux_1128_nl : STD_LOGIC;
  SIGNAL and_2140_nl : STD_LOGIC;
  SIGNAL nor_1898_nl : STD_LOGIC;
  SIGNAL and_1885_nl : STD_LOGIC;
  SIGNAL mux_1127_nl : STD_LOGIC;
  SIGNAL nor_1900_nl : STD_LOGIC;
  SIGNAL nor_1901_nl : STD_LOGIC;
  SIGNAL mux_1126_nl : STD_LOGIC;
  SIGNAL nor_1903_nl : STD_LOGIC;
  SIGNAL mux_1125_nl : STD_LOGIC;
  SIGNAL mux_1124_nl : STD_LOGIC;
  SIGNAL mux_1123_nl : STD_LOGIC;
  SIGNAL nand_430_nl : STD_LOGIC;
  SIGNAL or_1419_nl : STD_LOGIC;
  SIGNAL nor_1906_nl : STD_LOGIC;
  SIGNAL mux_1122_nl : STD_LOGIC;
  SIGNAL or_1416_nl : STD_LOGIC;
  SIGNAL or_1415_nl : STD_LOGIC;
  SIGNAL mux_1121_nl : STD_LOGIC;
  SIGNAL nand_68_nl : STD_LOGIC;
  SIGNAL mux_1119_nl : STD_LOGIC;
  SIGNAL mux_1118_nl : STD_LOGIC;
  SIGNAL and_1886_nl : STD_LOGIC;
  SIGNAL or_1411_nl : STD_LOGIC;
  SIGNAL mux_1117_nl : STD_LOGIC;
  SIGNAL nor_1907_nl : STD_LOGIC;
  SIGNAL or_1407_nl : STD_LOGIC;
  SIGNAL mux_1195_nl : STD_LOGIC;
  SIGNAL mux_1194_nl : STD_LOGIC;
  SIGNAL mux_1193_nl : STD_LOGIC;
  SIGNAL mux_1192_nl : STD_LOGIC;
  SIGNAL or_1488_nl : STD_LOGIC;
  SIGNAL or_1486_nl : STD_LOGIC;
  SIGNAL mux_1191_nl : STD_LOGIC;
  SIGNAL mux_1190_nl : STD_LOGIC;
  SIGNAL mux_1189_nl : STD_LOGIC;
  SIGNAL mux_1188_nl : STD_LOGIC;
  SIGNAL or_1485_nl : STD_LOGIC;
  SIGNAL mux_1187_nl : STD_LOGIC;
  SIGNAL or_1476_nl : STD_LOGIC;
  SIGNAL mux_1184_nl : STD_LOGIC;
  SIGNAL mux_1183_nl : STD_LOGIC;
  SIGNAL mux_1182_nl : STD_LOGIC;
  SIGNAL or_1475_nl : STD_LOGIC;
  SIGNAL mux_1181_nl : STD_LOGIC;
  SIGNAL or_1474_nl : STD_LOGIC;
  SIGNAL mux_1180_nl : STD_LOGIC;
  SIGNAL or_1473_nl : STD_LOGIC;
  SIGNAL mux_1178_nl : STD_LOGIC;
  SIGNAL mux_1177_nl : STD_LOGIC;
  SIGNAL or_1467_nl : STD_LOGIC;
  SIGNAL or_1466_nl : STD_LOGIC;
  SIGNAL mux_1176_nl : STD_LOGIC;
  SIGNAL or_1465_nl : STD_LOGIC;
  SIGNAL mux_1175_nl : STD_LOGIC;
  SIGNAL or_1463_nl : STD_LOGIC;
  SIGNAL nand_72_nl : STD_LOGIC;
  SIGNAL mux_1174_nl : STD_LOGIC;
  SIGNAL or_1462_nl : STD_LOGIC;
  SIGNAL mux_1173_nl : STD_LOGIC;
  SIGNAL mux_1172_nl : STD_LOGIC;
  SIGNAL or_1459_nl : STD_LOGIC;
  SIGNAL mux_1247_nl : STD_LOGIC;
  SIGNAL mux_1246_nl : STD_LOGIC;
  SIGNAL mux_1245_nl : STD_LOGIC;
  SIGNAL and_1862_nl : STD_LOGIC;
  SIGNAL mux_1244_nl : STD_LOGIC;
  SIGNAL and_2132_nl : STD_LOGIC;
  SIGNAL nor_1872_nl : STD_LOGIC;
  SIGNAL nor_1873_nl : STD_LOGIC;
  SIGNAL and_1863_nl : STD_LOGIC;
  SIGNAL mux_1242_nl : STD_LOGIC;
  SIGNAL nor_1874_nl : STD_LOGIC;
  SIGNAL nor_1875_nl : STD_LOGIC;
  SIGNAL mux_1241_nl : STD_LOGIC;
  SIGNAL mux_1240_nl : STD_LOGIC;
  SIGNAL mux_1239_nl : STD_LOGIC;
  SIGNAL mux_1238_nl : STD_LOGIC;
  SIGNAL or_1551_nl : STD_LOGIC;
  SIGNAL nor_1877_nl : STD_LOGIC;
  SIGNAL mux_1237_nl : STD_LOGIC;
  SIGNAL or_1548_nl : STD_LOGIC;
  SIGNAL mux_1236_nl : STD_LOGIC;
  SIGNAL or_1545_nl : STD_LOGIC;
  SIGNAL or_1543_nl : STD_LOGIC;
  SIGNAL mux_1235_nl : STD_LOGIC;
  SIGNAL nand_547_nl : STD_LOGIC;
  SIGNAL mux_1234_nl : STD_LOGIC;
  SIGNAL mux_1233_nl : STD_LOGIC;
  SIGNAL mux_1232_nl : STD_LOGIC;
  SIGNAL nor_1878_nl : STD_LOGIC;
  SIGNAL or_1534_nl : STD_LOGIC;
  SIGNAL mux_1231_nl : STD_LOGIC;
  SIGNAL nand_74_nl : STD_LOGIC;
  SIGNAL mux_1230_nl : STD_LOGIC;
  SIGNAL nor_1880_nl : STD_LOGIC;
  SIGNAL or_1530_nl : STD_LOGIC;
  SIGNAL mux_1280_nl : STD_LOGIC;
  SIGNAL mux_1279_nl : STD_LOGIC;
  SIGNAL mux_1276_nl : STD_LOGIC;
  SIGNAL or_1581_nl : STD_LOGIC;
  SIGNAL mux_1297_nl : STD_LOGIC;
  SIGNAL mux_1296_nl : STD_LOGIC;
  SIGNAL mux_1295_nl : STD_LOGIC;
  SIGNAL and_1851_nl : STD_LOGIC;
  SIGNAL mux_1294_nl : STD_LOGIC;
  SIGNAL and_2131_nl : STD_LOGIC;
  SIGNAL nor_1859_nl : STD_LOGIC;
  SIGNAL nor_1861_nl : STD_LOGIC;
  SIGNAL mux_1293_nl : STD_LOGIC;
  SIGNAL nor_1863_nl : STD_LOGIC;
  SIGNAL mux_1292_nl : STD_LOGIC;
  SIGNAL mux_1291_nl : STD_LOGIC;
  SIGNAL mux_1290_nl : STD_LOGIC;
  SIGNAL nand_419_nl : STD_LOGIC;
  SIGNAL or_1609_nl : STD_LOGIC;
  SIGNAL nor_1866_nl : STD_LOGIC;
  SIGNAL mux_1289_nl : STD_LOGIC;
  SIGNAL or_1606_nl : STD_LOGIC;
  SIGNAL mux_1288_nl : STD_LOGIC;
  SIGNAL or_1605_nl : STD_LOGIC;
  SIGNAL or_1600_nl : STD_LOGIC;
  SIGNAL or_1598_nl : STD_LOGIC;
  SIGNAL mux_1286_nl : STD_LOGIC;
  SIGNAL or_1597_nl : STD_LOGIC;
  SIGNAL nand_78_nl : STD_LOGIC;
  SIGNAL mux_1285_nl : STD_LOGIC;
  SIGNAL and_444_nl : STD_LOGIC;
  SIGNAL mux_1284_nl : STD_LOGIC;
  SIGNAL nor_1867_nl : STD_LOGIC;
  SIGNAL or_1591_nl : STD_LOGIC;
  SIGNAL mux_1349_nl : STD_LOGIC;
  SIGNAL mux_1348_nl : STD_LOGIC;
  SIGNAL mux_1347_nl : STD_LOGIC;
  SIGNAL and_1838_nl : STD_LOGIC;
  SIGNAL mux_1346_nl : STD_LOGIC;
  SIGNAL and_2139_nl : STD_LOGIC;
  SIGNAL nor_1843_nl : STD_LOGIC;
  SIGNAL and_1839_nl : STD_LOGIC;
  SIGNAL mux_1345_nl : STD_LOGIC;
  SIGNAL nor_1845_nl : STD_LOGIC;
  SIGNAL nor_1846_nl : STD_LOGIC;
  SIGNAL mux_1344_nl : STD_LOGIC;
  SIGNAL nor_1848_nl : STD_LOGIC;
  SIGNAL mux_1343_nl : STD_LOGIC;
  SIGNAL mux_1342_nl : STD_LOGIC;
  SIGNAL mux_1341_nl : STD_LOGIC;
  SIGNAL nand_411_nl : STD_LOGIC;
  SIGNAL nand_413_nl : STD_LOGIC;
  SIGNAL nor_1851_nl : STD_LOGIC;
  SIGNAL mux_1340_nl : STD_LOGIC;
  SIGNAL or_1663_nl : STD_LOGIC;
  SIGNAL or_1661_nl : STD_LOGIC;
  SIGNAL mux_1339_nl : STD_LOGIC;
  SIGNAL nand_81_nl : STD_LOGIC;
  SIGNAL mux_1337_nl : STD_LOGIC;
  SIGNAL mux_1336_nl : STD_LOGIC;
  SIGNAL and_1840_nl : STD_LOGIC;
  SIGNAL or_1655_nl : STD_LOGIC;
  SIGNAL mux_1335_nl : STD_LOGIC;
  SIGNAL nor_1852_nl : STD_LOGIC;
  SIGNAL nand_415_nl : STD_LOGIC;
  SIGNAL mux_1413_nl : STD_LOGIC;
  SIGNAL mux_1412_nl : STD_LOGIC;
  SIGNAL mux_1411_nl : STD_LOGIC;
  SIGNAL mux_1410_nl : STD_LOGIC;
  SIGNAL mux_1409_nl : STD_LOGIC;
  SIGNAL mux_1408_nl : STD_LOGIC;
  SIGNAL or_1740_nl : STD_LOGIC;
  SIGNAL mux_1407_nl : STD_LOGIC;
  SIGNAL mux_1406_nl : STD_LOGIC;
  SIGNAL mux_1405_nl : STD_LOGIC;
  SIGNAL or_1735_nl : STD_LOGIC;
  SIGNAL or_1732_nl : STD_LOGIC;
  SIGNAL or_1727_nl : STD_LOGIC;
  SIGNAL mux_1402_nl : STD_LOGIC;
  SIGNAL mux_1401_nl : STD_LOGIC;
  SIGNAL mux_1400_nl : STD_LOGIC;
  SIGNAL or_1726_nl : STD_LOGIC;
  SIGNAL mux_1399_nl : STD_LOGIC;
  SIGNAL or_1725_nl : STD_LOGIC;
  SIGNAL mux_1398_nl : STD_LOGIC;
  SIGNAL or_1724_nl : STD_LOGIC;
  SIGNAL mux_1396_nl : STD_LOGIC;
  SIGNAL mux_1395_nl : STD_LOGIC;
  SIGNAL or_1718_nl : STD_LOGIC;
  SIGNAL or_1717_nl : STD_LOGIC;
  SIGNAL mux_1394_nl : STD_LOGIC;
  SIGNAL or_1716_nl : STD_LOGIC;
  SIGNAL mux_1393_nl : STD_LOGIC;
  SIGNAL or_1714_nl : STD_LOGIC;
  SIGNAL nand_85_nl : STD_LOGIC;
  SIGNAL mux_1392_nl : STD_LOGIC;
  SIGNAL or_1713_nl : STD_LOGIC;
  SIGNAL mux_1391_nl : STD_LOGIC;
  SIGNAL mux_1390_nl : STD_LOGIC;
  SIGNAL and_1822_nl : STD_LOGIC;
  SIGNAL or_1710_nl : STD_LOGIC;
  SIGNAL mux_1464_nl : STD_LOGIC;
  SIGNAL mux_1463_nl : STD_LOGIC;
  SIGNAL mux_1462_nl : STD_LOGIC;
  SIGNAL and_1810_nl : STD_LOGIC;
  SIGNAL mux_1461_nl : STD_LOGIC;
  SIGNAL nor_1819_nl : STD_LOGIC;
  SIGNAL nor_1820_nl : STD_LOGIC;
  SIGNAL nor_1821_nl : STD_LOGIC;
  SIGNAL and_1811_nl : STD_LOGIC;
  SIGNAL mux_1459_nl : STD_LOGIC;
  SIGNAL nor_1823_nl : STD_LOGIC;
  SIGNAL mux_1458_nl : STD_LOGIC;
  SIGNAL mux_1457_nl : STD_LOGIC;
  SIGNAL mux_1456_nl : STD_LOGIC;
  SIGNAL mux_1455_nl : STD_LOGIC;
  SIGNAL nor_1824_nl : STD_LOGIC;
  SIGNAL or_1788_nl : STD_LOGIC;
  SIGNAL nor_1825_nl : STD_LOGIC;
  SIGNAL mux_1454_nl : STD_LOGIC;
  SIGNAL or_1785_nl : STD_LOGIC;
  SIGNAL mux_1453_nl : STD_LOGIC;
  SIGNAL or_1782_nl : STD_LOGIC;
  SIGNAL mux_1452_nl : STD_LOGIC;
  SIGNAL nand_401_nl : STD_LOGIC;
  SIGNAL mux_1451_nl : STD_LOGIC;
  SIGNAL mux_1450_nl : STD_LOGIC;
  SIGNAL mux_1449_nl : STD_LOGIC;
  SIGNAL nor_1826_nl : STD_LOGIC;
  SIGNAL or_1778_nl : STD_LOGIC;
  SIGNAL nand_87_nl : STD_LOGIC;
  SIGNAL mux_1448_nl : STD_LOGIC;
  SIGNAL and_2130_nl : STD_LOGIC;
  SIGNAL or_1774_nl : STD_LOGIC;
  SIGNAL or_1817_nl : STD_LOGIC;
  SIGNAL mux_1497_nl : STD_LOGIC;
  SIGNAL mux_1496_nl : STD_LOGIC;
  SIGNAL mux_1514_nl : STD_LOGIC;
  SIGNAL mux_1513_nl : STD_LOGIC;
  SIGNAL mux_1512_nl : STD_LOGIC;
  SIGNAL and_1797_nl : STD_LOGIC;
  SIGNAL mux_1511_nl : STD_LOGIC;
  SIGNAL nor_1808_nl : STD_LOGIC;
  SIGNAL nor_1809_nl : STD_LOGIC;
  SIGNAL and_1798_nl : STD_LOGIC;
  SIGNAL mux_1510_nl : STD_LOGIC;
  SIGNAL nor_1812_nl : STD_LOGIC;
  SIGNAL mux_1509_nl : STD_LOGIC;
  SIGNAL mux_1508_nl : STD_LOGIC;
  SIGNAL mux_1507_nl : STD_LOGIC;
  SIGNAL nand_392_nl : STD_LOGIC;
  SIGNAL or_1841_nl : STD_LOGIC;
  SIGNAL nor_1815_nl : STD_LOGIC;
  SIGNAL mux_1506_nl : STD_LOGIC;
  SIGNAL or_1838_nl : STD_LOGIC;
  SIGNAL mux_1505_nl : STD_LOGIC;
  SIGNAL or_1837_nl : STD_LOGIC;
  SIGNAL or_1833_nl : STD_LOGIC;
  SIGNAL mux_1503_nl : STD_LOGIC;
  SIGNAL nand_91_nl : STD_LOGIC;
  SIGNAL mux_1502_nl : STD_LOGIC;
  SIGNAL and_487_nl : STD_LOGIC;
  SIGNAL mux_1501_nl : STD_LOGIC;
  SIGNAL and_1800_nl : STD_LOGIC;
  SIGNAL or_1828_nl : STD_LOGIC;
  SIGNAL mux_1566_nl : STD_LOGIC;
  SIGNAL mux_1565_nl : STD_LOGIC;
  SIGNAL mux_1564_nl : STD_LOGIC;
  SIGNAL and_1784_nl : STD_LOGIC;
  SIGNAL mux_1563_nl : STD_LOGIC;
  SIGNAL nor_1792_nl : STD_LOGIC;
  SIGNAL nor_1793_nl : STD_LOGIC;
  SIGNAL and_1785_nl : STD_LOGIC;
  SIGNAL mux_1562_nl : STD_LOGIC;
  SIGNAL and_2144_nl : STD_LOGIC;
  SIGNAL nor_1796_nl : STD_LOGIC;
  SIGNAL mux_1561_nl : STD_LOGIC;
  SIGNAL nor_1798_nl : STD_LOGIC;
  SIGNAL mux_1560_nl : STD_LOGIC;
  SIGNAL mux_1559_nl : STD_LOGIC;
  SIGNAL mux_1558_nl : STD_LOGIC;
  SIGNAL nand_385_nl : STD_LOGIC;
  SIGNAL or_1895_nl : STD_LOGIC;
  SIGNAL nor_1801_nl : STD_LOGIC;
  SIGNAL mux_1557_nl : STD_LOGIC;
  SIGNAL or_1892_nl : STD_LOGIC;
  SIGNAL or_1890_nl : STD_LOGIC;
  SIGNAL mux_1556_nl : STD_LOGIC;
  SIGNAL nand_94_nl : STD_LOGIC;
  SIGNAL mux_1554_nl : STD_LOGIC;
  SIGNAL mux_1553_nl : STD_LOGIC;
  SIGNAL and_1787_nl : STD_LOGIC;
  SIGNAL or_1884_nl : STD_LOGIC;
  SIGNAL mux_1552_nl : STD_LOGIC;
  SIGNAL and_2129_nl : STD_LOGIC;
  SIGNAL or_1880_nl : STD_LOGIC;
  SIGNAL mux_1630_nl : STD_LOGIC;
  SIGNAL mux_1629_nl : STD_LOGIC;
  SIGNAL mux_1628_nl : STD_LOGIC;
  SIGNAL mux_1627_nl : STD_LOGIC;
  SIGNAL or_1967_nl : STD_LOGIC;
  SIGNAL or_1965_nl : STD_LOGIC;
  SIGNAL mux_1626_nl : STD_LOGIC;
  SIGNAL mux_1625_nl : STD_LOGIC;
  SIGNAL mux_1624_nl : STD_LOGIC;
  SIGNAL mux_1623_nl : STD_LOGIC;
  SIGNAL nand_550_nl : STD_LOGIC;
  SIGNAL mux_1622_nl : STD_LOGIC;
  SIGNAL or_1955_nl : STD_LOGIC;
  SIGNAL mux_1619_nl : STD_LOGIC;
  SIGNAL mux_1618_nl : STD_LOGIC;
  SIGNAL mux_1617_nl : STD_LOGIC;
  SIGNAL or_1954_nl : STD_LOGIC;
  SIGNAL mux_1616_nl : STD_LOGIC;
  SIGNAL or_1953_nl : STD_LOGIC;
  SIGNAL mux_1615_nl : STD_LOGIC;
  SIGNAL or_1952_nl : STD_LOGIC;
  SIGNAL mux_1613_nl : STD_LOGIC;
  SIGNAL mux_1612_nl : STD_LOGIC;
  SIGNAL or_1946_nl : STD_LOGIC;
  SIGNAL or_1945_nl : STD_LOGIC;
  SIGNAL mux_1611_nl : STD_LOGIC;
  SIGNAL or_1944_nl : STD_LOGIC;
  SIGNAL mux_1610_nl : STD_LOGIC;
  SIGNAL or_1942_nl : STD_LOGIC;
  SIGNAL nand_98_nl : STD_LOGIC;
  SIGNAL mux_1609_nl : STD_LOGIC;
  SIGNAL or_1941_nl : STD_LOGIC;
  SIGNAL mux_1608_nl : STD_LOGIC;
  SIGNAL mux_1607_nl : STD_LOGIC;
  SIGNAL and_1769_nl : STD_LOGIC;
  SIGNAL or_1938_nl : STD_LOGIC;
  SIGNAL mux_1681_nl : STD_LOGIC;
  SIGNAL mux_1680_nl : STD_LOGIC;
  SIGNAL mux_1679_nl : STD_LOGIC;
  SIGNAL and_1754_nl : STD_LOGIC;
  SIGNAL mux_1678_nl : STD_LOGIC;
  SIGNAL nor_1768_nl : STD_LOGIC;
  SIGNAL nor_1769_nl : STD_LOGIC;
  SIGNAL nor_1770_nl : STD_LOGIC;
  SIGNAL and_1755_nl : STD_LOGIC;
  SIGNAL mux_1676_nl : STD_LOGIC;
  SIGNAL nor_1772_nl : STD_LOGIC;
  SIGNAL mux_1675_nl : STD_LOGIC;
  SIGNAL mux_1674_nl : STD_LOGIC;
  SIGNAL mux_1673_nl : STD_LOGIC;
  SIGNAL mux_1672_nl : STD_LOGIC;
  SIGNAL nor_1773_nl : STD_LOGIC;
  SIGNAL and_1756_nl : STD_LOGIC;
  SIGNAL or_2016_nl : STD_LOGIC;
  SIGNAL nor_1774_nl : STD_LOGIC;
  SIGNAL mux_1671_nl : STD_LOGIC;
  SIGNAL or_2013_nl : STD_LOGIC;
  SIGNAL mux_1670_nl : STD_LOGIC;
  SIGNAL or_2012_nl : STD_LOGIC;
  SIGNAL or_2009_nl : STD_LOGIC;
  SIGNAL mux_1669_nl : STD_LOGIC;
  SIGNAL nand_362_nl : STD_LOGIC;
  SIGNAL mux_1668_nl : STD_LOGIC;
  SIGNAL mux_1667_nl : STD_LOGIC;
  SIGNAL mux_1666_nl : STD_LOGIC;
  SIGNAL nor_1775_nl : STD_LOGIC;
  SIGNAL nand_363_nl : STD_LOGIC;
  SIGNAL nand_100_nl : STD_LOGIC;
  SIGNAL mux_1665_nl : STD_LOGIC;
  SIGNAL and_2128_nl : STD_LOGIC;
  SIGNAL or_2003_nl : STD_LOGIC;
  SIGNAL mux_1714_nl : STD_LOGIC;
  SIGNAL mux_1713_nl : STD_LOGIC;
  SIGNAL mux_1710_nl : STD_LOGIC;
  SIGNAL or_2045_nl : STD_LOGIC;
  SIGNAL mux_1731_nl : STD_LOGIC;
  SIGNAL mux_1730_nl : STD_LOGIC;
  SIGNAL mux_1729_nl : STD_LOGIC;
  SIGNAL and_1733_nl : STD_LOGIC;
  SIGNAL mux_1728_nl : STD_LOGIC;
  SIGNAL nor_1756_nl : STD_LOGIC;
  SIGNAL nor_1757_nl : STD_LOGIC;
  SIGNAL nor_1759_nl : STD_LOGIC;
  SIGNAL mux_1727_nl : STD_LOGIC;
  SIGNAL nor_1761_nl : STD_LOGIC;
  SIGNAL mux_1726_nl : STD_LOGIC;
  SIGNAL mux_1725_nl : STD_LOGIC;
  SIGNAL mux_1724_nl : STD_LOGIC;
  SIGNAL nand_349_nl : STD_LOGIC;
  SIGNAL and_1734_nl : STD_LOGIC;
  SIGNAL nor_1764_nl : STD_LOGIC;
  SIGNAL mux_1723_nl : STD_LOGIC;
  SIGNAL or_2064_nl : STD_LOGIC;
  SIGNAL mux_1722_nl : STD_LOGIC;
  SIGNAL or_2063_nl : STD_LOGIC;
  SIGNAL or_2059_nl : STD_LOGIC;
  SIGNAL mux_1720_nl : STD_LOGIC;
  SIGNAL nand_104_nl : STD_LOGIC;
  SIGNAL mux_1719_nl : STD_LOGIC;
  SIGNAL and_529_nl : STD_LOGIC;
  SIGNAL mux_1718_nl : STD_LOGIC;
  SIGNAL and_1735_nl : STD_LOGIC;
  SIGNAL mux_1780_nl : STD_LOGIC;
  SIGNAL mux_1779_nl : STD_LOGIC;
  SIGNAL mux_1778_nl : STD_LOGIC;
  SIGNAL and_1707_nl : STD_LOGIC;
  SIGNAL mux_1777_nl : STD_LOGIC;
  SIGNAL and_1708_nl : STD_LOGIC;
  SIGNAL nor_1745_nl : STD_LOGIC;
  SIGNAL and_1709_nl : STD_LOGIC;
  SIGNAL mux_1776_nl : STD_LOGIC;
  SIGNAL and_1710_nl : STD_LOGIC;
  SIGNAL nor_1747_nl : STD_LOGIC;
  SIGNAL mux_1775_nl : STD_LOGIC;
  SIGNAL nor_1749_nl : STD_LOGIC;
  SIGNAL mux_1774_nl : STD_LOGIC;
  SIGNAL or_4557_nl : STD_LOGIC;
  SIGNAL mux_1773_nl : STD_LOGIC;
  SIGNAL nand_338_nl : STD_LOGIC;
  SIGNAL nor_1751_nl : STD_LOGIC;
  SIGNAL mux_1772_nl : STD_LOGIC;
  SIGNAL or_2108_nl : STD_LOGIC;
  SIGNAL or_2106_nl : STD_LOGIC;
  SIGNAL mux_1771_nl : STD_LOGIC;
  SIGNAL nand_339_nl : STD_LOGIC;
  SIGNAL mux_1769_nl : STD_LOGIC;
  SIGNAL or_2104_nl : STD_LOGIC;
  SIGNAL or_2103_nl : STD_LOGIC;
  SIGNAL mux_1842_nl : STD_LOGIC;
  SIGNAL mux_1841_nl : STD_LOGIC;
  SIGNAL mux_1840_nl : STD_LOGIC;
  SIGNAL or_2160_nl : STD_LOGIC;
  SIGNAL mux_1839_nl : STD_LOGIC;
  SIGNAL mux_1838_nl : STD_LOGIC;
  SIGNAL or_2159_nl : STD_LOGIC;
  SIGNAL or_2156_nl : STD_LOGIC;
  SIGNAL mux_1837_nl : STD_LOGIC;
  SIGNAL mux_1836_nl : STD_LOGIC;
  SIGNAL or_2155_nl : STD_LOGIC;
  SIGNAL or_2154_nl : STD_LOGIC;
  SIGNAL mux_1835_nl : STD_LOGIC;
  SIGNAL mux_1834_nl : STD_LOGIC;
  SIGNAL mux_1833_nl : STD_LOGIC;
  SIGNAL or_2151_nl : STD_LOGIC;
  SIGNAL mux_1831_nl : STD_LOGIC;
  SIGNAL or_2150_nl : STD_LOGIC;
  SIGNAL mux_1830_nl : STD_LOGIC;
  SIGNAL mux_1829_nl : STD_LOGIC;
  SIGNAL mux_1828_nl : STD_LOGIC;
  SIGNAL mux_1827_nl : STD_LOGIC;
  SIGNAL mux_1826_nl : STD_LOGIC;
  SIGNAL mux_1825_nl : STD_LOGIC;
  SIGNAL mux_1824_nl : STD_LOGIC;
  SIGNAL or_2146_nl : STD_LOGIC;
  SIGNAL or_2144_nl : STD_LOGIC;
  SIGNAL mux_1823_nl : STD_LOGIC;
  SIGNAL mux_1822_nl : STD_LOGIC;
  SIGNAL or_2137_nl : STD_LOGIC;
  SIGNAL mux_1876_nl : STD_LOGIC;
  SIGNAL and_1675_nl : STD_LOGIC;
  SIGNAL and_1677_nl : STD_LOGIC;
  SIGNAL mux_1867_nl : STD_LOGIC;
  SIGNAL and_1678_nl : STD_LOGIC;
  SIGNAL mux_1879_nl : STD_LOGIC;
  SIGNAL mux_1878_nl : STD_LOGIC;
  SIGNAL and_1676_nl : STD_LOGIC;
  SIGNAL mux_1875_nl : STD_LOGIC;
  SIGNAL mux_1874_nl : STD_LOGIC;
  SIGNAL mux_1873_nl : STD_LOGIC;
  SIGNAL or_2188_nl : STD_LOGIC;
  SIGNAL mux_1871_nl : STD_LOGIC;
  SIGNAL mux_1870_nl : STD_LOGIC;
  SIGNAL mux_1869_nl : STD_LOGIC;
  SIGNAL mux_1901_nl : STD_LOGIC;
  SIGNAL mux_1900_nl : STD_LOGIC;
  SIGNAL mux_1899_nl : STD_LOGIC;
  SIGNAL or_2217_nl : STD_LOGIC;
  SIGNAL mux_1898_nl : STD_LOGIC;
  SIGNAL mux_1897_nl : STD_LOGIC;
  SIGNAL mux_1896_nl : STD_LOGIC;
  SIGNAL nor_1727_nl : STD_LOGIC;
  SIGNAL nand_114_nl : STD_LOGIC;
  SIGNAL mux_1895_nl : STD_LOGIC;
  SIGNAL mux_1894_nl : STD_LOGIC;
  SIGNAL mux_1893_nl : STD_LOGIC;
  SIGNAL mux_1892_nl : STD_LOGIC;
  SIGNAL or_2213_nl : STD_LOGIC;
  SIGNAL nand_113_nl : STD_LOGIC;
  SIGNAL mux_1891_nl : STD_LOGIC;
  SIGNAL mux_1890_nl : STD_LOGIC;
  SIGNAL mux_1889_nl : STD_LOGIC;
  SIGNAL or_2211_nl : STD_LOGIC;
  SIGNAL mux_1888_nl : STD_LOGIC;
  SIGNAL nor_640_nl : STD_LOGIC;
  SIGNAL mux_1882_nl : STD_LOGIC;
  SIGNAL nand_111_nl : STD_LOGIC;
  SIGNAL mux_1881_nl : STD_LOGIC;
  SIGNAL nor_1728_nl : STD_LOGIC;
  SIGNAL nor_1729_nl : STD_LOGIC;
  SIGNAL mux_1926_nl : STD_LOGIC;
  SIGNAL mux_1925_nl : STD_LOGIC;
  SIGNAL or_2244_nl : STD_LOGIC;
  SIGNAL mux_1923_nl : STD_LOGIC;
  SIGNAL mux_1922_nl : STD_LOGIC;
  SIGNAL mux_1921_nl : STD_LOGIC;
  SIGNAL mux_1931_nl : STD_LOGIC;
  SIGNAL mux_1930_nl : STD_LOGIC;
  SIGNAL and_1670_nl : STD_LOGIC;
  SIGNAL mux_1949_nl : STD_LOGIC;
  SIGNAL mux_1948_nl : STD_LOGIC;
  SIGNAL mux_1947_nl : STD_LOGIC;
  SIGNAL mux_1946_nl : STD_LOGIC;
  SIGNAL mux_1945_nl : STD_LOGIC;
  SIGNAL mux_1944_nl : STD_LOGIC;
  SIGNAL or_2274_nl : STD_LOGIC;
  SIGNAL or_2270_nl : STD_LOGIC;
  SIGNAL mux_1943_nl : STD_LOGIC;
  SIGNAL mux_1942_nl : STD_LOGIC;
  SIGNAL mux_1941_nl : STD_LOGIC;
  SIGNAL or_2268_nl : STD_LOGIC;
  SIGNAL or_2267_nl : STD_LOGIC;
  SIGNAL mux_1940_nl : STD_LOGIC;
  SIGNAL mux_1939_nl : STD_LOGIC;
  SIGNAL or_2265_nl : STD_LOGIC;
  SIGNAL or_2263_nl : STD_LOGIC;
  SIGNAL mux_1933_nl : STD_LOGIC;
  SIGNAL or_2254_nl : STD_LOGIC;
  SIGNAL mux_1989_nl : STD_LOGIC;
  SIGNAL mux_1988_nl : STD_LOGIC;
  SIGNAL and_1659_nl : STD_LOGIC;
  SIGNAL mux_2009_nl : STD_LOGIC;
  SIGNAL mux_2008_nl : STD_LOGIC;
  SIGNAL mux_2007_nl : STD_LOGIC;
  SIGNAL or_2317_nl : STD_LOGIC;
  SIGNAL mux_2006_nl : STD_LOGIC;
  SIGNAL mux_2005_nl : STD_LOGIC;
  SIGNAL mux_2004_nl : STD_LOGIC;
  SIGNAL nor_1703_nl : STD_LOGIC;
  SIGNAL nand_119_nl : STD_LOGIC;
  SIGNAL mux_2003_nl : STD_LOGIC;
  SIGNAL mux_2002_nl : STD_LOGIC;
  SIGNAL mux_2001_nl : STD_LOGIC;
  SIGNAL or_2313_nl : STD_LOGIC;
  SIGNAL nand_118_nl : STD_LOGIC;
  SIGNAL mux_2000_nl : STD_LOGIC;
  SIGNAL or_2311_nl : STD_LOGIC;
  SIGNAL mux_1998_nl : STD_LOGIC;
  SIGNAL mux_1997_nl : STD_LOGIC;
  SIGNAL nor_664_nl : STD_LOGIC;
  SIGNAL mux_1992_nl : STD_LOGIC;
  SIGNAL or_4537_nl : STD_LOGIC;
  SIGNAL mux_1991_nl : STD_LOGIC;
  SIGNAL or_2303_nl : STD_LOGIC;
  SIGNAL mux_2050_nl : STD_LOGIC;
  SIGNAL mux_2049_nl : STD_LOGIC;
  SIGNAL and_1646_nl : STD_LOGIC;
  SIGNAL mux_2074_nl : STD_LOGIC;
  SIGNAL mux_2073_nl : STD_LOGIC;
  SIGNAL mux_2072_nl : STD_LOGIC;
  SIGNAL or_2368_nl : STD_LOGIC;
  SIGNAL mux_2071_nl : STD_LOGIC;
  SIGNAL mux_2070_nl : STD_LOGIC;
  SIGNAL or_2367_nl : STD_LOGIC;
  SIGNAL or_2364_nl : STD_LOGIC;
  SIGNAL mux_2069_nl : STD_LOGIC;
  SIGNAL mux_2068_nl : STD_LOGIC;
  SIGNAL or_2363_nl : STD_LOGIC;
  SIGNAL or_2362_nl : STD_LOGIC;
  SIGNAL mux_2067_nl : STD_LOGIC;
  SIGNAL mux_2066_nl : STD_LOGIC;
  SIGNAL mux_2065_nl : STD_LOGIC;
  SIGNAL or_2359_nl : STD_LOGIC;
  SIGNAL mux_2063_nl : STD_LOGIC;
  SIGNAL or_2358_nl : STD_LOGIC;
  SIGNAL mux_2062_nl : STD_LOGIC;
  SIGNAL mux_2061_nl : STD_LOGIC;
  SIGNAL or_2355_nl : STD_LOGIC;
  SIGNAL mux_2060_nl : STD_LOGIC;
  SIGNAL mux_2059_nl : STD_LOGIC;
  SIGNAL mux_2058_nl : STD_LOGIC;
  SIGNAL mux_2057_nl : STD_LOGIC;
  SIGNAL mux_2056_nl : STD_LOGIC;
  SIGNAL mux_2055_nl : STD_LOGIC;
  SIGNAL mux_2054_nl : STD_LOGIC;
  SIGNAL or_2352_nl : STD_LOGIC;
  SIGNAL or_2346_nl : STD_LOGIC;
  SIGNAL mux_2107_nl : STD_LOGIC;
  SIGNAL mux_2106_nl : STD_LOGIC;
  SIGNAL and_1636_nl : STD_LOGIC;
  SIGNAL mux_2103_nl : STD_LOGIC;
  SIGNAL mux_2102_nl : STD_LOGIC;
  SIGNAL mux_2101_nl : STD_LOGIC;
  SIGNAL or_2385_nl : STD_LOGIC;
  SIGNAL mux_2099_nl : STD_LOGIC;
  SIGNAL mux_2098_nl : STD_LOGIC;
  SIGNAL mux_2097_nl : STD_LOGIC;
  SIGNAL mux_2129_nl : STD_LOGIC;
  SIGNAL mux_2128_nl : STD_LOGIC;
  SIGNAL mux_2127_nl : STD_LOGIC;
  SIGNAL or_2422_nl : STD_LOGIC;
  SIGNAL mux_2126_nl : STD_LOGIC;
  SIGNAL mux_2125_nl : STD_LOGIC;
  SIGNAL mux_2124_nl : STD_LOGIC;
  SIGNAL nor_1683_nl : STD_LOGIC;
  SIGNAL nand_123_nl : STD_LOGIC;
  SIGNAL mux_2123_nl : STD_LOGIC;
  SIGNAL mux_2122_nl : STD_LOGIC;
  SIGNAL mux_2121_nl : STD_LOGIC;
  SIGNAL mux_2120_nl : STD_LOGIC;
  SIGNAL or_2418_nl : STD_LOGIC;
  SIGNAL nand_122_nl : STD_LOGIC;
  SIGNAL mux_2119_nl : STD_LOGIC;
  SIGNAL mux_2118_nl : STD_LOGIC;
  SIGNAL mux_2117_nl : STD_LOGIC;
  SIGNAL or_2415_nl : STD_LOGIC;
  SIGNAL mux_2116_nl : STD_LOGIC;
  SIGNAL nor_697_nl : STD_LOGIC;
  SIGNAL mux_2110_nl : STD_LOGIC;
  SIGNAL nand_120_nl : STD_LOGIC;
  SIGNAL mux_2109_nl : STD_LOGIC;
  SIGNAL nor_1684_nl : STD_LOGIC;
  SIGNAL nor_1685_nl : STD_LOGIC;
  SIGNAL mux_2151_nl : STD_LOGIC;
  SIGNAL mux_2150_nl : STD_LOGIC;
  SIGNAL or_2439_nl : STD_LOGIC;
  SIGNAL mux_2148_nl : STD_LOGIC;
  SIGNAL mux_2147_nl : STD_LOGIC;
  SIGNAL mux_2146_nl : STD_LOGIC;
  SIGNAL mux_2156_nl : STD_LOGIC;
  SIGNAL mux_2155_nl : STD_LOGIC;
  SIGNAL and_1630_nl : STD_LOGIC;
  SIGNAL mux_2174_nl : STD_LOGIC;
  SIGNAL mux_2173_nl : STD_LOGIC;
  SIGNAL mux_2172_nl : STD_LOGIC;
  SIGNAL mux_2171_nl : STD_LOGIC;
  SIGNAL mux_2170_nl : STD_LOGIC;
  SIGNAL mux_2169_nl : STD_LOGIC;
  SIGNAL or_2475_nl : STD_LOGIC;
  SIGNAL or_2471_nl : STD_LOGIC;
  SIGNAL mux_2168_nl : STD_LOGIC;
  SIGNAL mux_2167_nl : STD_LOGIC;
  SIGNAL mux_2166_nl : STD_LOGIC;
  SIGNAL or_2469_nl : STD_LOGIC;
  SIGNAL or_2468_nl : STD_LOGIC;
  SIGNAL mux_2165_nl : STD_LOGIC;
  SIGNAL mux_2164_nl : STD_LOGIC;
  SIGNAL or_2465_nl : STD_LOGIC;
  SIGNAL or_2463_nl : STD_LOGIC;
  SIGNAL mux_2158_nl : STD_LOGIC;
  SIGNAL or_2450_nl : STD_LOGIC;
  SIGNAL mux_2212_nl : STD_LOGIC;
  SIGNAL mux_2211_nl : STD_LOGIC;
  SIGNAL and_1619_nl : STD_LOGIC;
  SIGNAL mux_2232_nl : STD_LOGIC;
  SIGNAL mux_2231_nl : STD_LOGIC;
  SIGNAL mux_2230_nl : STD_LOGIC;
  SIGNAL or_2516_nl : STD_LOGIC;
  SIGNAL mux_2229_nl : STD_LOGIC;
  SIGNAL mux_2228_nl : STD_LOGIC;
  SIGNAL mux_2227_nl : STD_LOGIC;
  SIGNAL nor_1665_nl : STD_LOGIC;
  SIGNAL nand_128_nl : STD_LOGIC;
  SIGNAL mux_2226_nl : STD_LOGIC;
  SIGNAL mux_2225_nl : STD_LOGIC;
  SIGNAL mux_2224_nl : STD_LOGIC;
  SIGNAL or_2512_nl : STD_LOGIC;
  SIGNAL nand_127_nl : STD_LOGIC;
  SIGNAL mux_2223_nl : STD_LOGIC;
  SIGNAL or_2509_nl : STD_LOGIC;
  SIGNAL mux_2221_nl : STD_LOGIC;
  SIGNAL mux_2220_nl : STD_LOGIC;
  SIGNAL nor_724_nl : STD_LOGIC;
  SIGNAL mux_2215_nl : STD_LOGIC;
  SIGNAL or_4516_nl : STD_LOGIC;
  SIGNAL mux_2214_nl : STD_LOGIC;
  SIGNAL or_2497_nl : STD_LOGIC;
  SIGNAL mux_2270_nl : STD_LOGIC;
  SIGNAL mux_2269_nl : STD_LOGIC;
  SIGNAL and_1605_nl : STD_LOGIC;
  SIGNAL mux_2294_nl : STD_LOGIC;
  SIGNAL mux_2293_nl : STD_LOGIC;
  SIGNAL mux_2292_nl : STD_LOGIC;
  SIGNAL or_2558_nl : STD_LOGIC;
  SIGNAL mux_2291_nl : STD_LOGIC;
  SIGNAL mux_2290_nl : STD_LOGIC;
  SIGNAL or_2557_nl : STD_LOGIC;
  SIGNAL or_2554_nl : STD_LOGIC;
  SIGNAL mux_2289_nl : STD_LOGIC;
  SIGNAL mux_2288_nl : STD_LOGIC;
  SIGNAL or_2553_nl : STD_LOGIC;
  SIGNAL or_2552_nl : STD_LOGIC;
  SIGNAL mux_2287_nl : STD_LOGIC;
  SIGNAL mux_2286_nl : STD_LOGIC;
  SIGNAL mux_2285_nl : STD_LOGIC;
  SIGNAL or_2549_nl : STD_LOGIC;
  SIGNAL mux_2283_nl : STD_LOGIC;
  SIGNAL or_2548_nl : STD_LOGIC;
  SIGNAL mux_2282_nl : STD_LOGIC;
  SIGNAL mux_2281_nl : STD_LOGIC;
  SIGNAL mux_2280_nl : STD_LOGIC;
  SIGNAL mux_2279_nl : STD_LOGIC;
  SIGNAL mux_2278_nl : STD_LOGIC;
  SIGNAL mux_2277_nl : STD_LOGIC;
  SIGNAL mux_2276_nl : STD_LOGIC;
  SIGNAL or_2544_nl : STD_LOGIC;
  SIGNAL or_2542_nl : STD_LOGIC;
  SIGNAL mux_2275_nl : STD_LOGIC;
  SIGNAL mux_2274_nl : STD_LOGIC;
  SIGNAL or_2535_nl : STD_LOGIC;
  SIGNAL mux_2327_nl : STD_LOGIC;
  SIGNAL mux_2326_nl : STD_LOGIC;
  SIGNAL and_1595_nl : STD_LOGIC;
  SIGNAL mux_2323_nl : STD_LOGIC;
  SIGNAL mux_2322_nl : STD_LOGIC;
  SIGNAL mux_2321_nl : STD_LOGIC;
  SIGNAL or_2576_nl : STD_LOGIC;
  SIGNAL mux_2319_nl : STD_LOGIC;
  SIGNAL mux_2318_nl : STD_LOGIC;
  SIGNAL mux_2317_nl : STD_LOGIC;
  SIGNAL mux_2349_nl : STD_LOGIC;
  SIGNAL mux_2348_nl : STD_LOGIC;
  SIGNAL mux_2347_nl : STD_LOGIC;
  SIGNAL or_2603_nl : STD_LOGIC;
  SIGNAL mux_2346_nl : STD_LOGIC;
  SIGNAL mux_2345_nl : STD_LOGIC;
  SIGNAL mux_2344_nl : STD_LOGIC;
  SIGNAL nor_1650_nl : STD_LOGIC;
  SIGNAL nand_132_nl : STD_LOGIC;
  SIGNAL mux_2343_nl : STD_LOGIC;
  SIGNAL mux_2342_nl : STD_LOGIC;
  SIGNAL mux_2341_nl : STD_LOGIC;
  SIGNAL mux_2340_nl : STD_LOGIC;
  SIGNAL or_2599_nl : STD_LOGIC;
  SIGNAL nand_131_nl : STD_LOGIC;
  SIGNAL mux_2339_nl : STD_LOGIC;
  SIGNAL mux_2338_nl : STD_LOGIC;
  SIGNAL mux_2337_nl : STD_LOGIC;
  SIGNAL or_2597_nl : STD_LOGIC;
  SIGNAL mux_2336_nl : STD_LOGIC;
  SIGNAL nor_756_nl : STD_LOGIC;
  SIGNAL mux_2330_nl : STD_LOGIC;
  SIGNAL nand_129_nl : STD_LOGIC;
  SIGNAL mux_2329_nl : STD_LOGIC;
  SIGNAL nor_1651_nl : STD_LOGIC;
  SIGNAL nor_1652_nl : STD_LOGIC;
  SIGNAL mux_2371_nl : STD_LOGIC;
  SIGNAL mux_2370_nl : STD_LOGIC;
  SIGNAL or_2621_nl : STD_LOGIC;
  SIGNAL mux_2368_nl : STD_LOGIC;
  SIGNAL mux_2367_nl : STD_LOGIC;
  SIGNAL mux_2366_nl : STD_LOGIC;
  SIGNAL mux_2376_nl : STD_LOGIC;
  SIGNAL mux_2375_nl : STD_LOGIC;
  SIGNAL and_1589_nl : STD_LOGIC;
  SIGNAL mux_2394_nl : STD_LOGIC;
  SIGNAL mux_2393_nl : STD_LOGIC;
  SIGNAL mux_2392_nl : STD_LOGIC;
  SIGNAL mux_2391_nl : STD_LOGIC;
  SIGNAL mux_2390_nl : STD_LOGIC;
  SIGNAL mux_2389_nl : STD_LOGIC;
  SIGNAL or_2650_nl : STD_LOGIC;
  SIGNAL or_2646_nl : STD_LOGIC;
  SIGNAL mux_2388_nl : STD_LOGIC;
  SIGNAL mux_2387_nl : STD_LOGIC;
  SIGNAL mux_2386_nl : STD_LOGIC;
  SIGNAL or_2644_nl : STD_LOGIC;
  SIGNAL or_2643_nl : STD_LOGIC;
  SIGNAL mux_2385_nl : STD_LOGIC;
  SIGNAL mux_2384_nl : STD_LOGIC;
  SIGNAL or_2641_nl : STD_LOGIC;
  SIGNAL or_2639_nl : STD_LOGIC;
  SIGNAL mux_2378_nl : STD_LOGIC;
  SIGNAL or_2630_nl : STD_LOGIC;
  SIGNAL mux_2432_nl : STD_LOGIC;
  SIGNAL mux_2431_nl : STD_LOGIC;
  SIGNAL and_1578_nl : STD_LOGIC;
  SIGNAL mux_2452_nl : STD_LOGIC;
  SIGNAL mux_2451_nl : STD_LOGIC;
  SIGNAL mux_2450_nl : STD_LOGIC;
  SIGNAL or_2686_nl : STD_LOGIC;
  SIGNAL mux_2449_nl : STD_LOGIC;
  SIGNAL mux_2448_nl : STD_LOGIC;
  SIGNAL mux_2447_nl : STD_LOGIC;
  SIGNAL nor_1632_nl : STD_LOGIC;
  SIGNAL nand_137_nl : STD_LOGIC;
  SIGNAL mux_2446_nl : STD_LOGIC;
  SIGNAL mux_2445_nl : STD_LOGIC;
  SIGNAL mux_2444_nl : STD_LOGIC;
  SIGNAL or_2682_nl : STD_LOGIC;
  SIGNAL nand_136_nl : STD_LOGIC;
  SIGNAL mux_2443_nl : STD_LOGIC;
  SIGNAL or_2680_nl : STD_LOGIC;
  SIGNAL mux_2441_nl : STD_LOGIC;
  SIGNAL mux_2440_nl : STD_LOGIC;
  SIGNAL nor_780_nl : STD_LOGIC;
  SIGNAL mux_2435_nl : STD_LOGIC;
  SIGNAL or_4495_nl : STD_LOGIC;
  SIGNAL mux_2434_nl : STD_LOGIC;
  SIGNAL or_2672_nl : STD_LOGIC;
  SIGNAL mux_2490_nl : STD_LOGIC;
  SIGNAL mux_2489_nl : STD_LOGIC;
  SIGNAL and_1564_nl : STD_LOGIC;
  SIGNAL mux_2514_nl : STD_LOGIC;
  SIGNAL mux_2513_nl : STD_LOGIC;
  SIGNAL mux_2512_nl : STD_LOGIC;
  SIGNAL or_2729_nl : STD_LOGIC;
  SIGNAL mux_2511_nl : STD_LOGIC;
  SIGNAL mux_2510_nl : STD_LOGIC;
  SIGNAL or_2728_nl : STD_LOGIC;
  SIGNAL or_2725_nl : STD_LOGIC;
  SIGNAL mux_2509_nl : STD_LOGIC;
  SIGNAL mux_2508_nl : STD_LOGIC;
  SIGNAL or_2724_nl : STD_LOGIC;
  SIGNAL or_2723_nl : STD_LOGIC;
  SIGNAL mux_2507_nl : STD_LOGIC;
  SIGNAL mux_2506_nl : STD_LOGIC;
  SIGNAL mux_2505_nl : STD_LOGIC;
  SIGNAL or_2720_nl : STD_LOGIC;
  SIGNAL mux_2503_nl : STD_LOGIC;
  SIGNAL or_2719_nl : STD_LOGIC;
  SIGNAL mux_2502_nl : STD_LOGIC;
  SIGNAL mux_2501_nl : STD_LOGIC;
  SIGNAL or_2716_nl : STD_LOGIC;
  SIGNAL mux_2500_nl : STD_LOGIC;
  SIGNAL mux_2499_nl : STD_LOGIC;
  SIGNAL mux_2498_nl : STD_LOGIC;
  SIGNAL mux_2497_nl : STD_LOGIC;
  SIGNAL mux_2496_nl : STD_LOGIC;
  SIGNAL mux_2495_nl : STD_LOGIC;
  SIGNAL mux_2494_nl : STD_LOGIC;
  SIGNAL or_2713_nl : STD_LOGIC;
  SIGNAL or_2707_nl : STD_LOGIC;
  SIGNAL mux_2547_nl : STD_LOGIC;
  SIGNAL mux_2546_nl : STD_LOGIC;
  SIGNAL and_1554_nl : STD_LOGIC;
  SIGNAL mux_2543_nl : STD_LOGIC;
  SIGNAL mux_2542_nl : STD_LOGIC;
  SIGNAL mux_2541_nl : STD_LOGIC;
  SIGNAL or_2746_nl : STD_LOGIC;
  SIGNAL mux_2539_nl : STD_LOGIC;
  SIGNAL mux_2538_nl : STD_LOGIC;
  SIGNAL mux_2537_nl : STD_LOGIC;
  SIGNAL mux_2569_nl : STD_LOGIC;
  SIGNAL mux_2568_nl : STD_LOGIC;
  SIGNAL mux_2567_nl : STD_LOGIC;
  SIGNAL or_2782_nl : STD_LOGIC;
  SIGNAL mux_2566_nl : STD_LOGIC;
  SIGNAL mux_2565_nl : STD_LOGIC;
  SIGNAL mux_2564_nl : STD_LOGIC;
  SIGNAL nor_1617_nl : STD_LOGIC;
  SIGNAL nand_141_nl : STD_LOGIC;
  SIGNAL mux_2563_nl : STD_LOGIC;
  SIGNAL mux_2562_nl : STD_LOGIC;
  SIGNAL mux_2561_nl : STD_LOGIC;
  SIGNAL mux_2560_nl : STD_LOGIC;
  SIGNAL or_2778_nl : STD_LOGIC;
  SIGNAL nand_140_nl : STD_LOGIC;
  SIGNAL mux_2559_nl : STD_LOGIC;
  SIGNAL mux_2558_nl : STD_LOGIC;
  SIGNAL mux_2557_nl : STD_LOGIC;
  SIGNAL or_2775_nl : STD_LOGIC;
  SIGNAL mux_2556_nl : STD_LOGIC;
  SIGNAL nor_813_nl : STD_LOGIC;
  SIGNAL mux_2550_nl : STD_LOGIC;
  SIGNAL nand_138_nl : STD_LOGIC;
  SIGNAL mux_2549_nl : STD_LOGIC;
  SIGNAL nor_1618_nl : STD_LOGIC;
  SIGNAL nor_1619_nl : STD_LOGIC;
  SIGNAL mux_2591_nl : STD_LOGIC;
  SIGNAL mux_2590_nl : STD_LOGIC;
  SIGNAL or_2799_nl : STD_LOGIC;
  SIGNAL mux_2588_nl : STD_LOGIC;
  SIGNAL mux_2587_nl : STD_LOGIC;
  SIGNAL mux_2586_nl : STD_LOGIC;
  SIGNAL mux_2596_nl : STD_LOGIC;
  SIGNAL mux_2595_nl : STD_LOGIC;
  SIGNAL and_1547_nl : STD_LOGIC;
  SIGNAL mux_2614_nl : STD_LOGIC;
  SIGNAL mux_2613_nl : STD_LOGIC;
  SIGNAL mux_2612_nl : STD_LOGIC;
  SIGNAL mux_2611_nl : STD_LOGIC;
  SIGNAL mux_2610_nl : STD_LOGIC;
  SIGNAL mux_2609_nl : STD_LOGIC;
  SIGNAL or_2835_nl : STD_LOGIC;
  SIGNAL or_2831_nl : STD_LOGIC;
  SIGNAL mux_2608_nl : STD_LOGIC;
  SIGNAL mux_2607_nl : STD_LOGIC;
  SIGNAL mux_2606_nl : STD_LOGIC;
  SIGNAL or_2829_nl : STD_LOGIC;
  SIGNAL or_2828_nl : STD_LOGIC;
  SIGNAL mux_2605_nl : STD_LOGIC;
  SIGNAL mux_2604_nl : STD_LOGIC;
  SIGNAL or_2825_nl : STD_LOGIC;
  SIGNAL or_2823_nl : STD_LOGIC;
  SIGNAL mux_2598_nl : STD_LOGIC;
  SIGNAL or_2810_nl : STD_LOGIC;
  SIGNAL mux_2652_nl : STD_LOGIC;
  SIGNAL mux_2651_nl : STD_LOGIC;
  SIGNAL and_1534_nl : STD_LOGIC;
  SIGNAL mux_2672_nl : STD_LOGIC;
  SIGNAL mux_2671_nl : STD_LOGIC;
  SIGNAL mux_2670_nl : STD_LOGIC;
  SIGNAL or_2876_nl : STD_LOGIC;
  SIGNAL mux_2669_nl : STD_LOGIC;
  SIGNAL mux_2668_nl : STD_LOGIC;
  SIGNAL mux_2667_nl : STD_LOGIC;
  SIGNAL and_1531_nl : STD_LOGIC;
  SIGNAL nand_146_nl : STD_LOGIC;
  SIGNAL mux_2666_nl : STD_LOGIC;
  SIGNAL mux_2665_nl : STD_LOGIC;
  SIGNAL mux_2664_nl : STD_LOGIC;
  SIGNAL or_2872_nl : STD_LOGIC;
  SIGNAL nand_145_nl : STD_LOGIC;
  SIGNAL mux_2663_nl : STD_LOGIC;
  SIGNAL or_2869_nl : STD_LOGIC;
  SIGNAL mux_2661_nl : STD_LOGIC;
  SIGNAL mux_2660_nl : STD_LOGIC;
  SIGNAL mux_2655_nl : STD_LOGIC;
  SIGNAL or_4474_nl : STD_LOGIC;
  SIGNAL mux_2654_nl : STD_LOGIC;
  SIGNAL or_2857_nl : STD_LOGIC;
  SIGNAL mux_2710_nl : STD_LOGIC;
  SIGNAL mux_2709_nl : STD_LOGIC;
  SIGNAL and_1518_nl : STD_LOGIC;
  SIGNAL mux_2734_nl : STD_LOGIC;
  SIGNAL mux_2733_nl : STD_LOGIC;
  SIGNAL or_2930_nl : STD_LOGIC;
  SIGNAL or_2928_nl : STD_LOGIC;
  SIGNAL mux_2732_nl : STD_LOGIC;
  SIGNAL mux_2731_nl : STD_LOGIC;
  SIGNAL mux_2730_nl : STD_LOGIC;
  SIGNAL or_2927_nl : STD_LOGIC;
  SIGNAL mux_2729_nl : STD_LOGIC;
  SIGNAL or_2926_nl : STD_LOGIC;
  SIGNAL mux_2728_nl : STD_LOGIC;
  SIGNAL mux_2727_nl : STD_LOGIC;
  SIGNAL or_2923_nl : STD_LOGIC;
  SIGNAL mux_2726_nl : STD_LOGIC;
  SIGNAL mux_2725_nl : STD_LOGIC;
  SIGNAL or_2922_nl : STD_LOGIC;
  SIGNAL or_2918_nl : STD_LOGIC;
  SIGNAL mux_2724_nl : STD_LOGIC;
  SIGNAL mux_2722_nl : STD_LOGIC;
  SIGNAL mux_2721_nl : STD_LOGIC;
  SIGNAL mux_2720_nl : STD_LOGIC;
  SIGNAL mux_2719_nl : STD_LOGIC;
  SIGNAL mux_2718_nl : STD_LOGIC;
  SIGNAL mux_2717_nl : STD_LOGIC;
  SIGNAL mux_2716_nl : STD_LOGIC;
  SIGNAL or_2911_nl : STD_LOGIC;
  SIGNAL or_2908_nl : STD_LOGIC;
  SIGNAL mux_2715_nl : STD_LOGIC;
  SIGNAL mux_2714_nl : STD_LOGIC;
  SIGNAL or_2896_nl : STD_LOGIC;
  SIGNAL mux_2767_nl : STD_LOGIC;
  SIGNAL mux_2766_nl : STD_LOGIC;
  SIGNAL and_1507_nl : STD_LOGIC;
  SIGNAL mux_2763_nl : STD_LOGIC;
  SIGNAL mux_2762_nl : STD_LOGIC;
  SIGNAL mux_2761_nl : STD_LOGIC;
  SIGNAL or_2949_nl : STD_LOGIC;
  SIGNAL mux_2759_nl : STD_LOGIC;
  SIGNAL mux_2758_nl : STD_LOGIC;
  SIGNAL mux_2757_nl : STD_LOGIC;
  SIGNAL mux_2789_nl : STD_LOGIC;
  SIGNAL mux_2788_nl : STD_LOGIC;
  SIGNAL mux_2787_nl : STD_LOGIC;
  SIGNAL or_2980_nl : STD_LOGIC;
  SIGNAL nand_150_nl : STD_LOGIC;
  SIGNAL mux_2786_nl : STD_LOGIC;
  SIGNAL mux_2785_nl : STD_LOGIC;
  SIGNAL mux_2784_nl : STD_LOGIC;
  SIGNAL or_2978_nl : STD_LOGIC;
  SIGNAL mux_2783_nl : STD_LOGIC;
  SIGNAL nor_878_nl : STD_LOGIC;
  SIGNAL mux_2782_nl : STD_LOGIC;
  SIGNAL mux_2781_nl : STD_LOGIC;
  SIGNAL or_2976_nl : STD_LOGIC;
  SIGNAL mux_2780_nl : STD_LOGIC;
  SIGNAL mux_2779_nl : STD_LOGIC;
  SIGNAL mux_2778_nl : STD_LOGIC;
  SIGNAL nor_1587_nl : STD_LOGIC;
  SIGNAL nand_149_nl : STD_LOGIC;
  SIGNAL mux_2777_nl : STD_LOGIC;
  SIGNAL mux_2776_nl : STD_LOGIC;
  SIGNAL mux_2770_nl : STD_LOGIC;
  SIGNAL nand_147_nl : STD_LOGIC;
  SIGNAL mux_2769_nl : STD_LOGIC;
  SIGNAL nor_1588_nl : STD_LOGIC;
  SIGNAL nor_1589_nl : STD_LOGIC;
  SIGNAL mux_2811_nl : STD_LOGIC;
  SIGNAL mux_2810_nl : STD_LOGIC;
  SIGNAL or_3001_nl : STD_LOGIC;
  SIGNAL mux_2808_nl : STD_LOGIC;
  SIGNAL mux_2807_nl : STD_LOGIC;
  SIGNAL mux_2806_nl : STD_LOGIC;
  SIGNAL mux_2816_nl : STD_LOGIC;
  SIGNAL mux_2815_nl : STD_LOGIC;
  SIGNAL and_1501_nl : STD_LOGIC;
  SIGNAL mux_2834_nl : STD_LOGIC;
  SIGNAL mux_2833_nl : STD_LOGIC;
  SIGNAL mux_2832_nl : STD_LOGIC;
  SIGNAL or_3033_nl : STD_LOGIC;
  SIGNAL or_3031_nl : STD_LOGIC;
  SIGNAL mux_2831_nl : STD_LOGIC;
  SIGNAL mux_2830_nl : STD_LOGIC;
  SIGNAL or_3030_nl : STD_LOGIC;
  SIGNAL or_3028_nl : STD_LOGIC;
  SIGNAL mux_2829_nl : STD_LOGIC;
  SIGNAL mux_2828_nl : STD_LOGIC;
  SIGNAL mux_2827_nl : STD_LOGIC;
  SIGNAL mux_2826_nl : STD_LOGIC;
  SIGNAL mux_2825_nl : STD_LOGIC;
  SIGNAL or_3026_nl : STD_LOGIC;
  SIGNAL or_3021_nl : STD_LOGIC;
  SIGNAL mux_2824_nl : STD_LOGIC;
  SIGNAL mux_2818_nl : STD_LOGIC;
  SIGNAL or_3009_nl : STD_LOGIC;
  SIGNAL mux_2872_nl : STD_LOGIC;
  SIGNAL mux_2871_nl : STD_LOGIC;
  SIGNAL and_1490_nl : STD_LOGIC;
  SIGNAL mux_2892_nl : STD_LOGIC;
  SIGNAL mux_2891_nl : STD_LOGIC;
  SIGNAL mux_2890_nl : STD_LOGIC;
  SIGNAL or_3074_nl : STD_LOGIC;
  SIGNAL nand_155_nl : STD_LOGIC;
  SIGNAL mux_2889_nl : STD_LOGIC;
  SIGNAL or_3072_nl : STD_LOGIC;
  SIGNAL mux_2888_nl : STD_LOGIC;
  SIGNAL mux_2887_nl : STD_LOGIC;
  SIGNAL nor_906_nl : STD_LOGIC;
  SIGNAL mux_2886_nl : STD_LOGIC;
  SIGNAL mux_2885_nl : STD_LOGIC;
  SIGNAL or_3071_nl : STD_LOGIC;
  SIGNAL mux_2884_nl : STD_LOGIC;
  SIGNAL mux_2883_nl : STD_LOGIC;
  SIGNAL mux_2882_nl : STD_LOGIC;
  SIGNAL nor_1569_nl : STD_LOGIC;
  SIGNAL nand_154_nl : STD_LOGIC;
  SIGNAL mux_2881_nl : STD_LOGIC;
  SIGNAL mux_2875_nl : STD_LOGIC;
  SIGNAL or_4453_nl : STD_LOGIC;
  SIGNAL mux_2874_nl : STD_LOGIC;
  SIGNAL or_3057_nl : STD_LOGIC;
  SIGNAL mux_2930_nl : STD_LOGIC;
  SIGNAL mux_2929_nl : STD_LOGIC;
  SIGNAL and_1477_nl : STD_LOGIC;
  SIGNAL mux_2954_nl : STD_LOGIC;
  SIGNAL mux_2953_nl : STD_LOGIC;
  SIGNAL or_3131_nl : STD_LOGIC;
  SIGNAL or_3129_nl : STD_LOGIC;
  SIGNAL mux_2952_nl : STD_LOGIC;
  SIGNAL mux_2951_nl : STD_LOGIC;
  SIGNAL mux_2950_nl : STD_LOGIC;
  SIGNAL or_3128_nl : STD_LOGIC;
  SIGNAL mux_2949_nl : STD_LOGIC;
  SIGNAL or_3127_nl : STD_LOGIC;
  SIGNAL mux_2948_nl : STD_LOGIC;
  SIGNAL mux_2947_nl : STD_LOGIC;
  SIGNAL or_3124_nl : STD_LOGIC;
  SIGNAL mux_2946_nl : STD_LOGIC;
  SIGNAL mux_2945_nl : STD_LOGIC;
  SIGNAL or_3123_nl : STD_LOGIC;
  SIGNAL or_3119_nl : STD_LOGIC;
  SIGNAL mux_2944_nl : STD_LOGIC;
  SIGNAL mux_2942_nl : STD_LOGIC;
  SIGNAL mux_2941_nl : STD_LOGIC;
  SIGNAL or_3113_nl : STD_LOGIC;
  SIGNAL mux_2940_nl : STD_LOGIC;
  SIGNAL mux_2939_nl : STD_LOGIC;
  SIGNAL mux_2938_nl : STD_LOGIC;
  SIGNAL mux_2937_nl : STD_LOGIC;
  SIGNAL mux_2936_nl : STD_LOGIC;
  SIGNAL mux_2935_nl : STD_LOGIC;
  SIGNAL mux_2934_nl : STD_LOGIC;
  SIGNAL or_3109_nl : STD_LOGIC;
  SIGNAL or_3098_nl : STD_LOGIC;
  SIGNAL mux_2987_nl : STD_LOGIC;
  SIGNAL mux_2986_nl : STD_LOGIC;
  SIGNAL and_1467_nl : STD_LOGIC;
  SIGNAL mux_2983_nl : STD_LOGIC;
  SIGNAL mux_2982_nl : STD_LOGIC;
  SIGNAL mux_2981_nl : STD_LOGIC;
  SIGNAL or_3149_nl : STD_LOGIC;
  SIGNAL mux_2979_nl : STD_LOGIC;
  SIGNAL mux_2978_nl : STD_LOGIC;
  SIGNAL mux_2977_nl : STD_LOGIC;
  SIGNAL mux_3009_nl : STD_LOGIC;
  SIGNAL mux_3008_nl : STD_LOGIC;
  SIGNAL mux_3007_nl : STD_LOGIC;
  SIGNAL or_3189_nl : STD_LOGIC;
  SIGNAL nand_159_nl : STD_LOGIC;
  SIGNAL mux_3006_nl : STD_LOGIC;
  SIGNAL mux_3005_nl : STD_LOGIC;
  SIGNAL mux_3004_nl : STD_LOGIC;
  SIGNAL or_3187_nl : STD_LOGIC;
  SIGNAL mux_3003_nl : STD_LOGIC;
  SIGNAL nor_943_nl : STD_LOGIC;
  SIGNAL mux_3002_nl : STD_LOGIC;
  SIGNAL mux_3001_nl : STD_LOGIC;
  SIGNAL or_3185_nl : STD_LOGIC;
  SIGNAL mux_3000_nl : STD_LOGIC;
  SIGNAL mux_2999_nl : STD_LOGIC;
  SIGNAL mux_2998_nl : STD_LOGIC;
  SIGNAL nor_1553_nl : STD_LOGIC;
  SIGNAL nand_158_nl : STD_LOGIC;
  SIGNAL mux_2997_nl : STD_LOGIC;
  SIGNAL mux_2996_nl : STD_LOGIC;
  SIGNAL mux_2990_nl : STD_LOGIC;
  SIGNAL nand_156_nl : STD_LOGIC;
  SIGNAL mux_2989_nl : STD_LOGIC;
  SIGNAL nor_1554_nl : STD_LOGIC;
  SIGNAL nor_1555_nl : STD_LOGIC;
  SIGNAL mux_3031_nl : STD_LOGIC;
  SIGNAL mux_3030_nl : STD_LOGIC;
  SIGNAL or_3209_nl : STD_LOGIC;
  SIGNAL mux_3028_nl : STD_LOGIC;
  SIGNAL mux_3027_nl : STD_LOGIC;
  SIGNAL mux_3026_nl : STD_LOGIC;
  SIGNAL mux_3036_nl : STD_LOGIC;
  SIGNAL mux_3035_nl : STD_LOGIC;
  SIGNAL and_1461_nl : STD_LOGIC;
  SIGNAL mux_3054_nl : STD_LOGIC;
  SIGNAL mux_3053_nl : STD_LOGIC;
  SIGNAL mux_3052_nl : STD_LOGIC;
  SIGNAL or_3248_nl : STD_LOGIC;
  SIGNAL or_3246_nl : STD_LOGIC;
  SIGNAL mux_3051_nl : STD_LOGIC;
  SIGNAL mux_3050_nl : STD_LOGIC;
  SIGNAL or_3245_nl : STD_LOGIC;
  SIGNAL or_3243_nl : STD_LOGIC;
  SIGNAL mux_3049_nl : STD_LOGIC;
  SIGNAL mux_3048_nl : STD_LOGIC;
  SIGNAL mux_3047_nl : STD_LOGIC;
  SIGNAL mux_3046_nl : STD_LOGIC;
  SIGNAL mux_3045_nl : STD_LOGIC;
  SIGNAL or_3241_nl : STD_LOGIC;
  SIGNAL or_3236_nl : STD_LOGIC;
  SIGNAL mux_3044_nl : STD_LOGIC;
  SIGNAL mux_3038_nl : STD_LOGIC;
  SIGNAL or_3219_nl : STD_LOGIC;
  SIGNAL mux_3092_nl : STD_LOGIC;
  SIGNAL mux_3091_nl : STD_LOGIC;
  SIGNAL and_1449_nl : STD_LOGIC;
  SIGNAL mux_3112_nl : STD_LOGIC;
  SIGNAL mux_3111_nl : STD_LOGIC;
  SIGNAL mux_3110_nl : STD_LOGIC;
  SIGNAL or_3294_nl : STD_LOGIC;
  SIGNAL nand_164_nl : STD_LOGIC;
  SIGNAL mux_3109_nl : STD_LOGIC;
  SIGNAL or_3292_nl : STD_LOGIC;
  SIGNAL mux_3108_nl : STD_LOGIC;
  SIGNAL mux_3107_nl : STD_LOGIC;
  SIGNAL mux_3106_nl : STD_LOGIC;
  SIGNAL mux_3105_nl : STD_LOGIC;
  SIGNAL or_3291_nl : STD_LOGIC;
  SIGNAL mux_3104_nl : STD_LOGIC;
  SIGNAL mux_3103_nl : STD_LOGIC;
  SIGNAL mux_3102_nl : STD_LOGIC;
  SIGNAL and_2143_nl : STD_LOGIC;
  SIGNAL nand_163_nl : STD_LOGIC;
  SIGNAL mux_3101_nl : STD_LOGIC;
  SIGNAL mux_3095_nl : STD_LOGIC;
  SIGNAL or_4432_nl : STD_LOGIC;
  SIGNAL mux_3094_nl : STD_LOGIC;
  SIGNAL or_3272_nl : STD_LOGIC;
  SIGNAL mux_3150_nl : STD_LOGIC;
  SIGNAL mux_3149_nl : STD_LOGIC;
  SIGNAL and_1433_nl : STD_LOGIC;
  SIGNAL mux_3174_nl : STD_LOGIC;
  SIGNAL mux_3173_nl : STD_LOGIC;
  SIGNAL or_3350_nl : STD_LOGIC;
  SIGNAL or_3348_nl : STD_LOGIC;
  SIGNAL mux_3172_nl : STD_LOGIC;
  SIGNAL mux_3171_nl : STD_LOGIC;
  SIGNAL mux_3170_nl : STD_LOGIC;
  SIGNAL or_3347_nl : STD_LOGIC;
  SIGNAL mux_3169_nl : STD_LOGIC;
  SIGNAL or_3346_nl : STD_LOGIC;
  SIGNAL mux_3168_nl : STD_LOGIC;
  SIGNAL mux_3167_nl : STD_LOGIC;
  SIGNAL or_3343_nl : STD_LOGIC;
  SIGNAL mux_3166_nl : STD_LOGIC;
  SIGNAL mux_3165_nl : STD_LOGIC;
  SIGNAL or_3342_nl : STD_LOGIC;
  SIGNAL or_3338_nl : STD_LOGIC;
  SIGNAL mux_3164_nl : STD_LOGIC;
  SIGNAL mux_3162_nl : STD_LOGIC;
  SIGNAL mux_3161_nl : STD_LOGIC;
  SIGNAL mux_3160_nl : STD_LOGIC;
  SIGNAL mux_3159_nl : STD_LOGIC;
  SIGNAL mux_3158_nl : STD_LOGIC;
  SIGNAL mux_3157_nl : STD_LOGIC;
  SIGNAL mux_3156_nl : STD_LOGIC;
  SIGNAL or_3331_nl : STD_LOGIC;
  SIGNAL or_3328_nl : STD_LOGIC;
  SIGNAL mux_3155_nl : STD_LOGIC;
  SIGNAL mux_3154_nl : STD_LOGIC;
  SIGNAL or_3316_nl : STD_LOGIC;
  SIGNAL mux_3207_nl : STD_LOGIC;
  SIGNAL mux_3206_nl : STD_LOGIC;
  SIGNAL and_1423_nl : STD_LOGIC;
  SIGNAL mux_3203_nl : STD_LOGIC;
  SIGNAL mux_3202_nl : STD_LOGIC;
  SIGNAL mux_3201_nl : STD_LOGIC;
  SIGNAL or_3369_nl : STD_LOGIC;
  SIGNAL mux_3199_nl : STD_LOGIC;
  SIGNAL mux_3198_nl : STD_LOGIC;
  SIGNAL mux_3197_nl : STD_LOGIC;
  SIGNAL mux_3229_nl : STD_LOGIC;
  SIGNAL mux_3228_nl : STD_LOGIC;
  SIGNAL mux_3227_nl : STD_LOGIC;
  SIGNAL or_3399_nl : STD_LOGIC;
  SIGNAL nand_168_nl : STD_LOGIC;
  SIGNAL mux_3226_nl : STD_LOGIC;
  SIGNAL mux_3225_nl : STD_LOGIC;
  SIGNAL mux_3224_nl : STD_LOGIC;
  SIGNAL or_3397_nl : STD_LOGIC;
  SIGNAL mux_3223_nl : STD_LOGIC;
  SIGNAL nor_1016_nl : STD_LOGIC;
  SIGNAL mux_3222_nl : STD_LOGIC;
  SIGNAL mux_3221_nl : STD_LOGIC;
  SIGNAL or_3395_nl : STD_LOGIC;
  SIGNAL mux_3220_nl : STD_LOGIC;
  SIGNAL mux_3219_nl : STD_LOGIC;
  SIGNAL mux_3218_nl : STD_LOGIC;
  SIGNAL nor_1519_nl : STD_LOGIC;
  SIGNAL nand_167_nl : STD_LOGIC;
  SIGNAL mux_3217_nl : STD_LOGIC;
  SIGNAL mux_3216_nl : STD_LOGIC;
  SIGNAL mux_3210_nl : STD_LOGIC;
  SIGNAL nand_165_nl : STD_LOGIC;
  SIGNAL mux_3209_nl : STD_LOGIC;
  SIGNAL nor_1520_nl : STD_LOGIC;
  SIGNAL nor_1521_nl : STD_LOGIC;
  SIGNAL mux_3251_nl : STD_LOGIC;
  SIGNAL mux_3250_nl : STD_LOGIC;
  SIGNAL or_3420_nl : STD_LOGIC;
  SIGNAL mux_3248_nl : STD_LOGIC;
  SIGNAL mux_3247_nl : STD_LOGIC;
  SIGNAL mux_3246_nl : STD_LOGIC;
  SIGNAL mux_3256_nl : STD_LOGIC;
  SIGNAL mux_3255_nl : STD_LOGIC;
  SIGNAL and_1417_nl : STD_LOGIC;
  SIGNAL mux_3274_nl : STD_LOGIC;
  SIGNAL mux_3273_nl : STD_LOGIC;
  SIGNAL mux_3272_nl : STD_LOGIC;
  SIGNAL or_3452_nl : STD_LOGIC;
  SIGNAL or_3450_nl : STD_LOGIC;
  SIGNAL mux_3271_nl : STD_LOGIC;
  SIGNAL mux_3270_nl : STD_LOGIC;
  SIGNAL or_3449_nl : STD_LOGIC;
  SIGNAL or_3447_nl : STD_LOGIC;
  SIGNAL mux_3269_nl : STD_LOGIC;
  SIGNAL mux_3268_nl : STD_LOGIC;
  SIGNAL mux_3267_nl : STD_LOGIC;
  SIGNAL mux_3266_nl : STD_LOGIC;
  SIGNAL mux_3265_nl : STD_LOGIC;
  SIGNAL or_3445_nl : STD_LOGIC;
  SIGNAL or_3440_nl : STD_LOGIC;
  SIGNAL mux_3264_nl : STD_LOGIC;
  SIGNAL mux_3258_nl : STD_LOGIC;
  SIGNAL or_3428_nl : STD_LOGIC;
  SIGNAL mux_3312_nl : STD_LOGIC;
  SIGNAL mux_3311_nl : STD_LOGIC;
  SIGNAL and_1405_nl : STD_LOGIC;
  SIGNAL mux_3332_nl : STD_LOGIC;
  SIGNAL mux_3331_nl : STD_LOGIC;
  SIGNAL mux_3330_nl : STD_LOGIC;
  SIGNAL or_3493_nl : STD_LOGIC;
  SIGNAL nand_173_nl : STD_LOGIC;
  SIGNAL mux_3329_nl : STD_LOGIC;
  SIGNAL or_3491_nl : STD_LOGIC;
  SIGNAL mux_3328_nl : STD_LOGIC;
  SIGNAL mux_3327_nl : STD_LOGIC;
  SIGNAL mux_3326_nl : STD_LOGIC;
  SIGNAL mux_3325_nl : STD_LOGIC;
  SIGNAL or_3490_nl : STD_LOGIC;
  SIGNAL mux_3324_nl : STD_LOGIC;
  SIGNAL mux_3323_nl : STD_LOGIC;
  SIGNAL mux_3322_nl : STD_LOGIC;
  SIGNAL nor_1501_nl : STD_LOGIC;
  SIGNAL nand_172_nl : STD_LOGIC;
  SIGNAL mux_3321_nl : STD_LOGIC;
  SIGNAL mux_3315_nl : STD_LOGIC;
  SIGNAL or_4411_nl : STD_LOGIC;
  SIGNAL mux_3314_nl : STD_LOGIC;
  SIGNAL or_3476_nl : STD_LOGIC;
  SIGNAL mux_3370_nl : STD_LOGIC;
  SIGNAL mux_3369_nl : STD_LOGIC;
  SIGNAL and_1389_nl : STD_LOGIC;
  SIGNAL mux_3394_nl : STD_LOGIC;
  SIGNAL mux_3393_nl : STD_LOGIC;
  SIGNAL or_3547_nl : STD_LOGIC;
  SIGNAL or_3545_nl : STD_LOGIC;
  SIGNAL mux_3392_nl : STD_LOGIC;
  SIGNAL mux_3391_nl : STD_LOGIC;
  SIGNAL mux_3390_nl : STD_LOGIC;
  SIGNAL or_3544_nl : STD_LOGIC;
  SIGNAL mux_3389_nl : STD_LOGIC;
  SIGNAL or_3543_nl : STD_LOGIC;
  SIGNAL mux_3388_nl : STD_LOGIC;
  SIGNAL mux_3387_nl : STD_LOGIC;
  SIGNAL or_3540_nl : STD_LOGIC;
  SIGNAL mux_3386_nl : STD_LOGIC;
  SIGNAL mux_3385_nl : STD_LOGIC;
  SIGNAL or_3539_nl : STD_LOGIC;
  SIGNAL or_3535_nl : STD_LOGIC;
  SIGNAL mux_3384_nl : STD_LOGIC;
  SIGNAL mux_3382_nl : STD_LOGIC;
  SIGNAL mux_3381_nl : STD_LOGIC;
  SIGNAL or_3530_nl : STD_LOGIC;
  SIGNAL mux_3380_nl : STD_LOGIC;
  SIGNAL mux_3379_nl : STD_LOGIC;
  SIGNAL mux_3378_nl : STD_LOGIC;
  SIGNAL mux_3377_nl : STD_LOGIC;
  SIGNAL mux_3376_nl : STD_LOGIC;
  SIGNAL mux_3375_nl : STD_LOGIC;
  SIGNAL mux_3374_nl : STD_LOGIC;
  SIGNAL or_3526_nl : STD_LOGIC;
  SIGNAL or_3517_nl : STD_LOGIC;
  SIGNAL mux_3427_nl : STD_LOGIC;
  SIGNAL mux_3426_nl : STD_LOGIC;
  SIGNAL and_1376_nl : STD_LOGIC;
  SIGNAL mux_3423_nl : STD_LOGIC;
  SIGNAL mux_3422_nl : STD_LOGIC;
  SIGNAL mux_3421_nl : STD_LOGIC;
  SIGNAL or_3565_nl : STD_LOGIC;
  SIGNAL mux_3419_nl : STD_LOGIC;
  SIGNAL mux_3418_nl : STD_LOGIC;
  SIGNAL mux_3417_nl : STD_LOGIC;
  SIGNAL mux_3449_nl : STD_LOGIC;
  SIGNAL mux_3448_nl : STD_LOGIC;
  SIGNAL mux_3447_nl : STD_LOGIC;
  SIGNAL or_3599_nl : STD_LOGIC;
  SIGNAL nand_176_nl : STD_LOGIC;
  SIGNAL mux_3446_nl : STD_LOGIC;
  SIGNAL mux_3445_nl : STD_LOGIC;
  SIGNAL mux_3444_nl : STD_LOGIC;
  SIGNAL or_3597_nl : STD_LOGIC;
  SIGNAL mux_3443_nl : STD_LOGIC;
  SIGNAL mux_3442_nl : STD_LOGIC;
  SIGNAL mux_3441_nl : STD_LOGIC;
  SIGNAL or_3595_nl : STD_LOGIC;
  SIGNAL mux_3440_nl : STD_LOGIC;
  SIGNAL mux_3439_nl : STD_LOGIC;
  SIGNAL mux_3438_nl : STD_LOGIC;
  SIGNAL nor_1485_nl : STD_LOGIC;
  SIGNAL nand_175_nl : STD_LOGIC;
  SIGNAL mux_3437_nl : STD_LOGIC;
  SIGNAL mux_3436_nl : STD_LOGIC;
  SIGNAL mux_3430_nl : STD_LOGIC;
  SIGNAL nand_174_nl : STD_LOGIC;
  SIGNAL mux_3429_nl : STD_LOGIC;
  SIGNAL nor_1486_nl : STD_LOGIC;
  SIGNAL nor_1487_nl : STD_LOGIC;
  SIGNAL mux_3471_nl : STD_LOGIC;
  SIGNAL mux_3470_nl : STD_LOGIC;
  SIGNAL or_3619_nl : STD_LOGIC;
  SIGNAL mux_3468_nl : STD_LOGIC;
  SIGNAL mux_3467_nl : STD_LOGIC;
  SIGNAL mux_3466_nl : STD_LOGIC;
  SIGNAL mux_3476_nl : STD_LOGIC;
  SIGNAL mux_3475_nl : STD_LOGIC;
  SIGNAL and_1364_nl : STD_LOGIC;
  SIGNAL mux_3494_nl : STD_LOGIC;
  SIGNAL mux_3493_nl : STD_LOGIC;
  SIGNAL mux_3492_nl : STD_LOGIC;
  SIGNAL or_3656_nl : STD_LOGIC;
  SIGNAL or_3654_nl : STD_LOGIC;
  SIGNAL mux_3491_nl : STD_LOGIC;
  SIGNAL mux_3490_nl : STD_LOGIC;
  SIGNAL nand_513_nl : STD_LOGIC;
  SIGNAL or_3651_nl : STD_LOGIC;
  SIGNAL mux_3489_nl : STD_LOGIC;
  SIGNAL mux_3488_nl : STD_LOGIC;
  SIGNAL mux_3487_nl : STD_LOGIC;
  SIGNAL mux_3486_nl : STD_LOGIC;
  SIGNAL mux_3485_nl : STD_LOGIC;
  SIGNAL or_3649_nl : STD_LOGIC;
  SIGNAL or_3644_nl : STD_LOGIC;
  SIGNAL mux_3484_nl : STD_LOGIC;
  SIGNAL mux_3478_nl : STD_LOGIC;
  SIGNAL or_3629_nl : STD_LOGIC;
  SIGNAL mux_3532_nl : STD_LOGIC;
  SIGNAL mux_3531_nl : STD_LOGIC;
  SIGNAL and_1348_nl : STD_LOGIC;
  SIGNAL mux_3552_nl : STD_LOGIC;
  SIGNAL mux_3551_nl : STD_LOGIC;
  SIGNAL mux_3550_nl : STD_LOGIC;
  SIGNAL or_3696_nl : STD_LOGIC;
  SIGNAL nand_180_nl : STD_LOGIC;
  SIGNAL mux_3549_nl : STD_LOGIC;
  SIGNAL or_3694_nl : STD_LOGIC;
  SIGNAL mux_3548_nl : STD_LOGIC;
  SIGNAL mux_3547_nl : STD_LOGIC;
  SIGNAL mux_3546_nl : STD_LOGIC;
  SIGNAL mux_3545_nl : STD_LOGIC;
  SIGNAL or_3693_nl : STD_LOGIC;
  SIGNAL mux_3544_nl : STD_LOGIC;
  SIGNAL mux_3543_nl : STD_LOGIC;
  SIGNAL mux_3542_nl : STD_LOGIC;
  SIGNAL nand_179_nl : STD_LOGIC;
  SIGNAL mux_3541_nl : STD_LOGIC;
  SIGNAL mux_3535_nl : STD_LOGIC;
  SIGNAL or_4388_nl : STD_LOGIC;
  SIGNAL mux_3534_nl : STD_LOGIC;
  SIGNAL or_3680_nl : STD_LOGIC;
  SIGNAL mux_3590_nl : STD_LOGIC;
  SIGNAL mux_3589_nl : STD_LOGIC;
  SIGNAL and_1326_nl : STD_LOGIC;
  SIGNAL mux_3592_nl : STD_LOGIC;
  SIGNAL nor_1463_nl : STD_LOGIC;
  SIGNAL nor_1464_nl : STD_LOGIC;
  SIGNAL mux_3593_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_62_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_1_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_63_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_3_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_64_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_65_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_66_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_7_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_67_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_68_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_69_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_70_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_71_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_72_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_73_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_15_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_74_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_75_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_76_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_77_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_78_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_79_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_80_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_81_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_82_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_83_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_84_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_85_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_86_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_87_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_and_88_nl : STD_LOGIC;
  SIGNAL mux_3594_nl : STD_LOGIC;
  SIGNAL nor_1462_nl : STD_LOGIC;
  SIGNAL mux_3595_nl : STD_LOGIC;
  SIGNAL mux_3596_nl : STD_LOGIC;
  SIGNAL nor_1459_nl : STD_LOGIC;
  SIGNAL nor_1460_nl : STD_LOGIC;
  SIGNAL mux_3597_nl : STD_LOGIC;
  SIGNAL mux_3598_nl : STD_LOGIC;
  SIGNAL nor_1457_nl : STD_LOGIC;
  SIGNAL nor_1458_nl : STD_LOGIC;
  SIGNAL mux_3599_nl : STD_LOGIC;
  SIGNAL mux_3600_nl : STD_LOGIC;
  SIGNAL nor_1455_nl : STD_LOGIC;
  SIGNAL nor_1456_nl : STD_LOGIC;
  SIGNAL mux_3601_nl : STD_LOGIC;
  SIGNAL mux_3602_nl : STD_LOGIC;
  SIGNAL nor_1453_nl : STD_LOGIC;
  SIGNAL nor_1454_nl : STD_LOGIC;
  SIGNAL mux_3603_nl : STD_LOGIC;
  SIGNAL mux_3604_nl : STD_LOGIC;
  SIGNAL nor_1451_nl : STD_LOGIC;
  SIGNAL nor_1452_nl : STD_LOGIC;
  SIGNAL mux_3605_nl : STD_LOGIC;
  SIGNAL mux_3606_nl : STD_LOGIC;
  SIGNAL nor_1449_nl : STD_LOGIC;
  SIGNAL nor_1450_nl : STD_LOGIC;
  SIGNAL mux_3607_nl : STD_LOGIC;
  SIGNAL mux_3608_nl : STD_LOGIC;
  SIGNAL nor_1447_nl : STD_LOGIC;
  SIGNAL nor_1448_nl : STD_LOGIC;
  SIGNAL mux_3609_nl : STD_LOGIC;
  SIGNAL mux_3610_nl : STD_LOGIC;
  SIGNAL nor_1446_nl : STD_LOGIC;
  SIGNAL mux_3611_nl : STD_LOGIC;
  SIGNAL mux_3612_nl : STD_LOGIC;
  SIGNAL nor_1443_nl : STD_LOGIC;
  SIGNAL nor_1444_nl : STD_LOGIC;
  SIGNAL mux_3613_nl : STD_LOGIC;
  SIGNAL mux_3614_nl : STD_LOGIC;
  SIGNAL nor_1441_nl : STD_LOGIC;
  SIGNAL nor_1442_nl : STD_LOGIC;
  SIGNAL mux_3615_nl : STD_LOGIC;
  SIGNAL mux_3616_nl : STD_LOGIC;
  SIGNAL nor_1439_nl : STD_LOGIC;
  SIGNAL nor_1440_nl : STD_LOGIC;
  SIGNAL mux_3617_nl : STD_LOGIC;
  SIGNAL mux_3618_nl : STD_LOGIC;
  SIGNAL nor_1437_nl : STD_LOGIC;
  SIGNAL nor_1438_nl : STD_LOGIC;
  SIGNAL mux_3619_nl : STD_LOGIC;
  SIGNAL mux_3620_nl : STD_LOGIC;
  SIGNAL nor_1435_nl : STD_LOGIC;
  SIGNAL nor_1436_nl : STD_LOGIC;
  SIGNAL mux_3621_nl : STD_LOGIC;
  SIGNAL mux_3622_nl : STD_LOGIC;
  SIGNAL nor_1433_nl : STD_LOGIC;
  SIGNAL nor_1434_nl : STD_LOGIC;
  SIGNAL mux_3623_nl : STD_LOGIC;
  SIGNAL mux_3624_nl : STD_LOGIC;
  SIGNAL nor_1431_nl : STD_LOGIC;
  SIGNAL nor_1432_nl : STD_LOGIC;
  SIGNAL mux_3625_nl : STD_LOGIC;
  SIGNAL or_1283_nl : STD_LOGIC;
  SIGNAL mux_3626_nl : STD_LOGIC;
  SIGNAL nor_1430_nl : STD_LOGIC;
  SIGNAL mux_3627_nl : STD_LOGIC;
  SIGNAL or_1340_nl : STD_LOGIC;
  SIGNAL mux_3628_nl : STD_LOGIC;
  SIGNAL nor_1427_nl : STD_LOGIC;
  SIGNAL nor_1428_nl : STD_LOGIC;
  SIGNAL mux_3629_nl : STD_LOGIC;
  SIGNAL or_1393_nl : STD_LOGIC;
  SIGNAL mux_3630_nl : STD_LOGIC;
  SIGNAL nor_1425_nl : STD_LOGIC;
  SIGNAL nor_1426_nl : STD_LOGIC;
  SIGNAL mux_3631_nl : STD_LOGIC;
  SIGNAL or_1445_nl : STD_LOGIC;
  SIGNAL mux_3632_nl : STD_LOGIC;
  SIGNAL nor_1423_nl : STD_LOGIC;
  SIGNAL nor_1424_nl : STD_LOGIC;
  SIGNAL mux_3633_nl : STD_LOGIC;
  SIGNAL or_1510_nl : STD_LOGIC;
  SIGNAL mux_3634_nl : STD_LOGIC;
  SIGNAL nor_1421_nl : STD_LOGIC;
  SIGNAL nor_1422_nl : STD_LOGIC;
  SIGNAL mux_3635_nl : STD_LOGIC;
  SIGNAL or_1578_nl : STD_LOGIC;
  SIGNAL mux_3636_nl : STD_LOGIC;
  SIGNAL nor_1419_nl : STD_LOGIC;
  SIGNAL nor_1420_nl : STD_LOGIC;
  SIGNAL mux_3637_nl : STD_LOGIC;
  SIGNAL or_1638_nl : STD_LOGIC;
  SIGNAL mux_3638_nl : STD_LOGIC;
  SIGNAL nor_1417_nl : STD_LOGIC;
  SIGNAL nor_1418_nl : STD_LOGIC;
  SIGNAL mux_3639_nl : STD_LOGIC;
  SIGNAL or_1697_nl : STD_LOGIC;
  SIGNAL mux_3640_nl : STD_LOGIC;
  SIGNAL nor_1415_nl : STD_LOGIC;
  SIGNAL nor_1416_nl : STD_LOGIC;
  SIGNAL mux_3641_nl : STD_LOGIC;
  SIGNAL or_1758_nl : STD_LOGIC;
  SIGNAL mux_3642_nl : STD_LOGIC;
  SIGNAL nor_1413_nl : STD_LOGIC;
  SIGNAL nor_1414_nl : STD_LOGIC;
  SIGNAL mux_3643_nl : STD_LOGIC;
  SIGNAL or_1814_nl : STD_LOGIC;
  SIGNAL mux_3644_nl : STD_LOGIC;
  SIGNAL nor_1411_nl : STD_LOGIC;
  SIGNAL nor_1412_nl : STD_LOGIC;
  SIGNAL mux_3645_nl : STD_LOGIC;
  SIGNAL or_1867_nl : STD_LOGIC;
  SIGNAL mux_3646_nl : STD_LOGIC;
  SIGNAL and_2133_nl : STD_LOGIC;
  SIGNAL nor_1410_nl : STD_LOGIC;
  SIGNAL mux_3647_nl : STD_LOGIC;
  SIGNAL nand_378_nl : STD_LOGIC;
  SIGNAL mux_3648_nl : STD_LOGIC;
  SIGNAL nor_1407_nl : STD_LOGIC;
  SIGNAL nor_1408_nl : STD_LOGIC;
  SIGNAL mux_3649_nl : STD_LOGIC;
  SIGNAL or_1988_nl : STD_LOGIC;
  SIGNAL mux_3650_nl : STD_LOGIC;
  SIGNAL nor_1405_nl : STD_LOGIC;
  SIGNAL nor_1406_nl : STD_LOGIC;
  SIGNAL mux_3651_nl : STD_LOGIC;
  SIGNAL or_2042_nl : STD_LOGIC;
  SIGNAL mux_3652_nl : STD_LOGIC;
  SIGNAL nor_1403_nl : STD_LOGIC;
  SIGNAL nor_1404_nl : STD_LOGIC;
  SIGNAL mux_3653_nl : STD_LOGIC;
  SIGNAL or_2091_nl : STD_LOGIC;
  SIGNAL mux_3654_nl : STD_LOGIC;
  SIGNAL and_1324_nl : STD_LOGIC;
  SIGNAL and_1325_nl : STD_LOGIC;
  SIGNAL mux_3655_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_tf_mux_1_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL not_10627_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_k_mux_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL not_nl : STD_LOGIC;
  SIGNAL and_1112_nl : STD_LOGIC;
  SIGNAL mux_3668_nl : STD_LOGIC;
  SIGNAL mux_3667_nl : STD_LOGIC;
  SIGNAL mux_3666_nl : STD_LOGIC;
  SIGNAL mux_3665_nl : STD_LOGIC;
  SIGNAL and_1322_nl : STD_LOGIC;
  SIGNAL mux_3664_nl : STD_LOGIC;
  SIGNAL or_3820_nl : STD_LOGIC;
  SIGNAL mux_3663_nl : STD_LOGIC;
  SIGNAL mux_3662_nl : STD_LOGIC;
  SIGNAL mux_3661_nl : STD_LOGIC;
  SIGNAL or_3817_nl : STD_LOGIC;
  SIGNAL mux_3660_nl : STD_LOGIC;
  SIGNAL nand_530_nl : STD_LOGIC;
  SIGNAL mux_3658_nl : STD_LOGIC;
  SIGNAL mux_3657_nl : STD_LOGIC;
  SIGNAL mux_3656_nl : STD_LOGIC;
  SIGNAL nor_1393_nl : STD_LOGIC;
  SIGNAL mux_3677_nl : STD_LOGIC;
  SIGNAL mux_3676_nl : STD_LOGIC;
  SIGNAL and_1319_nl : STD_LOGIC;
  SIGNAL mux_3675_nl : STD_LOGIC;
  SIGNAL nor_1394_nl : STD_LOGIC;
  SIGNAL nor_1396_nl : STD_LOGIC;
  SIGNAL nor_1397_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_k_mux1h_1_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL S2_INNER_LOOP1_r_S2_INNER_LOOP1_r_and_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL not_9789_nl : STD_LOGIC;
  SIGNAL mux_4109_nl : STD_LOGIC;
  SIGNAL mux_4108_nl : STD_LOGIC;
  SIGNAL mux_4107_nl : STD_LOGIC;
  SIGNAL nor_1262_nl : STD_LOGIC;
  SIGNAL mux_4106_nl : STD_LOGIC;
  SIGNAL mux_4105_nl : STD_LOGIC;
  SIGNAL mux_4104_nl : STD_LOGIC;
  SIGNAL mux_4103_nl : STD_LOGIC;
  SIGNAL mux_4102_nl : STD_LOGIC;
  SIGNAL and_1270_nl : STD_LOGIC;
  SIGNAL mux_4101_nl : STD_LOGIC;
  SIGNAL nor_1263_nl : STD_LOGIC;
  SIGNAL mux_4100_nl : STD_LOGIC;
  SIGNAL mux_4099_nl : STD_LOGIC;
  SIGNAL mux_4098_nl : STD_LOGIC;
  SIGNAL mux_4097_nl : STD_LOGIC;
  SIGNAL mux_4096_nl : STD_LOGIC;
  SIGNAL mux_4095_nl : STD_LOGIC;
  SIGNAL mux_4093_nl : STD_LOGIC;
  SIGNAL mux_4092_nl : STD_LOGIC;
  SIGNAL and_1172_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_k_or_nl : STD_LOGIC;
  SIGNAL and_1179_nl : STD_LOGIC;
  SIGNAL mux_3729_nl : STD_LOGIC;
  SIGNAL mux_3728_nl : STD_LOGIC;
  SIGNAL nor_2306_nl : STD_LOGIC;
  SIGNAL nor_2308_nl : STD_LOGIC;
  SIGNAL mux_3741_nl : STD_LOGIC;
  SIGNAL mux_3740_nl : STD_LOGIC;
  SIGNAL mux_3739_nl : STD_LOGIC;
  SIGNAL mux_3738_nl : STD_LOGIC;
  SIGNAL or_3906_nl : STD_LOGIC;
  SIGNAL and_1307_nl : STD_LOGIC;
  SIGNAL mux_3736_nl : STD_LOGIC;
  SIGNAL mux_3735_nl : STD_LOGIC;
  SIGNAL mux_3734_nl : STD_LOGIC;
  SIGNAL mux_3733_nl : STD_LOGIC;
  SIGNAL mux_3732_nl : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_p_or_nl : STD_LOGIC;
  SIGNAL mux_3727_nl : STD_LOGIC;
  SIGNAL or_4690_nl : STD_LOGIC;
  SIGNAL nand_534_nl : STD_LOGIC;
  SIGNAL mux_3726_nl : STD_LOGIC;
  SIGNAL and_1312_nl : STD_LOGIC;
  SIGNAL and_1313_nl : STD_LOGIC;
  SIGNAL mux_3724_nl : STD_LOGIC;
  SIGNAL nor_1362_nl : STD_LOGIC;
  SIGNAL nor_1363_nl : STD_LOGIC;
  SIGNAL mux_4278_nl : STD_LOGIC;
  SIGNAL mux_4277_nl : STD_LOGIC;
  SIGNAL mux_4276_nl : STD_LOGIC;
  SIGNAL mux_4275_nl : STD_LOGIC;
  SIGNAL mux_4274_nl : STD_LOGIC;
  SIGNAL mux_4273_nl : STD_LOGIC;
  SIGNAL mux_4272_nl : STD_LOGIC;
  SIGNAL mux_4271_nl : STD_LOGIC;
  SIGNAL mux_4268_nl : STD_LOGIC;
  SIGNAL mux_4267_nl : STD_LOGIC;
  SIGNAL mux_4266_nl : STD_LOGIC;
  SIGNAL and_2894_nl : STD_LOGIC;
  SIGNAL mux_4265_nl : STD_LOGIC;
  SIGNAL mux_4264_nl : STD_LOGIC;
  SIGNAL mux_nl : STD_LOGIC;
  SIGNAL and_2895_nl : STD_LOGIC;
  SIGNAL mux_4293_nl : STD_LOGIC;
  SIGNAL mux_4292_nl : STD_LOGIC;
  SIGNAL mux_4291_nl : STD_LOGIC;
  SIGNAL or_4766_nl : STD_LOGIC;
  SIGNAL mux_4290_nl : STD_LOGIC;
  SIGNAL mux_4289_nl : STD_LOGIC;
  SIGNAL or_4764_nl : STD_LOGIC;
  SIGNAL mux_4288_nl : STD_LOGIC;
  SIGNAL mux_4287_nl : STD_LOGIC;
  SIGNAL or_4762_nl : STD_LOGIC;
  SIGNAL or_4761_nl : STD_LOGIC;
  SIGNAL mux_4286_nl : STD_LOGIC;
  SIGNAL mux_4285_nl : STD_LOGIC;
  SIGNAL mux_4284_nl : STD_LOGIC;
  SIGNAL or_4758_nl : STD_LOGIC;
  SIGNAL mux_4283_nl : STD_LOGIC;
  SIGNAL mux_4282_nl : STD_LOGIC;
  SIGNAL or_4755_nl : STD_LOGIC;
  SIGNAL mux_4281_nl : STD_LOGIC;
  SIGNAL mux_4280_nl : STD_LOGIC;
  SIGNAL or_4753_nl : STD_LOGIC;
  SIGNAL mux_4279_nl : STD_LOGIC;
  SIGNAL or_115_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_k_asn_S2_COPY_LOOP_for_i_5_0_sva_2_4_S1_OUTER_LOOP_k_and_nl
      : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL S1_OUTER_LOOP_k_mux1h_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL and_67_nl : STD_LOGIC;
  SIGNAL and_74_nl : STD_LOGIC;
  SIGNAL and_77_nl : STD_LOGIC;
  SIGNAL mux_94_nl : STD_LOGIC;
  SIGNAL mux_93_nl : STD_LOGIC;
  SIGNAL nor_nl : STD_LOGIC;
  SIGNAL mux_92_nl : STD_LOGIC;
  SIGNAL or_271_nl : STD_LOGIC;
  SIGNAL nand_535_nl : STD_LOGIC;
  SIGNAL and_2150_nl : STD_LOGIC;
  SIGNAL and_2151_nl : STD_LOGIC;
  SIGNAL mux_91_nl : STD_LOGIC;
  SIGNAL nor_2184_nl : STD_LOGIC;
  SIGNAL nor_2185_nl : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_for_p_S2_INNER_LOOP1_for_p_and_nl : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL not_9788_nl : STD_LOGIC;
  SIGNAL mux_3757_nl : STD_LOGIC;
  SIGNAL mux_3756_nl : STD_LOGIC;
  SIGNAL mux_3755_nl : STD_LOGIC;
  SIGNAL nor_1347_nl : STD_LOGIC;
  SIGNAL mux_3754_nl : STD_LOGIC;
  SIGNAL and_2138_nl : STD_LOGIC;
  SIGNAL and_1301_nl : STD_LOGIC;
  SIGNAL and_1302_nl : STD_LOGIC;
  SIGNAL mux_3753_nl : STD_LOGIC;
  SIGNAL nor_1352_nl : STD_LOGIC;
  SIGNAL mux_3776_nl : STD_LOGIC;
  SIGNAL mux_3775_nl : STD_LOGIC;
  SIGNAL mux_3774_nl : STD_LOGIC;
  SIGNAL mux_3773_nl : STD_LOGIC;
  SIGNAL mux_3772_nl : STD_LOGIC;
  SIGNAL mux_3771_nl : STD_LOGIC;
  SIGNAL mux_3770_nl : STD_LOGIC;
  SIGNAL mux_3768_nl : STD_LOGIC;
  SIGNAL mux_3767_nl : STD_LOGIC;
  SIGNAL mux_3766_nl : STD_LOGIC;
  SIGNAL mux_3765_nl : STD_LOGIC;
  SIGNAL mux_3764_nl : STD_LOGIC;
  SIGNAL mux_3763_nl : STD_LOGIC;
  SIGNAL mux_3762_nl : STD_LOGIC;
  SIGNAL or_3935_nl : STD_LOGIC;
  SIGNAL mux_3761_nl : STD_LOGIC;
  SIGNAL mux_3760_nl : STD_LOGIC;
  SIGNAL mux_3759_nl : STD_LOGIC;
  SIGNAL mux_3758_nl : STD_LOGIC;
  SIGNAL mux_4303_nl : STD_LOGIC;
  SIGNAL mux_4302_nl : STD_LOGIC;
  SIGNAL mux_4301_nl : STD_LOGIC;
  SIGNAL mux_4300_nl : STD_LOGIC;
  SIGNAL mux_4299_nl : STD_LOGIC;
  SIGNAL or_4853_nl : STD_LOGIC;
  SIGNAL mux_4298_nl : STD_LOGIC;
  SIGNAL mux_4297_nl : STD_LOGIC;
  SIGNAL nand_562_nl : STD_LOGIC;
  SIGNAL nor_2422_nl : STD_LOGIC;
  SIGNAL mux_4296_nl : STD_LOGIC;
  SIGNAL nor_2423_nl : STD_LOGIC;
  SIGNAL and_2866_nl : STD_LOGIC;
  SIGNAL mux_4295_nl : STD_LOGIC;
  SIGNAL mux_4294_nl : STD_LOGIC;
  SIGNAL or_4768_nl : STD_LOGIC;
  SIGNAL mux_4318_nl : STD_LOGIC;
  SIGNAL mux_4317_nl : STD_LOGIC;
  SIGNAL mux_4316_nl : STD_LOGIC;
  SIGNAL mux_4315_nl : STD_LOGIC;
  SIGNAL mux_4314_nl : STD_LOGIC;
  SIGNAL mux_4313_nl : STD_LOGIC;
  SIGNAL mux_4312_nl : STD_LOGIC;
  SIGNAL mux_4311_nl : STD_LOGIC;
  SIGNAL mux_4310_nl : STD_LOGIC;
  SIGNAL or_4782_nl : STD_LOGIC;
  SIGNAL mux_4309_nl : STD_LOGIC;
  SIGNAL mux_4411_nl : STD_LOGIC;
  SIGNAL nor_2420_nl : STD_LOGIC;
  SIGNAL mux_4308_nl : STD_LOGIC;
  SIGNAL nor_2421_nl : STD_LOGIC;
  SIGNAL mux_4307_nl : STD_LOGIC;
  SIGNAL mux_4306_nl : STD_LOGIC;
  SIGNAL and_2889_nl : STD_LOGIC;
  SIGNAL mux_4305_nl : STD_LOGIC;
  SIGNAL mux_4304_nl : STD_LOGIC;
  SIGNAL or_4776_nl : STD_LOGIC;
  SIGNAL mux_4334_nl : STD_LOGIC;
  SIGNAL mux_4333_nl : STD_LOGIC;
  SIGNAL mux_4332_nl : STD_LOGIC;
  SIGNAL mux_4331_nl : STD_LOGIC;
  SIGNAL or_4796_nl : STD_LOGIC;
  SIGNAL mux_4330_nl : STD_LOGIC;
  SIGNAL or_4795_nl : STD_LOGIC;
  SIGNAL mux_4329_nl : STD_LOGIC;
  SIGNAL or_4793_nl : STD_LOGIC;
  SIGNAL or_4792_nl : STD_LOGIC;
  SIGNAL mux_4328_nl : STD_LOGIC;
  SIGNAL mux_4327_nl : STD_LOGIC;
  SIGNAL mux_4326_nl : STD_LOGIC;
  SIGNAL mux_4325_nl : STD_LOGIC;
  SIGNAL or_4790_nl : STD_LOGIC;
  SIGNAL or_4789_nl : STD_LOGIC;
  SIGNAL or_4788_nl : STD_LOGIC;
  SIGNAL mux_4324_nl : STD_LOGIC;
  SIGNAL or_4787_nl : STD_LOGIC;
  SIGNAL mux_4323_nl : STD_LOGIC;
  SIGNAL mux_4322_nl : STD_LOGIC;
  SIGNAL mux_4321_nl : STD_LOGIC;
  SIGNAL or_4786_nl : STD_LOGIC;
  SIGNAL mux_4320_nl : STD_LOGIC;
  SIGNAL mux_4319_nl : STD_LOGIC;
  SIGNAL S2_INNER_LOOP1_S2_INNER_LOOP1_and_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL nor_2209_nl : STD_LOGIC;
  SIGNAL mux_106_nl : STD_LOGIC;
  SIGNAL or_4683_nl : STD_LOGIC;
  SIGNAL mux_105_nl : STD_LOGIC;
  SIGNAL or_290_nl : STD_LOGIC;
  SIGNAL or_289_nl : STD_LOGIC;
  SIGNAL or_4684_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_mux1h_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL S5_COPY_LOOP_for_acc_6_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL operator_20_true_1_acc_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL and_1193_nl : STD_LOGIC;
  SIGNAL mux_3828_nl : STD_LOGIC;
  SIGNAL mux_3827_nl : STD_LOGIC;
  SIGNAL mux_3826_nl : STD_LOGIC;
  SIGNAL mux_3825_nl : STD_LOGIC;
  SIGNAL mux_48_nl : STD_LOGIC;
  SIGNAL mux_47_nl : STD_LOGIC;
  SIGNAL mux_3822_nl : STD_LOGIC;
  SIGNAL mux_3820_nl : STD_LOGIC;
  SIGNAL mux_3818_nl : STD_LOGIC;
  SIGNAL mux_3817_nl : STD_LOGIC;
  SIGNAL or_3984_nl : STD_LOGIC;
  SIGNAL mux_3816_nl : STD_LOGIC;
  SIGNAL mux_3815_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_nand_nl : STD_LOGIC;
  SIGNAL mux_3814_nl : STD_LOGIC;
  SIGNAL mux_3813_nl : STD_LOGIC;
  SIGNAL or_3982_nl : STD_LOGIC;
  SIGNAL or_3981_nl : STD_LOGIC;
  SIGNAL mux_4361_nl : STD_LOGIC;
  SIGNAL mux_4360_nl : STD_LOGIC;
  SIGNAL mux_4359_nl : STD_LOGIC;
  SIGNAL mux_4358_nl : STD_LOGIC;
  SIGNAL mux_4357_nl : STD_LOGIC;
  SIGNAL mux_4356_nl : STD_LOGIC;
  SIGNAL mux_4355_nl : STD_LOGIC;
  SIGNAL mux_4354_nl : STD_LOGIC;
  SIGNAL mux_4353_nl : STD_LOGIC;
  SIGNAL mux_4352_nl : STD_LOGIC;
  SIGNAL mux_4351_nl : STD_LOGIC;
  SIGNAL mux_4350_nl : STD_LOGIC;
  SIGNAL and_2885_nl : STD_LOGIC;
  SIGNAL mux_4349_nl : STD_LOGIC;
  SIGNAL mux_4348_nl : STD_LOGIC;
  SIGNAL mux_4347_nl : STD_LOGIC;
  SIGNAL mux_4346_nl : STD_LOGIC;
  SIGNAL mux_4345_nl : STD_LOGIC;
  SIGNAL mux_4344_nl : STD_LOGIC;
  SIGNAL mux_4343_nl : STD_LOGIC;
  SIGNAL mux_4342_nl : STD_LOGIC;
  SIGNAL nor_2417_nl : STD_LOGIC;
  SIGNAL mux_4341_nl : STD_LOGIC;
  SIGNAL mux_4340_nl : STD_LOGIC;
  SIGNAL mux_4339_nl : STD_LOGIC;
  SIGNAL mux_4338_nl : STD_LOGIC;
  SIGNAL mux_4337_nl : STD_LOGIC;
  SIGNAL nor_2418_nl : STD_LOGIC;
  SIGNAL mux_4335_nl : STD_LOGIC;
  SIGNAL mux_4373_nl : STD_LOGIC;
  SIGNAL mux_4372_nl : STD_LOGIC;
  SIGNAL mux_4371_nl : STD_LOGIC;
  SIGNAL mux_4370_nl : STD_LOGIC;
  SIGNAL nor_2410_nl : STD_LOGIC;
  SIGNAL mux_4369_nl : STD_LOGIC;
  SIGNAL mux_4368_nl : STD_LOGIC;
  SIGNAL mux_4367_nl : STD_LOGIC;
  SIGNAL mux_4366_nl : STD_LOGIC;
  SIGNAL mux_4365_nl : STD_LOGIC;
  SIGNAL mux_4364_nl : STD_LOGIC;
  SIGNAL nor_2413_nl : STD_LOGIC;
  SIGNAL nor_2414_nl : STD_LOGIC;
  SIGNAL mux_4363_nl : STD_LOGIC;
  SIGNAL nor_2415_nl : STD_LOGIC;
  SIGNAL mux_4362_nl : STD_LOGIC;
  SIGNAL or_4810_nl : STD_LOGIC;
  SIGNAL or_4808_nl : STD_LOGIC;
  SIGNAL nor_2416_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_25_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_26_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_nor_3_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_28_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_nor_7_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_32_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_45_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_39_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_53_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_57_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_59_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_60_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_nor_nl : STD_LOGIC;
  SIGNAL mux_3854_nl : STD_LOGIC;
  SIGNAL mux_3853_nl : STD_LOGIC;
  SIGNAL or_4691_nl : STD_LOGIC;
  SIGNAL or_4692_nl : STD_LOGIC;
  SIGNAL or_4693_nl : STD_LOGIC;
  SIGNAL mux_3852_nl : STD_LOGIC;
  SIGNAL or_4020_nl : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_nor_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_nl : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_nor_1_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_1_nl : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_nor_3_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_3_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_6_nl : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_nor_7_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_7_nl : STD_LOGIC;
  SIGNAL butterFly_7_f1_butterFly_7_f1_nor_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_10_nl : STD_LOGIC;
  SIGNAL butterFly_7_f1_butterFly_7_f1_and_4_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_12_nl : STD_LOGIC;
  SIGNAL butterFly_7_f1_butterFly_7_f1_and_5_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_13_nl : STD_LOGIC;
  SIGNAL S2_COPY_LOOP_for_nor_14_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_nor_14_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_18_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_20_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_21_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_24_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_25_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_27_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_2_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_4_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_5_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_8_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_9_nl : STD_LOGIC;
  SIGNAL butterFly_7_f1_butterFly_7_f1_and_2_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_11_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_16_nl : STD_LOGIC;
  SIGNAL butterFly_4_f1_butterFly_4_f1_and_2_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_17_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_19_nl : STD_LOGIC;
  SIGNAL S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_23_nl : STD_LOGIC;
  SIGNAL and_1222_nl : STD_LOGIC;
  SIGNAL mux_3910_nl : STD_LOGIC;
  SIGNAL and_1287_nl : STD_LOGIC;
  SIGNAL mux_3909_nl : STD_LOGIC;
  SIGNAL and_1225_nl : STD_LOGIC;
  SIGNAL mux_3912_nl : STD_LOGIC;
  SIGNAL mux_3911_nl : STD_LOGIC;
  SIGNAL nor_1309_nl : STD_LOGIC;
  SIGNAL nor_1310_nl : STD_LOGIC;
  SIGNAL and_1286_nl : STD_LOGIC;
  SIGNAL and_1229_nl : STD_LOGIC;
  SIGNAL mux_3913_nl : STD_LOGIC;
  SIGNAL nor_1307_nl : STD_LOGIC;
  SIGNAL and_1231_nl : STD_LOGIC;
  SIGNAL mux_3914_nl : STD_LOGIC;
  SIGNAL and_1285_nl : STD_LOGIC;
  SIGNAL nor_1306_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_25_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_26_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_27_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_28_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_29_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_82_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_83_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_30_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_31_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_32_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_33_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_34_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_35_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_36_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_37_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_38_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_39_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_84_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_40_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_41_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_42_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_43_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_44_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_45_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_46_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_47_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_48_nl : STD_LOGIC;
  SIGNAL S1_OUTER_LOOP_for_mux_49_nl : STD_LOGIC;
  SIGNAL mux_4081_nl : STD_LOGIC;
  SIGNAL mux_4080_nl : STD_LOGIC;
  SIGNAL mux_4079_nl : STD_LOGIC;
  SIGNAL mux_4078_nl : STD_LOGIC;
  SIGNAL or_4296_nl : STD_LOGIC;
  SIGNAL mux_4077_nl : STD_LOGIC;
  SIGNAL mux_4076_nl : STD_LOGIC;
  SIGNAL mux_4072_nl : STD_LOGIC;
  SIGNAL mux_4071_nl : STD_LOGIC;
  SIGNAL mux_4070_nl : STD_LOGIC;
  SIGNAL mux_4391_nl : STD_LOGIC;
  SIGNAL mux_4390_nl : STD_LOGIC;
  SIGNAL mux_4389_nl : STD_LOGIC;
  SIGNAL mux_4388_nl : STD_LOGIC;
  SIGNAL mux_4387_nl : STD_LOGIC;
  SIGNAL or_4824_nl : STD_LOGIC;
  SIGNAL mux_4386_nl : STD_LOGIC;
  SIGNAL nor_2402_nl : STD_LOGIC;
  SIGNAL mux_4385_nl : STD_LOGIC;
  SIGNAL mux_4384_nl : STD_LOGIC;
  SIGNAL mux_4383_nl : STD_LOGIC;
  SIGNAL mux_4382_nl : STD_LOGIC;
  SIGNAL mux_4381_nl : STD_LOGIC;
  SIGNAL mux_4380_nl : STD_LOGIC;
  SIGNAL or_4821_nl : STD_LOGIC;
  SIGNAL nor_2403_nl : STD_LOGIC;
  SIGNAL mux_4379_nl : STD_LOGIC;
  SIGNAL mux_4378_nl : STD_LOGIC;
  SIGNAL mux_4377_nl : STD_LOGIC;
  SIGNAL and_2882_nl : STD_LOGIC;
  SIGNAL mux_4374_nl : STD_LOGIC;
  SIGNAL mux_4397_nl : STD_LOGIC;
  SIGNAL mux_4396_nl : STD_LOGIC;
  SIGNAL mux_4395_nl : STD_LOGIC;
  SIGNAL mux_4394_nl : STD_LOGIC;
  SIGNAL nor_2404_nl : STD_LOGIC;
  SIGNAL mux_4393_nl : STD_LOGIC;
  SIGNAL nor_2405_nl : STD_LOGIC;
  SIGNAL nor_2406_nl : STD_LOGIC;
  SIGNAL nor_2407_nl : STD_LOGIC;
  SIGNAL mux_4392_nl : STD_LOGIC;
  SIGNAL or_4831_nl : STD_LOGIC;
  SIGNAL or_4830_nl : STD_LOGIC;
  SIGNAL nor_2408_nl : STD_LOGIC;
  SIGNAL nor_2409_nl : STD_LOGIC;
  SIGNAL mux_4091_nl : STD_LOGIC;
  SIGNAL mux_4404_nl : STD_LOGIC;
  SIGNAL mux_4403_nl : STD_LOGIC;
  SIGNAL mux_4402_nl : STD_LOGIC;
  SIGNAL mux_4401_nl : STD_LOGIC;
  SIGNAL and_2879_nl : STD_LOGIC;
  SIGNAL or_4842_nl : STD_LOGIC;
  SIGNAL or_4841_nl : STD_LOGIC;
  SIGNAL mux_4400_nl : STD_LOGIC;
  SIGNAL or_4839_nl : STD_LOGIC;
  SIGNAL mux_4399_nl : STD_LOGIC;
  SIGNAL mux_4410_nl : STD_LOGIC;
  SIGNAL or_4849_nl : STD_LOGIC;
  SIGNAL mux_4409_nl : STD_LOGIC;
  SIGNAL mux_4408_nl : STD_LOGIC;
  SIGNAL and_2875_nl : STD_LOGIC;
  SIGNAL and_2877_nl : STD_LOGIC;
  SIGNAL mux_4407_nl : STD_LOGIC;
  SIGNAL mux_4406_nl : STD_LOGIC;
  SIGNAL or_4846_nl : STD_LOGIC;
  SIGNAL mux_4405_nl : STD_LOGIC;
  SIGNAL or_4845_nl : STD_LOGIC;
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_3_res_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mux_4413_nl : STD_LOGIC;
  SIGNAL and_2897_nl : STD_LOGIC;
  SIGNAL mux_4414_nl : STD_LOGIC;
  SIGNAL mux_4415_nl : STD_LOGIC;
  SIGNAL mux_4416_nl : STD_LOGIC;
  SIGNAL nor_2426_nl : STD_LOGIC;
  SIGNAL nor_2427_nl : STD_LOGIC;
  SIGNAL nor_2428_nl : STD_LOGIC;
  SIGNAL mux_4417_nl : STD_LOGIC;
  SIGNAL or_4856_nl : STD_LOGIC;
  SIGNAL nand_573_nl : STD_LOGIC;
  SIGNAL nor_2429_nl : STD_LOGIC;
  SIGNAL mux_4418_nl : STD_LOGIC;
  SIGNAL nor_2430_nl : STD_LOGIC;
  SIGNAL mux_4419_nl : STD_LOGIC;
  SIGNAL or_4857_nl : STD_LOGIC;
  SIGNAL and_2898_nl : STD_LOGIC;
  SIGNAL mux_4420_nl : STD_LOGIC;
  SIGNAL mux_4421_nl : STD_LOGIC;
  SIGNAL mux_4422_nl : STD_LOGIC;
  SIGNAL nand_574_nl : STD_LOGIC;
  SIGNAL nand_575_nl : STD_LOGIC;
  SIGNAL mux_4423_nl : STD_LOGIC;
  SIGNAL or_4858_nl : STD_LOGIC;
  SIGNAL or_4859_nl : STD_LOGIC;
  SIGNAL mux_4424_nl : STD_LOGIC;
  SIGNAL nor_2431_nl : STD_LOGIC;
  SIGNAL mux_4425_nl : STD_LOGIC;
  SIGNAL or_4860_nl : STD_LOGIC;
  SIGNAL or_4861_nl : STD_LOGIC;
  SIGNAL mux_4426_nl : STD_LOGIC;
  SIGNAL mux_4427_nl : STD_LOGIC;
  SIGNAL nor_2432_nl : STD_LOGIC;
  SIGNAL mux_4428_nl : STD_LOGIC;
  SIGNAL nor_2433_nl : STD_LOGIC;
  SIGNAL nor_2434_nl : STD_LOGIC;
  SIGNAL nor_2435_nl : STD_LOGIC;
  SIGNAL acc_15_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_3_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2918_nl : STD_LOGIC;
  SIGNAL acc_17_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_2_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2925_nl : STD_LOGIC;
  SIGNAL acc_19_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_1_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2929_nl : STD_LOGIC;
  SIGNAL and_2930_nl : STD_LOGIC;
  SIGNAL and_2931_nl : STD_LOGIC;
  SIGNAL and_2932_nl : STD_LOGIC;
  SIGNAL acc_20_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_7_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_21_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_6_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2934_nl : STD_LOGIC;
  SIGNAL and_2935_nl : STD_LOGIC;
  SIGNAL and_2936_nl : STD_LOGIC;
  SIGNAL and_2937_nl : STD_LOGIC;
  SIGNAL acc_18_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_5_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2926_nl : STD_LOGIC;
  SIGNAL and_2927_nl : STD_LOGIC;
  SIGNAL and_2928_nl : STD_LOGIC;
  SIGNAL acc_22_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_11_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2938_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_1_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_15_nl : STD_LOGIC;
  SIGNAL modulo_add_13_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_sub_18_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL nor_2169_nl : STD_LOGIC;
  SIGNAL or_4688_nl : STD_LOGIC;
  SIGNAL or_4689_nl : STD_LOGIC;
  SIGNAL mux_112_nl : STD_LOGIC;
  SIGNAL nor_2165_nl : STD_LOGIC;
  SIGNAL nor_2166_nl : STD_LOGIC;
  SIGNAL mux_113_nl : STD_LOGIC;
  SIGNAL or_4696_nl : STD_LOGIC;
  SIGNAL or_4697_nl : STD_LOGIC;
  SIGNAL and_2095_nl : STD_LOGIC;
  SIGNAL nor_2162_nl : STD_LOGIC;
  SIGNAL or_320_nl : STD_LOGIC;
  SIGNAL or_318_nl : STD_LOGIC;
  SIGNAL or_331_nl : STD_LOGIC;
  SIGNAL mux_127_nl : STD_LOGIC;
  SIGNAL or_329_nl : STD_LOGIC;
  SIGNAL or_341_nl : STD_LOGIC;
  SIGNAL mux_141_nl : STD_LOGIC;
  SIGNAL nand_502_nl : STD_LOGIC;
  SIGNAL nand_501_nl : STD_LOGIC;
  SIGNAL mux_155_nl : STD_LOGIC;
  SIGNAL nor_2154_nl : STD_LOGIC;
  SIGNAL nor_2150_nl : STD_LOGIC;
  SIGNAL nor_2151_nl : STD_LOGIC;
  SIGNAL or_405_nl : STD_LOGIC;
  SIGNAL and_2134_nl : STD_LOGIC;
  SIGNAL nor_2135_nl : STD_LOGIC;
  SIGNAL mux_211_nl : STD_LOGIC;
  SIGNAL or_452_nl : STD_LOGIC;
  SIGNAL mux_243_nl : STD_LOGIC;
  SIGNAL nor_2120_nl : STD_LOGIC;
  SIGNAL nor_2121_nl : STD_LOGIC;
  SIGNAL nor_2117_nl : STD_LOGIC;
  SIGNAL nor_2118_nl : STD_LOGIC;
  SIGNAL mux_262_nl : STD_LOGIC;
  SIGNAL or_483_nl : STD_LOGIC;
  SIGNAL mux_301_nl : STD_LOGIC;
  SIGNAL and_2057_nl : STD_LOGIC;
  SIGNAL and_2058_nl : STD_LOGIC;
  SIGNAL mux_300_nl : STD_LOGIC;
  SIGNAL or_527_nl : STD_LOGIC;
  SIGNAL and_2054_nl : STD_LOGIC;
  SIGNAL nor_2101_nl : STD_LOGIC;
  SIGNAL mux_316_nl : STD_LOGIC;
  SIGNAL or_534_nl : STD_LOGIC;
  SIGNAL or_560_nl : STD_LOGIC;
  SIGNAL or_558_nl : STD_LOGIC;
  SIGNAL or_571_nl : STD_LOGIC;
  SIGNAL mux_346_nl : STD_LOGIC;
  SIGNAL or_569_nl : STD_LOGIC;
  SIGNAL or_625_nl : STD_LOGIC;
  SIGNAL or_623_nl : STD_LOGIC;
  SIGNAL or_648_nl : STD_LOGIC;
  SIGNAL or_693_nl : STD_LOGIC;
  SIGNAL mux_515_nl : STD_LOGIC;
  SIGNAL and_2014_nl : STD_LOGIC;
  SIGNAL and_2015_nl : STD_LOGIC;
  SIGNAL mux_514_nl : STD_LOGIC;
  SIGNAL or_767_nl : STD_LOGIC;
  SIGNAL or_800_nl : STD_LOGIC;
  SIGNAL or_798_nl : STD_LOGIC;
  SIGNAL or_811_nl : STD_LOGIC;
  SIGNAL mux_555_nl : STD_LOGIC;
  SIGNAL or_809_nl : STD_LOGIC;
  SIGNAL or_874_nl : STD_LOGIC;
  SIGNAL or_915_nl : STD_LOGIC;
  SIGNAL mux_718_nl : STD_LOGIC;
  SIGNAL and_1972_nl : STD_LOGIC;
  SIGNAL and_1973_nl : STD_LOGIC;
  SIGNAL mux_717_nl : STD_LOGIC;
  SIGNAL or_988_nl : STD_LOGIC;
  SIGNAL or_1017_nl : STD_LOGIC;
  SIGNAL or_1015_nl : STD_LOGIC;
  SIGNAL or_1028_nl : STD_LOGIC;
  SIGNAL mux_761_nl : STD_LOGIC;
  SIGNAL or_1026_nl : STD_LOGIC;
  SIGNAL or_1097_nl : STD_LOGIC;
  SIGNAL or_1142_nl : STD_LOGIC;
  SIGNAL or_1140_nl : STD_LOGIC;
  SIGNAL mux_927_nl : STD_LOGIC;
  SIGNAL and_1923_nl : STD_LOGIC;
  SIGNAL and_1925_nl : STD_LOGIC;
  SIGNAL mux_926_nl : STD_LOGIC;
  SIGNAL nand_442_nl : STD_LOGIC;
  SIGNAL or_1245_nl : STD_LOGIC;
  SIGNAL or_1243_nl : STD_LOGIC;
  SIGNAL or_1255_nl : STD_LOGIC;
  SIGNAL mux_968_nl : STD_LOGIC;
  SIGNAL or_1253_nl : STD_LOGIC;
  SIGNAL or_1322_nl : STD_LOGIC;
  SIGNAL or_1362_nl : STD_LOGIC;
  SIGNAL mux_1141_nl : STD_LOGIC;
  SIGNAL and_1879_nl : STD_LOGIC;
  SIGNAL and_1880_nl : STD_LOGIC;
  SIGNAL mux_1140_nl : STD_LOGIC;
  SIGNAL or_1439_nl : STD_LOGIC;
  SIGNAL or_1470_nl : STD_LOGIC;
  SIGNAL or_1468_nl : STD_LOGIC;
  SIGNAL or_1480_nl : STD_LOGIC;
  SIGNAL mux_1185_nl : STD_LOGIC;
  SIGNAL or_1478_nl : STD_LOGIC;
  SIGNAL nand_546_nl : STD_LOGIC;
  SIGNAL or_1559_nl : STD_LOGIC;
  SIGNAL or_1604_nl : STD_LOGIC;
  SIGNAL or_1602_nl : STD_LOGIC;
  SIGNAL mux_1362_nl : STD_LOGIC;
  SIGNAL and_1831_nl : STD_LOGIC;
  SIGNAL and_1833_nl : STD_LOGIC;
  SIGNAL mux_1361_nl : STD_LOGIC;
  SIGNAL nand_408_nl : STD_LOGIC;
  SIGNAL or_1721_nl : STD_LOGIC;
  SIGNAL or_1719_nl : STD_LOGIC;
  SIGNAL or_1731_nl : STD_LOGIC;
  SIGNAL mux_1403_nl : STD_LOGIC;
  SIGNAL or_1729_nl : STD_LOGIC;
  SIGNAL or_1796_nl : STD_LOGIC;
  SIGNAL nand_396_nl : STD_LOGIC;
  SIGNAL mux_1576_nl : STD_LOGIC;
  SIGNAL and_1777_nl : STD_LOGIC;
  SIGNAL and_1779_nl : STD_LOGIC;
  SIGNAL mux_1575_nl : STD_LOGIC;
  SIGNAL nand_380_nl : STD_LOGIC;
  SIGNAL or_1949_nl : STD_LOGIC;
  SIGNAL or_1947_nl : STD_LOGIC;
  SIGNAL nand_518_nl : STD_LOGIC;
  SIGNAL mux_1620_nl : STD_LOGIC;
  SIGNAL or_1957_nl : STD_LOGIC;
  SIGNAL or_2025_nl : STD_LOGIC;
  SIGNAL nand_353_nl : STD_LOGIC;
  SIGNAL or_2062_nl : STD_LOGIC;
  SIGNAL mux_1792_nl : STD_LOGIC;
  SIGNAL and_1699_nl : STD_LOGIC;
  SIGNAL and_1701_nl : STD_LOGIC;
  SIGNAL mux_1791_nl : STD_LOGIC;
  SIGNAL nand_335_nl : STD_LOGIC;
  SIGNAL or_2140_nl : STD_LOGIC;
  SIGNAL or_2139_nl : STD_LOGIC;
  SIGNAL or_2142_nl : STD_LOGIC;
  SIGNAL or_2141_nl : STD_LOGIC;
  SIGNAL nor_1740_nl : STD_LOGIC;
  SIGNAL nor_1741_nl : STD_LOGIC;
  SIGNAL mux_1845_nl : STD_LOGIC;
  SIGNAL nor_1732_nl : STD_LOGIC;
  SIGNAL mux_1863_nl : STD_LOGIC;
  SIGNAL or_2184_nl : STD_LOGIC;
  SIGNAL or_2182_nl : STD_LOGIC;
  SIGNAL nor_1733_nl : STD_LOGIC;
  SIGNAL or_2209_nl : STD_LOGIC;
  SIGNAL mux_1886_nl : STD_LOGIC;
  SIGNAL or_2208_nl : STD_LOGIC;
  SIGNAL or_2207_nl : STD_LOGIC;
  SIGNAL mux_1885_nl : STD_LOGIC;
  SIGNAL mux_1884_nl : STD_LOGIC;
  SIGNAL or_2206_nl : STD_LOGIC;
  SIGNAL nand_112_nl : STD_LOGIC;
  SIGNAL mux_1883_nl : STD_LOGIC;
  SIGNAL or_2203_nl : STD_LOGIC;
  SIGNAL mux_1903_nl : STD_LOGIC;
  SIGNAL or_4685_nl : STD_LOGIC;
  SIGNAL or_4686_nl : STD_LOGIC;
  SIGNAL nor_1717_nl : STD_LOGIC;
  SIGNAL mux_1915_nl : STD_LOGIC;
  SIGNAL nand_532_nl : STD_LOGIC;
  SIGNAL or_2238_nl : STD_LOGIC;
  SIGNAL nor_1718_nl : STD_LOGIC;
  SIGNAL mux_1937_nl : STD_LOGIC;
  SIGNAL or_2262_nl : STD_LOGIC;
  SIGNAL or_2261_nl : STD_LOGIC;
  SIGNAL mux_1936_nl : STD_LOGIC;
  SIGNAL mux_1935_nl : STD_LOGIC;
  SIGNAL or_2259_nl : STD_LOGIC;
  SIGNAL or_2258_nl : STD_LOGIC;
  SIGNAL nand_115_nl : STD_LOGIC;
  SIGNAL mux_1934_nl : STD_LOGIC;
  SIGNAL nor_1713_nl : STD_LOGIC;
  SIGNAL nor_1714_nl : STD_LOGIC;
  SIGNAL and_1666_nl : STD_LOGIC;
  SIGNAL mux_1957_nl : STD_LOGIC;
  SIGNAL mux_1956_nl : STD_LOGIC;
  SIGNAL or_2277_nl : STD_LOGIC;
  SIGNAL mux_1955_nl : STD_LOGIC;
  SIGNAL or_2276_nl : STD_LOGIC;
  SIGNAL nor_1706_nl : STD_LOGIC;
  SIGNAL mux_1973_nl : STD_LOGIC;
  SIGNAL or_2289_nl : STD_LOGIC;
  SIGNAL or_2287_nl : STD_LOGIC;
  SIGNAL nor_1707_nl : STD_LOGIC;
  SIGNAL mux_1995_nl : STD_LOGIC;
  SIGNAL nand_117_nl : STD_LOGIC;
  SIGNAL mux_1994_nl : STD_LOGIC;
  SIGNAL mux_1993_nl : STD_LOGIC;
  SIGNAL or_2306_nl : STD_LOGIC;
  SIGNAL or_2312_nl : STD_LOGIC;
  SIGNAL mux_2011_nl : STD_LOGIC;
  SIGNAL nor_1701_nl : STD_LOGIC;
  SIGNAL nor_1702_nl : STD_LOGIC;
  SIGNAL and_1656_nl : STD_LOGIC;
  SIGNAL mux_2018_nl : STD_LOGIC;
  SIGNAL mux_2017_nl : STD_LOGIC;
  SIGNAL or_2323_nl : STD_LOGIC;
  SIGNAL mux_2016_nl : STD_LOGIC;
  SIGNAL or_2322_nl : STD_LOGIC;
  SIGNAL nor_1695_nl : STD_LOGIC;
  SIGNAL mux_2034_nl : STD_LOGIC;
  SIGNAL or_2333_nl : STD_LOGIC;
  SIGNAL nor_1696_nl : STD_LOGIC;
  SIGNAL or_2349_nl : STD_LOGIC;
  SIGNAL or_2348_nl : STD_LOGIC;
  SIGNAL or_2351_nl : STD_LOGIC;
  SIGNAL or_2350_nl : STD_LOGIC;
  SIGNAL or_2412_nl : STD_LOGIC;
  SIGNAL mux_2114_nl : STD_LOGIC;
  SIGNAL or_2411_nl : STD_LOGIC;
  SIGNAL or_2409_nl : STD_LOGIC;
  SIGNAL mux_2113_nl : STD_LOGIC;
  SIGNAL mux_2112_nl : STD_LOGIC;
  SIGNAL or_2407_nl : STD_LOGIC;
  SIGNAL nand_121_nl : STD_LOGIC;
  SIGNAL mux_2111_nl : STD_LOGIC;
  SIGNAL or_2403_nl : STD_LOGIC;
  SIGNAL mux_2162_nl : STD_LOGIC;
  SIGNAL or_2462_nl : STD_LOGIC;
  SIGNAL or_2460_nl : STD_LOGIC;
  SIGNAL mux_2161_nl : STD_LOGIC;
  SIGNAL mux_2160_nl : STD_LOGIC;
  SIGNAL or_2457_nl : STD_LOGIC;
  SIGNAL or_2455_nl : STD_LOGIC;
  SIGNAL nand_124_nl : STD_LOGIC;
  SIGNAL mux_2159_nl : STD_LOGIC;
  SIGNAL nor_1673_nl : STD_LOGIC;
  SIGNAL nor_1674_nl : STD_LOGIC;
  SIGNAL and_1626_nl : STD_LOGIC;
  SIGNAL mux_2186_nl : STD_LOGIC;
  SIGNAL mux_2185_nl : STD_LOGIC;
  SIGNAL or_2480_nl : STD_LOGIC;
  SIGNAL mux_2184_nl : STD_LOGIC;
  SIGNAL or_2479_nl : STD_LOGIC;
  SIGNAL mux_2218_nl : STD_LOGIC;
  SIGNAL nand_126_nl : STD_LOGIC;
  SIGNAL mux_2217_nl : STD_LOGIC;
  SIGNAL mux_2216_nl : STD_LOGIC;
  SIGNAL or_2502_nl : STD_LOGIC;
  SIGNAL or_2511_nl : STD_LOGIC;
  SIGNAL and_1615_nl : STD_LOGIC;
  SIGNAL mux_2244_nl : STD_LOGIC;
  SIGNAL mux_2243_nl : STD_LOGIC;
  SIGNAL or_2521_nl : STD_LOGIC;
  SIGNAL mux_2242_nl : STD_LOGIC;
  SIGNAL or_2520_nl : STD_LOGIC;
  SIGNAL or_2538_nl : STD_LOGIC;
  SIGNAL or_2537_nl : STD_LOGIC;
  SIGNAL or_2540_nl : STD_LOGIC;
  SIGNAL or_2539_nl : STD_LOGIC;
  SIGNAL or_2595_nl : STD_LOGIC;
  SIGNAL mux_2334_nl : STD_LOGIC;
  SIGNAL or_2594_nl : STD_LOGIC;
  SIGNAL or_2593_nl : STD_LOGIC;
  SIGNAL mux_2333_nl : STD_LOGIC;
  SIGNAL mux_2332_nl : STD_LOGIC;
  SIGNAL or_2592_nl : STD_LOGIC;
  SIGNAL nand_130_nl : STD_LOGIC;
  SIGNAL mux_2331_nl : STD_LOGIC;
  SIGNAL or_2589_nl : STD_LOGIC;
  SIGNAL mux_2382_nl : STD_LOGIC;
  SIGNAL or_2638_nl : STD_LOGIC;
  SIGNAL or_2637_nl : STD_LOGIC;
  SIGNAL mux_2381_nl : STD_LOGIC;
  SIGNAL mux_2380_nl : STD_LOGIC;
  SIGNAL or_2635_nl : STD_LOGIC;
  SIGNAL or_2634_nl : STD_LOGIC;
  SIGNAL nand_133_nl : STD_LOGIC;
  SIGNAL mux_2379_nl : STD_LOGIC;
  SIGNAL nor_1640_nl : STD_LOGIC;
  SIGNAL nor_1641_nl : STD_LOGIC;
  SIGNAL and_1585_nl : STD_LOGIC;
  SIGNAL mux_2402_nl : STD_LOGIC;
  SIGNAL mux_2401_nl : STD_LOGIC;
  SIGNAL or_2653_nl : STD_LOGIC;
  SIGNAL mux_2400_nl : STD_LOGIC;
  SIGNAL or_2652_nl : STD_LOGIC;
  SIGNAL mux_2438_nl : STD_LOGIC;
  SIGNAL nand_135_nl : STD_LOGIC;
  SIGNAL mux_2437_nl : STD_LOGIC;
  SIGNAL mux_2436_nl : STD_LOGIC;
  SIGNAL or_2675_nl : STD_LOGIC;
  SIGNAL or_2681_nl : STD_LOGIC;
  SIGNAL and_1574_nl : STD_LOGIC;
  SIGNAL mux_2460_nl : STD_LOGIC;
  SIGNAL mux_2459_nl : STD_LOGIC;
  SIGNAL or_2689_nl : STD_LOGIC;
  SIGNAL mux_2458_nl : STD_LOGIC;
  SIGNAL or_2688_nl : STD_LOGIC;
  SIGNAL or_2710_nl : STD_LOGIC;
  SIGNAL or_2709_nl : STD_LOGIC;
  SIGNAL or_2712_nl : STD_LOGIC;
  SIGNAL or_2711_nl : STD_LOGIC;
  SIGNAL or_2772_nl : STD_LOGIC;
  SIGNAL mux_2554_nl : STD_LOGIC;
  SIGNAL or_2771_nl : STD_LOGIC;
  SIGNAL or_2769_nl : STD_LOGIC;
  SIGNAL mux_2553_nl : STD_LOGIC;
  SIGNAL mux_2552_nl : STD_LOGIC;
  SIGNAL or_2767_nl : STD_LOGIC;
  SIGNAL nand_139_nl : STD_LOGIC;
  SIGNAL mux_2551_nl : STD_LOGIC;
  SIGNAL or_2763_nl : STD_LOGIC;
  SIGNAL mux_2602_nl : STD_LOGIC;
  SIGNAL or_2822_nl : STD_LOGIC;
  SIGNAL or_2820_nl : STD_LOGIC;
  SIGNAL mux_2601_nl : STD_LOGIC;
  SIGNAL mux_2600_nl : STD_LOGIC;
  SIGNAL or_2817_nl : STD_LOGIC;
  SIGNAL or_2815_nl : STD_LOGIC;
  SIGNAL nand_142_nl : STD_LOGIC;
  SIGNAL mux_2599_nl : STD_LOGIC;
  SIGNAL nor_1608_nl : STD_LOGIC;
  SIGNAL nor_1609_nl : STD_LOGIC;
  SIGNAL and_1542_nl : STD_LOGIC;
  SIGNAL mux_2626_nl : STD_LOGIC;
  SIGNAL mux_2625_nl : STD_LOGIC;
  SIGNAL or_2840_nl : STD_LOGIC;
  SIGNAL mux_2624_nl : STD_LOGIC;
  SIGNAL or_2839_nl : STD_LOGIC;
  SIGNAL mux_2658_nl : STD_LOGIC;
  SIGNAL nand_144_nl : STD_LOGIC;
  SIGNAL mux_2657_nl : STD_LOGIC;
  SIGNAL mux_2656_nl : STD_LOGIC;
  SIGNAL or_2862_nl : STD_LOGIC;
  SIGNAL or_2871_nl : STD_LOGIC;
  SIGNAL and_1528_nl : STD_LOGIC;
  SIGNAL mux_2684_nl : STD_LOGIC;
  SIGNAL mux_2683_nl : STD_LOGIC;
  SIGNAL or_2881_nl : STD_LOGIC;
  SIGNAL mux_2682_nl : STD_LOGIC;
  SIGNAL or_2880_nl : STD_LOGIC;
  SIGNAL or_2901_nl : STD_LOGIC;
  SIGNAL or_2899_nl : STD_LOGIC;
  SIGNAL or_2905_nl : STD_LOGIC;
  SIGNAL or_2903_nl : STD_LOGIC;
  SIGNAL or_2969_nl : STD_LOGIC;
  SIGNAL mux_2774_nl : STD_LOGIC;
  SIGNAL or_2968_nl : STD_LOGIC;
  SIGNAL or_2967_nl : STD_LOGIC;
  SIGNAL mux_2773_nl : STD_LOGIC;
  SIGNAL mux_2772_nl : STD_LOGIC;
  SIGNAL or_2966_nl : STD_LOGIC;
  SIGNAL nand_148_nl : STD_LOGIC;
  SIGNAL mux_2771_nl : STD_LOGIC;
  SIGNAL or_2961_nl : STD_LOGIC;
  SIGNAL mux_2822_nl : STD_LOGIC;
  SIGNAL or_3018_nl : STD_LOGIC;
  SIGNAL or_3017_nl : STD_LOGIC;
  SIGNAL mux_2821_nl : STD_LOGIC;
  SIGNAL mux_2820_nl : STD_LOGIC;
  SIGNAL or_3015_nl : STD_LOGIC;
  SIGNAL or_3014_nl : STD_LOGIC;
  SIGNAL nand_151_nl : STD_LOGIC;
  SIGNAL mux_2819_nl : STD_LOGIC;
  SIGNAL nor_1577_nl : STD_LOGIC;
  SIGNAL nor_1578_nl : STD_LOGIC;
  SIGNAL and_1498_nl : STD_LOGIC;
  SIGNAL mux_2842_nl : STD_LOGIC;
  SIGNAL mux_2841_nl : STD_LOGIC;
  SIGNAL or_3036_nl : STD_LOGIC;
  SIGNAL mux_2840_nl : STD_LOGIC;
  SIGNAL or_3035_nl : STD_LOGIC;
  SIGNAL mux_2878_nl : STD_LOGIC;
  SIGNAL nand_153_nl : STD_LOGIC;
  SIGNAL mux_2877_nl : STD_LOGIC;
  SIGNAL mux_2876_nl : STD_LOGIC;
  SIGNAL or_3059_nl : STD_LOGIC;
  SIGNAL or_3067_nl : STD_LOGIC;
  SIGNAL and_1487_nl : STD_LOGIC;
  SIGNAL mux_2900_nl : STD_LOGIC;
  SIGNAL mux_2899_nl : STD_LOGIC;
  SIGNAL or_3077_nl : STD_LOGIC;
  SIGNAL mux_2898_nl : STD_LOGIC;
  SIGNAL or_3076_nl : STD_LOGIC;
  SIGNAL or_3103_nl : STD_LOGIC;
  SIGNAL or_3101_nl : STD_LOGIC;
  SIGNAL or_3107_nl : STD_LOGIC;
  SIGNAL or_3105_nl : STD_LOGIC;
  SIGNAL or_3176_nl : STD_LOGIC;
  SIGNAL mux_2994_nl : STD_LOGIC;
  SIGNAL or_3175_nl : STD_LOGIC;
  SIGNAL or_3173_nl : STD_LOGIC;
  SIGNAL mux_2993_nl : STD_LOGIC;
  SIGNAL mux_2992_nl : STD_LOGIC;
  SIGNAL or_3171_nl : STD_LOGIC;
  SIGNAL nand_157_nl : STD_LOGIC;
  SIGNAL mux_2991_nl : STD_LOGIC;
  SIGNAL or_3165_nl : STD_LOGIC;
  SIGNAL mux_3042_nl : STD_LOGIC;
  SIGNAL or_3232_nl : STD_LOGIC;
  SIGNAL or_3230_nl : STD_LOGIC;
  SIGNAL mux_3041_nl : STD_LOGIC;
  SIGNAL mux_3040_nl : STD_LOGIC;
  SIGNAL or_3227_nl : STD_LOGIC;
  SIGNAL or_3225_nl : STD_LOGIC;
  SIGNAL nand_160_nl : STD_LOGIC;
  SIGNAL mux_3039_nl : STD_LOGIC;
  SIGNAL nor_1543_nl : STD_LOGIC;
  SIGNAL nor_1544_nl : STD_LOGIC;
  SIGNAL and_1457_nl : STD_LOGIC;
  SIGNAL mux_3066_nl : STD_LOGIC;
  SIGNAL mux_3065_nl : STD_LOGIC;
  SIGNAL or_3253_nl : STD_LOGIC;
  SIGNAL mux_3064_nl : STD_LOGIC;
  SIGNAL or_3252_nl : STD_LOGIC;
  SIGNAL mux_3098_nl : STD_LOGIC;
  SIGNAL nand_162_nl : STD_LOGIC;
  SIGNAL mux_3097_nl : STD_LOGIC;
  SIGNAL mux_3096_nl : STD_LOGIC;
  SIGNAL or_3276_nl : STD_LOGIC;
  SIGNAL or_3287_nl : STD_LOGIC;
  SIGNAL and_1444_nl : STD_LOGIC;
  SIGNAL mux_3124_nl : STD_LOGIC;
  SIGNAL mux_3123_nl : STD_LOGIC;
  SIGNAL or_3299_nl : STD_LOGIC;
  SIGNAL mux_3122_nl : STD_LOGIC;
  SIGNAL or_3298_nl : STD_LOGIC;
  SIGNAL or_3321_nl : STD_LOGIC;
  SIGNAL or_3319_nl : STD_LOGIC;
  SIGNAL or_3325_nl : STD_LOGIC;
  SIGNAL or_3323_nl : STD_LOGIC;
  SIGNAL or_3388_nl : STD_LOGIC;
  SIGNAL mux_3214_nl : STD_LOGIC;
  SIGNAL or_3387_nl : STD_LOGIC;
  SIGNAL or_3386_nl : STD_LOGIC;
  SIGNAL mux_3213_nl : STD_LOGIC;
  SIGNAL mux_3212_nl : STD_LOGIC;
  SIGNAL or_3385_nl : STD_LOGIC;
  SIGNAL nand_166_nl : STD_LOGIC;
  SIGNAL mux_3211_nl : STD_LOGIC;
  SIGNAL or_3380_nl : STD_LOGIC;
  SIGNAL mux_3262_nl : STD_LOGIC;
  SIGNAL or_3437_nl : STD_LOGIC;
  SIGNAL or_3436_nl : STD_LOGIC;
  SIGNAL mux_3261_nl : STD_LOGIC;
  SIGNAL mux_3260_nl : STD_LOGIC;
  SIGNAL or_3434_nl : STD_LOGIC;
  SIGNAL or_3433_nl : STD_LOGIC;
  SIGNAL nand_169_nl : STD_LOGIC;
  SIGNAL mux_3259_nl : STD_LOGIC;
  SIGNAL nor_1509_nl : STD_LOGIC;
  SIGNAL nor_1510_nl : STD_LOGIC;
  SIGNAL and_1413_nl : STD_LOGIC;
  SIGNAL mux_3282_nl : STD_LOGIC;
  SIGNAL mux_3281_nl : STD_LOGIC;
  SIGNAL or_3455_nl : STD_LOGIC;
  SIGNAL mux_3280_nl : STD_LOGIC;
  SIGNAL or_3454_nl : STD_LOGIC;
  SIGNAL mux_3318_nl : STD_LOGIC;
  SIGNAL nand_171_nl : STD_LOGIC;
  SIGNAL mux_3317_nl : STD_LOGIC;
  SIGNAL mux_3316_nl : STD_LOGIC;
  SIGNAL or_3478_nl : STD_LOGIC;
  SIGNAL or_3486_nl : STD_LOGIC;
  SIGNAL and_1400_nl : STD_LOGIC;
  SIGNAL mux_3340_nl : STD_LOGIC;
  SIGNAL mux_3339_nl : STD_LOGIC;
  SIGNAL or_3496_nl : STD_LOGIC;
  SIGNAL mux_3338_nl : STD_LOGIC;
  SIGNAL or_3495_nl : STD_LOGIC;
  SIGNAL or_3522_nl : STD_LOGIC;
  SIGNAL or_3520_nl : STD_LOGIC;
  SIGNAL or_3525_nl : STD_LOGIC;
  SIGNAL or_3524_nl : STD_LOGIC;
  SIGNAL or_3588_nl : STD_LOGIC;
  SIGNAL mux_3434_nl : STD_LOGIC;
  SIGNAL or_3587_nl : STD_LOGIC;
  SIGNAL or_3586_nl : STD_LOGIC;
  SIGNAL mux_3433_nl : STD_LOGIC;
  SIGNAL mux_3432_nl : STD_LOGIC;
  SIGNAL or_4398_nl : STD_LOGIC;
  SIGNAL nand_277_nl : STD_LOGIC;
  SIGNAL mux_3431_nl : STD_LOGIC;
  SIGNAL or_3580_nl : STD_LOGIC;
  SIGNAL mux_3482_nl : STD_LOGIC;
  SIGNAL or_3642_nl : STD_LOGIC;
  SIGNAL or_3640_nl : STD_LOGIC;
  SIGNAL mux_3481_nl : STD_LOGIC;
  SIGNAL mux_3480_nl : STD_LOGIC;
  SIGNAL or_3637_nl : STD_LOGIC;
  SIGNAL or_3635_nl : STD_LOGIC;
  SIGNAL nand_177_nl : STD_LOGIC;
  SIGNAL mux_3479_nl : STD_LOGIC;
  SIGNAL nor_1476_nl : STD_LOGIC;
  SIGNAL nor_1477_nl : STD_LOGIC;
  SIGNAL and_1359_nl : STD_LOGIC;
  SIGNAL mux_3506_nl : STD_LOGIC;
  SIGNAL mux_3505_nl : STD_LOGIC;
  SIGNAL or_3661_nl : STD_LOGIC;
  SIGNAL mux_3504_nl : STD_LOGIC;
  SIGNAL or_3660_nl : STD_LOGIC;
  SIGNAL mux_3538_nl : STD_LOGIC;
  SIGNAL or_4389_nl : STD_LOGIC;
  SIGNAL nand_259_nl : STD_LOGIC;
  SIGNAL mux_3537_nl : STD_LOGIC;
  SIGNAL mux_3536_nl : STD_LOGIC;
  SIGNAL or_3684_nl : STD_LOGIC;
  SIGNAL or_3691_nl : STD_LOGIC;
  SIGNAL and_1341_nl : STD_LOGIC;
  SIGNAL mux_3564_nl : STD_LOGIC;
  SIGNAL mux_3563_nl : STD_LOGIC;
  SIGNAL nand_256_nl : STD_LOGIC;
  SIGNAL mux_3562_nl : STD_LOGIC;
  SIGNAL nand_257_nl : STD_LOGIC;
  SIGNAL mux_3683_nl : STD_LOGIC;
  SIGNAL mux_3682_nl : STD_LOGIC;
  SIGNAL nor_1388_nl : STD_LOGIC;
  SIGNAL nor_1389_nl : STD_LOGIC;
  SIGNAL nor_1390_nl : STD_LOGIC;
  SIGNAL mux_3681_nl : STD_LOGIC;
  SIGNAL or_3846_nl : STD_LOGIC;
  SIGNAL or_3844_nl : STD_LOGIC;
  SIGNAL nor_1391_nl : STD_LOGIC;
  SIGNAL mux_3680_nl : STD_LOGIC;
  SIGNAL or_3841_nl : STD_LOGIC;
  SIGNAL or_3839_nl : STD_LOGIC;
  SIGNAL mux_3798_nl : STD_LOGIC;
  SIGNAL nor_1343_nl : STD_LOGIC;
  SIGNAL nor_1344_nl : STD_LOGIC;
  SIGNAL or_3980_nl : STD_LOGIC;
  SIGNAL or_3979_nl : STD_LOGIC;
  SIGNAL mux_3856_nl : STD_LOGIC;
  SIGNAL mux_3855_nl : STD_LOGIC;
  SIGNAL nor_1326_nl : STD_LOGIC;
  SIGNAL nor_1327_nl : STD_LOGIC;
  SIGNAL nor_1328_nl : STD_LOGIC;
  SIGNAL nor_1323_nl : STD_LOGIC;
  SIGNAL mux_3860_nl : STD_LOGIC;
  SIGNAL nand_197_nl : STD_LOGIC;
  SIGNAL mux_3859_nl : STD_LOGIC;
  SIGNAL mux_3858_nl : STD_LOGIC;
  SIGNAL or_99_nl : STD_LOGIC;
  SIGNAL or_100_nl : STD_LOGIC;
  SIGNAL mux_3857_nl : STD_LOGIC;
  SIGNAL nor_1324_nl : STD_LOGIC;
  SIGNAL nor_1325_nl : STD_LOGIC;
  SIGNAL mux_3875_nl : STD_LOGIC;
  SIGNAL mux_3874_nl : STD_LOGIC;
  SIGNAL nor_1321_nl : STD_LOGIC;
  SIGNAL and_1289_nl : STD_LOGIC;
  SIGNAL nor_1322_nl : STD_LOGIC;
  SIGNAL mux_3898_nl : STD_LOGIC;
  SIGNAL mux_3897_nl : STD_LOGIC;
  SIGNAL mux_3896_nl : STD_LOGIC;
  SIGNAL or_4095_nl : STD_LOGIC;
  SIGNAL mux_3895_nl : STD_LOGIC;
  SIGNAL or_4092_nl : STD_LOGIC;
  SIGNAL mux_3894_nl : STD_LOGIC;
  SIGNAL or_4090_nl : STD_LOGIC;
  SIGNAL mux_3907_nl : STD_LOGIC;
  SIGNAL nor_1312_nl : STD_LOGIC;
  SIGNAL nor_1313_nl : STD_LOGIC;
  SIGNAL mux_3908_nl : STD_LOGIC;
  SIGNAL or_4112_nl : STD_LOGIC;
  SIGNAL nor_1269_nl : STD_LOGIC;
  SIGNAL mux_4056_nl : STD_LOGIC;
  SIGNAL or_4288_nl : STD_LOGIC;
  SIGNAL mux_4055_nl : STD_LOGIC;
  SIGNAL or_4287_nl : STD_LOGIC;
  SIGNAL or_4286_nl : STD_LOGIC;
  SIGNAL and_1275_nl : STD_LOGIC;
  SIGNAL mux_4054_nl : STD_LOGIC;
  SIGNAL nor_1270_nl : STD_LOGIC;
  SIGNAL nor_1271_nl : STD_LOGIC;
  SIGNAL mux_4053_nl : STD_LOGIC;
  SIGNAL mux_73_nl : STD_LOGIC;
  SIGNAL nor_1268_nl : STD_LOGIC;
  SIGNAL mux_4068_nl : STD_LOGIC;
  SIGNAL mux_4067_nl : STD_LOGIC;
  SIGNAL mux_4066_nl : STD_LOGIC;
  SIGNAL mux_4065_nl : STD_LOGIC;
  SIGNAL mux_4064_nl : STD_LOGIC;
  SIGNAL mux_4063_nl : STD_LOGIC;
  SIGNAL mux_4061_nl : STD_LOGIC;
  SIGNAL mux_4060_nl : STD_LOGIC;
  SIGNAL or_4291_nl : STD_LOGIC;
  SIGNAL mux_4059_nl : STD_LOGIC;
  SIGNAL mux_4074_nl : STD_LOGIC;
  SIGNAL mux_4073_nl : STD_LOGIC;
  SIGNAL nor_1339_nl : STD_LOGIC;
  SIGNAL mux_3802_nl : STD_LOGIC;
  SIGNAL or_3962_nl : STD_LOGIC;
  SIGNAL mux_3809_nl : STD_LOGIC;
  SIGNAL or_3971_nl : STD_LOGIC;
  SIGNAL or_3969_nl : STD_LOGIC;
  SIGNAL mux_3800_nl : STD_LOGIC;
  SIGNAL and_1294_nl : STD_LOGIC;
  SIGNAL mux_3799_nl : STD_LOGIC;
  SIGNAL nor_1340_nl : STD_LOGIC;
  SIGNAL nor_1251_nl : STD_LOGIC;
  SIGNAL nor_1342_nl : STD_LOGIC;
  SIGNAL nor_1304_nl : STD_LOGIC;
  SIGNAL nor_1305_nl : STD_LOGIC;
  SIGNAL mux_3918_nl : STD_LOGIC;
  SIGNAL or_4127_nl : STD_LOGIC;
  SIGNAL mux_3917_nl : STD_LOGIC;
  SIGNAL mux_3916_nl : STD_LOGIC;
  SIGNAL or_4125_nl : STD_LOGIC;
  SIGNAL or_4087_nl : STD_LOGIC;
  SIGNAL or_4123_nl : STD_LOGIC;
  SIGNAL mux_3915_nl : STD_LOGIC;
  SIGNAL nor_1299_nl : STD_LOGIC;
  SIGNAL and_1282_nl : STD_LOGIC;
  SIGNAL mux_3949_nl : STD_LOGIC;
  SIGNAL nor_1300_nl : STD_LOGIC;
  SIGNAL mux_3948_nl : STD_LOGIC;
  SIGNAL mux_3947_nl : STD_LOGIC;
  SIGNAL and_1283_nl : STD_LOGIC;
  SIGNAL mux_3946_nl : STD_LOGIC;
  SIGNAL nor_2195_nl : STD_LOGIC;
  SIGNAL nor_1302_nl : STD_LOGIC;
  SIGNAL nor_1298_nl : STD_LOGIC;
  SIGNAL nor_1289_nl : STD_LOGIC;
  SIGNAL mux_3991_nl : STD_LOGIC;
  SIGNAL mux_3990_nl : STD_LOGIC;
  SIGNAL nor_1290_nl : STD_LOGIC;
  SIGNAL nor_1291_nl : STD_LOGIC;
  SIGNAL mux_3989_nl : STD_LOGIC;
  SIGNAL or_4198_nl : STD_LOGIC;
  SIGNAL nor_1292_nl : STD_LOGIC;
  SIGNAL mux_3988_nl : STD_LOGIC;
  SIGNAL or_4195_nl : STD_LOGIC;
  SIGNAL or_4194_nl : STD_LOGIC;
  SIGNAL mux_4008_nl : STD_LOGIC;
  SIGNAL and_1279_nl : STD_LOGIC;
  SIGNAL mux_4007_nl : STD_LOGIC;
  SIGNAL nor_1283_nl : STD_LOGIC;
  SIGNAL nor_1284_nl : STD_LOGIC;
  SIGNAL nor_1285_nl : STD_LOGIC;
  SIGNAL mux_4006_nl : STD_LOGIC;
  SIGNAL nor_1287_nl : STD_LOGIC;
  SIGNAL mux_4005_nl : STD_LOGIC;
  SIGNAL or_4220_nl : STD_LOGIC;
  SIGNAL or_4219_nl : STD_LOGIC;
  SIGNAL mux_4025_nl : STD_LOGIC;
  SIGNAL nor_1278_nl : STD_LOGIC;
  SIGNAL mux_4024_nl : STD_LOGIC;
  SIGNAL mux_4023_nl : STD_LOGIC;
  SIGNAL nor_1279_nl : STD_LOGIC;
  SIGNAL nor_1280_nl : STD_LOGIC;
  SIGNAL nor_1281_nl : STD_LOGIC;
  SIGNAL mux_4022_nl : STD_LOGIC;
  SIGNAL or_4243_nl : STD_LOGIC;
  SIGNAL or_4131_nl : STD_LOGIC;
  SIGNAL nor_1282_nl : STD_LOGIC;
  SIGNAL mux_4043_nl : STD_LOGIC;
  SIGNAL mux_4042_nl : STD_LOGIC;
  SIGNAL and_1277_nl : STD_LOGIC;
  SIGNAL mux_4041_nl : STD_LOGIC;
  SIGNAL nor_1274_nl : STD_LOGIC;
  SIGNAL nor_1275_nl : STD_LOGIC;
  SIGNAL and_1278_nl : STD_LOGIC;
  SIGNAL mux_4040_nl : STD_LOGIC;
  SIGNAL nor_1276_nl : STD_LOGIC;
  SIGNAL nor_1277_nl : STD_LOGIC;
  SIGNAL mux_140_nl : STD_LOGIC;
  SIGNAL or_345_nl : STD_LOGIC;
  SIGNAL mux_192_nl : STD_LOGIC;
  SIGNAL or_412_nl : STD_LOGIC;
  SIGNAL mux_242_nl : STD_LOGIC;
  SIGNAL or_470_nl : STD_LOGIC;
  SIGNAL mux_294_nl : STD_LOGIC;
  SIGNAL or_525_nl : STD_LOGIC;
  SIGNAL mux_358_nl : STD_LOGIC;
  SIGNAL or_581_nl : STD_LOGIC;
  SIGNAL mux_409_nl : STD_LOGIC;
  SIGNAL or_657_nl : STD_LOGIC;
  SIGNAL mux_456_nl : STD_LOGIC;
  SIGNAL or_713_nl : STD_LOGIC;
  SIGNAL mux_505_nl : STD_LOGIC;
  SIGNAL or_766_nl : STD_LOGIC;
  SIGNAL mux_567_nl : STD_LOGIC;
  SIGNAL or_822_nl : STD_LOGIC;
  SIGNAL mux_615_nl : STD_LOGIC;
  SIGNAL or_881_nl : STD_LOGIC;
  SIGNAL mux_662_nl : STD_LOGIC;
  SIGNAL or_933_nl : STD_LOGIC;
  SIGNAL mux_711_nl : STD_LOGIC;
  SIGNAL or_986_nl : STD_LOGIC;
  SIGNAL mux_773_nl : STD_LOGIC;
  SIGNAL or_1038_nl : STD_LOGIC;
  SIGNAL mux_821_nl : STD_LOGIC;
  SIGNAL or_1105_nl : STD_LOGIC;
  SIGNAL mux_868_nl : STD_LOGIC;
  SIGNAL or_1162_nl : STD_LOGIC;
  SIGNAL mux_917_nl : STD_LOGIC;
  SIGNAL or_1212_nl : STD_LOGIC;
  SIGNAL mux_981_nl : STD_LOGIC;
  SIGNAL or_1267_nl : STD_LOGIC;
  SIGNAL mux_980_nl : STD_LOGIC;
  SIGNAL or_1265_nl : STD_LOGIC;
  SIGNAL mux_1032_nl : STD_LOGIC;
  SIGNAL or_1331_nl : STD_LOGIC;
  SIGNAL mux_1031_nl : STD_LOGIC;
  SIGNAL or_1330_nl : STD_LOGIC;
  SIGNAL mux_1082_nl : STD_LOGIC;
  SIGNAL or_1384_nl : STD_LOGIC;
  SIGNAL mux_1081_nl : STD_LOGIC;
  SIGNAL or_1383_nl : STD_LOGIC;
  SIGNAL mux_1134_nl : STD_LOGIC;
  SIGNAL or_1437_nl : STD_LOGIC;
  SIGNAL mux_1133_nl : STD_LOGIC;
  SIGNAL or_1436_nl : STD_LOGIC;
  SIGNAL mux_1198_nl : STD_LOGIC;
  SIGNAL or_1491_nl : STD_LOGIC;
  SIGNAL mux_1197_nl : STD_LOGIC;
  SIGNAL or_1489_nl : STD_LOGIC;
  SIGNAL mux_1250_nl : STD_LOGIC;
  SIGNAL or_1569_nl : STD_LOGIC;
  SIGNAL mux_1249_nl : STD_LOGIC;
  SIGNAL or_1568_nl : STD_LOGIC;
  SIGNAL mux_1300_nl : STD_LOGIC;
  SIGNAL or_1629_nl : STD_LOGIC;
  SIGNAL mux_1299_nl : STD_LOGIC;
  SIGNAL or_1627_nl : STD_LOGIC;
  SIGNAL mux_1352_nl : STD_LOGIC;
  SIGNAL or_1687_nl : STD_LOGIC;
  SIGNAL mux_1351_nl : STD_LOGIC;
  SIGNAL or_1686_nl : STD_LOGIC;
  SIGNAL mux_1416_nl : STD_LOGIC;
  SIGNAL or_1742_nl : STD_LOGIC;
  SIGNAL mux_1415_nl : STD_LOGIC;
  SIGNAL or_1741_nl : STD_LOGIC;
  SIGNAL mux_1467_nl : STD_LOGIC;
  SIGNAL or_1805_nl : STD_LOGIC;
  SIGNAL mux_1466_nl : STD_LOGIC;
  SIGNAL or_1804_nl : STD_LOGIC;
  SIGNAL mux_1517_nl : STD_LOGIC;
  SIGNAL or_1858_nl : STD_LOGIC;
  SIGNAL mux_1516_nl : STD_LOGIC;
  SIGNAL or_1857_nl : STD_LOGIC;
  SIGNAL mux_1569_nl : STD_LOGIC;
  SIGNAL or_1916_nl : STD_LOGIC;
  SIGNAL mux_1568_nl : STD_LOGIC;
  SIGNAL nand_382_nl : STD_LOGIC;
  SIGNAL mux_1633_nl : STD_LOGIC;
  SIGNAL or_1969_nl : STD_LOGIC;
  SIGNAL mux_1632_nl : STD_LOGIC;
  SIGNAL or_1968_nl : STD_LOGIC;
  SIGNAL mux_1684_nl : STD_LOGIC;
  SIGNAL or_2033_nl : STD_LOGIC;
  SIGNAL mux_1683_nl : STD_LOGIC;
  SIGNAL or_2032_nl : STD_LOGIC;
  SIGNAL mux_1734_nl : STD_LOGIC;
  SIGNAL or_2084_nl : STD_LOGIC;
  SIGNAL mux_1733_nl : STD_LOGIC;
  SIGNAL and_2137_nl : STD_LOGIC;
  SIGNAL mux_1782_nl : STD_LOGIC;
  SIGNAL nand_109_nl : STD_LOGIC;
  SIGNAL mux_145_nl : STD_LOGIC;
  SIGNAL nor_2160_nl : STD_LOGIC;
  SIGNAL and_2091_nl : STD_LOGIC;
  SIGNAL or_352_nl : STD_LOGIC;
  SIGNAL mux_144_nl : STD_LOGIC;
  SIGNAL mux_143_nl : STD_LOGIC;
  SIGNAL mux_142_nl : STD_LOGIC;
  SIGNAL and_2092_nl : STD_LOGIC;
  SIGNAL mux_151_nl : STD_LOGIC;
  SIGNAL mux_150_nl : STD_LOGIC;
  SIGNAL mux_149_nl : STD_LOGIC;
  SIGNAL mux_148_nl : STD_LOGIC;
  SIGNAL nor_2158_nl : STD_LOGIC;
  SIGNAL nor_2159_nl : STD_LOGIC;
  SIGNAL mux_147_nl : STD_LOGIC;
  SIGNAL mux_207_nl : STD_LOGIC;
  SIGNAL mux_206_nl : STD_LOGIC;
  SIGNAL mux_205_nl : STD_LOGIC;
  SIGNAL mux_204_nl : STD_LOGIC;
  SIGNAL mux_203_nl : STD_LOGIC;
  SIGNAL or_420_nl : STD_LOGIC;
  SIGNAL mux_201_nl : STD_LOGIC;
  SIGNAL mux_200_nl : STD_LOGIC;
  SIGNAL and_2078_nl : STD_LOGIC;
  SIGNAL and_2079_nl : STD_LOGIC;
  SIGNAL mux_199_nl : STD_LOGIC;
  SIGNAL mux_198_nl : STD_LOGIC;
  SIGNAL or_415_nl : STD_LOGIC;
  SIGNAL mux_197_nl : STD_LOGIC;
  SIGNAL mux_196_nl : STD_LOGIC;
  SIGNAL mux_195_nl : STD_LOGIC;
  SIGNAL mux_258_nl : STD_LOGIC;
  SIGNAL mux_257_nl : STD_LOGIC;
  SIGNAL mux_256_nl : STD_LOGIC;
  SIGNAL or_478_nl : STD_LOGIC;
  SIGNAL mux_255_nl : STD_LOGIC;
  SIGNAL mux_254_nl : STD_LOGIC;
  SIGNAL and_2069_nl : STD_LOGIC;
  SIGNAL and_2070_nl : STD_LOGIC;
  SIGNAL mux_253_nl : STD_LOGIC;
  SIGNAL or_475_nl : STD_LOGIC;
  SIGNAL mux_252_nl : STD_LOGIC;
  SIGNAL mux_251_nl : STD_LOGIC;
  SIGNAL or_474_nl : STD_LOGIC;
  SIGNAL mux_250_nl : STD_LOGIC;
  SIGNAL mux_249_nl : STD_LOGIC;
  SIGNAL mux_248_nl : STD_LOGIC;
  SIGNAL mux_247_nl : STD_LOGIC;
  SIGNAL or_473_nl : STD_LOGIC;
  SIGNAL or_530_nl : STD_LOGIC;
  SIGNAL mux_307_nl : STD_LOGIC;
  SIGNAL mux_306_nl : STD_LOGIC;
  SIGNAL nor_78_nl : STD_LOGIC;
  SIGNAL mux_305_nl : STD_LOGIC;
  SIGNAL mux_312_nl : STD_LOGIC;
  SIGNAL mux_311_nl : STD_LOGIC;
  SIGNAL mux_310_nl : STD_LOGIC;
  SIGNAL mux_304_nl : STD_LOGIC;
  SIGNAL mux_303_nl : STD_LOGIC;
  SIGNAL mux_368_nl : STD_LOGIC;
  SIGNAL mux_367_nl : STD_LOGIC;
  SIGNAL mux_366_nl : STD_LOGIC;
  SIGNAL mux_365_nl : STD_LOGIC;
  SIGNAL nor_2094_nl : STD_LOGIC;
  SIGNAL nor_2095_nl : STD_LOGIC;
  SIGNAL mux_364_nl : STD_LOGIC;
  SIGNAL mux_423_nl : STD_LOGIC;
  SIGNAL mux_422_nl : STD_LOGIC;
  SIGNAL mux_421_nl : STD_LOGIC;
  SIGNAL mux_420_nl : STD_LOGIC;
  SIGNAL mux_419_nl : STD_LOGIC;
  SIGNAL or_663_nl : STD_LOGIC;
  SIGNAL mux_417_nl : STD_LOGIC;
  SIGNAL mux_416_nl : STD_LOGIC;
  SIGNAL and_2036_nl : STD_LOGIC;
  SIGNAL and_2037_nl : STD_LOGIC;
  SIGNAL mux_415_nl : STD_LOGIC;
  SIGNAL mux_414_nl : STD_LOGIC;
  SIGNAL nor_105_nl : STD_LOGIC;
  SIGNAL mux_413_nl : STD_LOGIC;
  SIGNAL mux_412_nl : STD_LOGIC;
  SIGNAL mux_411_nl : STD_LOGIC;
  SIGNAL mux_471_nl : STD_LOGIC;
  SIGNAL mux_470_nl : STD_LOGIC;
  SIGNAL mux_469_nl : STD_LOGIC;
  SIGNAL nor_126_nl : STD_LOGIC;
  SIGNAL mux_468_nl : STD_LOGIC;
  SIGNAL mux_467_nl : STD_LOGIC;
  SIGNAL and_2027_nl : STD_LOGIC;
  SIGNAL and_2028_nl : STD_LOGIC;
  SIGNAL mux_466_nl : STD_LOGIC;
  SIGNAL or_714_nl : STD_LOGIC;
  SIGNAL mux_465_nl : STD_LOGIC;
  SIGNAL mux_464_nl : STD_LOGIC;
  SIGNAL nor_121_nl : STD_LOGIC;
  SIGNAL mux_463_nl : STD_LOGIC;
  SIGNAL mux_462_nl : STD_LOGIC;
  SIGNAL mux_461_nl : STD_LOGIC;
  SIGNAL mux_460_nl : STD_LOGIC;
  SIGNAL nor_120_nl : STD_LOGIC;
  SIGNAL mux_523_nl : STD_LOGIC;
  SIGNAL mux_522_nl : STD_LOGIC;
  SIGNAL mux_520_nl : STD_LOGIC;
  SIGNAL mux_519_nl : STD_LOGIC;
  SIGNAL mux_518_nl : STD_LOGIC;
  SIGNAL mux_577_nl : STD_LOGIC;
  SIGNAL mux_576_nl : STD_LOGIC;
  SIGNAL mux_575_nl : STD_LOGIC;
  SIGNAL mux_574_nl : STD_LOGIC;
  SIGNAL nor_2043_nl : STD_LOGIC;
  SIGNAL nor_2044_nl : STD_LOGIC;
  SIGNAL mux_573_nl : STD_LOGIC;
  SIGNAL mux_629_nl : STD_LOGIC;
  SIGNAL mux_628_nl : STD_LOGIC;
  SIGNAL mux_627_nl : STD_LOGIC;
  SIGNAL mux_626_nl : STD_LOGIC;
  SIGNAL mux_625_nl : STD_LOGIC;
  SIGNAL or_889_nl : STD_LOGIC;
  SIGNAL mux_623_nl : STD_LOGIC;
  SIGNAL mux_622_nl : STD_LOGIC;
  SIGNAL and_1994_nl : STD_LOGIC;
  SIGNAL and_1995_nl : STD_LOGIC;
  SIGNAL mux_621_nl : STD_LOGIC;
  SIGNAL mux_620_nl : STD_LOGIC;
  SIGNAL or_884_nl : STD_LOGIC;
  SIGNAL mux_619_nl : STD_LOGIC;
  SIGNAL mux_618_nl : STD_LOGIC;
  SIGNAL mux_617_nl : STD_LOGIC;
  SIGNAL mux_677_nl : STD_LOGIC;
  SIGNAL mux_676_nl : STD_LOGIC;
  SIGNAL mux_675_nl : STD_LOGIC;
  SIGNAL or_939_nl : STD_LOGIC;
  SIGNAL mux_674_nl : STD_LOGIC;
  SIGNAL mux_673_nl : STD_LOGIC;
  SIGNAL and_1985_nl : STD_LOGIC;
  SIGNAL and_1986_nl : STD_LOGIC;
  SIGNAL mux_672_nl : STD_LOGIC;
  SIGNAL or_936_nl : STD_LOGIC;
  SIGNAL mux_671_nl : STD_LOGIC;
  SIGNAL mux_670_nl : STD_LOGIC;
  SIGNAL or_935_nl : STD_LOGIC;
  SIGNAL mux_669_nl : STD_LOGIC;
  SIGNAL mux_668_nl : STD_LOGIC;
  SIGNAL mux_667_nl : STD_LOGIC;
  SIGNAL mux_666_nl : STD_LOGIC;
  SIGNAL or_934_nl : STD_LOGIC;
  SIGNAL mux_729_nl : STD_LOGIC;
  SIGNAL mux_728_nl : STD_LOGIC;
  SIGNAL mux_727_nl : STD_LOGIC;
  SIGNAL mux_721_nl : STD_LOGIC;
  SIGNAL mux_720_nl : STD_LOGIC;
  SIGNAL mux_783_nl : STD_LOGIC;
  SIGNAL mux_782_nl : STD_LOGIC;
  SIGNAL mux_781_nl : STD_LOGIC;
  SIGNAL mux_780_nl : STD_LOGIC;
  SIGNAL nor_1991_nl : STD_LOGIC;
  SIGNAL nor_1992_nl : STD_LOGIC;
  SIGNAL mux_779_nl : STD_LOGIC;
  SIGNAL mux_835_nl : STD_LOGIC;
  SIGNAL mux_834_nl : STD_LOGIC;
  SIGNAL mux_833_nl : STD_LOGIC;
  SIGNAL mux_832_nl : STD_LOGIC;
  SIGNAL mux_831_nl : STD_LOGIC;
  SIGNAL or_1111_nl : STD_LOGIC;
  SIGNAL mux_829_nl : STD_LOGIC;
  SIGNAL mux_828_nl : STD_LOGIC;
  SIGNAL and_1950_nl : STD_LOGIC;
  SIGNAL and_1951_nl : STD_LOGIC;
  SIGNAL mux_827_nl : STD_LOGIC;
  SIGNAL mux_826_nl : STD_LOGIC;
  SIGNAL and_1952_nl : STD_LOGIC;
  SIGNAL mux_825_nl : STD_LOGIC;
  SIGNAL mux_824_nl : STD_LOGIC;
  SIGNAL mux_823_nl : STD_LOGIC;
  SIGNAL mux_883_nl : STD_LOGIC;
  SIGNAL mux_882_nl : STD_LOGIC;
  SIGNAL mux_881_nl : STD_LOGIC;
  SIGNAL nor_257_nl : STD_LOGIC;
  SIGNAL mux_880_nl : STD_LOGIC;
  SIGNAL mux_879_nl : STD_LOGIC;
  SIGNAL and_1939_nl : STD_LOGIC;
  SIGNAL and_1940_nl : STD_LOGIC;
  SIGNAL mux_878_nl : STD_LOGIC;
  SIGNAL or_1163_nl : STD_LOGIC;
  SIGNAL mux_877_nl : STD_LOGIC;
  SIGNAL mux_876_nl : STD_LOGIC;
  SIGNAL nor_252_nl : STD_LOGIC;
  SIGNAL mux_875_nl : STD_LOGIC;
  SIGNAL mux_874_nl : STD_LOGIC;
  SIGNAL mux_873_nl : STD_LOGIC;
  SIGNAL mux_872_nl : STD_LOGIC;
  SIGNAL and_1941_nl : STD_LOGIC;
  SIGNAL mux_935_nl : STD_LOGIC;
  SIGNAL mux_934_nl : STD_LOGIC;
  SIGNAL mux_932_nl : STD_LOGIC;
  SIGNAL mux_931_nl : STD_LOGIC;
  SIGNAL mux_930_nl : STD_LOGIC;
  SIGNAL mux_991_nl : STD_LOGIC;
  SIGNAL mux_990_nl : STD_LOGIC;
  SIGNAL nor_1940_nl : STD_LOGIC;
  SIGNAL mux_989_nl : STD_LOGIC;
  SIGNAL mux_988_nl : STD_LOGIC;
  SIGNAL nor_1943_nl : STD_LOGIC;
  SIGNAL nor_296_nl : STD_LOGIC;
  SIGNAL mux_987_nl : STD_LOGIC;
  SIGNAL mux_1046_nl : STD_LOGIC;
  SIGNAL mux_1045_nl : STD_LOGIC;
  SIGNAL mux_1044_nl : STD_LOGIC;
  SIGNAL mux_1043_nl : STD_LOGIC;
  SIGNAL mux_1042_nl : STD_LOGIC;
  SIGNAL nor_310_nl : STD_LOGIC;
  SIGNAL mux_1040_nl : STD_LOGIC;
  SIGNAL mux_1039_nl : STD_LOGIC;
  SIGNAL and_1900_nl : STD_LOGIC;
  SIGNAL and_1901_nl : STD_LOGIC;
  SIGNAL mux_1038_nl : STD_LOGIC;
  SIGNAL mux_1037_nl : STD_LOGIC;
  SIGNAL or_1334_nl : STD_LOGIC;
  SIGNAL mux_1036_nl : STD_LOGIC;
  SIGNAL mux_1035_nl : STD_LOGIC;
  SIGNAL mux_1034_nl : STD_LOGIC;
  SIGNAL mux_1097_nl : STD_LOGIC;
  SIGNAL mux_1096_nl : STD_LOGIC;
  SIGNAL mux_1095_nl : STD_LOGIC;
  SIGNAL or_1390_nl : STD_LOGIC;
  SIGNAL mux_1094_nl : STD_LOGIC;
  SIGNAL mux_1093_nl : STD_LOGIC;
  SIGNAL and_1891_nl : STD_LOGIC;
  SIGNAL and_1892_nl : STD_LOGIC;
  SIGNAL mux_1092_nl : STD_LOGIC;
  SIGNAL or_1387_nl : STD_LOGIC;
  SIGNAL mux_1091_nl : STD_LOGIC;
  SIGNAL mux_1090_nl : STD_LOGIC;
  SIGNAL or_1386_nl : STD_LOGIC;
  SIGNAL mux_1089_nl : STD_LOGIC;
  SIGNAL mux_1088_nl : STD_LOGIC;
  SIGNAL mux_1087_nl : STD_LOGIC;
  SIGNAL mux_1086_nl : STD_LOGIC;
  SIGNAL or_1385_nl : STD_LOGIC;
  SIGNAL mux_1152_nl : STD_LOGIC;
  SIGNAL mux_1151_nl : STD_LOGIC;
  SIGNAL mux_1150_nl : STD_LOGIC;
  SIGNAL mux_1144_nl : STD_LOGIC;
  SIGNAL mux_1143_nl : STD_LOGIC;
  SIGNAL mux_1208_nl : STD_LOGIC;
  SIGNAL mux_1207_nl : STD_LOGIC;
  SIGNAL nor_1887_nl : STD_LOGIC;
  SIGNAL mux_1206_nl : STD_LOGIC;
  SIGNAL mux_1205_nl : STD_LOGIC;
  SIGNAL nor_1890_nl : STD_LOGIC;
  SIGNAL nor_361_nl : STD_LOGIC;
  SIGNAL mux_1204_nl : STD_LOGIC;
  SIGNAL mux_1264_nl : STD_LOGIC;
  SIGNAL mux_1263_nl : STD_LOGIC;
  SIGNAL mux_1262_nl : STD_LOGIC;
  SIGNAL mux_1261_nl : STD_LOGIC;
  SIGNAL mux_1260_nl : STD_LOGIC;
  SIGNAL nor_381_nl : STD_LOGIC;
  SIGNAL mux_1258_nl : STD_LOGIC;
  SIGNAL mux_1257_nl : STD_LOGIC;
  SIGNAL and_1856_nl : STD_LOGIC;
  SIGNAL and_1857_nl : STD_LOGIC;
  SIGNAL mux_1256_nl : STD_LOGIC;
  SIGNAL mux_1255_nl : STD_LOGIC;
  SIGNAL and_1858_nl : STD_LOGIC;
  SIGNAL mux_1254_nl : STD_LOGIC;
  SIGNAL mux_1253_nl : STD_LOGIC;
  SIGNAL mux_1252_nl : STD_LOGIC;
  SIGNAL mux_1315_nl : STD_LOGIC;
  SIGNAL mux_1314_nl : STD_LOGIC;
  SIGNAL mux_1313_nl : STD_LOGIC;
  SIGNAL nor_401_nl : STD_LOGIC;
  SIGNAL mux_1312_nl : STD_LOGIC;
  SIGNAL mux_1311_nl : STD_LOGIC;
  SIGNAL and_1845_nl : STD_LOGIC;
  SIGNAL and_1846_nl : STD_LOGIC;
  SIGNAL mux_1310_nl : STD_LOGIC;
  SIGNAL or_1630_nl : STD_LOGIC;
  SIGNAL mux_1309_nl : STD_LOGIC;
  SIGNAL mux_1308_nl : STD_LOGIC;
  SIGNAL nor_396_nl : STD_LOGIC;
  SIGNAL mux_1307_nl : STD_LOGIC;
  SIGNAL mux_1306_nl : STD_LOGIC;
  SIGNAL mux_1305_nl : STD_LOGIC;
  SIGNAL mux_1304_nl : STD_LOGIC;
  SIGNAL and_1847_nl : STD_LOGIC;
  SIGNAL mux_1370_nl : STD_LOGIC;
  SIGNAL mux_1369_nl : STD_LOGIC;
  SIGNAL mux_1367_nl : STD_LOGIC;
  SIGNAL mux_1366_nl : STD_LOGIC;
  SIGNAL mux_1365_nl : STD_LOGIC;
  SIGNAL mux_1426_nl : STD_LOGIC;
  SIGNAL mux_1425_nl : STD_LOGIC;
  SIGNAL nor_1834_nl : STD_LOGIC;
  SIGNAL mux_1424_nl : STD_LOGIC;
  SIGNAL mux_1423_nl : STD_LOGIC;
  SIGNAL nor_1837_nl : STD_LOGIC;
  SIGNAL nor_442_nl : STD_LOGIC;
  SIGNAL mux_1422_nl : STD_LOGIC;
  SIGNAL mux_1481_nl : STD_LOGIC;
  SIGNAL mux_1480_nl : STD_LOGIC;
  SIGNAL mux_1479_nl : STD_LOGIC;
  SIGNAL mux_1478_nl : STD_LOGIC;
  SIGNAL mux_1477_nl : STD_LOGIC;
  SIGNAL nor_460_nl : STD_LOGIC;
  SIGNAL mux_1475_nl : STD_LOGIC;
  SIGNAL mux_1474_nl : STD_LOGIC;
  SIGNAL and_1805_nl : STD_LOGIC;
  SIGNAL and_1806_nl : STD_LOGIC;
  SIGNAL mux_1473_nl : STD_LOGIC;
  SIGNAL mux_1472_nl : STD_LOGIC;
  SIGNAL nand_399_nl : STD_LOGIC;
  SIGNAL mux_1471_nl : STD_LOGIC;
  SIGNAL mux_1470_nl : STD_LOGIC;
  SIGNAL mux_1469_nl : STD_LOGIC;
  SIGNAL mux_1532_nl : STD_LOGIC;
  SIGNAL mux_1531_nl : STD_LOGIC;
  SIGNAL mux_1530_nl : STD_LOGIC;
  SIGNAL or_1864_nl : STD_LOGIC;
  SIGNAL mux_1529_nl : STD_LOGIC;
  SIGNAL mux_1528_nl : STD_LOGIC;
  SIGNAL and_1793_nl : STD_LOGIC;
  SIGNAL and_1794_nl : STD_LOGIC;
  SIGNAL mux_1527_nl : STD_LOGIC;
  SIGNAL or_1861_nl : STD_LOGIC;
  SIGNAL mux_1526_nl : STD_LOGIC;
  SIGNAL mux_1525_nl : STD_LOGIC;
  SIGNAL or_1860_nl : STD_LOGIC;
  SIGNAL mux_1524_nl : STD_LOGIC;
  SIGNAL mux_1523_nl : STD_LOGIC;
  SIGNAL mux_1522_nl : STD_LOGIC;
  SIGNAL mux_1521_nl : STD_LOGIC;
  SIGNAL nand_390_nl : STD_LOGIC;
  SIGNAL mux_1587_nl : STD_LOGIC;
  SIGNAL mux_1586_nl : STD_LOGIC;
  SIGNAL mux_1585_nl : STD_LOGIC;
  SIGNAL mux_1579_nl : STD_LOGIC;
  SIGNAL mux_1578_nl : STD_LOGIC;
  SIGNAL mux_1643_nl : STD_LOGIC;
  SIGNAL mux_1642_nl : STD_LOGIC;
  SIGNAL nor_1783_nl : STD_LOGIC;
  SIGNAL mux_1641_nl : STD_LOGIC;
  SIGNAL mux_1640_nl : STD_LOGIC;
  SIGNAL nor_1786_nl : STD_LOGIC;
  SIGNAL nor_520_nl : STD_LOGIC;
  SIGNAL mux_1639_nl : STD_LOGIC;
  SIGNAL mux_1698_nl : STD_LOGIC;
  SIGNAL mux_1697_nl : STD_LOGIC;
  SIGNAL mux_1696_nl : STD_LOGIC;
  SIGNAL mux_1695_nl : STD_LOGIC;
  SIGNAL mux_1694_nl : STD_LOGIC;
  SIGNAL and_1744_nl : STD_LOGIC;
  SIGNAL mux_1692_nl : STD_LOGIC;
  SIGNAL mux_1691_nl : STD_LOGIC;
  SIGNAL and_1745_nl : STD_LOGIC;
  SIGNAL and_1747_nl : STD_LOGIC;
  SIGNAL mux_1690_nl : STD_LOGIC;
  SIGNAL mux_1689_nl : STD_LOGIC;
  SIGNAL and_1749_nl : STD_LOGIC;
  SIGNAL mux_1688_nl : STD_LOGIC;
  SIGNAL mux_1687_nl : STD_LOGIC;
  SIGNAL mux_1686_nl : STD_LOGIC;
  SIGNAL mux_1749_nl : STD_LOGIC;
  SIGNAL mux_1748_nl : STD_LOGIC;
  SIGNAL mux_1747_nl : STD_LOGIC;
  SIGNAL nor_574_nl : STD_LOGIC;
  SIGNAL mux_1746_nl : STD_LOGIC;
  SIGNAL mux_1745_nl : STD_LOGIC;
  SIGNAL and_1724_nl : STD_LOGIC;
  SIGNAL and_1726_nl : STD_LOGIC;
  SIGNAL mux_1744_nl : STD_LOGIC;
  SIGNAL nand_346_nl : STD_LOGIC;
  SIGNAL mux_1743_nl : STD_LOGIC;
  SIGNAL mux_1742_nl : STD_LOGIC;
  SIGNAL and_1728_nl : STD_LOGIC;
  SIGNAL mux_1741_nl : STD_LOGIC;
  SIGNAL mux_1740_nl : STD_LOGIC;
  SIGNAL mux_1739_nl : STD_LOGIC;
  SIGNAL mux_1738_nl : STD_LOGIC;
  SIGNAL and_1729_nl : STD_LOGIC;
  SIGNAL mux_1800_nl : STD_LOGIC;
  SIGNAL mux_1799_nl : STD_LOGIC;
  SIGNAL mux_1797_nl : STD_LOGIC;
  SIGNAL mux_1796_nl : STD_LOGIC;
  SIGNAL mux_1795_nl : STD_LOGIC;
  SIGNAL and_1680_nl : STD_LOGIC;
  SIGNAL mux_1856_nl : STD_LOGIC;
  SIGNAL nor_630_nl : STD_LOGIC;
  SIGNAL or_2175_nl : STD_LOGIC;
  SIGNAL mux_1846_nl : STD_LOGIC;
  SIGNAL and_1683_nl : STD_LOGIC;
  SIGNAL mux_1859_nl : STD_LOGIC;
  SIGNAL mux_1858_nl : STD_LOGIC;
  SIGNAL mux_1855_nl : STD_LOGIC;
  SIGNAL and_1681_nl : STD_LOGIC;
  SIGNAL and_1682_nl : STD_LOGIC;
  SIGNAL mux_1853_nl : STD_LOGIC;
  SIGNAL mux_1852_nl : STD_LOGIC;
  SIGNAL mux_1851_nl : STD_LOGIC;
  SIGNAL mux_1850_nl : STD_LOGIC;
  SIGNAL or_2169_nl : STD_LOGIC;
  SIGNAL mux_1849_nl : STD_LOGIC;
  SIGNAL or_2168_nl : STD_LOGIC;
  SIGNAL mux_1911_nl : STD_LOGIC;
  SIGNAL nor_1722_nl : STD_LOGIC;
  SIGNAL mux_1910_nl : STD_LOGIC;
  SIGNAL mux_1909_nl : STD_LOGIC;
  SIGNAL mux_1908_nl : STD_LOGIC;
  SIGNAL or_2231_nl : STD_LOGIC;
  SIGNAL or_2230_nl : STD_LOGIC;
  SIGNAL or_2229_nl : STD_LOGIC;
  SIGNAL or_2228_nl : STD_LOGIC;
  SIGNAL nor_1723_nl : STD_LOGIC;
  SIGNAL mux_1907_nl : STD_LOGIC;
  SIGNAL mux_1906_nl : STD_LOGIC;
  SIGNAL mux_1905_nl : STD_LOGIC;
  SIGNAL mux_1904_nl : STD_LOGIC;
  SIGNAL or_2223_nl : STD_LOGIC;
  SIGNAL mux_1952_nl : STD_LOGIC;
  SIGNAL mux_1951_nl : STD_LOGIC;
  SIGNAL or_2281_nl : STD_LOGIC;
  SIGNAL mux_1965_nl : STD_LOGIC;
  SIGNAL mux_1964_nl : STD_LOGIC;
  SIGNAL and_1663_nl : STD_LOGIC;
  SIGNAL mux_1963_nl : STD_LOGIC;
  SIGNAL mux_1962_nl : STD_LOGIC;
  SIGNAL nor_655_nl : STD_LOGIC;
  SIGNAL mux_1969_nl : STD_LOGIC;
  SIGNAL mux_1968_nl : STD_LOGIC;
  SIGNAL mux_1960_nl : STD_LOGIC;
  SIGNAL mux_1959_nl : STD_LOGIC;
  SIGNAL or_2327_nl : STD_LOGIC;
  SIGNAL mux_2026_nl : STD_LOGIC;
  SIGNAL mux_2025_nl : STD_LOGIC;
  SIGNAL mux_2023_nl : STD_LOGIC;
  SIGNAL and_1652_nl : STD_LOGIC;
  SIGNAL mux_2030_nl : STD_LOGIC;
  SIGNAL mux_2029_nl : STD_LOGIC;
  SIGNAL mux_2021_nl : STD_LOGIC;
  SIGNAL mux_2020_nl : STD_LOGIC;
  SIGNAL mux_2089_nl : STD_LOGIC;
  SIGNAL mux_2088_nl : STD_LOGIC;
  SIGNAL mux_2085_nl : STD_LOGIC;
  SIGNAL and_1641_nl : STD_LOGIC;
  SIGNAL and_1642_nl : STD_LOGIC;
  SIGNAL mux_2083_nl : STD_LOGIC;
  SIGNAL mux_2082_nl : STD_LOGIC;
  SIGNAL mux_2081_nl : STD_LOGIC;
  SIGNAL mux_2080_nl : STD_LOGIC;
  SIGNAL or_2373_nl : STD_LOGIC;
  SIGNAL mux_2079_nl : STD_LOGIC;
  SIGNAL or_2372_nl : STD_LOGIC;
  SIGNAL mux_2138_nl : STD_LOGIC;
  SIGNAL nor_1680_nl : STD_LOGIC;
  SIGNAL mux_2137_nl : STD_LOGIC;
  SIGNAL mux_2136_nl : STD_LOGIC;
  SIGNAL mux_2135_nl : STD_LOGIC;
  SIGNAL or_2433_nl : STD_LOGIC;
  SIGNAL or_2432_nl : STD_LOGIC;
  SIGNAL or_2431_nl : STD_LOGIC;
  SIGNAL or_2430_nl : STD_LOGIC;
  SIGNAL nor_1681_nl : STD_LOGIC;
  SIGNAL mux_2134_nl : STD_LOGIC;
  SIGNAL mux_2133_nl : STD_LOGIC;
  SIGNAL mux_2132_nl : STD_LOGIC;
  SIGNAL mux_2131_nl : STD_LOGIC;
  SIGNAL or_2425_nl : STD_LOGIC;
  SIGNAL mux_2194_nl : STD_LOGIC;
  SIGNAL mux_2193_nl : STD_LOGIC;
  SIGNAL mux_2189_nl : STD_LOGIC;
  SIGNAL mux_2188_nl : STD_LOGIC;
  SIGNAL mux_2252_nl : STD_LOGIC;
  SIGNAL mux_2251_nl : STD_LOGIC;
  SIGNAL mux_2247_nl : STD_LOGIC;
  SIGNAL mux_2246_nl : STD_LOGIC;
  SIGNAL mux_2309_nl : STD_LOGIC;
  SIGNAL mux_2308_nl : STD_LOGIC;
  SIGNAL mux_2305_nl : STD_LOGIC;
  SIGNAL and_1600_nl : STD_LOGIC;
  SIGNAL and_1601_nl : STD_LOGIC;
  SIGNAL mux_2303_nl : STD_LOGIC;
  SIGNAL mux_2302_nl : STD_LOGIC;
  SIGNAL mux_2301_nl : STD_LOGIC;
  SIGNAL mux_2300_nl : STD_LOGIC;
  SIGNAL or_2563_nl : STD_LOGIC;
  SIGNAL mux_2299_nl : STD_LOGIC;
  SIGNAL or_2562_nl : STD_LOGIC;
  SIGNAL mux_2358_nl : STD_LOGIC;
  SIGNAL nor_1647_nl : STD_LOGIC;
  SIGNAL mux_2357_nl : STD_LOGIC;
  SIGNAL mux_2356_nl : STD_LOGIC;
  SIGNAL mux_2355_nl : STD_LOGIC;
  SIGNAL or_2614_nl : STD_LOGIC;
  SIGNAL or_2613_nl : STD_LOGIC;
  SIGNAL or_2612_nl : STD_LOGIC;
  SIGNAL or_2611_nl : STD_LOGIC;
  SIGNAL nor_1648_nl : STD_LOGIC;
  SIGNAL mux_2354_nl : STD_LOGIC;
  SIGNAL mux_2353_nl : STD_LOGIC;
  SIGNAL mux_2352_nl : STD_LOGIC;
  SIGNAL mux_2351_nl : STD_LOGIC;
  SIGNAL or_2606_nl : STD_LOGIC;
  SIGNAL mux_2414_nl : STD_LOGIC;
  SIGNAL mux_2413_nl : STD_LOGIC;
  SIGNAL mux_2405_nl : STD_LOGIC;
  SIGNAL mux_2404_nl : STD_LOGIC;
  SIGNAL mux_2472_nl : STD_LOGIC;
  SIGNAL mux_2471_nl : STD_LOGIC;
  SIGNAL mux_2463_nl : STD_LOGIC;
  SIGNAL mux_2462_nl : STD_LOGIC;
  SIGNAL mux_2529_nl : STD_LOGIC;
  SIGNAL mux_2528_nl : STD_LOGIC;
  SIGNAL mux_2525_nl : STD_LOGIC;
  SIGNAL and_1559_nl : STD_LOGIC;
  SIGNAL and_1560_nl : STD_LOGIC;
  SIGNAL mux_2523_nl : STD_LOGIC;
  SIGNAL mux_2522_nl : STD_LOGIC;
  SIGNAL mux_2521_nl : STD_LOGIC;
  SIGNAL mux_2520_nl : STD_LOGIC;
  SIGNAL or_2734_nl : STD_LOGIC;
  SIGNAL mux_2519_nl : STD_LOGIC;
  SIGNAL or_2733_nl : STD_LOGIC;
  SIGNAL mux_2578_nl : STD_LOGIC;
  SIGNAL nor_1614_nl : STD_LOGIC;
  SIGNAL mux_2577_nl : STD_LOGIC;
  SIGNAL mux_2576_nl : STD_LOGIC;
  SIGNAL mux_2575_nl : STD_LOGIC;
  SIGNAL or_2793_nl : STD_LOGIC;
  SIGNAL or_2792_nl : STD_LOGIC;
  SIGNAL or_2791_nl : STD_LOGIC;
  SIGNAL or_2790_nl : STD_LOGIC;
  SIGNAL nor_1615_nl : STD_LOGIC;
  SIGNAL mux_2574_nl : STD_LOGIC;
  SIGNAL mux_2573_nl : STD_LOGIC;
  SIGNAL mux_2572_nl : STD_LOGIC;
  SIGNAL mux_2571_nl : STD_LOGIC;
  SIGNAL or_2785_nl : STD_LOGIC;
  SIGNAL mux_2634_nl : STD_LOGIC;
  SIGNAL mux_2633_nl : STD_LOGIC;
  SIGNAL mux_2629_nl : STD_LOGIC;
  SIGNAL mux_2628_nl : STD_LOGIC;
  SIGNAL mux_2692_nl : STD_LOGIC;
  SIGNAL mux_2691_nl : STD_LOGIC;
  SIGNAL mux_2687_nl : STD_LOGIC;
  SIGNAL mux_2686_nl : STD_LOGIC;
  SIGNAL mux_2749_nl : STD_LOGIC;
  SIGNAL and_1512_nl : STD_LOGIC;
  SIGNAL mux_2748_nl : STD_LOGIC;
  SIGNAL mux_2745_nl : STD_LOGIC;
  SIGNAL and_1514_nl : STD_LOGIC;
  SIGNAL mux_2743_nl : STD_LOGIC;
  SIGNAL mux_2742_nl : STD_LOGIC;
  SIGNAL mux_2741_nl : STD_LOGIC;
  SIGNAL mux_2740_nl : STD_LOGIC;
  SIGNAL or_2934_nl : STD_LOGIC;
  SIGNAL mux_2739_nl : STD_LOGIC;
  SIGNAL or_2933_nl : STD_LOGIC;
  SIGNAL mux_2798_nl : STD_LOGIC;
  SIGNAL nor_1584_nl : STD_LOGIC;
  SIGNAL mux_2797_nl : STD_LOGIC;
  SIGNAL mux_2796_nl : STD_LOGIC;
  SIGNAL mux_2795_nl : STD_LOGIC;
  SIGNAL or_2991_nl : STD_LOGIC;
  SIGNAL or_2990_nl : STD_LOGIC;
  SIGNAL or_2989_nl : STD_LOGIC;
  SIGNAL or_2988_nl : STD_LOGIC;
  SIGNAL nor_1585_nl : STD_LOGIC;
  SIGNAL mux_2794_nl : STD_LOGIC;
  SIGNAL mux_2793_nl : STD_LOGIC;
  SIGNAL mux_2792_nl : STD_LOGIC;
  SIGNAL mux_2791_nl : STD_LOGIC;
  SIGNAL or_2983_nl : STD_LOGIC;
  SIGNAL mux_2854_nl : STD_LOGIC;
  SIGNAL mux_2853_nl : STD_LOGIC;
  SIGNAL mux_2845_nl : STD_LOGIC;
  SIGNAL mux_2844_nl : STD_LOGIC;
  SIGNAL mux_2912_nl : STD_LOGIC;
  SIGNAL mux_2911_nl : STD_LOGIC;
  SIGNAL mux_2903_nl : STD_LOGIC;
  SIGNAL mux_2902_nl : STD_LOGIC;
  SIGNAL mux_2969_nl : STD_LOGIC;
  SIGNAL and_1472_nl : STD_LOGIC;
  SIGNAL mux_2968_nl : STD_LOGIC;
  SIGNAL mux_2965_nl : STD_LOGIC;
  SIGNAL and_1474_nl : STD_LOGIC;
  SIGNAL mux_2963_nl : STD_LOGIC;
  SIGNAL mux_2962_nl : STD_LOGIC;
  SIGNAL mux_2961_nl : STD_LOGIC;
  SIGNAL mux_2960_nl : STD_LOGIC;
  SIGNAL or_3135_nl : STD_LOGIC;
  SIGNAL mux_2959_nl : STD_LOGIC;
  SIGNAL or_3134_nl : STD_LOGIC;
  SIGNAL mux_3018_nl : STD_LOGIC;
  SIGNAL nor_1550_nl : STD_LOGIC;
  SIGNAL mux_3017_nl : STD_LOGIC;
  SIGNAL mux_3016_nl : STD_LOGIC;
  SIGNAL mux_3015_nl : STD_LOGIC;
  SIGNAL or_3200_nl : STD_LOGIC;
  SIGNAL or_3199_nl : STD_LOGIC;
  SIGNAL or_3198_nl : STD_LOGIC;
  SIGNAL or_3197_nl : STD_LOGIC;
  SIGNAL nor_1551_nl : STD_LOGIC;
  SIGNAL mux_3014_nl : STD_LOGIC;
  SIGNAL mux_3013_nl : STD_LOGIC;
  SIGNAL mux_3012_nl : STD_LOGIC;
  SIGNAL mux_3011_nl : STD_LOGIC;
  SIGNAL or_3192_nl : STD_LOGIC;
  SIGNAL mux_3074_nl : STD_LOGIC;
  SIGNAL mux_3073_nl : STD_LOGIC;
  SIGNAL mux_3069_nl : STD_LOGIC;
  SIGNAL mux_3068_nl : STD_LOGIC;
  SIGNAL mux_3132_nl : STD_LOGIC;
  SIGNAL mux_3131_nl : STD_LOGIC;
  SIGNAL mux_3127_nl : STD_LOGIC;
  SIGNAL mux_3126_nl : STD_LOGIC;
  SIGNAL mux_3189_nl : STD_LOGIC;
  SIGNAL and_1428_nl : STD_LOGIC;
  SIGNAL mux_3188_nl : STD_LOGIC;
  SIGNAL mux_3185_nl : STD_LOGIC;
  SIGNAL and_1430_nl : STD_LOGIC;
  SIGNAL mux_3183_nl : STD_LOGIC;
  SIGNAL mux_3182_nl : STD_LOGIC;
  SIGNAL mux_3181_nl : STD_LOGIC;
  SIGNAL mux_3180_nl : STD_LOGIC;
  SIGNAL or_3354_nl : STD_LOGIC;
  SIGNAL mux_3179_nl : STD_LOGIC;
  SIGNAL or_3353_nl : STD_LOGIC;
  SIGNAL mux_3238_nl : STD_LOGIC;
  SIGNAL nor_1516_nl : STD_LOGIC;
  SIGNAL mux_3237_nl : STD_LOGIC;
  SIGNAL mux_3236_nl : STD_LOGIC;
  SIGNAL mux_3235_nl : STD_LOGIC;
  SIGNAL or_3410_nl : STD_LOGIC;
  SIGNAL or_3409_nl : STD_LOGIC;
  SIGNAL or_3408_nl : STD_LOGIC;
  SIGNAL or_3407_nl : STD_LOGIC;
  SIGNAL nor_1517_nl : STD_LOGIC;
  SIGNAL mux_3234_nl : STD_LOGIC;
  SIGNAL mux_3233_nl : STD_LOGIC;
  SIGNAL mux_3232_nl : STD_LOGIC;
  SIGNAL mux_3231_nl : STD_LOGIC;
  SIGNAL or_3402_nl : STD_LOGIC;
  SIGNAL mux_3294_nl : STD_LOGIC;
  SIGNAL mux_3293_nl : STD_LOGIC;
  SIGNAL mux_3285_nl : STD_LOGIC;
  SIGNAL mux_3284_nl : STD_LOGIC;
  SIGNAL mux_3352_nl : STD_LOGIC;
  SIGNAL mux_3351_nl : STD_LOGIC;
  SIGNAL mux_3343_nl : STD_LOGIC;
  SIGNAL mux_3342_nl : STD_LOGIC;
  SIGNAL mux_3409_nl : STD_LOGIC;
  SIGNAL and_1382_nl : STD_LOGIC;
  SIGNAL mux_3408_nl : STD_LOGIC;
  SIGNAL mux_3405_nl : STD_LOGIC;
  SIGNAL and_1384_nl : STD_LOGIC;
  SIGNAL mux_3403_nl : STD_LOGIC;
  SIGNAL mux_3402_nl : STD_LOGIC;
  SIGNAL mux_3401_nl : STD_LOGIC;
  SIGNAL mux_3400_nl : STD_LOGIC;
  SIGNAL or_3551_nl : STD_LOGIC;
  SIGNAL mux_3399_nl : STD_LOGIC;
  SIGNAL or_3550_nl : STD_LOGIC;
  SIGNAL mux_3458_nl : STD_LOGIC;
  SIGNAL nor_1483_nl : STD_LOGIC;
  SIGNAL mux_3457_nl : STD_LOGIC;
  SIGNAL mux_3456_nl : STD_LOGIC;
  SIGNAL mux_3455_nl : STD_LOGIC;
  SIGNAL nand_271_nl : STD_LOGIC;
  SIGNAL nand_272_nl : STD_LOGIC;
  SIGNAL or_3608_nl : STD_LOGIC;
  SIGNAL nand_273_nl : STD_LOGIC;
  SIGNAL nor_1484_nl : STD_LOGIC;
  SIGNAL mux_3454_nl : STD_LOGIC;
  SIGNAL mux_3453_nl : STD_LOGIC;
  SIGNAL mux_3452_nl : STD_LOGIC;
  SIGNAL mux_3451_nl : STD_LOGIC;
  SIGNAL or_3602_nl : STD_LOGIC;
  SIGNAL mux_3514_nl : STD_LOGIC;
  SIGNAL mux_3513_nl : STD_LOGIC;
  SIGNAL mux_3509_nl : STD_LOGIC;
  SIGNAL mux_3508_nl : STD_LOGIC;
  SIGNAL mux_3572_nl : STD_LOGIC;
  SIGNAL mux_3571_nl : STD_LOGIC;
  SIGNAL mux_3567_nl : STD_LOGIC;
  SIGNAL mux_3566_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_168_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_31_nl : STD_LOGIC;
  SIGNAL mux1h_62_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2274_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_191_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_93_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_72_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_230_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_169_nl : STD_LOGIC;
  SIGNAL mux1h_63_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_202_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_264_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_1_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_or_38_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_39_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_167_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_and_149_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_150_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_1_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_311_nl : STD_LOGIC;
  SIGNAL mux_173_nl : STD_LOGIC;
  SIGNAL mux_172_nl : STD_LOGIC;
  SIGNAL or_373_nl : STD_LOGIC;
  SIGNAL mux_166_nl : STD_LOGIC;
  SIGNAL mux_165_nl : STD_LOGIC;
  SIGNAL mux_164_nl : STD_LOGIC;
  SIGNAL mux_161_nl : STD_LOGIC;
  SIGNAL mux_160_nl : STD_LOGIC;
  SIGNAL mux_159_nl : STD_LOGIC;
  SIGNAL mux_158_nl : STD_LOGIC;
  SIGNAL or_370_nl : STD_LOGIC;
  SIGNAL or_368_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_165_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_30_nl : STD_LOGIC;
  SIGNAL mux1h_60_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2275_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_190_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_92_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_71_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_228_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_170_nl : STD_LOGIC;
  SIGNAL mux1h_61_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_205_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_265_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_or_36_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_37_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_166_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_and_143_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_144_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_3_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_312_nl : STD_LOGIC;
  SIGNAL mux_227_nl : STD_LOGIC;
  SIGNAL mux_219_nl : STD_LOGIC;
  SIGNAL mux_218_nl : STD_LOGIC;
  SIGNAL and_2075_nl : STD_LOGIC;
  SIGNAL mux_217_nl : STD_LOGIC;
  SIGNAL mux_216_nl : STD_LOGIC;
  SIGNAL mux_215_nl : STD_LOGIC;
  SIGNAL nor_49_nl : STD_LOGIC;
  SIGNAL or_432_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_162_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_29_nl : STD_LOGIC;
  SIGNAL mux1h_58_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2276_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_189_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_91_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_70_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_226_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_171_nl : STD_LOGIC;
  SIGNAL mux1h_59_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_208_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_266_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_9_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_or_34_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_35_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_165_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_and_137_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_138_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_5_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_313_nl : STD_LOGIC;
  SIGNAL mux_278_nl : STD_LOGIC;
  SIGNAL mux_270_nl : STD_LOGIC;
  SIGNAL mux_269_nl : STD_LOGIC;
  SIGNAL and_2066_nl : STD_LOGIC;
  SIGNAL mux_268_nl : STD_LOGIC;
  SIGNAL mux_267_nl : STD_LOGIC;
  SIGNAL mux_266_nl : STD_LOGIC;
  SIGNAL nor_62_nl : STD_LOGIC;
  SIGNAL or_489_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_159_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_28_nl : STD_LOGIC;
  SIGNAL mux1h_56_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2277_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_188_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_90_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_69_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_224_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_172_nl : STD_LOGIC;
  SIGNAL mux1h_57_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_211_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_267_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_13_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_or_32_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_33_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_164_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_7_and_131_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_132_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_7_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_314_nl : STD_LOGIC;
  SIGNAL mux_332_nl : STD_LOGIC;
  SIGNAL mux_324_nl : STD_LOGIC;
  SIGNAL mux_323_nl : STD_LOGIC;
  SIGNAL and_2052_nl : STD_LOGIC;
  SIGNAL mux_322_nl : STD_LOGIC;
  SIGNAL mux_321_nl : STD_LOGIC;
  SIGNAL mux_320_nl : STD_LOGIC;
  SIGNAL nor_82_nl : STD_LOGIC;
  SIGNAL or_537_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_156_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_27_nl : STD_LOGIC;
  SIGNAL mux1h_54_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2278_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_187_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_89_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_68_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_222_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_173_nl : STD_LOGIC;
  SIGNAL mux1h_55_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_214_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_268_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_9_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_315_nl : STD_LOGIC;
  SIGNAL mux_388_nl : STD_LOGIC;
  SIGNAL mux_387_nl : STD_LOGIC;
  SIGNAL nor_97_nl : STD_LOGIC;
  SIGNAL mux_381_nl : STD_LOGIC;
  SIGNAL mux_380_nl : STD_LOGIC;
  SIGNAL mux_379_nl : STD_LOGIC;
  SIGNAL mux_376_nl : STD_LOGIC;
  SIGNAL mux_375_nl : STD_LOGIC;
  SIGNAL mux_374_nl : STD_LOGIC;
  SIGNAL mux_373_nl : STD_LOGIC;
  SIGNAL or_605_nl : STD_LOGIC;
  SIGNAL or_603_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_153_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_26_nl : STD_LOGIC;
  SIGNAL mux1h_52_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2279_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_186_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_88_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_67_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_220_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_174_nl : STD_LOGIC;
  SIGNAL mux1h_53_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_217_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_269_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_11_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_316_nl : STD_LOGIC;
  SIGNAL mux_441_nl : STD_LOGIC;
  SIGNAL mux_433_nl : STD_LOGIC;
  SIGNAL mux_432_nl : STD_LOGIC;
  SIGNAL and_2033_nl : STD_LOGIC;
  SIGNAL mux_431_nl : STD_LOGIC;
  SIGNAL mux_430_nl : STD_LOGIC;
  SIGNAL mux_429_nl : STD_LOGIC;
  SIGNAL nor_113_nl : STD_LOGIC;
  SIGNAL or_670_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_150_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_25_nl : STD_LOGIC;
  SIGNAL mux1h_50_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2280_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_185_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_87_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_66_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_218_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_175_nl : STD_LOGIC;
  SIGNAL mux1h_51_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_220_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_270_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_13_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_317_nl : STD_LOGIC;
  SIGNAL mux_489_nl : STD_LOGIC;
  SIGNAL mux_488_nl : STD_LOGIC;
  SIGNAL mux_487_nl : STD_LOGIC;
  SIGNAL mux_486_nl : STD_LOGIC;
  SIGNAL mux_481_nl : STD_LOGIC;
  SIGNAL mux_480_nl : STD_LOGIC;
  SIGNAL and_2024_nl : STD_LOGIC;
  SIGNAL mux_479_nl : STD_LOGIC;
  SIGNAL mux_478_nl : STD_LOGIC;
  SIGNAL mux_477_nl : STD_LOGIC;
  SIGNAL nor_129_nl : STD_LOGIC;
  SIGNAL or_724_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_147_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_24_nl : STD_LOGIC;
  SIGNAL mux1h_48_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2281_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_184_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_86_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_65_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_216_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_176_nl : STD_LOGIC;
  SIGNAL mux1h_49_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_223_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_271_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_15_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_318_nl : STD_LOGIC;
  SIGNAL mux_541_nl : STD_LOGIC;
  SIGNAL mux_533_nl : STD_LOGIC;
  SIGNAL mux_532_nl : STD_LOGIC;
  SIGNAL and_2010_nl : STD_LOGIC;
  SIGNAL mux_531_nl : STD_LOGIC;
  SIGNAL mux_530_nl : STD_LOGIC;
  SIGNAL mux_529_nl : STD_LOGIC;
  SIGNAL nor_152_nl : STD_LOGIC;
  SIGNAL or_777_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_144_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_23_nl : STD_LOGIC;
  SIGNAL mux1h_46_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2282_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_183_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_85_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_64_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_214_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_177_nl : STD_LOGIC;
  SIGNAL mux1h_47_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_226_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_272_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_17_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_319_nl : STD_LOGIC;
  SIGNAL mux_597_nl : STD_LOGIC;
  SIGNAL mux_596_nl : STD_LOGIC;
  SIGNAL or_846_nl : STD_LOGIC;
  SIGNAL mux_590_nl : STD_LOGIC;
  SIGNAL mux_589_nl : STD_LOGIC;
  SIGNAL mux_588_nl : STD_LOGIC;
  SIGNAL mux_585_nl : STD_LOGIC;
  SIGNAL mux_584_nl : STD_LOGIC;
  SIGNAL mux_583_nl : STD_LOGIC;
  SIGNAL mux_582_nl : STD_LOGIC;
  SIGNAL or_843_nl : STD_LOGIC;
  SIGNAL or_841_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_141_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_22_nl : STD_LOGIC;
  SIGNAL mux1h_44_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2283_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_182_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_84_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_63_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_212_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_178_nl : STD_LOGIC;
  SIGNAL mux1h_45_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_229_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_273_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_19_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_320_nl : STD_LOGIC;
  SIGNAL mux_647_nl : STD_LOGIC;
  SIGNAL mux_639_nl : STD_LOGIC;
  SIGNAL mux_638_nl : STD_LOGIC;
  SIGNAL and_1991_nl : STD_LOGIC;
  SIGNAL mux_637_nl : STD_LOGIC;
  SIGNAL mux_636_nl : STD_LOGIC;
  SIGNAL mux_635_nl : STD_LOGIC;
  SIGNAL nor_177_nl : STD_LOGIC;
  SIGNAL or_895_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_138_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_21_nl : STD_LOGIC;
  SIGNAL mux1h_42_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2284_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_181_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_83_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_62_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_210_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_179_nl : STD_LOGIC;
  SIGNAL mux1h_43_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_232_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_274_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_21_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_321_nl : STD_LOGIC;
  SIGNAL mux_695_nl : STD_LOGIC;
  SIGNAL mux_687_nl : STD_LOGIC;
  SIGNAL mux_686_nl : STD_LOGIC;
  SIGNAL and_1982_nl : STD_LOGIC;
  SIGNAL mux_685_nl : STD_LOGIC;
  SIGNAL mux_684_nl : STD_LOGIC;
  SIGNAL mux_683_nl : STD_LOGIC;
  SIGNAL nor_190_nl : STD_LOGIC;
  SIGNAL or_944_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_135_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_20_nl : STD_LOGIC;
  SIGNAL mux1h_40_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2285_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_180_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_82_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_61_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_208_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_180_nl : STD_LOGIC;
  SIGNAL mux1h_41_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_235_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_275_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_23_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_322_nl : STD_LOGIC;
  SIGNAL mux_747_nl : STD_LOGIC;
  SIGNAL mux_746_nl : STD_LOGIC;
  SIGNAL mux_745_nl : STD_LOGIC;
  SIGNAL mux_744_nl : STD_LOGIC;
  SIGNAL nor_213_nl : STD_LOGIC;
  SIGNAL mux_739_nl : STD_LOGIC;
  SIGNAL mux_738_nl : STD_LOGIC;
  SIGNAL and_1968_nl : STD_LOGIC;
  SIGNAL mux_737_nl : STD_LOGIC;
  SIGNAL mux_736_nl : STD_LOGIC;
  SIGNAL mux_735_nl : STD_LOGIC;
  SIGNAL nor_210_nl : STD_LOGIC;
  SIGNAL or_995_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_132_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_19_nl : STD_LOGIC;
  SIGNAL mux1h_38_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2286_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_179_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_81_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_60_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_206_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_181_nl : STD_LOGIC;
  SIGNAL mux1h_39_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_238_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_276_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_25_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_323_nl : STD_LOGIC;
  SIGNAL mux_803_nl : STD_LOGIC;
  SIGNAL mux_802_nl : STD_LOGIC;
  SIGNAL nor_226_nl : STD_LOGIC;
  SIGNAL mux_796_nl : STD_LOGIC;
  SIGNAL mux_795_nl : STD_LOGIC;
  SIGNAL mux_794_nl : STD_LOGIC;
  SIGNAL mux_791_nl : STD_LOGIC;
  SIGNAL mux_790_nl : STD_LOGIC;
  SIGNAL mux_789_nl : STD_LOGIC;
  SIGNAL mux_788_nl : STD_LOGIC;
  SIGNAL or_1062_nl : STD_LOGIC;
  SIGNAL or_1060_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_129_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_18_nl : STD_LOGIC;
  SIGNAL mux1h_36_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2287_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_178_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_80_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_59_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_204_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_182_nl : STD_LOGIC;
  SIGNAL mux1h_37_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_241_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_277_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_27_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_324_nl : STD_LOGIC;
  SIGNAL mux_853_nl : STD_LOGIC;
  SIGNAL mux_845_nl : STD_LOGIC;
  SIGNAL mux_844_nl : STD_LOGIC;
  SIGNAL and_1947_nl : STD_LOGIC;
  SIGNAL mux_843_nl : STD_LOGIC;
  SIGNAL mux_842_nl : STD_LOGIC;
  SIGNAL mux_841_nl : STD_LOGIC;
  SIGNAL nor_242_nl : STD_LOGIC;
  SIGNAL or_1119_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_126_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_17_nl : STD_LOGIC;
  SIGNAL mux1h_34_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2288_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_177_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_79_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_58_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_202_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_183_nl : STD_LOGIC;
  SIGNAL mux1h_35_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_244_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_278_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_29_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_325_nl : STD_LOGIC;
  SIGNAL mux_901_nl : STD_LOGIC;
  SIGNAL mux_893_nl : STD_LOGIC;
  SIGNAL mux_892_nl : STD_LOGIC;
  SIGNAL and_1936_nl : STD_LOGIC;
  SIGNAL mux_891_nl : STD_LOGIC;
  SIGNAL mux_890_nl : STD_LOGIC;
  SIGNAL mux_889_nl : STD_LOGIC;
  SIGNAL nor_260_nl : STD_LOGIC;
  SIGNAL or_1173_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_123_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_16_nl : STD_LOGIC;
  SIGNAL mux1h_32_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2289_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_176_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_78_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_57_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_200_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_184_nl : STD_LOGIC;
  SIGNAL mux1h_33_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_247_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_279_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_31_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_326_nl : STD_LOGIC;
  SIGNAL mux_953_nl : STD_LOGIC;
  SIGNAL mux_952_nl : STD_LOGIC;
  SIGNAL mux_951_nl : STD_LOGIC;
  SIGNAL mux_950_nl : STD_LOGIC;
  SIGNAL or_1226_nl : STD_LOGIC;
  SIGNAL mux_945_nl : STD_LOGIC;
  SIGNAL mux_944_nl : STD_LOGIC;
  SIGNAL and_1917_nl : STD_LOGIC;
  SIGNAL mux_943_nl : STD_LOGIC;
  SIGNAL mux_942_nl : STD_LOGIC;
  SIGNAL mux_941_nl : STD_LOGIC;
  SIGNAL and_1918_nl : STD_LOGIC;
  SIGNAL or_1223_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_120_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_15_nl : STD_LOGIC;
  SIGNAL mux1h_30_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2290_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_175_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_77_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_56_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_198_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_185_nl : STD_LOGIC;
  SIGNAL mux1h_31_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_250_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_280_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_33_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_327_nl : STD_LOGIC;
  SIGNAL mux_1011_nl : STD_LOGIC;
  SIGNAL mux_1010_nl : STD_LOGIC;
  SIGNAL or_1289_nl : STD_LOGIC;
  SIGNAL mux_1004_nl : STD_LOGIC;
  SIGNAL mux_1003_nl : STD_LOGIC;
  SIGNAL mux_1002_nl : STD_LOGIC;
  SIGNAL mux_999_nl : STD_LOGIC;
  SIGNAL mux_998_nl : STD_LOGIC;
  SIGNAL mux_997_nl : STD_LOGIC;
  SIGNAL mux_996_nl : STD_LOGIC;
  SIGNAL or_1286_nl : STD_LOGIC;
  SIGNAL or_1284_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_117_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_14_nl : STD_LOGIC;
  SIGNAL mux1h_28_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2291_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_174_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_76_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_55_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_196_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_186_nl : STD_LOGIC;
  SIGNAL mux1h_29_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_253_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_281_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_35_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_328_nl : STD_LOGIC;
  SIGNAL mux_1064_nl : STD_LOGIC;
  SIGNAL mux_1056_nl : STD_LOGIC;
  SIGNAL mux_1055_nl : STD_LOGIC;
  SIGNAL and_1897_nl : STD_LOGIC;
  SIGNAL mux_1054_nl : STD_LOGIC;
  SIGNAL mux_1053_nl : STD_LOGIC;
  SIGNAL mux_1052_nl : STD_LOGIC;
  SIGNAL nor_314_nl : STD_LOGIC;
  SIGNAL or_1341_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_114_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_13_nl : STD_LOGIC;
  SIGNAL mux1h_26_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2292_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_173_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_75_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_54_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_194_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_187_nl : STD_LOGIC;
  SIGNAL mux1h_27_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_256_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_282_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_37_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_329_nl : STD_LOGIC;
  SIGNAL mux_1115_nl : STD_LOGIC;
  SIGNAL mux_1107_nl : STD_LOGIC;
  SIGNAL mux_1106_nl : STD_LOGIC;
  SIGNAL and_1888_nl : STD_LOGIC;
  SIGNAL mux_1105_nl : STD_LOGIC;
  SIGNAL mux_1104_nl : STD_LOGIC;
  SIGNAL mux_1103_nl : STD_LOGIC;
  SIGNAL nor_327_nl : STD_LOGIC;
  SIGNAL or_1394_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_111_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_12_nl : STD_LOGIC;
  SIGNAL mux1h_24_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2293_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_172_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_74_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_53_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_192_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_188_nl : STD_LOGIC;
  SIGNAL mux1h_25_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_259_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_283_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_39_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_330_nl : STD_LOGIC;
  SIGNAL mux_1170_nl : STD_LOGIC;
  SIGNAL mux_1162_nl : STD_LOGIC;
  SIGNAL mux_1161_nl : STD_LOGIC;
  SIGNAL and_1875_nl : STD_LOGIC;
  SIGNAL mux_1160_nl : STD_LOGIC;
  SIGNAL mux_1159_nl : STD_LOGIC;
  SIGNAL mux_1158_nl : STD_LOGIC;
  SIGNAL nor_347_nl : STD_LOGIC;
  SIGNAL or_1446_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_108_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_11_nl : STD_LOGIC;
  SIGNAL mux1h_22_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2294_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_171_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_73_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_52_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_190_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_189_nl : STD_LOGIC;
  SIGNAL mux1h_23_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_262_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_284_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_41_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_331_nl : STD_LOGIC;
  SIGNAL mux_1228_nl : STD_LOGIC;
  SIGNAL mux_1227_nl : STD_LOGIC;
  SIGNAL nor_367_nl : STD_LOGIC;
  SIGNAL mux_1221_nl : STD_LOGIC;
  SIGNAL mux_1220_nl : STD_LOGIC;
  SIGNAL mux_1219_nl : STD_LOGIC;
  SIGNAL mux_1216_nl : STD_LOGIC;
  SIGNAL mux_1215_nl : STD_LOGIC;
  SIGNAL mux_1214_nl : STD_LOGIC;
  SIGNAL mux_1213_nl : STD_LOGIC;
  SIGNAL or_1513_nl : STD_LOGIC;
  SIGNAL or_1511_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_105_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_10_nl : STD_LOGIC;
  SIGNAL mux1h_20_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2295_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_170_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_72_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_51_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_188_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_190_nl : STD_LOGIC;
  SIGNAL mux1h_21_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_265_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_285_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_43_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_332_nl : STD_LOGIC;
  SIGNAL mux_1282_nl : STD_LOGIC;
  SIGNAL mux_1274_nl : STD_LOGIC;
  SIGNAL mux_1273_nl : STD_LOGIC;
  SIGNAL and_1853_nl : STD_LOGIC;
  SIGNAL mux_1272_nl : STD_LOGIC;
  SIGNAL mux_1271_nl : STD_LOGIC;
  SIGNAL mux_1270_nl : STD_LOGIC;
  SIGNAL nor_386_nl : STD_LOGIC;
  SIGNAL or_1579_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_102_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_9_nl : STD_LOGIC;
  SIGNAL mux1h_18_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2296_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_169_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_71_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_50_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_186_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_191_nl : STD_LOGIC;
  SIGNAL mux1h_19_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_268_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_286_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_45_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_333_nl : STD_LOGIC;
  SIGNAL mux_1333_nl : STD_LOGIC;
  SIGNAL mux_1325_nl : STD_LOGIC;
  SIGNAL mux_1324_nl : STD_LOGIC;
  SIGNAL and_1842_nl : STD_LOGIC;
  SIGNAL mux_1323_nl : STD_LOGIC;
  SIGNAL mux_1322_nl : STD_LOGIC;
  SIGNAL mux_1321_nl : STD_LOGIC;
  SIGNAL nor_405_nl : STD_LOGIC;
  SIGNAL or_1639_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_99_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_8_nl : STD_LOGIC;
  SIGNAL mux1h_16_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2297_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_168_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_70_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_49_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_184_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_192_nl : STD_LOGIC;
  SIGNAL mux1h_17_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_271_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_287_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_47_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_334_nl : STD_LOGIC;
  SIGNAL mux_1388_nl : STD_LOGIC;
  SIGNAL mux_1380_nl : STD_LOGIC;
  SIGNAL mux_1379_nl : STD_LOGIC;
  SIGNAL and_1825_nl : STD_LOGIC;
  SIGNAL mux_1378_nl : STD_LOGIC;
  SIGNAL mux_1377_nl : STD_LOGIC;
  SIGNAL mux_1376_nl : STD_LOGIC;
  SIGNAL and_1826_nl : STD_LOGIC;
  SIGNAL or_1698_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_96_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_7_nl : STD_LOGIC;
  SIGNAL mux1h_14_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2298_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_167_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_69_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_48_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_182_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_193_nl : STD_LOGIC;
  SIGNAL mux1h_15_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_274_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_288_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_49_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_335_nl : STD_LOGIC;
  SIGNAL mux_1446_nl : STD_LOGIC;
  SIGNAL mux_1445_nl : STD_LOGIC;
  SIGNAL or_1764_nl : STD_LOGIC;
  SIGNAL mux_1439_nl : STD_LOGIC;
  SIGNAL mux_1438_nl : STD_LOGIC;
  SIGNAL mux_1437_nl : STD_LOGIC;
  SIGNAL mux_1434_nl : STD_LOGIC;
  SIGNAL mux_1433_nl : STD_LOGIC;
  SIGNAL mux_1432_nl : STD_LOGIC;
  SIGNAL mux_1431_nl : STD_LOGIC;
  SIGNAL or_1761_nl : STD_LOGIC;
  SIGNAL or_1759_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_93_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_6_nl : STD_LOGIC;
  SIGNAL mux1h_12_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2299_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_166_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_68_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_47_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_180_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_194_nl : STD_LOGIC;
  SIGNAL mux1h_13_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_277_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_289_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_51_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_336_nl : STD_LOGIC;
  SIGNAL mux_1499_nl : STD_LOGIC;
  SIGNAL mux_1491_nl : STD_LOGIC;
  SIGNAL mux_1490_nl : STD_LOGIC;
  SIGNAL and_1802_nl : STD_LOGIC;
  SIGNAL mux_1489_nl : STD_LOGIC;
  SIGNAL mux_1488_nl : STD_LOGIC;
  SIGNAL mux_1487_nl : STD_LOGIC;
  SIGNAL nor_464_nl : STD_LOGIC;
  SIGNAL or_1815_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_90_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_5_nl : STD_LOGIC;
  SIGNAL mux1h_10_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2300_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_165_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_67_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_46_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_178_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_195_nl : STD_LOGIC;
  SIGNAL mux1h_11_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_280_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_290_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_53_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_337_nl : STD_LOGIC;
  SIGNAL mux_1550_nl : STD_LOGIC;
  SIGNAL mux_1549_nl : STD_LOGIC;
  SIGNAL mux_1548_nl : STD_LOGIC;
  SIGNAL mux_1547_nl : STD_LOGIC;
  SIGNAL nor_483_nl : STD_LOGIC;
  SIGNAL mux_1542_nl : STD_LOGIC;
  SIGNAL mux_1541_nl : STD_LOGIC;
  SIGNAL and_1790_nl : STD_LOGIC;
  SIGNAL mux_1540_nl : STD_LOGIC;
  SIGNAL mux_1539_nl : STD_LOGIC;
  SIGNAL mux_1538_nl : STD_LOGIC;
  SIGNAL nor_480_nl : STD_LOGIC;
  SIGNAL or_1869_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_87_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_4_nl : STD_LOGIC;
  SIGNAL mux1h_8_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2301_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_164_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_66_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_45_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_176_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_196_nl : STD_LOGIC;
  SIGNAL mux1h_9_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_283_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_291_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_55_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_338_nl : STD_LOGIC;
  SIGNAL mux_1605_nl : STD_LOGIC;
  SIGNAL mux_1597_nl : STD_LOGIC;
  SIGNAL mux_1596_nl : STD_LOGIC;
  SIGNAL and_1771_nl : STD_LOGIC;
  SIGNAL mux_1595_nl : STD_LOGIC;
  SIGNAL mux_1594_nl : STD_LOGIC;
  SIGNAL mux_1593_nl : STD_LOGIC;
  SIGNAL and_1772_nl : STD_LOGIC;
  SIGNAL or_1925_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_84_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_3_nl : STD_LOGIC;
  SIGNAL mux1h_6_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2302_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_163_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_65_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_44_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_174_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_197_nl : STD_LOGIC;
  SIGNAL mux1h_7_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_286_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_292_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_57_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_339_nl : STD_LOGIC;
  SIGNAL mux_1663_nl : STD_LOGIC;
  SIGNAL mux_1662_nl : STD_LOGIC;
  SIGNAL and_1759_nl : STD_LOGIC;
  SIGNAL mux_1656_nl : STD_LOGIC;
  SIGNAL mux_1655_nl : STD_LOGIC;
  SIGNAL mux_1654_nl : STD_LOGIC;
  SIGNAL mux_1651_nl : STD_LOGIC;
  SIGNAL mux_1650_nl : STD_LOGIC;
  SIGNAL mux_1649_nl : STD_LOGIC;
  SIGNAL mux_1648_nl : STD_LOGIC;
  SIGNAL or_1991_nl : STD_LOGIC;
  SIGNAL or_1989_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_81_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_2_nl : STD_LOGIC;
  SIGNAL mux1h_4_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2303_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_162_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_64_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_43_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_172_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_198_nl : STD_LOGIC;
  SIGNAL mux1h_5_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_289_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_293_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_59_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_340_nl : STD_LOGIC;
  SIGNAL mux_1716_nl : STD_LOGIC;
  SIGNAL mux_1708_nl : STD_LOGIC;
  SIGNAL mux_1707_nl : STD_LOGIC;
  SIGNAL and_1738_nl : STD_LOGIC;
  SIGNAL mux_1706_nl : STD_LOGIC;
  SIGNAL mux_1705_nl : STD_LOGIC;
  SIGNAL mux_1704_nl : STD_LOGIC;
  SIGNAL and_1739_nl : STD_LOGIC;
  SIGNAL or_2043_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_78_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_1_nl : STD_LOGIC;
  SIGNAL mux1h_2_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2304_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_161_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_63_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_42_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_170_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_199_nl : STD_LOGIC;
  SIGNAL mux1h_3_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_292_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_294_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_61_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_341_nl : STD_LOGIC;
  SIGNAL mux_1767_nl : STD_LOGIC;
  SIGNAL mux_1759_nl : STD_LOGIC;
  SIGNAL mux_1758_nl : STD_LOGIC;
  SIGNAL and_1719_nl : STD_LOGIC;
  SIGNAL mux_1757_nl : STD_LOGIC;
  SIGNAL mux_1756_nl : STD_LOGIC;
  SIGNAL mux_1755_nl : STD_LOGIC;
  SIGNAL and_1720_nl : STD_LOGIC;
  SIGNAL or_2092_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_75_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_mux_nl : STD_LOGIC;
  SIGNAL mux1h_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL nor_2305_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_160_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_41_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_168_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_200_nl : STD_LOGIC;
  SIGNAL mux1h_1_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_7_or_295_nl : STD_LOGIC;
  SIGNAL butterFly_7_mux1h_295_nl : STD_LOGIC;
  SIGNAL butterFly_7_butterFly_7_or_63_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_342_nl : STD_LOGIC;
  SIGNAL mux_1818_nl : STD_LOGIC;
  SIGNAL mux_1810_nl : STD_LOGIC;
  SIGNAL mux_1809_nl : STD_LOGIC;
  SIGNAL and_1689_nl : STD_LOGIC;
  SIGNAL mux_1808_nl : STD_LOGIC;
  SIGNAL mux_1807_nl : STD_LOGIC;
  SIGNAL mux_1806_nl : STD_LOGIC;
  SIGNAL and_1691_nl : STD_LOGIC;
  SIGNAL or_2130_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_70_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_1_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_137_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_134_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_103_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_135_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_298_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_136_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_1_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_and_18_nl : STD_LOGIC;
  SIGNAL butterFly_3_and_19_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_39_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_or_6_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_7_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_343_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_68_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_3_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_139_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_132_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_101_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_134_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_303_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_137_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_and_12_nl : STD_LOGIC;
  SIGNAL butterFly_3_and_13_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_38_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_or_4_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_5_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_1_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_344_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_66_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_5_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_141_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_130_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_99_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_133_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_308_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_138_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_5_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_and_6_nl : STD_LOGIC;
  SIGNAL butterFly_3_and_7_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_37_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_or_2_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_3_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_2_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_345_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_64_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_7_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_143_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_128_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_97_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_132_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_313_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_139_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_and_nl : STD_LOGIC;
  SIGNAL butterFly_3_and_1_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_36_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly_3_or_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_1_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_3_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_346_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_62_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_9_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_145_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_126_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_95_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_131_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_318_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_140_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_4_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_347_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_60_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_11_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_147_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_124_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_93_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_130_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_323_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_141_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_5_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_348_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_58_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_13_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_149_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_122_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_91_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_129_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_328_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_142_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_6_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_349_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_56_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_15_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_151_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_120_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_89_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_128_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_333_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_143_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_7_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_350_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_54_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_17_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_153_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_118_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_87_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_127_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_338_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_144_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_8_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_351_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_52_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_19_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_155_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_116_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_85_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_126_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_343_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_145_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_9_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_352_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_50_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_21_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_157_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_114_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_83_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_125_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_348_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_146_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_10_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_353_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_48_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_23_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_159_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_112_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_81_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_124_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_353_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_147_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_11_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_354_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_46_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_25_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_161_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_110_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_79_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_123_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_358_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_148_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_12_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_355_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_44_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_27_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_163_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_108_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_77_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_122_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_363_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_149_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_13_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_356_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_42_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_29_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_165_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_106_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_75_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_121_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_368_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_150_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_14_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_357_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_40_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_31_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_167_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_104_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_73_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_120_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_373_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_151_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_15_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_358_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_38_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_33_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_169_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_102_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_71_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_119_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_378_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_152_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_16_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_359_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_36_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_35_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_171_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_100_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_69_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_118_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_383_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_153_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_17_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_360_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_34_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_37_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_173_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_98_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_67_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_117_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_388_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_154_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_18_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_361_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_32_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_39_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_175_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_96_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_65_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_116_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_393_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_155_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_19_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_362_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_30_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_41_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_177_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_94_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_63_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_115_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_398_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_156_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_20_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_363_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_28_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_43_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_179_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_92_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_61_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_114_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_403_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_157_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_21_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_364_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_26_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_45_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_181_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_90_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_59_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_113_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_408_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_158_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_22_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_365_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_24_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_47_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_183_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_88_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_57_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_112_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_413_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_159_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_23_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_366_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_22_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_49_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_185_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_86_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_55_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_111_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_418_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_160_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_24_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_367_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_20_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_51_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_187_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_84_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_53_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_110_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_423_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_161_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_25_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_368_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_18_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_53_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_189_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_82_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_51_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_109_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_428_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_162_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_26_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_369_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_16_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_55_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_191_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_80_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_49_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_108_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_433_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_163_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_27_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_370_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_14_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_57_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_193_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_78_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_47_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_107_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_438_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_164_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_28_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_371_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_12_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_59_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_195_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_76_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_45_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_106_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_443_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_165_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_29_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_372_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_10_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_61_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_197_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_74_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_43_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_105_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_448_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_166_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_30_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_373_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_8_nl : STD_LOGIC;
  SIGNAL butterFly_3_butterFly_3_mux_63_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_199_nl : STD_LOGIC;
  SIGNAL butterFly_3_or_72_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_41_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_104_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL butterFly_3_or_453_nl : STD_LOGIC;
  SIGNAL butterFly_3_mux1h_167_nl : STD_LOGIC;
  SIGNAL butterFly_7_or_31_nl : STD_LOGIC;
  SIGNAL butterFly_7_and_374_nl : STD_LOGIC;
  SIGNAL mux_4244_nl : STD_LOGIC;
  SIGNAL nor_2367_nl : STD_LOGIC;
  SIGNAL nor_2368_nl : STD_LOGIC;
  SIGNAL mux_4241_nl : STD_LOGIC;
  SIGNAL nor_2338_nl : STD_LOGIC;
  SIGNAL mux_4240_nl : STD_LOGIC;
  SIGNAL nor_2340_nl : STD_LOGIC;
  SIGNAL S5_COPY_LOOP_for_mux_3_nl : STD_LOGIC;
  SIGNAL S5_COPY_LOOP_for_mux_4_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL acc_2_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_3_if_mux_1_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_if_or_4_nl : STD_LOGIC;
  SIGNAL acc_3_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_sub_3_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL and_2906_nl : STD_LOGIC;
  SIGNAL and_2907_nl : STD_LOGIC;
  SIGNAL modulo_sub_2_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL nor_2436_nl : STD_LOGIC;
  SIGNAL and_2908_nl : STD_LOGIC;
  SIGNAL modulo_sub_1_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL nor_2437_nl : STD_LOGIC;
  SIGNAL and_2909_nl : STD_LOGIC;
  SIGNAL and_2910_nl : STD_LOGIC;
  SIGNAL and_2911_nl : STD_LOGIC;
  SIGNAL modulo_sub_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL and_2912_nl : STD_LOGIC;
  SIGNAL modulo_sub_7_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL and_2914_nl : STD_LOGIC;
  SIGNAL acc_9_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly_18_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL and_2915_nl : STD_LOGIC;
  SIGNAL modulo_sub_5_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL and_2916_nl : STD_LOGIC;
  SIGNAL modulo_sub_12_qif_mux1h_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL nor_2438_nl : STD_LOGIC;
  SIGNAL and_2917_nl : STD_LOGIC;
  SIGNAL operator_20_true_15_acc_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL acc_14_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL acc_16_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_1_if_mult_1_if_mux_1_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_if_or_2_nl : STD_LOGIC;
  SIGNAL S34_OUTER_LOOP_for_mux_3_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL and_2939_nl : STD_LOGIC;
  SIGNAL m_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL m_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_12_z_mul_cmp_a : STD_LOGIC_VECTOR (19 DOWNTO 0);
  SIGNAL mult_12_z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_mul_cmp_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL operator_33_true_1_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_z : STD_LOGIC_VECTOR (3 DOWNTO 0);

  COMPONENT hybrid_core_twiddle_rsci_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsci_oswt : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsci_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_adrb_d : STD_LOGIC_VECTOR (4
      DOWNTO 0);
  SIGNAL hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_qb_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_adrb_d_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_qb_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      xx_rsc_0_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_1_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_2_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_3_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_4_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_5_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_6_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_7_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_8_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_9_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_10_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_11_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_12_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_13_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_14_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_15_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_16_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_17_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_18_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_19_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_20_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_21_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_22_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_23_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_24_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_25_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_26_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_27_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_28_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_29_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_30_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_31_0_cgo_iro : IN STD_LOGIC;
      xx_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_0_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_1_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_2_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_3_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_4_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_5_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_6_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_7_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_8_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_9_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_10_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_11_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_12_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_13_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_14_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_15_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_16_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_17_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_18_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_19_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_20_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_21_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_22_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_23_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_24_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_25_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_26_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_27_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_28_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_29_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_30_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_31_0_cgo_iro : IN STD_LOGIC;
      yy_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
      ensig_cgo_iro : IN STD_LOGIC;
      S34_OUTER_LOOP_for_tf_mul_cmp_z : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      ensig_cgo_iro_1 : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      xx_rsc_0_0_cgo : IN STD_LOGIC;
      xx_rsc_1_0_cgo : IN STD_LOGIC;
      xx_rsc_2_0_cgo : IN STD_LOGIC;
      xx_rsc_3_0_cgo : IN STD_LOGIC;
      xx_rsc_4_0_cgo : IN STD_LOGIC;
      xx_rsc_5_0_cgo : IN STD_LOGIC;
      xx_rsc_6_0_cgo : IN STD_LOGIC;
      xx_rsc_7_0_cgo : IN STD_LOGIC;
      xx_rsc_8_0_cgo : IN STD_LOGIC;
      xx_rsc_9_0_cgo : IN STD_LOGIC;
      xx_rsc_10_0_cgo : IN STD_LOGIC;
      xx_rsc_11_0_cgo : IN STD_LOGIC;
      xx_rsc_12_0_cgo : IN STD_LOGIC;
      xx_rsc_13_0_cgo : IN STD_LOGIC;
      xx_rsc_14_0_cgo : IN STD_LOGIC;
      xx_rsc_15_0_cgo : IN STD_LOGIC;
      xx_rsc_16_0_cgo : IN STD_LOGIC;
      xx_rsc_17_0_cgo : IN STD_LOGIC;
      xx_rsc_18_0_cgo : IN STD_LOGIC;
      xx_rsc_19_0_cgo : IN STD_LOGIC;
      xx_rsc_20_0_cgo : IN STD_LOGIC;
      xx_rsc_21_0_cgo : IN STD_LOGIC;
      xx_rsc_22_0_cgo : IN STD_LOGIC;
      xx_rsc_23_0_cgo : IN STD_LOGIC;
      xx_rsc_24_0_cgo : IN STD_LOGIC;
      xx_rsc_25_0_cgo : IN STD_LOGIC;
      xx_rsc_26_0_cgo : IN STD_LOGIC;
      xx_rsc_27_0_cgo : IN STD_LOGIC;
      xx_rsc_28_0_cgo : IN STD_LOGIC;
      xx_rsc_29_0_cgo : IN STD_LOGIC;
      xx_rsc_30_0_cgo : IN STD_LOGIC;
      xx_rsc_31_0_cgo : IN STD_LOGIC;
      yy_rsc_0_0_cgo : IN STD_LOGIC;
      yy_rsc_1_0_cgo : IN STD_LOGIC;
      yy_rsc_2_0_cgo : IN STD_LOGIC;
      yy_rsc_3_0_cgo : IN STD_LOGIC;
      yy_rsc_4_0_cgo : IN STD_LOGIC;
      yy_rsc_5_0_cgo : IN STD_LOGIC;
      yy_rsc_6_0_cgo : IN STD_LOGIC;
      yy_rsc_7_0_cgo : IN STD_LOGIC;
      yy_rsc_8_0_cgo : IN STD_LOGIC;
      yy_rsc_9_0_cgo : IN STD_LOGIC;
      yy_rsc_10_0_cgo : IN STD_LOGIC;
      yy_rsc_11_0_cgo : IN STD_LOGIC;
      yy_rsc_12_0_cgo : IN STD_LOGIC;
      yy_rsc_13_0_cgo : IN STD_LOGIC;
      yy_rsc_14_0_cgo : IN STD_LOGIC;
      yy_rsc_15_0_cgo : IN STD_LOGIC;
      yy_rsc_16_0_cgo : IN STD_LOGIC;
      yy_rsc_17_0_cgo : IN STD_LOGIC;
      yy_rsc_18_0_cgo : IN STD_LOGIC;
      yy_rsc_19_0_cgo : IN STD_LOGIC;
      yy_rsc_20_0_cgo : IN STD_LOGIC;
      yy_rsc_21_0_cgo : IN STD_LOGIC;
      yy_rsc_22_0_cgo : IN STD_LOGIC;
      yy_rsc_23_0_cgo : IN STD_LOGIC;
      yy_rsc_24_0_cgo : IN STD_LOGIC;
      yy_rsc_25_0_cgo : IN STD_LOGIC;
      yy_rsc_26_0_cgo : IN STD_LOGIC;
      yy_rsc_27_0_cgo : IN STD_LOGIC;
      yy_rsc_28_0_cgo : IN STD_LOGIC;
      yy_rsc_29_0_cgo : IN STD_LOGIC;
      yy_rsc_30_0_cgo : IN STD_LOGIC;
      yy_rsc_31_0_cgo : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      mult_12_z_mul_cmp_en : OUT STD_LOGIC;
      S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      ensig_cgo_1 : IN STD_LOGIC;
      mult_z_mul_cmp_en : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_0_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_4_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_8_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_12_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_16_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_20_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_24_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_xx_rsc_28_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_0_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_1_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_2_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_3_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_4_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_5_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_6_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_7_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_8_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_9_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_10_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_11_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_12_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_13_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_14_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_15_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_16_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_17_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_18_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_19_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_20_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_21_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_22_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_23_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_24_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_25_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_26_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_27_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_28_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_29_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_30_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_yy_rsc_31_0_cgo_iro : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z : STD_LOGIC_VECTOR
      (9 DOWNTO 0);
  SIGNAL hybrid_core_wait_dp_inst_ensig_cgo_iro_1 : STD_LOGIC;
  SIGNAL hybrid_core_wait_dp_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg : STD_LOGIC_VECTOR
      (9 DOWNTO 0);

  COMPONENT hybrid_core_twiddle_h_rsci_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_h_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsci_oswt : IN STD_LOGIC;
      twiddle_h_rsci_adrb_d_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_h_rsci_qb_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsci_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_adrb_d : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_qb_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_adrb_d_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_qb_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_revArr_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      revArr_rsc_s_tdone : IN STD_LOGIC;
      revArr_rsc_tr_write_done : IN STD_LOGIC;
      revArr_rsc_RREADY : IN STD_LOGIC;
      revArr_rsc_RVALID : OUT STD_LOGIC;
      revArr_rsc_RUSER : OUT STD_LOGIC;
      revArr_rsc_RLAST : OUT STD_LOGIC;
      revArr_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      revArr_rsc_RID : OUT STD_LOGIC;
      revArr_rsc_ARREADY : OUT STD_LOGIC;
      revArr_rsc_ARVALID : IN STD_LOGIC;
      revArr_rsc_ARUSER : IN STD_LOGIC;
      revArr_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_ARLOCK : IN STD_LOGIC;
      revArr_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      revArr_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      revArr_rsc_ARID : IN STD_LOGIC;
      revArr_rsc_BREADY : IN STD_LOGIC;
      revArr_rsc_BVALID : OUT STD_LOGIC;
      revArr_rsc_BUSER : OUT STD_LOGIC;
      revArr_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_BID : OUT STD_LOGIC;
      revArr_rsc_WREADY : OUT STD_LOGIC;
      revArr_rsc_WVALID : IN STD_LOGIC;
      revArr_rsc_WUSER : IN STD_LOGIC;
      revArr_rsc_WLAST : IN STD_LOGIC;
      revArr_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      revArr_rsc_AWREADY : OUT STD_LOGIC;
      revArr_rsc_AWVALID : IN STD_LOGIC;
      revArr_rsc_AWUSER : IN STD_LOGIC;
      revArr_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_AWLOCK : IN STD_LOGIC;
      revArr_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      revArr_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      revArr_rsc_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      revArr_rsci_oswt : IN STD_LOGIC;
      revArr_rsci_wen_comp : OUT STD_LOGIC;
      revArr_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      revArr_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (9 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsc_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsci_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_revArr_rsci_inst_revArr_rsci_s_din_mxwt : STD_LOGIC_VECTOR (9
      DOWNTO 0);

  COMPONENT hybrid_core_tw_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      tw_rsc_s_tdone : IN STD_LOGIC;
      tw_rsc_tr_write_done : IN STD_LOGIC;
      tw_rsc_RREADY : IN STD_LOGIC;
      tw_rsc_RVALID : OUT STD_LOGIC;
      tw_rsc_RUSER : OUT STD_LOGIC;
      tw_rsc_RLAST : OUT STD_LOGIC;
      tw_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_rsc_RID : OUT STD_LOGIC;
      tw_rsc_ARREADY : OUT STD_LOGIC;
      tw_rsc_ARVALID : IN STD_LOGIC;
      tw_rsc_ARUSER : IN STD_LOGIC;
      tw_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_ARLOCK : IN STD_LOGIC;
      tw_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_rsc_ARID : IN STD_LOGIC;
      tw_rsc_BREADY : IN STD_LOGIC;
      tw_rsc_BVALID : OUT STD_LOGIC;
      tw_rsc_BUSER : OUT STD_LOGIC;
      tw_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_BID : OUT STD_LOGIC;
      tw_rsc_WREADY : OUT STD_LOGIC;
      tw_rsc_WVALID : IN STD_LOGIC;
      tw_rsc_WUSER : IN STD_LOGIC;
      tw_rsc_WLAST : IN STD_LOGIC;
      tw_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_rsc_AWREADY : OUT STD_LOGIC;
      tw_rsc_AWVALID : IN STD_LOGIC;
      tw_rsc_AWUSER : IN STD_LOGIC;
      tw_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_AWLOCK : IN STD_LOGIC;
      tw_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_rsc_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      tw_rsci_oswt : IN STD_LOGIC;
      tw_rsci_wen_comp : OUT STD_LOGIC;
      tw_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      tw_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsc_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsci_s_raddr_core : STD_LOGIC_VECTOR (9 DOWNTO
      0);
  SIGNAL hybrid_core_tw_rsci_inst_tw_rsci_s_din_mxwt : STD_LOGIC_VECTOR (19 DOWNTO
      0);

  COMPONENT hybrid_core_tw_h_rsci
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      tw_h_rsc_s_tdone : IN STD_LOGIC;
      tw_h_rsc_tr_write_done : IN STD_LOGIC;
      tw_h_rsc_RREADY : IN STD_LOGIC;
      tw_h_rsc_RVALID : OUT STD_LOGIC;
      tw_h_rsc_RUSER : OUT STD_LOGIC;
      tw_h_rsc_RLAST : OUT STD_LOGIC;
      tw_h_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_h_rsc_RID : OUT STD_LOGIC;
      tw_h_rsc_ARREADY : OUT STD_LOGIC;
      tw_h_rsc_ARVALID : IN STD_LOGIC;
      tw_h_rsc_ARUSER : IN STD_LOGIC;
      tw_h_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_ARLOCK : IN STD_LOGIC;
      tw_h_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_h_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_h_rsc_ARID : IN STD_LOGIC;
      tw_h_rsc_BREADY : IN STD_LOGIC;
      tw_h_rsc_BVALID : OUT STD_LOGIC;
      tw_h_rsc_BUSER : OUT STD_LOGIC;
      tw_h_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_BID : OUT STD_LOGIC;
      tw_h_rsc_WREADY : OUT STD_LOGIC;
      tw_h_rsc_WVALID : IN STD_LOGIC;
      tw_h_rsc_WUSER : IN STD_LOGIC;
      tw_h_rsc_WLAST : IN STD_LOGIC;
      tw_h_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_h_rsc_AWREADY : OUT STD_LOGIC;
      tw_h_rsc_AWVALID : IN STD_LOGIC;
      tw_h_rsc_AWUSER : IN STD_LOGIC;
      tw_h_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_AWLOCK : IN STD_LOGIC;
      tw_h_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_h_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_h_rsc_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      tw_h_rsci_oswt : IN STD_LOGIC;
      tw_h_rsci_wen_comp : OUT STD_LOGIC;
      tw_h_rsci_s_raddr_core : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      tw_h_rsci_s_din_mxwt : OUT STD_LOGIC_VECTOR (19 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsci_s_raddr_core : STD_LOGIC_VECTOR (9
      DOWNTO 0);
  SIGNAL hybrid_core_tw_h_rsci_inst_tw_h_rsci_s_din_mxwt : STD_LOGIC_VECTOR (19 DOWNTO
      0);

  COMPONENT hybrid_core_x_rsc_0_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_0_0_s_tdone : IN STD_LOGIC;
      x_rsc_0_0_tr_write_done : IN STD_LOGIC;
      x_rsc_0_0_RREADY : IN STD_LOGIC;
      x_rsc_0_0_RVALID : OUT STD_LOGIC;
      x_rsc_0_0_RUSER : OUT STD_LOGIC;
      x_rsc_0_0_RLAST : OUT STD_LOGIC;
      x_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_RID : OUT STD_LOGIC;
      x_rsc_0_0_ARREADY : OUT STD_LOGIC;
      x_rsc_0_0_ARVALID : IN STD_LOGIC;
      x_rsc_0_0_ARUSER : IN STD_LOGIC;
      x_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_ARLOCK : IN STD_LOGIC;
      x_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_0_0_ARID : IN STD_LOGIC;
      x_rsc_0_0_BREADY : IN STD_LOGIC;
      x_rsc_0_0_BVALID : OUT STD_LOGIC;
      x_rsc_0_0_BUSER : OUT STD_LOGIC;
      x_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_BID : OUT STD_LOGIC;
      x_rsc_0_0_WREADY : OUT STD_LOGIC;
      x_rsc_0_0_WVALID : IN STD_LOGIC;
      x_rsc_0_0_WUSER : IN STD_LOGIC;
      x_rsc_0_0_WLAST : IN STD_LOGIC;
      x_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_AWREADY : OUT STD_LOGIC;
      x_rsc_0_0_AWVALID : IN STD_LOGIC;
      x_rsc_0_0_AWUSER : IN STD_LOGIC;
      x_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_AWLOCK : IN STD_LOGIC;
      x_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_0_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_0_0_i_oswt : IN STD_LOGIC;
      x_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_0_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_0_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_0_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_1_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_1_0_s_tdone : IN STD_LOGIC;
      x_rsc_1_0_tr_write_done : IN STD_LOGIC;
      x_rsc_1_0_RREADY : IN STD_LOGIC;
      x_rsc_1_0_RVALID : OUT STD_LOGIC;
      x_rsc_1_0_RUSER : OUT STD_LOGIC;
      x_rsc_1_0_RLAST : OUT STD_LOGIC;
      x_rsc_1_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_RID : OUT STD_LOGIC;
      x_rsc_1_0_ARREADY : OUT STD_LOGIC;
      x_rsc_1_0_ARVALID : IN STD_LOGIC;
      x_rsc_1_0_ARUSER : IN STD_LOGIC;
      x_rsc_1_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_ARLOCK : IN STD_LOGIC;
      x_rsc_1_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_1_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_1_0_ARID : IN STD_LOGIC;
      x_rsc_1_0_BREADY : IN STD_LOGIC;
      x_rsc_1_0_BVALID : OUT STD_LOGIC;
      x_rsc_1_0_BUSER : OUT STD_LOGIC;
      x_rsc_1_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_BID : OUT STD_LOGIC;
      x_rsc_1_0_WREADY : OUT STD_LOGIC;
      x_rsc_1_0_WVALID : IN STD_LOGIC;
      x_rsc_1_0_WUSER : IN STD_LOGIC;
      x_rsc_1_0_WLAST : IN STD_LOGIC;
      x_rsc_1_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_AWREADY : OUT STD_LOGIC;
      x_rsc_1_0_AWVALID : IN STD_LOGIC;
      x_rsc_1_0_AWUSER : IN STD_LOGIC;
      x_rsc_1_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_AWLOCK : IN STD_LOGIC;
      x_rsc_1_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_1_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_1_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_1_0_i_oswt : IN STD_LOGIC;
      x_rsc_1_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_1_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_1_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_1_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_1_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_1_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_2_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_2_0_s_tdone : IN STD_LOGIC;
      x_rsc_2_0_tr_write_done : IN STD_LOGIC;
      x_rsc_2_0_RREADY : IN STD_LOGIC;
      x_rsc_2_0_RVALID : OUT STD_LOGIC;
      x_rsc_2_0_RUSER : OUT STD_LOGIC;
      x_rsc_2_0_RLAST : OUT STD_LOGIC;
      x_rsc_2_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_RID : OUT STD_LOGIC;
      x_rsc_2_0_ARREADY : OUT STD_LOGIC;
      x_rsc_2_0_ARVALID : IN STD_LOGIC;
      x_rsc_2_0_ARUSER : IN STD_LOGIC;
      x_rsc_2_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_ARLOCK : IN STD_LOGIC;
      x_rsc_2_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_2_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_2_0_ARID : IN STD_LOGIC;
      x_rsc_2_0_BREADY : IN STD_LOGIC;
      x_rsc_2_0_BVALID : OUT STD_LOGIC;
      x_rsc_2_0_BUSER : OUT STD_LOGIC;
      x_rsc_2_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_BID : OUT STD_LOGIC;
      x_rsc_2_0_WREADY : OUT STD_LOGIC;
      x_rsc_2_0_WVALID : IN STD_LOGIC;
      x_rsc_2_0_WUSER : IN STD_LOGIC;
      x_rsc_2_0_WLAST : IN STD_LOGIC;
      x_rsc_2_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_AWREADY : OUT STD_LOGIC;
      x_rsc_2_0_AWVALID : IN STD_LOGIC;
      x_rsc_2_0_AWUSER : IN STD_LOGIC;
      x_rsc_2_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_AWLOCK : IN STD_LOGIC;
      x_rsc_2_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_2_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_2_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_2_0_i_oswt : IN STD_LOGIC;
      x_rsc_2_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_2_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_2_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_2_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_2_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_2_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_3_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_3_0_s_tdone : IN STD_LOGIC;
      x_rsc_3_0_tr_write_done : IN STD_LOGIC;
      x_rsc_3_0_RREADY : IN STD_LOGIC;
      x_rsc_3_0_RVALID : OUT STD_LOGIC;
      x_rsc_3_0_RUSER : OUT STD_LOGIC;
      x_rsc_3_0_RLAST : OUT STD_LOGIC;
      x_rsc_3_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_RID : OUT STD_LOGIC;
      x_rsc_3_0_ARREADY : OUT STD_LOGIC;
      x_rsc_3_0_ARVALID : IN STD_LOGIC;
      x_rsc_3_0_ARUSER : IN STD_LOGIC;
      x_rsc_3_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_ARLOCK : IN STD_LOGIC;
      x_rsc_3_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_3_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_3_0_ARID : IN STD_LOGIC;
      x_rsc_3_0_BREADY : IN STD_LOGIC;
      x_rsc_3_0_BVALID : OUT STD_LOGIC;
      x_rsc_3_0_BUSER : OUT STD_LOGIC;
      x_rsc_3_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_BID : OUT STD_LOGIC;
      x_rsc_3_0_WREADY : OUT STD_LOGIC;
      x_rsc_3_0_WVALID : IN STD_LOGIC;
      x_rsc_3_0_WUSER : IN STD_LOGIC;
      x_rsc_3_0_WLAST : IN STD_LOGIC;
      x_rsc_3_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_AWREADY : OUT STD_LOGIC;
      x_rsc_3_0_AWVALID : IN STD_LOGIC;
      x_rsc_3_0_AWUSER : IN STD_LOGIC;
      x_rsc_3_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_AWLOCK : IN STD_LOGIC;
      x_rsc_3_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_3_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_3_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_3_0_i_oswt : IN STD_LOGIC;
      x_rsc_3_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_3_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_3_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_3_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_3_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_3_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_4_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_4_0_s_tdone : IN STD_LOGIC;
      x_rsc_4_0_tr_write_done : IN STD_LOGIC;
      x_rsc_4_0_RREADY : IN STD_LOGIC;
      x_rsc_4_0_RVALID : OUT STD_LOGIC;
      x_rsc_4_0_RUSER : OUT STD_LOGIC;
      x_rsc_4_0_RLAST : OUT STD_LOGIC;
      x_rsc_4_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_RID : OUT STD_LOGIC;
      x_rsc_4_0_ARREADY : OUT STD_LOGIC;
      x_rsc_4_0_ARVALID : IN STD_LOGIC;
      x_rsc_4_0_ARUSER : IN STD_LOGIC;
      x_rsc_4_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_ARLOCK : IN STD_LOGIC;
      x_rsc_4_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_4_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_4_0_ARID : IN STD_LOGIC;
      x_rsc_4_0_BREADY : IN STD_LOGIC;
      x_rsc_4_0_BVALID : OUT STD_LOGIC;
      x_rsc_4_0_BUSER : OUT STD_LOGIC;
      x_rsc_4_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_BID : OUT STD_LOGIC;
      x_rsc_4_0_WREADY : OUT STD_LOGIC;
      x_rsc_4_0_WVALID : IN STD_LOGIC;
      x_rsc_4_0_WUSER : IN STD_LOGIC;
      x_rsc_4_0_WLAST : IN STD_LOGIC;
      x_rsc_4_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_AWREADY : OUT STD_LOGIC;
      x_rsc_4_0_AWVALID : IN STD_LOGIC;
      x_rsc_4_0_AWUSER : IN STD_LOGIC;
      x_rsc_4_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_AWLOCK : IN STD_LOGIC;
      x_rsc_4_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_4_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_4_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_4_0_i_oswt : IN STD_LOGIC;
      x_rsc_4_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_4_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_4_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_4_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_4_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_4_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_5_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_5_0_s_tdone : IN STD_LOGIC;
      x_rsc_5_0_tr_write_done : IN STD_LOGIC;
      x_rsc_5_0_RREADY : IN STD_LOGIC;
      x_rsc_5_0_RVALID : OUT STD_LOGIC;
      x_rsc_5_0_RUSER : OUT STD_LOGIC;
      x_rsc_5_0_RLAST : OUT STD_LOGIC;
      x_rsc_5_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_RID : OUT STD_LOGIC;
      x_rsc_5_0_ARREADY : OUT STD_LOGIC;
      x_rsc_5_0_ARVALID : IN STD_LOGIC;
      x_rsc_5_0_ARUSER : IN STD_LOGIC;
      x_rsc_5_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_ARLOCK : IN STD_LOGIC;
      x_rsc_5_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_5_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_5_0_ARID : IN STD_LOGIC;
      x_rsc_5_0_BREADY : IN STD_LOGIC;
      x_rsc_5_0_BVALID : OUT STD_LOGIC;
      x_rsc_5_0_BUSER : OUT STD_LOGIC;
      x_rsc_5_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_BID : OUT STD_LOGIC;
      x_rsc_5_0_WREADY : OUT STD_LOGIC;
      x_rsc_5_0_WVALID : IN STD_LOGIC;
      x_rsc_5_0_WUSER : IN STD_LOGIC;
      x_rsc_5_0_WLAST : IN STD_LOGIC;
      x_rsc_5_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_AWREADY : OUT STD_LOGIC;
      x_rsc_5_0_AWVALID : IN STD_LOGIC;
      x_rsc_5_0_AWUSER : IN STD_LOGIC;
      x_rsc_5_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_AWLOCK : IN STD_LOGIC;
      x_rsc_5_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_5_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_5_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_5_0_i_oswt : IN STD_LOGIC;
      x_rsc_5_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_5_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_5_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_5_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_5_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_5_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_6_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_6_0_s_tdone : IN STD_LOGIC;
      x_rsc_6_0_tr_write_done : IN STD_LOGIC;
      x_rsc_6_0_RREADY : IN STD_LOGIC;
      x_rsc_6_0_RVALID : OUT STD_LOGIC;
      x_rsc_6_0_RUSER : OUT STD_LOGIC;
      x_rsc_6_0_RLAST : OUT STD_LOGIC;
      x_rsc_6_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_RID : OUT STD_LOGIC;
      x_rsc_6_0_ARREADY : OUT STD_LOGIC;
      x_rsc_6_0_ARVALID : IN STD_LOGIC;
      x_rsc_6_0_ARUSER : IN STD_LOGIC;
      x_rsc_6_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_ARLOCK : IN STD_LOGIC;
      x_rsc_6_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_6_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_6_0_ARID : IN STD_LOGIC;
      x_rsc_6_0_BREADY : IN STD_LOGIC;
      x_rsc_6_0_BVALID : OUT STD_LOGIC;
      x_rsc_6_0_BUSER : OUT STD_LOGIC;
      x_rsc_6_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_BID : OUT STD_LOGIC;
      x_rsc_6_0_WREADY : OUT STD_LOGIC;
      x_rsc_6_0_WVALID : IN STD_LOGIC;
      x_rsc_6_0_WUSER : IN STD_LOGIC;
      x_rsc_6_0_WLAST : IN STD_LOGIC;
      x_rsc_6_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_AWREADY : OUT STD_LOGIC;
      x_rsc_6_0_AWVALID : IN STD_LOGIC;
      x_rsc_6_0_AWUSER : IN STD_LOGIC;
      x_rsc_6_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_AWLOCK : IN STD_LOGIC;
      x_rsc_6_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_6_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_6_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_6_0_i_oswt : IN STD_LOGIC;
      x_rsc_6_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_6_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_6_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_6_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_6_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_6_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_7_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_7_0_s_tdone : IN STD_LOGIC;
      x_rsc_7_0_tr_write_done : IN STD_LOGIC;
      x_rsc_7_0_RREADY : IN STD_LOGIC;
      x_rsc_7_0_RVALID : OUT STD_LOGIC;
      x_rsc_7_0_RUSER : OUT STD_LOGIC;
      x_rsc_7_0_RLAST : OUT STD_LOGIC;
      x_rsc_7_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_RID : OUT STD_LOGIC;
      x_rsc_7_0_ARREADY : OUT STD_LOGIC;
      x_rsc_7_0_ARVALID : IN STD_LOGIC;
      x_rsc_7_0_ARUSER : IN STD_LOGIC;
      x_rsc_7_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_ARLOCK : IN STD_LOGIC;
      x_rsc_7_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_7_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_7_0_ARID : IN STD_LOGIC;
      x_rsc_7_0_BREADY : IN STD_LOGIC;
      x_rsc_7_0_BVALID : OUT STD_LOGIC;
      x_rsc_7_0_BUSER : OUT STD_LOGIC;
      x_rsc_7_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_BID : OUT STD_LOGIC;
      x_rsc_7_0_WREADY : OUT STD_LOGIC;
      x_rsc_7_0_WVALID : IN STD_LOGIC;
      x_rsc_7_0_WUSER : IN STD_LOGIC;
      x_rsc_7_0_WLAST : IN STD_LOGIC;
      x_rsc_7_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_AWREADY : OUT STD_LOGIC;
      x_rsc_7_0_AWVALID : IN STD_LOGIC;
      x_rsc_7_0_AWUSER : IN STD_LOGIC;
      x_rsc_7_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_AWLOCK : IN STD_LOGIC;
      x_rsc_7_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_7_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_7_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_7_0_i_oswt : IN STD_LOGIC;
      x_rsc_7_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_7_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_7_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_7_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_7_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_7_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_8_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_8_0_s_tdone : IN STD_LOGIC;
      x_rsc_8_0_tr_write_done : IN STD_LOGIC;
      x_rsc_8_0_RREADY : IN STD_LOGIC;
      x_rsc_8_0_RVALID : OUT STD_LOGIC;
      x_rsc_8_0_RUSER : OUT STD_LOGIC;
      x_rsc_8_0_RLAST : OUT STD_LOGIC;
      x_rsc_8_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_RID : OUT STD_LOGIC;
      x_rsc_8_0_ARREADY : OUT STD_LOGIC;
      x_rsc_8_0_ARVALID : IN STD_LOGIC;
      x_rsc_8_0_ARUSER : IN STD_LOGIC;
      x_rsc_8_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_ARLOCK : IN STD_LOGIC;
      x_rsc_8_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_8_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_8_0_ARID : IN STD_LOGIC;
      x_rsc_8_0_BREADY : IN STD_LOGIC;
      x_rsc_8_0_BVALID : OUT STD_LOGIC;
      x_rsc_8_0_BUSER : OUT STD_LOGIC;
      x_rsc_8_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_BID : OUT STD_LOGIC;
      x_rsc_8_0_WREADY : OUT STD_LOGIC;
      x_rsc_8_0_WVALID : IN STD_LOGIC;
      x_rsc_8_0_WUSER : IN STD_LOGIC;
      x_rsc_8_0_WLAST : IN STD_LOGIC;
      x_rsc_8_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_AWREADY : OUT STD_LOGIC;
      x_rsc_8_0_AWVALID : IN STD_LOGIC;
      x_rsc_8_0_AWUSER : IN STD_LOGIC;
      x_rsc_8_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_AWLOCK : IN STD_LOGIC;
      x_rsc_8_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_8_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_8_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_8_0_i_oswt : IN STD_LOGIC;
      x_rsc_8_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_8_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_8_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_8_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_8_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_8_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_9_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_9_0_s_tdone : IN STD_LOGIC;
      x_rsc_9_0_tr_write_done : IN STD_LOGIC;
      x_rsc_9_0_RREADY : IN STD_LOGIC;
      x_rsc_9_0_RVALID : OUT STD_LOGIC;
      x_rsc_9_0_RUSER : OUT STD_LOGIC;
      x_rsc_9_0_RLAST : OUT STD_LOGIC;
      x_rsc_9_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_RID : OUT STD_LOGIC;
      x_rsc_9_0_ARREADY : OUT STD_LOGIC;
      x_rsc_9_0_ARVALID : IN STD_LOGIC;
      x_rsc_9_0_ARUSER : IN STD_LOGIC;
      x_rsc_9_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_ARLOCK : IN STD_LOGIC;
      x_rsc_9_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_9_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_9_0_ARID : IN STD_LOGIC;
      x_rsc_9_0_BREADY : IN STD_LOGIC;
      x_rsc_9_0_BVALID : OUT STD_LOGIC;
      x_rsc_9_0_BUSER : OUT STD_LOGIC;
      x_rsc_9_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_BID : OUT STD_LOGIC;
      x_rsc_9_0_WREADY : OUT STD_LOGIC;
      x_rsc_9_0_WVALID : IN STD_LOGIC;
      x_rsc_9_0_WUSER : IN STD_LOGIC;
      x_rsc_9_0_WLAST : IN STD_LOGIC;
      x_rsc_9_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_AWREADY : OUT STD_LOGIC;
      x_rsc_9_0_AWVALID : IN STD_LOGIC;
      x_rsc_9_0_AWUSER : IN STD_LOGIC;
      x_rsc_9_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_AWLOCK : IN STD_LOGIC;
      x_rsc_9_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_9_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_9_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_9_0_i_oswt : IN STD_LOGIC;
      x_rsc_9_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_9_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_9_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_9_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_9_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_9_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_10_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_10_0_s_tdone : IN STD_LOGIC;
      x_rsc_10_0_tr_write_done : IN STD_LOGIC;
      x_rsc_10_0_RREADY : IN STD_LOGIC;
      x_rsc_10_0_RVALID : OUT STD_LOGIC;
      x_rsc_10_0_RUSER : OUT STD_LOGIC;
      x_rsc_10_0_RLAST : OUT STD_LOGIC;
      x_rsc_10_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_RID : OUT STD_LOGIC;
      x_rsc_10_0_ARREADY : OUT STD_LOGIC;
      x_rsc_10_0_ARVALID : IN STD_LOGIC;
      x_rsc_10_0_ARUSER : IN STD_LOGIC;
      x_rsc_10_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_ARLOCK : IN STD_LOGIC;
      x_rsc_10_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_10_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_10_0_ARID : IN STD_LOGIC;
      x_rsc_10_0_BREADY : IN STD_LOGIC;
      x_rsc_10_0_BVALID : OUT STD_LOGIC;
      x_rsc_10_0_BUSER : OUT STD_LOGIC;
      x_rsc_10_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_BID : OUT STD_LOGIC;
      x_rsc_10_0_WREADY : OUT STD_LOGIC;
      x_rsc_10_0_WVALID : IN STD_LOGIC;
      x_rsc_10_0_WUSER : IN STD_LOGIC;
      x_rsc_10_0_WLAST : IN STD_LOGIC;
      x_rsc_10_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_AWREADY : OUT STD_LOGIC;
      x_rsc_10_0_AWVALID : IN STD_LOGIC;
      x_rsc_10_0_AWUSER : IN STD_LOGIC;
      x_rsc_10_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_AWLOCK : IN STD_LOGIC;
      x_rsc_10_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_10_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_10_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_10_0_i_oswt : IN STD_LOGIC;
      x_rsc_10_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_10_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_10_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_10_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_10_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_10_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_11_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_11_0_s_tdone : IN STD_LOGIC;
      x_rsc_11_0_tr_write_done : IN STD_LOGIC;
      x_rsc_11_0_RREADY : IN STD_LOGIC;
      x_rsc_11_0_RVALID : OUT STD_LOGIC;
      x_rsc_11_0_RUSER : OUT STD_LOGIC;
      x_rsc_11_0_RLAST : OUT STD_LOGIC;
      x_rsc_11_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_RID : OUT STD_LOGIC;
      x_rsc_11_0_ARREADY : OUT STD_LOGIC;
      x_rsc_11_0_ARVALID : IN STD_LOGIC;
      x_rsc_11_0_ARUSER : IN STD_LOGIC;
      x_rsc_11_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_ARLOCK : IN STD_LOGIC;
      x_rsc_11_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_11_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_11_0_ARID : IN STD_LOGIC;
      x_rsc_11_0_BREADY : IN STD_LOGIC;
      x_rsc_11_0_BVALID : OUT STD_LOGIC;
      x_rsc_11_0_BUSER : OUT STD_LOGIC;
      x_rsc_11_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_BID : OUT STD_LOGIC;
      x_rsc_11_0_WREADY : OUT STD_LOGIC;
      x_rsc_11_0_WVALID : IN STD_LOGIC;
      x_rsc_11_0_WUSER : IN STD_LOGIC;
      x_rsc_11_0_WLAST : IN STD_LOGIC;
      x_rsc_11_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_AWREADY : OUT STD_LOGIC;
      x_rsc_11_0_AWVALID : IN STD_LOGIC;
      x_rsc_11_0_AWUSER : IN STD_LOGIC;
      x_rsc_11_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_AWLOCK : IN STD_LOGIC;
      x_rsc_11_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_11_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_11_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_11_0_i_oswt : IN STD_LOGIC;
      x_rsc_11_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_11_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_11_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_11_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_11_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_11_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_12_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_12_0_s_tdone : IN STD_LOGIC;
      x_rsc_12_0_tr_write_done : IN STD_LOGIC;
      x_rsc_12_0_RREADY : IN STD_LOGIC;
      x_rsc_12_0_RVALID : OUT STD_LOGIC;
      x_rsc_12_0_RUSER : OUT STD_LOGIC;
      x_rsc_12_0_RLAST : OUT STD_LOGIC;
      x_rsc_12_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_RID : OUT STD_LOGIC;
      x_rsc_12_0_ARREADY : OUT STD_LOGIC;
      x_rsc_12_0_ARVALID : IN STD_LOGIC;
      x_rsc_12_0_ARUSER : IN STD_LOGIC;
      x_rsc_12_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_ARLOCK : IN STD_LOGIC;
      x_rsc_12_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_12_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_12_0_ARID : IN STD_LOGIC;
      x_rsc_12_0_BREADY : IN STD_LOGIC;
      x_rsc_12_0_BVALID : OUT STD_LOGIC;
      x_rsc_12_0_BUSER : OUT STD_LOGIC;
      x_rsc_12_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_BID : OUT STD_LOGIC;
      x_rsc_12_0_WREADY : OUT STD_LOGIC;
      x_rsc_12_0_WVALID : IN STD_LOGIC;
      x_rsc_12_0_WUSER : IN STD_LOGIC;
      x_rsc_12_0_WLAST : IN STD_LOGIC;
      x_rsc_12_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_AWREADY : OUT STD_LOGIC;
      x_rsc_12_0_AWVALID : IN STD_LOGIC;
      x_rsc_12_0_AWUSER : IN STD_LOGIC;
      x_rsc_12_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_AWLOCK : IN STD_LOGIC;
      x_rsc_12_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_12_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_12_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_12_0_i_oswt : IN STD_LOGIC;
      x_rsc_12_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_12_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_12_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_12_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_12_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_12_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_13_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_13_0_s_tdone : IN STD_LOGIC;
      x_rsc_13_0_tr_write_done : IN STD_LOGIC;
      x_rsc_13_0_RREADY : IN STD_LOGIC;
      x_rsc_13_0_RVALID : OUT STD_LOGIC;
      x_rsc_13_0_RUSER : OUT STD_LOGIC;
      x_rsc_13_0_RLAST : OUT STD_LOGIC;
      x_rsc_13_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_RID : OUT STD_LOGIC;
      x_rsc_13_0_ARREADY : OUT STD_LOGIC;
      x_rsc_13_0_ARVALID : IN STD_LOGIC;
      x_rsc_13_0_ARUSER : IN STD_LOGIC;
      x_rsc_13_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_ARLOCK : IN STD_LOGIC;
      x_rsc_13_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_13_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_13_0_ARID : IN STD_LOGIC;
      x_rsc_13_0_BREADY : IN STD_LOGIC;
      x_rsc_13_0_BVALID : OUT STD_LOGIC;
      x_rsc_13_0_BUSER : OUT STD_LOGIC;
      x_rsc_13_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_BID : OUT STD_LOGIC;
      x_rsc_13_0_WREADY : OUT STD_LOGIC;
      x_rsc_13_0_WVALID : IN STD_LOGIC;
      x_rsc_13_0_WUSER : IN STD_LOGIC;
      x_rsc_13_0_WLAST : IN STD_LOGIC;
      x_rsc_13_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_AWREADY : OUT STD_LOGIC;
      x_rsc_13_0_AWVALID : IN STD_LOGIC;
      x_rsc_13_0_AWUSER : IN STD_LOGIC;
      x_rsc_13_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_AWLOCK : IN STD_LOGIC;
      x_rsc_13_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_13_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_13_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_13_0_i_oswt : IN STD_LOGIC;
      x_rsc_13_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_13_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_13_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_13_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_13_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_13_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_14_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_14_0_s_tdone : IN STD_LOGIC;
      x_rsc_14_0_tr_write_done : IN STD_LOGIC;
      x_rsc_14_0_RREADY : IN STD_LOGIC;
      x_rsc_14_0_RVALID : OUT STD_LOGIC;
      x_rsc_14_0_RUSER : OUT STD_LOGIC;
      x_rsc_14_0_RLAST : OUT STD_LOGIC;
      x_rsc_14_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_RID : OUT STD_LOGIC;
      x_rsc_14_0_ARREADY : OUT STD_LOGIC;
      x_rsc_14_0_ARVALID : IN STD_LOGIC;
      x_rsc_14_0_ARUSER : IN STD_LOGIC;
      x_rsc_14_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_ARLOCK : IN STD_LOGIC;
      x_rsc_14_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_14_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_14_0_ARID : IN STD_LOGIC;
      x_rsc_14_0_BREADY : IN STD_LOGIC;
      x_rsc_14_0_BVALID : OUT STD_LOGIC;
      x_rsc_14_0_BUSER : OUT STD_LOGIC;
      x_rsc_14_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_BID : OUT STD_LOGIC;
      x_rsc_14_0_WREADY : OUT STD_LOGIC;
      x_rsc_14_0_WVALID : IN STD_LOGIC;
      x_rsc_14_0_WUSER : IN STD_LOGIC;
      x_rsc_14_0_WLAST : IN STD_LOGIC;
      x_rsc_14_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_AWREADY : OUT STD_LOGIC;
      x_rsc_14_0_AWVALID : IN STD_LOGIC;
      x_rsc_14_0_AWUSER : IN STD_LOGIC;
      x_rsc_14_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_AWLOCK : IN STD_LOGIC;
      x_rsc_14_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_14_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_14_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_14_0_i_oswt : IN STD_LOGIC;
      x_rsc_14_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_14_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_14_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_14_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_14_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_14_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_15_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_15_0_s_tdone : IN STD_LOGIC;
      x_rsc_15_0_tr_write_done : IN STD_LOGIC;
      x_rsc_15_0_RREADY : IN STD_LOGIC;
      x_rsc_15_0_RVALID : OUT STD_LOGIC;
      x_rsc_15_0_RUSER : OUT STD_LOGIC;
      x_rsc_15_0_RLAST : OUT STD_LOGIC;
      x_rsc_15_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_RID : OUT STD_LOGIC;
      x_rsc_15_0_ARREADY : OUT STD_LOGIC;
      x_rsc_15_0_ARVALID : IN STD_LOGIC;
      x_rsc_15_0_ARUSER : IN STD_LOGIC;
      x_rsc_15_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_ARLOCK : IN STD_LOGIC;
      x_rsc_15_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_15_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_15_0_ARID : IN STD_LOGIC;
      x_rsc_15_0_BREADY : IN STD_LOGIC;
      x_rsc_15_0_BVALID : OUT STD_LOGIC;
      x_rsc_15_0_BUSER : OUT STD_LOGIC;
      x_rsc_15_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_BID : OUT STD_LOGIC;
      x_rsc_15_0_WREADY : OUT STD_LOGIC;
      x_rsc_15_0_WVALID : IN STD_LOGIC;
      x_rsc_15_0_WUSER : IN STD_LOGIC;
      x_rsc_15_0_WLAST : IN STD_LOGIC;
      x_rsc_15_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_AWREADY : OUT STD_LOGIC;
      x_rsc_15_0_AWVALID : IN STD_LOGIC;
      x_rsc_15_0_AWUSER : IN STD_LOGIC;
      x_rsc_15_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_AWLOCK : IN STD_LOGIC;
      x_rsc_15_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_15_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_15_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_15_0_i_oswt : IN STD_LOGIC;
      x_rsc_15_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_15_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_15_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_15_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_15_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_15_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_16_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_16_0_s_tdone : IN STD_LOGIC;
      x_rsc_16_0_tr_write_done : IN STD_LOGIC;
      x_rsc_16_0_RREADY : IN STD_LOGIC;
      x_rsc_16_0_RVALID : OUT STD_LOGIC;
      x_rsc_16_0_RUSER : OUT STD_LOGIC;
      x_rsc_16_0_RLAST : OUT STD_LOGIC;
      x_rsc_16_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_RID : OUT STD_LOGIC;
      x_rsc_16_0_ARREADY : OUT STD_LOGIC;
      x_rsc_16_0_ARVALID : IN STD_LOGIC;
      x_rsc_16_0_ARUSER : IN STD_LOGIC;
      x_rsc_16_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_ARLOCK : IN STD_LOGIC;
      x_rsc_16_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_16_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_16_0_ARID : IN STD_LOGIC;
      x_rsc_16_0_BREADY : IN STD_LOGIC;
      x_rsc_16_0_BVALID : OUT STD_LOGIC;
      x_rsc_16_0_BUSER : OUT STD_LOGIC;
      x_rsc_16_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_BID : OUT STD_LOGIC;
      x_rsc_16_0_WREADY : OUT STD_LOGIC;
      x_rsc_16_0_WVALID : IN STD_LOGIC;
      x_rsc_16_0_WUSER : IN STD_LOGIC;
      x_rsc_16_0_WLAST : IN STD_LOGIC;
      x_rsc_16_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_AWREADY : OUT STD_LOGIC;
      x_rsc_16_0_AWVALID : IN STD_LOGIC;
      x_rsc_16_0_AWUSER : IN STD_LOGIC;
      x_rsc_16_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_AWLOCK : IN STD_LOGIC;
      x_rsc_16_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_16_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_16_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_16_0_i_oswt : IN STD_LOGIC;
      x_rsc_16_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_16_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_16_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_16_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_16_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_16_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_17_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_17_0_s_tdone : IN STD_LOGIC;
      x_rsc_17_0_tr_write_done : IN STD_LOGIC;
      x_rsc_17_0_RREADY : IN STD_LOGIC;
      x_rsc_17_0_RVALID : OUT STD_LOGIC;
      x_rsc_17_0_RUSER : OUT STD_LOGIC;
      x_rsc_17_0_RLAST : OUT STD_LOGIC;
      x_rsc_17_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_RID : OUT STD_LOGIC;
      x_rsc_17_0_ARREADY : OUT STD_LOGIC;
      x_rsc_17_0_ARVALID : IN STD_LOGIC;
      x_rsc_17_0_ARUSER : IN STD_LOGIC;
      x_rsc_17_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_ARLOCK : IN STD_LOGIC;
      x_rsc_17_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_17_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_17_0_ARID : IN STD_LOGIC;
      x_rsc_17_0_BREADY : IN STD_LOGIC;
      x_rsc_17_0_BVALID : OUT STD_LOGIC;
      x_rsc_17_0_BUSER : OUT STD_LOGIC;
      x_rsc_17_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_BID : OUT STD_LOGIC;
      x_rsc_17_0_WREADY : OUT STD_LOGIC;
      x_rsc_17_0_WVALID : IN STD_LOGIC;
      x_rsc_17_0_WUSER : IN STD_LOGIC;
      x_rsc_17_0_WLAST : IN STD_LOGIC;
      x_rsc_17_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_AWREADY : OUT STD_LOGIC;
      x_rsc_17_0_AWVALID : IN STD_LOGIC;
      x_rsc_17_0_AWUSER : IN STD_LOGIC;
      x_rsc_17_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_AWLOCK : IN STD_LOGIC;
      x_rsc_17_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_17_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_17_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_17_0_i_oswt : IN STD_LOGIC;
      x_rsc_17_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_17_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_17_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_17_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_17_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_17_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_18_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_18_0_s_tdone : IN STD_LOGIC;
      x_rsc_18_0_tr_write_done : IN STD_LOGIC;
      x_rsc_18_0_RREADY : IN STD_LOGIC;
      x_rsc_18_0_RVALID : OUT STD_LOGIC;
      x_rsc_18_0_RUSER : OUT STD_LOGIC;
      x_rsc_18_0_RLAST : OUT STD_LOGIC;
      x_rsc_18_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_RID : OUT STD_LOGIC;
      x_rsc_18_0_ARREADY : OUT STD_LOGIC;
      x_rsc_18_0_ARVALID : IN STD_LOGIC;
      x_rsc_18_0_ARUSER : IN STD_LOGIC;
      x_rsc_18_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_ARLOCK : IN STD_LOGIC;
      x_rsc_18_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_18_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_18_0_ARID : IN STD_LOGIC;
      x_rsc_18_0_BREADY : IN STD_LOGIC;
      x_rsc_18_0_BVALID : OUT STD_LOGIC;
      x_rsc_18_0_BUSER : OUT STD_LOGIC;
      x_rsc_18_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_BID : OUT STD_LOGIC;
      x_rsc_18_0_WREADY : OUT STD_LOGIC;
      x_rsc_18_0_WVALID : IN STD_LOGIC;
      x_rsc_18_0_WUSER : IN STD_LOGIC;
      x_rsc_18_0_WLAST : IN STD_LOGIC;
      x_rsc_18_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_AWREADY : OUT STD_LOGIC;
      x_rsc_18_0_AWVALID : IN STD_LOGIC;
      x_rsc_18_0_AWUSER : IN STD_LOGIC;
      x_rsc_18_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_AWLOCK : IN STD_LOGIC;
      x_rsc_18_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_18_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_18_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_18_0_i_oswt : IN STD_LOGIC;
      x_rsc_18_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_18_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_18_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_18_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_18_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_18_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_19_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_19_0_s_tdone : IN STD_LOGIC;
      x_rsc_19_0_tr_write_done : IN STD_LOGIC;
      x_rsc_19_0_RREADY : IN STD_LOGIC;
      x_rsc_19_0_RVALID : OUT STD_LOGIC;
      x_rsc_19_0_RUSER : OUT STD_LOGIC;
      x_rsc_19_0_RLAST : OUT STD_LOGIC;
      x_rsc_19_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_RID : OUT STD_LOGIC;
      x_rsc_19_0_ARREADY : OUT STD_LOGIC;
      x_rsc_19_0_ARVALID : IN STD_LOGIC;
      x_rsc_19_0_ARUSER : IN STD_LOGIC;
      x_rsc_19_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_ARLOCK : IN STD_LOGIC;
      x_rsc_19_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_19_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_19_0_ARID : IN STD_LOGIC;
      x_rsc_19_0_BREADY : IN STD_LOGIC;
      x_rsc_19_0_BVALID : OUT STD_LOGIC;
      x_rsc_19_0_BUSER : OUT STD_LOGIC;
      x_rsc_19_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_BID : OUT STD_LOGIC;
      x_rsc_19_0_WREADY : OUT STD_LOGIC;
      x_rsc_19_0_WVALID : IN STD_LOGIC;
      x_rsc_19_0_WUSER : IN STD_LOGIC;
      x_rsc_19_0_WLAST : IN STD_LOGIC;
      x_rsc_19_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_AWREADY : OUT STD_LOGIC;
      x_rsc_19_0_AWVALID : IN STD_LOGIC;
      x_rsc_19_0_AWUSER : IN STD_LOGIC;
      x_rsc_19_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_AWLOCK : IN STD_LOGIC;
      x_rsc_19_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_19_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_19_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_19_0_i_oswt : IN STD_LOGIC;
      x_rsc_19_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_19_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_19_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_19_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_19_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_19_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_20_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_20_0_s_tdone : IN STD_LOGIC;
      x_rsc_20_0_tr_write_done : IN STD_LOGIC;
      x_rsc_20_0_RREADY : IN STD_LOGIC;
      x_rsc_20_0_RVALID : OUT STD_LOGIC;
      x_rsc_20_0_RUSER : OUT STD_LOGIC;
      x_rsc_20_0_RLAST : OUT STD_LOGIC;
      x_rsc_20_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_RID : OUT STD_LOGIC;
      x_rsc_20_0_ARREADY : OUT STD_LOGIC;
      x_rsc_20_0_ARVALID : IN STD_LOGIC;
      x_rsc_20_0_ARUSER : IN STD_LOGIC;
      x_rsc_20_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_ARLOCK : IN STD_LOGIC;
      x_rsc_20_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_20_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_20_0_ARID : IN STD_LOGIC;
      x_rsc_20_0_BREADY : IN STD_LOGIC;
      x_rsc_20_0_BVALID : OUT STD_LOGIC;
      x_rsc_20_0_BUSER : OUT STD_LOGIC;
      x_rsc_20_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_BID : OUT STD_LOGIC;
      x_rsc_20_0_WREADY : OUT STD_LOGIC;
      x_rsc_20_0_WVALID : IN STD_LOGIC;
      x_rsc_20_0_WUSER : IN STD_LOGIC;
      x_rsc_20_0_WLAST : IN STD_LOGIC;
      x_rsc_20_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_AWREADY : OUT STD_LOGIC;
      x_rsc_20_0_AWVALID : IN STD_LOGIC;
      x_rsc_20_0_AWUSER : IN STD_LOGIC;
      x_rsc_20_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_AWLOCK : IN STD_LOGIC;
      x_rsc_20_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_20_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_20_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_20_0_i_oswt : IN STD_LOGIC;
      x_rsc_20_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_20_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_20_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_20_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_20_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_20_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_21_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_21_0_s_tdone : IN STD_LOGIC;
      x_rsc_21_0_tr_write_done : IN STD_LOGIC;
      x_rsc_21_0_RREADY : IN STD_LOGIC;
      x_rsc_21_0_RVALID : OUT STD_LOGIC;
      x_rsc_21_0_RUSER : OUT STD_LOGIC;
      x_rsc_21_0_RLAST : OUT STD_LOGIC;
      x_rsc_21_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_RID : OUT STD_LOGIC;
      x_rsc_21_0_ARREADY : OUT STD_LOGIC;
      x_rsc_21_0_ARVALID : IN STD_LOGIC;
      x_rsc_21_0_ARUSER : IN STD_LOGIC;
      x_rsc_21_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_ARLOCK : IN STD_LOGIC;
      x_rsc_21_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_21_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_21_0_ARID : IN STD_LOGIC;
      x_rsc_21_0_BREADY : IN STD_LOGIC;
      x_rsc_21_0_BVALID : OUT STD_LOGIC;
      x_rsc_21_0_BUSER : OUT STD_LOGIC;
      x_rsc_21_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_BID : OUT STD_LOGIC;
      x_rsc_21_0_WREADY : OUT STD_LOGIC;
      x_rsc_21_0_WVALID : IN STD_LOGIC;
      x_rsc_21_0_WUSER : IN STD_LOGIC;
      x_rsc_21_0_WLAST : IN STD_LOGIC;
      x_rsc_21_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_AWREADY : OUT STD_LOGIC;
      x_rsc_21_0_AWVALID : IN STD_LOGIC;
      x_rsc_21_0_AWUSER : IN STD_LOGIC;
      x_rsc_21_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_AWLOCK : IN STD_LOGIC;
      x_rsc_21_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_21_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_21_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_21_0_i_oswt : IN STD_LOGIC;
      x_rsc_21_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_21_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_21_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_21_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_21_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_21_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_22_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_22_0_s_tdone : IN STD_LOGIC;
      x_rsc_22_0_tr_write_done : IN STD_LOGIC;
      x_rsc_22_0_RREADY : IN STD_LOGIC;
      x_rsc_22_0_RVALID : OUT STD_LOGIC;
      x_rsc_22_0_RUSER : OUT STD_LOGIC;
      x_rsc_22_0_RLAST : OUT STD_LOGIC;
      x_rsc_22_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_RID : OUT STD_LOGIC;
      x_rsc_22_0_ARREADY : OUT STD_LOGIC;
      x_rsc_22_0_ARVALID : IN STD_LOGIC;
      x_rsc_22_0_ARUSER : IN STD_LOGIC;
      x_rsc_22_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_ARLOCK : IN STD_LOGIC;
      x_rsc_22_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_22_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_22_0_ARID : IN STD_LOGIC;
      x_rsc_22_0_BREADY : IN STD_LOGIC;
      x_rsc_22_0_BVALID : OUT STD_LOGIC;
      x_rsc_22_0_BUSER : OUT STD_LOGIC;
      x_rsc_22_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_BID : OUT STD_LOGIC;
      x_rsc_22_0_WREADY : OUT STD_LOGIC;
      x_rsc_22_0_WVALID : IN STD_LOGIC;
      x_rsc_22_0_WUSER : IN STD_LOGIC;
      x_rsc_22_0_WLAST : IN STD_LOGIC;
      x_rsc_22_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_AWREADY : OUT STD_LOGIC;
      x_rsc_22_0_AWVALID : IN STD_LOGIC;
      x_rsc_22_0_AWUSER : IN STD_LOGIC;
      x_rsc_22_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_AWLOCK : IN STD_LOGIC;
      x_rsc_22_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_22_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_22_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_22_0_i_oswt : IN STD_LOGIC;
      x_rsc_22_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_22_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_22_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_22_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_22_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_22_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_23_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_23_0_s_tdone : IN STD_LOGIC;
      x_rsc_23_0_tr_write_done : IN STD_LOGIC;
      x_rsc_23_0_RREADY : IN STD_LOGIC;
      x_rsc_23_0_RVALID : OUT STD_LOGIC;
      x_rsc_23_0_RUSER : OUT STD_LOGIC;
      x_rsc_23_0_RLAST : OUT STD_LOGIC;
      x_rsc_23_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_RID : OUT STD_LOGIC;
      x_rsc_23_0_ARREADY : OUT STD_LOGIC;
      x_rsc_23_0_ARVALID : IN STD_LOGIC;
      x_rsc_23_0_ARUSER : IN STD_LOGIC;
      x_rsc_23_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_ARLOCK : IN STD_LOGIC;
      x_rsc_23_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_23_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_23_0_ARID : IN STD_LOGIC;
      x_rsc_23_0_BREADY : IN STD_LOGIC;
      x_rsc_23_0_BVALID : OUT STD_LOGIC;
      x_rsc_23_0_BUSER : OUT STD_LOGIC;
      x_rsc_23_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_BID : OUT STD_LOGIC;
      x_rsc_23_0_WREADY : OUT STD_LOGIC;
      x_rsc_23_0_WVALID : IN STD_LOGIC;
      x_rsc_23_0_WUSER : IN STD_LOGIC;
      x_rsc_23_0_WLAST : IN STD_LOGIC;
      x_rsc_23_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_AWREADY : OUT STD_LOGIC;
      x_rsc_23_0_AWVALID : IN STD_LOGIC;
      x_rsc_23_0_AWUSER : IN STD_LOGIC;
      x_rsc_23_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_AWLOCK : IN STD_LOGIC;
      x_rsc_23_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_23_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_23_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_23_0_i_oswt : IN STD_LOGIC;
      x_rsc_23_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_23_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_23_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_23_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_23_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_23_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_24_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_24_0_s_tdone : IN STD_LOGIC;
      x_rsc_24_0_tr_write_done : IN STD_LOGIC;
      x_rsc_24_0_RREADY : IN STD_LOGIC;
      x_rsc_24_0_RVALID : OUT STD_LOGIC;
      x_rsc_24_0_RUSER : OUT STD_LOGIC;
      x_rsc_24_0_RLAST : OUT STD_LOGIC;
      x_rsc_24_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_RID : OUT STD_LOGIC;
      x_rsc_24_0_ARREADY : OUT STD_LOGIC;
      x_rsc_24_0_ARVALID : IN STD_LOGIC;
      x_rsc_24_0_ARUSER : IN STD_LOGIC;
      x_rsc_24_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_ARLOCK : IN STD_LOGIC;
      x_rsc_24_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_24_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_24_0_ARID : IN STD_LOGIC;
      x_rsc_24_0_BREADY : IN STD_LOGIC;
      x_rsc_24_0_BVALID : OUT STD_LOGIC;
      x_rsc_24_0_BUSER : OUT STD_LOGIC;
      x_rsc_24_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_BID : OUT STD_LOGIC;
      x_rsc_24_0_WREADY : OUT STD_LOGIC;
      x_rsc_24_0_WVALID : IN STD_LOGIC;
      x_rsc_24_0_WUSER : IN STD_LOGIC;
      x_rsc_24_0_WLAST : IN STD_LOGIC;
      x_rsc_24_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_AWREADY : OUT STD_LOGIC;
      x_rsc_24_0_AWVALID : IN STD_LOGIC;
      x_rsc_24_0_AWUSER : IN STD_LOGIC;
      x_rsc_24_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_AWLOCK : IN STD_LOGIC;
      x_rsc_24_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_24_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_24_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_24_0_i_oswt : IN STD_LOGIC;
      x_rsc_24_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_24_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_24_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_24_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_24_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_24_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_25_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_25_0_s_tdone : IN STD_LOGIC;
      x_rsc_25_0_tr_write_done : IN STD_LOGIC;
      x_rsc_25_0_RREADY : IN STD_LOGIC;
      x_rsc_25_0_RVALID : OUT STD_LOGIC;
      x_rsc_25_0_RUSER : OUT STD_LOGIC;
      x_rsc_25_0_RLAST : OUT STD_LOGIC;
      x_rsc_25_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_RID : OUT STD_LOGIC;
      x_rsc_25_0_ARREADY : OUT STD_LOGIC;
      x_rsc_25_0_ARVALID : IN STD_LOGIC;
      x_rsc_25_0_ARUSER : IN STD_LOGIC;
      x_rsc_25_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_ARLOCK : IN STD_LOGIC;
      x_rsc_25_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_25_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_25_0_ARID : IN STD_LOGIC;
      x_rsc_25_0_BREADY : IN STD_LOGIC;
      x_rsc_25_0_BVALID : OUT STD_LOGIC;
      x_rsc_25_0_BUSER : OUT STD_LOGIC;
      x_rsc_25_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_BID : OUT STD_LOGIC;
      x_rsc_25_0_WREADY : OUT STD_LOGIC;
      x_rsc_25_0_WVALID : IN STD_LOGIC;
      x_rsc_25_0_WUSER : IN STD_LOGIC;
      x_rsc_25_0_WLAST : IN STD_LOGIC;
      x_rsc_25_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_AWREADY : OUT STD_LOGIC;
      x_rsc_25_0_AWVALID : IN STD_LOGIC;
      x_rsc_25_0_AWUSER : IN STD_LOGIC;
      x_rsc_25_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_AWLOCK : IN STD_LOGIC;
      x_rsc_25_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_25_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_25_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_25_0_i_oswt : IN STD_LOGIC;
      x_rsc_25_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_25_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_25_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_25_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_25_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_25_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_26_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_26_0_s_tdone : IN STD_LOGIC;
      x_rsc_26_0_tr_write_done : IN STD_LOGIC;
      x_rsc_26_0_RREADY : IN STD_LOGIC;
      x_rsc_26_0_RVALID : OUT STD_LOGIC;
      x_rsc_26_0_RUSER : OUT STD_LOGIC;
      x_rsc_26_0_RLAST : OUT STD_LOGIC;
      x_rsc_26_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_RID : OUT STD_LOGIC;
      x_rsc_26_0_ARREADY : OUT STD_LOGIC;
      x_rsc_26_0_ARVALID : IN STD_LOGIC;
      x_rsc_26_0_ARUSER : IN STD_LOGIC;
      x_rsc_26_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_ARLOCK : IN STD_LOGIC;
      x_rsc_26_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_26_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_26_0_ARID : IN STD_LOGIC;
      x_rsc_26_0_BREADY : IN STD_LOGIC;
      x_rsc_26_0_BVALID : OUT STD_LOGIC;
      x_rsc_26_0_BUSER : OUT STD_LOGIC;
      x_rsc_26_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_BID : OUT STD_LOGIC;
      x_rsc_26_0_WREADY : OUT STD_LOGIC;
      x_rsc_26_0_WVALID : IN STD_LOGIC;
      x_rsc_26_0_WUSER : IN STD_LOGIC;
      x_rsc_26_0_WLAST : IN STD_LOGIC;
      x_rsc_26_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_AWREADY : OUT STD_LOGIC;
      x_rsc_26_0_AWVALID : IN STD_LOGIC;
      x_rsc_26_0_AWUSER : IN STD_LOGIC;
      x_rsc_26_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_AWLOCK : IN STD_LOGIC;
      x_rsc_26_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_26_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_26_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_26_0_i_oswt : IN STD_LOGIC;
      x_rsc_26_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_26_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_26_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_26_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_26_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_26_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_27_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_27_0_s_tdone : IN STD_LOGIC;
      x_rsc_27_0_tr_write_done : IN STD_LOGIC;
      x_rsc_27_0_RREADY : IN STD_LOGIC;
      x_rsc_27_0_RVALID : OUT STD_LOGIC;
      x_rsc_27_0_RUSER : OUT STD_LOGIC;
      x_rsc_27_0_RLAST : OUT STD_LOGIC;
      x_rsc_27_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_RID : OUT STD_LOGIC;
      x_rsc_27_0_ARREADY : OUT STD_LOGIC;
      x_rsc_27_0_ARVALID : IN STD_LOGIC;
      x_rsc_27_0_ARUSER : IN STD_LOGIC;
      x_rsc_27_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_ARLOCK : IN STD_LOGIC;
      x_rsc_27_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_27_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_27_0_ARID : IN STD_LOGIC;
      x_rsc_27_0_BREADY : IN STD_LOGIC;
      x_rsc_27_0_BVALID : OUT STD_LOGIC;
      x_rsc_27_0_BUSER : OUT STD_LOGIC;
      x_rsc_27_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_BID : OUT STD_LOGIC;
      x_rsc_27_0_WREADY : OUT STD_LOGIC;
      x_rsc_27_0_WVALID : IN STD_LOGIC;
      x_rsc_27_0_WUSER : IN STD_LOGIC;
      x_rsc_27_0_WLAST : IN STD_LOGIC;
      x_rsc_27_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_AWREADY : OUT STD_LOGIC;
      x_rsc_27_0_AWVALID : IN STD_LOGIC;
      x_rsc_27_0_AWUSER : IN STD_LOGIC;
      x_rsc_27_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_AWLOCK : IN STD_LOGIC;
      x_rsc_27_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_27_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_27_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_27_0_i_oswt : IN STD_LOGIC;
      x_rsc_27_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_27_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_27_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_27_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_27_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_27_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_28_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_28_0_s_tdone : IN STD_LOGIC;
      x_rsc_28_0_tr_write_done : IN STD_LOGIC;
      x_rsc_28_0_RREADY : IN STD_LOGIC;
      x_rsc_28_0_RVALID : OUT STD_LOGIC;
      x_rsc_28_0_RUSER : OUT STD_LOGIC;
      x_rsc_28_0_RLAST : OUT STD_LOGIC;
      x_rsc_28_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_RID : OUT STD_LOGIC;
      x_rsc_28_0_ARREADY : OUT STD_LOGIC;
      x_rsc_28_0_ARVALID : IN STD_LOGIC;
      x_rsc_28_0_ARUSER : IN STD_LOGIC;
      x_rsc_28_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_ARLOCK : IN STD_LOGIC;
      x_rsc_28_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_28_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_28_0_ARID : IN STD_LOGIC;
      x_rsc_28_0_BREADY : IN STD_LOGIC;
      x_rsc_28_0_BVALID : OUT STD_LOGIC;
      x_rsc_28_0_BUSER : OUT STD_LOGIC;
      x_rsc_28_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_BID : OUT STD_LOGIC;
      x_rsc_28_0_WREADY : OUT STD_LOGIC;
      x_rsc_28_0_WVALID : IN STD_LOGIC;
      x_rsc_28_0_WUSER : IN STD_LOGIC;
      x_rsc_28_0_WLAST : IN STD_LOGIC;
      x_rsc_28_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_AWREADY : OUT STD_LOGIC;
      x_rsc_28_0_AWVALID : IN STD_LOGIC;
      x_rsc_28_0_AWUSER : IN STD_LOGIC;
      x_rsc_28_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_AWLOCK : IN STD_LOGIC;
      x_rsc_28_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_28_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_28_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_28_0_i_oswt : IN STD_LOGIC;
      x_rsc_28_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_28_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_28_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_28_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_28_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_28_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_29_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_29_0_s_tdone : IN STD_LOGIC;
      x_rsc_29_0_tr_write_done : IN STD_LOGIC;
      x_rsc_29_0_RREADY : IN STD_LOGIC;
      x_rsc_29_0_RVALID : OUT STD_LOGIC;
      x_rsc_29_0_RUSER : OUT STD_LOGIC;
      x_rsc_29_0_RLAST : OUT STD_LOGIC;
      x_rsc_29_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_RID : OUT STD_LOGIC;
      x_rsc_29_0_ARREADY : OUT STD_LOGIC;
      x_rsc_29_0_ARVALID : IN STD_LOGIC;
      x_rsc_29_0_ARUSER : IN STD_LOGIC;
      x_rsc_29_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_ARLOCK : IN STD_LOGIC;
      x_rsc_29_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_29_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_29_0_ARID : IN STD_LOGIC;
      x_rsc_29_0_BREADY : IN STD_LOGIC;
      x_rsc_29_0_BVALID : OUT STD_LOGIC;
      x_rsc_29_0_BUSER : OUT STD_LOGIC;
      x_rsc_29_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_BID : OUT STD_LOGIC;
      x_rsc_29_0_WREADY : OUT STD_LOGIC;
      x_rsc_29_0_WVALID : IN STD_LOGIC;
      x_rsc_29_0_WUSER : IN STD_LOGIC;
      x_rsc_29_0_WLAST : IN STD_LOGIC;
      x_rsc_29_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_AWREADY : OUT STD_LOGIC;
      x_rsc_29_0_AWVALID : IN STD_LOGIC;
      x_rsc_29_0_AWUSER : IN STD_LOGIC;
      x_rsc_29_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_AWLOCK : IN STD_LOGIC;
      x_rsc_29_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_29_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_29_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_29_0_i_oswt : IN STD_LOGIC;
      x_rsc_29_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_29_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_29_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_29_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_29_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_29_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_30_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_30_0_s_tdone : IN STD_LOGIC;
      x_rsc_30_0_tr_write_done : IN STD_LOGIC;
      x_rsc_30_0_RREADY : IN STD_LOGIC;
      x_rsc_30_0_RVALID : OUT STD_LOGIC;
      x_rsc_30_0_RUSER : OUT STD_LOGIC;
      x_rsc_30_0_RLAST : OUT STD_LOGIC;
      x_rsc_30_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_RID : OUT STD_LOGIC;
      x_rsc_30_0_ARREADY : OUT STD_LOGIC;
      x_rsc_30_0_ARVALID : IN STD_LOGIC;
      x_rsc_30_0_ARUSER : IN STD_LOGIC;
      x_rsc_30_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_ARLOCK : IN STD_LOGIC;
      x_rsc_30_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_30_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_30_0_ARID : IN STD_LOGIC;
      x_rsc_30_0_BREADY : IN STD_LOGIC;
      x_rsc_30_0_BVALID : OUT STD_LOGIC;
      x_rsc_30_0_BUSER : OUT STD_LOGIC;
      x_rsc_30_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_BID : OUT STD_LOGIC;
      x_rsc_30_0_WREADY : OUT STD_LOGIC;
      x_rsc_30_0_WVALID : IN STD_LOGIC;
      x_rsc_30_0_WUSER : IN STD_LOGIC;
      x_rsc_30_0_WLAST : IN STD_LOGIC;
      x_rsc_30_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_AWREADY : OUT STD_LOGIC;
      x_rsc_30_0_AWVALID : IN STD_LOGIC;
      x_rsc_30_0_AWUSER : IN STD_LOGIC;
      x_rsc_30_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_AWLOCK : IN STD_LOGIC;
      x_rsc_30_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_30_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_30_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_30_0_i_oswt : IN STD_LOGIC;
      x_rsc_30_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_30_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_30_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_30_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_30_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_30_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_31_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_31_0_s_tdone : IN STD_LOGIC;
      x_rsc_31_0_tr_write_done : IN STD_LOGIC;
      x_rsc_31_0_RREADY : IN STD_LOGIC;
      x_rsc_31_0_RVALID : OUT STD_LOGIC;
      x_rsc_31_0_RUSER : OUT STD_LOGIC;
      x_rsc_31_0_RLAST : OUT STD_LOGIC;
      x_rsc_31_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_RID : OUT STD_LOGIC;
      x_rsc_31_0_ARREADY : OUT STD_LOGIC;
      x_rsc_31_0_ARVALID : IN STD_LOGIC;
      x_rsc_31_0_ARUSER : IN STD_LOGIC;
      x_rsc_31_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_ARLOCK : IN STD_LOGIC;
      x_rsc_31_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_31_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_31_0_ARID : IN STD_LOGIC;
      x_rsc_31_0_BREADY : IN STD_LOGIC;
      x_rsc_31_0_BVALID : OUT STD_LOGIC;
      x_rsc_31_0_BUSER : OUT STD_LOGIC;
      x_rsc_31_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_BID : OUT STD_LOGIC;
      x_rsc_31_0_WREADY : OUT STD_LOGIC;
      x_rsc_31_0_WVALID : IN STD_LOGIC;
      x_rsc_31_0_WUSER : IN STD_LOGIC;
      x_rsc_31_0_WLAST : IN STD_LOGIC;
      x_rsc_31_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_AWREADY : OUT STD_LOGIC;
      x_rsc_31_0_AWVALID : IN STD_LOGIC;
      x_rsc_31_0_AWUSER : IN STD_LOGIC;
      x_rsc_31_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_AWLOCK : IN STD_LOGIC;
      x_rsc_31_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_31_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_31_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      x_rsc_31_0_i_oswt : IN STD_LOGIC;
      x_rsc_31_0_i_wen_comp : OUT STD_LOGIC;
      x_rsc_31_0_i_oswt_1 : IN STD_LOGIC;
      x_rsc_31_0_i_wen_comp_1 : OUT STD_LOGIC;
      x_rsc_31_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_31_0_i_s_waddr_core : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      x_rsc_31_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_i_s_dout_core : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWREGION : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_waddr_core : STD_LOGIC_VECTOR
      (4 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_dout_core : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT hybrid_core_x_rsc_triosy_31_0_obj
    PORT(
      x_rsc_triosy_31_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_31_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_30_0_obj
    PORT(
      x_rsc_triosy_30_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_30_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_29_0_obj
    PORT(
      x_rsc_triosy_29_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_29_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_28_0_obj
    PORT(
      x_rsc_triosy_28_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_28_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_27_0_obj
    PORT(
      x_rsc_triosy_27_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_27_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_26_0_obj
    PORT(
      x_rsc_triosy_26_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_26_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_25_0_obj
    PORT(
      x_rsc_triosy_25_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_25_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_24_0_obj
    PORT(
      x_rsc_triosy_24_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_24_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_23_0_obj
    PORT(
      x_rsc_triosy_23_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_23_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_22_0_obj
    PORT(
      x_rsc_triosy_22_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_22_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_21_0_obj
    PORT(
      x_rsc_triosy_21_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_21_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_20_0_obj
    PORT(
      x_rsc_triosy_20_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_20_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_19_0_obj
    PORT(
      x_rsc_triosy_19_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_19_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_18_0_obj
    PORT(
      x_rsc_triosy_18_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_18_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_17_0_obj
    PORT(
      x_rsc_triosy_17_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_17_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_16_0_obj
    PORT(
      x_rsc_triosy_16_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_16_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_15_0_obj
    PORT(
      x_rsc_triosy_15_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_15_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_14_0_obj
    PORT(
      x_rsc_triosy_14_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_14_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_13_0_obj
    PORT(
      x_rsc_triosy_13_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_13_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_12_0_obj
    PORT(
      x_rsc_triosy_12_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_12_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_11_0_obj
    PORT(
      x_rsc_triosy_11_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_11_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_10_0_obj
    PORT(
      x_rsc_triosy_10_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_10_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_9_0_obj
    PORT(
      x_rsc_triosy_9_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_9_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_8_0_obj
    PORT(
      x_rsc_triosy_8_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_8_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_7_0_obj
    PORT(
      x_rsc_triosy_7_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_7_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_6_0_obj
    PORT(
      x_rsc_triosy_6_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_6_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_5_0_obj
    PORT(
      x_rsc_triosy_5_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_5_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_4_0_obj
    PORT(
      x_rsc_triosy_4_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_4_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_3_0_obj
    PORT(
      x_rsc_triosy_3_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_3_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_2_0_obj
    PORT(
      x_rsc_triosy_2_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_2_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_1_0_obj
    PORT(
      x_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_x_rsc_triosy_0_0_obj
    PORT(
      x_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      x_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_m_rsc_triosy_obj
    PORT(
      m_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      m_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_twiddle_rsc_triosy_obj
    PORT(
      twiddle_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_twiddle_h_rsc_triosy_obj
    PORT(
      twiddle_h_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_revArr_rsc_triosy_obj
    PORT(
      revArr_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      revArr_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_tw_rsc_triosy_obj
    PORT(
      tw_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      tw_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_tw_h_rsc_triosy_obj
    PORT(
      tw_h_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      tw_h_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_staller
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      core_wen : OUT STD_LOGIC;
      core_wten : OUT STD_LOGIC;
      revArr_rsci_wen_comp : IN STD_LOGIC;
      tw_rsci_wen_comp : IN STD_LOGIC;
      tw_h_rsci_wen_comp : IN STD_LOGIC;
      x_rsc_0_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_0_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_1_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_1_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_2_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_2_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_3_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_3_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_4_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_4_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_5_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_5_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_6_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_6_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_7_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_7_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_8_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_8_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_9_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_9_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_10_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_10_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_11_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_11_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_12_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_12_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_13_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_13_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_14_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_14_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_15_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_15_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_16_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_16_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_17_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_17_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_18_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_18_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_19_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_19_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_20_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_20_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_21_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_21_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_22_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_22_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_23_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_23_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_24_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_24_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_25_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_25_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_26_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_26_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_27_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_27_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_28_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_28_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_29_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_29_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_30_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_30_0_i_wen_comp_1 : IN STD_LOGIC;
      x_rsc_31_0_i_wen_comp : IN STD_LOGIC;
      x_rsc_31_0_i_wen_comp_1 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT hybrid_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
      S1_OUTER_LOOP_for_C_5_tr0 : IN STD_LOGIC;
      S1_OUTER_LOOP_C_0_tr0 : IN STD_LOGIC;
      S2_COPY_LOOP_for_C_4_tr0 : IN STD_LOGIC;
      S2_COPY_LOOP_C_0_tr0 : IN STD_LOGIC;
      S2_INNER_LOOP1_for_C_20_tr0 : IN STD_LOGIC;
      S2_INNER_LOOP1_C_2_tr0 : IN STD_LOGIC;
      S2_INNER_LOOP2_for_C_20_tr0 : IN STD_LOGIC;
      S2_INNER_LOOP2_C_2_tr0 : IN STD_LOGIC;
      S2_INNER_LOOP2_C_2_tr1 : IN STD_LOGIC;
      S2_INNER_LOOP3_for_C_20_tr0 : IN STD_LOGIC;
      S2_INNER_LOOP3_C_2_tr0 : IN STD_LOGIC;
      S34_OUTER_LOOP_for_C_12_tr0 : IN STD_LOGIC;
      S34_OUTER_LOOP_C_0_tr0 : IN STD_LOGIC;
      S5_COPY_LOOP_for_C_4_tr0 : IN STD_LOGIC;
      S5_COPY_LOOP_C_0_tr0 : IN STD_LOGIC;
      S5_INNER_LOOP1_for_C_20_tr0 : IN STD_LOGIC;
      S5_INNER_LOOP1_C_2_tr0 : IN STD_LOGIC;
      S5_INNER_LOOP2_for_C_20_tr0 : IN STD_LOGIC;
      S5_INNER_LOOP2_C_2_tr0 : IN STD_LOGIC;
      S5_INNER_LOOP2_C_2_tr1 : IN STD_LOGIC;
      S5_INNER_LOOP3_for_C_20_tr0 : IN STD_LOGIC;
      S5_INNER_LOOP3_C_2_tr0 : IN STD_LOGIC;
      S6_OUTER_LOOP_for_C_4_tr0 : IN STD_LOGIC;
      S6_OUTER_LOOP_C_0_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL hybrid_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_core_fsm_inst_S1_OUTER_LOOP_for_C_5_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S1_OUTER_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_COPY_LOOP_for_C_4_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_COPY_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP1_for_C_20_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP1_C_2_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP2_for_C_20_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP2_C_2_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP2_C_2_tr1 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP3_for_C_20_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S2_INNER_LOOP3_C_2_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S34_OUTER_LOOP_for_C_12_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S34_OUTER_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_COPY_LOOP_for_C_4_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_COPY_LOOP_C_0_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP1_for_C_20_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP1_C_2_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP2_for_C_20_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP2_C_2_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP2_C_2_tr1 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP3_for_C_20_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S5_INNER_LOOP3_C_2_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S6_OUTER_LOOP_for_C_4_tr0 : STD_LOGIC;
  SIGNAL hybrid_core_core_fsm_inst_S6_OUTER_LOOP_C_0_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_3_2(input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_s_1_5_2(input_4 : STD_LOGIC;
  input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
      tmp := sel(4);
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_31_3_2(input_2 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_31_4_2(input_3 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_10_2(input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(9 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_11_2(input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(10 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_32_2(input_31 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(31 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_33_2(input_32 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(32 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_34_2(input_33 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_32 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_31 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_30 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_29 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_28 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_27 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_26 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_25 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_24 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_23 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_22 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_21 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_20 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_19 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_18 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_17 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_16 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_15 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_14 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_13 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_12 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(33 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
      tmp := (OTHERS=>sel( 12));
      result := result or ( input_12 and tmp);
      tmp := (OTHERS=>sel( 13));
      result := result or ( input_13 and tmp);
      tmp := (OTHERS=>sel( 14));
      result := result or ( input_14 and tmp);
      tmp := (OTHERS=>sel( 15));
      result := result or ( input_15 and tmp);
      tmp := (OTHERS=>sel( 16));
      result := result or ( input_16 and tmp);
      tmp := (OTHERS=>sel( 17));
      result := result or ( input_17 and tmp);
      tmp := (OTHERS=>sel( 18));
      result := result or ( input_18 and tmp);
      tmp := (OTHERS=>sel( 19));
      result := result or ( input_19 and tmp);
      tmp := (OTHERS=>sel( 20));
      result := result or ( input_20 and tmp);
      tmp := (OTHERS=>sel( 21));
      result := result or ( input_21 and tmp);
      tmp := (OTHERS=>sel( 22));
      result := result or ( input_22 and tmp);
      tmp := (OTHERS=>sel( 23));
      result := result or ( input_23 and tmp);
      tmp := (OTHERS=>sel( 24));
      result := result or ( input_24 and tmp);
      tmp := (OTHERS=>sel( 25));
      result := result or ( input_25 and tmp);
      tmp := (OTHERS=>sel( 26));
      result := result or ( input_26 and tmp);
      tmp := (OTHERS=>sel( 27));
      result := result or ( input_27 and tmp);
      tmp := (OTHERS=>sel( 28));
      result := result or ( input_28 and tmp);
      tmp := (OTHERS=>sel( 29));
      result := result or ( input_29 and tmp);
      tmp := (OTHERS=>sel( 30));
      result := result or ( input_30 and tmp);
      tmp := (OTHERS=>sel( 31));
      result := result or ( input_31 and tmp);
      tmp := (OTHERS=>sel( 32));
      result := result or ( input_32 and tmp);
      tmp := (OTHERS=>sel( 33));
      result := result or ( input_33 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_3_2(input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_4_2(input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_5_2(input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_6_2(input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_7_2(input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(6 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_8_2(input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_9_2(input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_5_2(input_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_3_2(input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_4_2(input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_5_5_2(input_4 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_6_3_2(input_2 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_15_2_2(input_0 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(14 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(14 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_20_2_2(input_0 : STD_LOGIC_VECTOR(19 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(19 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(19 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  m_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 32
      )
    PORT MAP(
      dat => m_rsci_dat,
      idat => m_rsci_idat_1
    );
  m_rsci_dat <= m_rsc_dat;
  m_rsci_idat <= m_rsci_idat_1;

  mult_12_z_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 20,
      signd_a => 1,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_12_z_mul_cmp_a,
      b => mult_12_z_mul_cmp_b,
      clk => clk,
      en => mult_12_z_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_12_z_mul_cmp_z_1
    );
  mult_12_z_mul_cmp_a <= MUX_v_20_2_2(tw_rsci_s_din_mxwt, S34_OUTER_LOOP_for_tf_sva,
      and_dcpl_1007);
  mult_12_z_mul_cmp_b <= MUX_v_32_2_2(tmp_37_lpi_3_dfm_mx0w0, tmp_36_lpi_3_dfm, and_dcpl_1007);
  mult_12_z_mul_cmp_z <= mult_12_z_mul_cmp_z_1;

  mult_z_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_a,
      b => mult_z_mul_cmp_b,
      clk => clk,
      en => mult_z_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_z_1
    );
  mult_z_mul_cmp_a <= MUX1HOT_v_32_32_2(tmp_7_lpi_4_dfm_mx0w0, tmp_5_lpi_4_dfm, tmp_3_lpi_4_dfm,
      tmp_1_lpi_4_dfm, tmp_7_lpi_4_dfm, operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm,
      mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm, operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm,
      operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm, tmp_33_lpi_4_dfm,
      tmp_31_lpi_4_dfm, tmp_29_lpi_4_dfm, tmp_35_lpi_4_dfm, tmp_13_lpi_3_dfm, tmp_11_lpi_3_dfm,
      tmp_9_lpi_3_dfm, tmp_15_lpi_3_dfm, tmp_37_lpi_3_dfm_mx0w0, tmp_36_lpi_3_dfm,
      (mult_z_mul_cmp_z(51 DOWNTO 20)), tmp_43_lpi_4_dfm, tmp_41_lpi_4_dfm, tmp_39_lpi_4_dfm,
      tmp_45_lpi_4_dfm, tmp_22_lpi_4_dfm, tmp_20_lpi_4_dfm, tmp_18_lpi_4_dfm, tmp_24_lpi_4_dfm,
      tmp_51_lpi_3_dfm, tmp_49_lpi_3_dfm, tmp_47_lpi_3_dfm, tmp_53_lpi_3_dfm, STD_LOGIC_VECTOR'(
      (MUX_s_1_2_2((MUX_s_1_2_2((NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(5)))
      OR (fsm_output(7)) OR (NOT (fsm_output(2))) OR (fsm_output(0)) OR (fsm_output(4)))),
      (NOT((fsm_output(3)) OR (MUX_s_1_2_2(((fsm_output(7)) OR (NOT (fsm_output(2)))
      OR (fsm_output(0)) OR (fsm_output(4))), or_tmp_3550, fsm_output(5))))), fsm_output(6))),
      (NOT((fsm_output(6)) OR (MUX_s_1_2_2((MUX_s_1_2_2(or_tmp_3550, ((NOT (fsm_output(7)))
      OR (fsm_output(2)) OR (fsm_output(0)) OR (fsm_output(4))), fsm_output(5))),
      ((fsm_output(5)) OR (NOT (fsm_output(7))) OR (fsm_output(2)) OR (fsm_output(0))
      OR (fsm_output(4))), fsm_output(3))))), fsm_output(1))) & (and_dcpl_1014 AND
      and_dcpl_1013) & (and_dcpl_1014 AND and_dcpl_1000 AND and_dcpl_1011) & (nor_tmp_3
      AND xor_dcpl_1 AND and_dcpl_1013) & (and_dcpl_76 AND and_dcpl_70) & (MUX_s_1_2_2((NOT((NOT
      (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(2)) OR (NOT (fsm_output(4)))
      OR (fsm_output(7)) OR not_tmp_1345)), mux_3678_cse, fsm_output(0))) & not_tmp_1349
      & ((MUX_s_1_2_2((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(6))) OR (fsm_output(7))
      OR (NOT (fsm_output(4))) OR (NOT (fsm_output(3))) OR (fsm_output(1)))), (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((NOT((NOT
      (fsm_output(4))) OR (NOT (fsm_output(3))) OR (fsm_output(1)))), (NOT((NOT (fsm_output(4)))
      OR (fsm_output(3)) OR (fsm_output(1)))), fsm_output(7))), (NOT((fsm_output(7))
      OR (fsm_output(4)) OR (NOT (fsm_output(3))) OR (fsm_output(1)))), fsm_output(6))),
      (NOT((fsm_output(6)) OR (MUX_s_1_2_2(((NOT (fsm_output(4))) OR (fsm_output(3))
      OR (NOT (fsm_output(1)))), or_3852_cse, fsm_output(7))))), fsm_output(5))),
      fsm_output(0))) AND (fsm_output(2))) & (MUX_s_1_2_2(((fsm_output(5)) AND (MUX_s_1_2_2((NOT((NOT
      (fsm_output(4))) OR (fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(0)) OR
      (NOT (fsm_output(2))))), (NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(6)))
      OR (fsm_output(7)) OR (NOT (fsm_output(0))) OR (fsm_output(2)))), fsm_output(3)))),
      (MUX_s_1_2_2((MUX_s_1_2_2((NOT((NOT (fsm_output(4))) OR (fsm_output(6)) OR
      (NOT (fsm_output(7))) OR (fsm_output(0)) OR (fsm_output(2)))), (MUX_s_1_2_2((NOT((NOT
      (fsm_output(6))) OR (fsm_output(7)) OR (fsm_output(0)) OR (NOT (fsm_output(2))))),
      (NOT((fsm_output(6)) OR (fsm_output(7)) OR (fsm_output(0)) OR (NOT (fsm_output(2))))),
      fsm_output(4))), fsm_output(3))), (NOT((NOT (fsm_output(3))) OR (fsm_output(4))
      OR (fsm_output(6)) OR (NOT (fsm_output(7))) OR (fsm_output(0)) OR (fsm_output(2)))),
      fsm_output(5))), fsm_output(1))) & (and_dcpl_1024 AND and_dcpl_1023) & (and_dcpl_1027
      AND and_dcpl_1012 AND and_dcpl_1022) & (and_dcpl_1027 AND and_dcpl_1023) &
      (and_dcpl_130 AND and_dcpl_478) & (and_dcpl_1033 AND and_dcpl_1032) & (and_dcpl_1037
      AND and_dcpl_1035 AND and_dcpl_1011) & (and_dcpl_1037 AND and_dcpl_1032) &
      (and_dcpl_72 AND and_dcpl_90) & and_dcpl_1041 & and_dcpl_1007 & (nor_tmp_4
      AND ((fsm_output(1)) XOR (fsm_output(0))) AND and_dcpl_90) & (nor_tmp_3 AND
      and_dcpl_1035 AND and_dcpl_1044) & (nor_tmp_674 AND and_dcpl_1044) & (and_dcpl_1014
      AND and_dcpl_1035 AND and_dcpl_1022) & (and_dcpl_148 AND and_dcpl_108) & (and_dcpl_1052
      AND and_dcpl_460 AND (fsm_output(7))) & (and_dcpl_1024 AND and_dcpl_1012 AND
      and_dcpl_1054) & (and_dcpl_1024 AND and_dcpl_1000 AND and_dcpl_1054) & (and_dcpl_111
      AND and_dcpl_115) & (and_dcpl_1052 AND and_dcpl_117) & (and_dcpl_1033 AND and_dcpl_1012
      AND and_2112_cse) & (and_dcpl_1033 AND and_dcpl_1000 AND and_2112_cse) & (and_dcpl_111
      AND and_dcpl_75)));
  mult_z_mul_cmp_b <= MUX1HOT_v_32_5_2(S2_INNER_LOOP1_tfh_sva, S2_INNER_LOOP1_tf_sva,
      m_sva, STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tw_h_rsci_s_din_mxwt),32)), STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(S34_OUTER_LOOP_for_tf_h_sva),32)),
      STD_LOGIC_VECTOR'( (NOT (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((NOT
      nor_tmp_4), mux_tmp_3698, fsm_output(0))), or_2273_cse, fsm_output(6))), (NOT((fsm_output(6))
      AND (NOT (MUX_s_1_2_2(mux_tmp_3698, or_119_cse, fsm_output(0)))))), fsm_output(5))),
      ((NOT (fsm_output(5))) OR (fsm_output(6)) OR (NOT (fsm_output(2))) OR (fsm_output(4))),
      fsm_output(3))), (MUX_s_1_2_2((CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01"))
      OR mux_37_cse), (CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"))
      OR mux_37_cse), fsm_output(3))), fsm_output(7)))) & (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2((NOT((NOT
      (fsm_output(4))) OR (fsm_output(1)) OR (NOT (fsm_output(7))) OR (fsm_output(6)))),
      (NOT((NOT (fsm_output(4))) OR (fsm_output(7)) OR (fsm_output(6)))), fsm_output(5))),
      (MUX_s_1_2_2((MUX_s_1_2_2(nor_1368_cse, (NOT(and_1317_cse OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("00")))), fsm_output(4))), (MUX_s_1_2_2((NOT((fsm_output(1))
      OR (NOT (fsm_output(7))) OR (fsm_output(6)))), (NOT((fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(7)) OR (NOT (fsm_output(6))))), fsm_output(4))), fsm_output(5))),
      fsm_output(3))), (MUX_s_1_2_2((MUX_s_1_2_2((NOT((NOT (fsm_output(4))) OR (NOT
      (fsm_output(0))) OR (NOT (fsm_output(1))) OR (fsm_output(7)) OR (fsm_output(6)))),
      (MUX_s_1_2_2((NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(7))) OR (fsm_output(6)))),
      (NOT(nor_1375_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01")))),
      fsm_output(4))), fsm_output(5))), (NOT((fsm_output(5)) OR (fsm_output(4)) OR
      (NOT (fsm_output(1))) OR (NOT (fsm_output(7))) OR (fsm_output(6)))), fsm_output(3))),
      fsm_output(2))) & (MUX_s_1_2_2((MUX_s_1_2_2((MUX_s_1_2_2(((fsm_output(5)) AND
      (fsm_output(4)) AND (fsm_output(2))), (NOT(CONV_SL_1_1(fsm_output(5 DOWNTO
      4)/=STD_LOGIC_VECTOR'("01")) OR (MUX_s_1_2_2((NOT (fsm_output(2))), (fsm_output(2)),
      and_1317_cse)))), fsm_output(3))), ((fsm_output(3)) AND (MUX_s_1_2_2((MUX_s_1_2_2((fsm_output(2)),
      (MUX_s_1_2_2(and_2141_cse, nor_2247_cse, fsm_output(0))), fsm_output(4))),
      ((fsm_output(4)) AND (MUX_s_1_2_2((fsm_output(2)), (NOT (fsm_output(2))), or_3894_cse))),
      fsm_output(5)))), fsm_output(6))), (NOT((fsm_output(6)) OR (MUX_s_1_2_2((CONV_SL_1_1(fsm_output(5
      DOWNTO 4)/=STD_LOGIC_VECTOR'("01")) OR mux_tmp_3714), (CONV_SL_1_1(fsm_output(5
      DOWNTO 4)/=STD_LOGIC_VECTOR'("10")) OR mux_tmp_3714), fsm_output(3))))), fsm_output(7)))
      & and_dcpl_1041 & and_dcpl_1007));
  mult_z_mul_cmp_z <= mult_z_mul_cmp_z_1;

  operator_33_true_1_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_bl_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 4,
      width_z => 4
      )
    PORT MAP(
      a => operator_33_true_1_lshift_rg_a,
      s => operator_33_true_1_lshift_rg_s,
      z => operator_33_true_1_lshift_rg_z
    );
  operator_33_true_1_lshift_rg_a(0) <= '1';
  operator_33_true_1_lshift_rg_s <= STD_LOGIC_VECTOR'( '0' & (S2_OUTER_LOOP_c_2_sva
      AND (NOT and_2383_ssc)) & (MUX_s_1_2_2(S2_OUTER_LOOP_c_1_sva, (NOT S2_OUTER_LOOP_c_1_sva),
      and_2383_ssc)) & and_2383_ssc);
  z_out_3 <= operator_33_true_1_lshift_rg_z;

  hybrid_core_twiddle_rsci_1_inst : hybrid_core_twiddle_rsci_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsci_adrb_d => hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_adrb_d,
      twiddle_rsci_qb_d => hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_qb_d,
      twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      twiddle_rsci_oswt => reg_twiddle_rsci_oswt_cse,
      core_wten => core_wten,
      twiddle_rsci_adrb_d_core => hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_adrb_d_core,
      twiddle_rsci_qb_d_mxwt => hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_qb_d_mxwt,
      twiddle_rsci_oswt_pff => mux_111_rmff
    );
  twiddle_rsci_adrb_d_reg <= hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_adrb_d;
  hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_qb_d <= twiddle_rsci_qb_d;
  hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_adrb_d_core <= '0' & S2_INNER_LOOP1_tfh_S2_INNER_LOOP1_tfh_mux_rmff
      & S2_INNER_LOOP1_tfh_mux1h_rmff;
  twiddle_rsci_qb_d_mxwt <= hybrid_core_twiddle_rsci_1_inst_twiddle_rsci_qb_d_mxwt;

  hybrid_core_wait_dp_inst : hybrid_core_wait_dp
    PORT MAP(
      clk => clk,
      xx_rsc_0_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_0_0_cgo_iro,
      xx_rsc_0_0_i_clka_en_d => xx_rsc_0_0_i_clka_en_d,
      xx_rsc_1_0_cgo_iro => mux_191_rmff,
      xx_rsc_1_0_i_clka_en_d => xx_rsc_1_0_i_clka_en_d,
      xx_rsc_2_0_cgo_iro => mux_241_rmff,
      xx_rsc_2_0_i_clka_en_d => xx_rsc_2_0_i_clka_en_d,
      xx_rsc_3_0_cgo_iro => mux_293_rmff,
      xx_rsc_3_0_i_clka_en_d => xx_rsc_3_0_i_clka_en_d,
      xx_rsc_4_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_4_0_cgo_iro,
      xx_rsc_4_0_i_clka_en_d => xx_rsc_4_0_i_clka_en_d,
      xx_rsc_5_0_cgo_iro => mux_408_rmff,
      xx_rsc_5_0_i_clka_en_d => xx_rsc_5_0_i_clka_en_d,
      xx_rsc_6_0_cgo_iro => mux_455_rmff,
      xx_rsc_6_0_i_clka_en_d => xx_rsc_6_0_i_clka_en_d,
      xx_rsc_7_0_cgo_iro => mux_504_rmff,
      xx_rsc_7_0_i_clka_en_d => xx_rsc_7_0_i_clka_en_d,
      xx_rsc_8_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_8_0_cgo_iro,
      xx_rsc_8_0_i_clka_en_d => xx_rsc_8_0_i_clka_en_d,
      xx_rsc_9_0_cgo_iro => mux_614_rmff,
      xx_rsc_9_0_i_clka_en_d => xx_rsc_9_0_i_clka_en_d,
      xx_rsc_10_0_cgo_iro => mux_661_rmff,
      xx_rsc_10_0_i_clka_en_d => xx_rsc_10_0_i_clka_en_d,
      xx_rsc_11_0_cgo_iro => mux_710_rmff,
      xx_rsc_11_0_i_clka_en_d => xx_rsc_11_0_i_clka_en_d,
      xx_rsc_12_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_12_0_cgo_iro,
      xx_rsc_12_0_i_clka_en_d => xx_rsc_12_0_i_clka_en_d,
      xx_rsc_13_0_cgo_iro => mux_820_rmff,
      xx_rsc_13_0_i_clka_en_d => xx_rsc_13_0_i_clka_en_d,
      xx_rsc_14_0_cgo_iro => mux_867_rmff,
      xx_rsc_14_0_i_clka_en_d => xx_rsc_14_0_i_clka_en_d,
      xx_rsc_15_0_cgo_iro => mux_916_rmff,
      xx_rsc_15_0_i_clka_en_d => xx_rsc_15_0_i_clka_en_d,
      xx_rsc_16_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_16_0_cgo_iro,
      xx_rsc_16_0_i_clka_en_d => xx_rsc_16_0_i_clka_en_d,
      xx_rsc_17_0_cgo_iro => mux_1030_rmff,
      xx_rsc_17_0_i_clka_en_d => xx_rsc_17_0_i_clka_en_d,
      xx_rsc_18_0_cgo_iro => mux_1080_rmff,
      xx_rsc_18_0_i_clka_en_d => xx_rsc_18_0_i_clka_en_d,
      xx_rsc_19_0_cgo_iro => mux_1132_rmff,
      xx_rsc_19_0_i_clka_en_d => xx_rsc_19_0_i_clka_en_d,
      xx_rsc_20_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_20_0_cgo_iro,
      xx_rsc_20_0_i_clka_en_d => xx_rsc_20_0_i_clka_en_d,
      xx_rsc_21_0_cgo_iro => mux_1248_rmff,
      xx_rsc_21_0_i_clka_en_d => xx_rsc_21_0_i_clka_en_d,
      xx_rsc_22_0_cgo_iro => mux_1298_rmff,
      xx_rsc_22_0_i_clka_en_d => xx_rsc_22_0_i_clka_en_d,
      xx_rsc_23_0_cgo_iro => mux_1350_rmff,
      xx_rsc_23_0_i_clka_en_d => xx_rsc_23_0_i_clka_en_d,
      xx_rsc_24_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_24_0_cgo_iro,
      xx_rsc_24_0_i_clka_en_d => xx_rsc_24_0_i_clka_en_d,
      xx_rsc_25_0_cgo_iro => mux_1465_rmff,
      xx_rsc_25_0_i_clka_en_d => xx_rsc_25_0_i_clka_en_d,
      xx_rsc_26_0_cgo_iro => mux_1515_rmff,
      xx_rsc_26_0_i_clka_en_d => xx_rsc_26_0_i_clka_en_d,
      xx_rsc_27_0_cgo_iro => mux_1567_rmff,
      xx_rsc_27_0_i_clka_en_d => xx_rsc_27_0_i_clka_en_d,
      xx_rsc_28_0_cgo_iro => hybrid_core_wait_dp_inst_xx_rsc_28_0_cgo_iro,
      xx_rsc_28_0_i_clka_en_d => xx_rsc_28_0_i_clka_en_d,
      xx_rsc_29_0_cgo_iro => mux_1682_rmff,
      xx_rsc_29_0_i_clka_en_d => xx_rsc_29_0_i_clka_en_d,
      xx_rsc_30_0_cgo_iro => mux_1732_rmff,
      xx_rsc_30_0_i_clka_en_d => xx_rsc_30_0_i_clka_en_d,
      xx_rsc_31_0_cgo_iro => mux_1781_rmff,
      xx_rsc_31_0_i_clka_en_d => xx_rsc_31_0_i_clka_en_d,
      yy_rsc_0_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_0_0_cgo_iro,
      yy_rsc_0_0_i_clka_en_d => yy_rsc_0_0_i_clka_en_d,
      yy_rsc_1_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_1_0_cgo_iro,
      yy_rsc_1_0_i_clka_en_d => yy_rsc_1_0_i_clka_en_d,
      yy_rsc_2_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_2_0_cgo_iro,
      yy_rsc_2_0_i_clka_en_d => yy_rsc_2_0_i_clka_en_d,
      yy_rsc_3_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_3_0_cgo_iro,
      yy_rsc_3_0_i_clka_en_d => yy_rsc_3_0_i_clka_en_d,
      yy_rsc_4_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_4_0_cgo_iro,
      yy_rsc_4_0_i_clka_en_d => yy_rsc_4_0_i_clka_en_d,
      yy_rsc_5_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_5_0_cgo_iro,
      yy_rsc_5_0_i_clka_en_d => yy_rsc_5_0_i_clka_en_d,
      yy_rsc_6_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_6_0_cgo_iro,
      yy_rsc_6_0_i_clka_en_d => yy_rsc_6_0_i_clka_en_d,
      yy_rsc_7_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_7_0_cgo_iro,
      yy_rsc_7_0_i_clka_en_d => yy_rsc_7_0_i_clka_en_d,
      yy_rsc_8_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_8_0_cgo_iro,
      yy_rsc_8_0_i_clka_en_d => yy_rsc_8_0_i_clka_en_d,
      yy_rsc_9_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_9_0_cgo_iro,
      yy_rsc_9_0_i_clka_en_d => yy_rsc_9_0_i_clka_en_d,
      yy_rsc_10_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_10_0_cgo_iro,
      yy_rsc_10_0_i_clka_en_d => yy_rsc_10_0_i_clka_en_d,
      yy_rsc_11_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_11_0_cgo_iro,
      yy_rsc_11_0_i_clka_en_d => yy_rsc_11_0_i_clka_en_d,
      yy_rsc_12_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_12_0_cgo_iro,
      yy_rsc_12_0_i_clka_en_d => yy_rsc_12_0_i_clka_en_d,
      yy_rsc_13_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_13_0_cgo_iro,
      yy_rsc_13_0_i_clka_en_d => yy_rsc_13_0_i_clka_en_d,
      yy_rsc_14_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_14_0_cgo_iro,
      yy_rsc_14_0_i_clka_en_d => yy_rsc_14_0_i_clka_en_d,
      yy_rsc_15_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_15_0_cgo_iro,
      yy_rsc_15_0_i_clka_en_d => yy_rsc_15_0_i_clka_en_d,
      yy_rsc_16_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_16_0_cgo_iro,
      yy_rsc_16_0_i_clka_en_d => yy_rsc_16_0_i_clka_en_d,
      yy_rsc_17_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_17_0_cgo_iro,
      yy_rsc_17_0_i_clka_en_d => yy_rsc_17_0_i_clka_en_d,
      yy_rsc_18_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_18_0_cgo_iro,
      yy_rsc_18_0_i_clka_en_d => yy_rsc_18_0_i_clka_en_d,
      yy_rsc_19_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_19_0_cgo_iro,
      yy_rsc_19_0_i_clka_en_d => yy_rsc_19_0_i_clka_en_d,
      yy_rsc_20_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_20_0_cgo_iro,
      yy_rsc_20_0_i_clka_en_d => yy_rsc_20_0_i_clka_en_d,
      yy_rsc_21_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_21_0_cgo_iro,
      yy_rsc_21_0_i_clka_en_d => yy_rsc_21_0_i_clka_en_d,
      yy_rsc_22_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_22_0_cgo_iro,
      yy_rsc_22_0_i_clka_en_d => yy_rsc_22_0_i_clka_en_d,
      yy_rsc_23_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_23_0_cgo_iro,
      yy_rsc_23_0_i_clka_en_d => yy_rsc_23_0_i_clka_en_d,
      yy_rsc_24_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_24_0_cgo_iro,
      yy_rsc_24_0_i_clka_en_d => yy_rsc_24_0_i_clka_en_d,
      yy_rsc_25_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_25_0_cgo_iro,
      yy_rsc_25_0_i_clka_en_d => yy_rsc_25_0_i_clka_en_d,
      yy_rsc_26_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_26_0_cgo_iro,
      yy_rsc_26_0_i_clka_en_d => yy_rsc_26_0_i_clka_en_d,
      yy_rsc_27_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_27_0_cgo_iro,
      yy_rsc_27_0_i_clka_en_d => yy_rsc_27_0_i_clka_en_d,
      yy_rsc_28_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_28_0_cgo_iro,
      yy_rsc_28_0_i_clka_en_d => yy_rsc_28_0_i_clka_en_d,
      yy_rsc_29_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_29_0_cgo_iro,
      yy_rsc_29_0_i_clka_en_d => yy_rsc_29_0_i_clka_en_d,
      yy_rsc_30_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_30_0_cgo_iro,
      yy_rsc_30_0_i_clka_en_d => yy_rsc_30_0_i_clka_en_d,
      yy_rsc_31_0_cgo_iro => hybrid_core_wait_dp_inst_yy_rsc_31_0_cgo_iro,
      yy_rsc_31_0_i_clka_en_d => yy_rsc_31_0_i_clka_en_d,
      ensig_cgo_iro => and_1109_rmff,
      S34_OUTER_LOOP_for_tf_mul_cmp_z => hybrid_core_wait_dp_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z,
      ensig_cgo_iro_1 => hybrid_core_wait_dp_inst_ensig_cgo_iro_1,
      core_wen => core_wen,
      xx_rsc_0_0_cgo => reg_xx_rsc_0_0_cgo_cse,
      xx_rsc_1_0_cgo => reg_xx_rsc_1_0_cgo_cse,
      xx_rsc_2_0_cgo => reg_xx_rsc_2_0_cgo_cse,
      xx_rsc_3_0_cgo => reg_xx_rsc_3_0_cgo_cse,
      xx_rsc_4_0_cgo => reg_xx_rsc_4_0_cgo_cse,
      xx_rsc_5_0_cgo => reg_xx_rsc_5_0_cgo_cse,
      xx_rsc_6_0_cgo => reg_xx_rsc_6_0_cgo_cse,
      xx_rsc_7_0_cgo => reg_xx_rsc_7_0_cgo_cse,
      xx_rsc_8_0_cgo => reg_xx_rsc_8_0_cgo_cse,
      xx_rsc_9_0_cgo => reg_xx_rsc_9_0_cgo_cse,
      xx_rsc_10_0_cgo => reg_xx_rsc_10_0_cgo_cse,
      xx_rsc_11_0_cgo => reg_xx_rsc_11_0_cgo_cse,
      xx_rsc_12_0_cgo => reg_xx_rsc_12_0_cgo_cse,
      xx_rsc_13_0_cgo => reg_xx_rsc_13_0_cgo_cse,
      xx_rsc_14_0_cgo => reg_xx_rsc_14_0_cgo_cse,
      xx_rsc_15_0_cgo => reg_xx_rsc_15_0_cgo_cse,
      xx_rsc_16_0_cgo => reg_xx_rsc_16_0_cgo_cse,
      xx_rsc_17_0_cgo => reg_xx_rsc_17_0_cgo_cse,
      xx_rsc_18_0_cgo => reg_xx_rsc_18_0_cgo_cse,
      xx_rsc_19_0_cgo => reg_xx_rsc_19_0_cgo_cse,
      xx_rsc_20_0_cgo => reg_xx_rsc_20_0_cgo_cse,
      xx_rsc_21_0_cgo => reg_xx_rsc_21_0_cgo_cse,
      xx_rsc_22_0_cgo => reg_xx_rsc_22_0_cgo_cse,
      xx_rsc_23_0_cgo => reg_xx_rsc_23_0_cgo_cse,
      xx_rsc_24_0_cgo => reg_xx_rsc_24_0_cgo_cse,
      xx_rsc_25_0_cgo => reg_xx_rsc_25_0_cgo_cse,
      xx_rsc_26_0_cgo => reg_xx_rsc_26_0_cgo_cse,
      xx_rsc_27_0_cgo => reg_xx_rsc_27_0_cgo_cse,
      xx_rsc_28_0_cgo => reg_xx_rsc_28_0_cgo_cse,
      xx_rsc_29_0_cgo => reg_xx_rsc_29_0_cgo_cse,
      xx_rsc_30_0_cgo => reg_xx_rsc_30_0_cgo_cse,
      xx_rsc_31_0_cgo => reg_xx_rsc_31_0_cgo_cse,
      yy_rsc_0_0_cgo => reg_yy_rsc_0_0_cgo_cse,
      yy_rsc_1_0_cgo => reg_yy_rsc_1_0_cgo_cse,
      yy_rsc_2_0_cgo => reg_yy_rsc_2_0_cgo_cse,
      yy_rsc_3_0_cgo => reg_yy_rsc_3_0_cgo_cse,
      yy_rsc_4_0_cgo => reg_yy_rsc_4_0_cgo_cse,
      yy_rsc_5_0_cgo => reg_yy_rsc_5_0_cgo_cse,
      yy_rsc_6_0_cgo => reg_yy_rsc_6_0_cgo_cse,
      yy_rsc_7_0_cgo => reg_yy_rsc_7_0_cgo_cse,
      yy_rsc_8_0_cgo => reg_yy_rsc_8_0_cgo_cse,
      yy_rsc_9_0_cgo => reg_yy_rsc_9_0_cgo_cse,
      yy_rsc_10_0_cgo => reg_yy_rsc_10_0_cgo_cse,
      yy_rsc_11_0_cgo => reg_yy_rsc_11_0_cgo_cse,
      yy_rsc_12_0_cgo => reg_yy_rsc_12_0_cgo_cse,
      yy_rsc_13_0_cgo => reg_yy_rsc_13_0_cgo_cse,
      yy_rsc_14_0_cgo => reg_yy_rsc_14_0_cgo_cse,
      yy_rsc_15_0_cgo => reg_yy_rsc_15_0_cgo_cse,
      yy_rsc_16_0_cgo => reg_yy_rsc_16_0_cgo_cse,
      yy_rsc_17_0_cgo => reg_yy_rsc_17_0_cgo_cse,
      yy_rsc_18_0_cgo => reg_yy_rsc_18_0_cgo_cse,
      yy_rsc_19_0_cgo => reg_yy_rsc_19_0_cgo_cse,
      yy_rsc_20_0_cgo => reg_yy_rsc_20_0_cgo_cse,
      yy_rsc_21_0_cgo => reg_yy_rsc_21_0_cgo_cse,
      yy_rsc_22_0_cgo => reg_yy_rsc_22_0_cgo_cse,
      yy_rsc_23_0_cgo => reg_yy_rsc_23_0_cgo_cse,
      yy_rsc_24_0_cgo => reg_yy_rsc_24_0_cgo_cse,
      yy_rsc_25_0_cgo => reg_yy_rsc_25_0_cgo_cse,
      yy_rsc_26_0_cgo => reg_yy_rsc_26_0_cgo_cse,
      yy_rsc_27_0_cgo => reg_yy_rsc_27_0_cgo_cse,
      yy_rsc_28_0_cgo => reg_yy_rsc_28_0_cgo_cse,
      yy_rsc_29_0_cgo => reg_yy_rsc_29_0_cgo_cse,
      yy_rsc_30_0_cgo => reg_yy_rsc_30_0_cgo_cse,
      yy_rsc_31_0_cgo => reg_yy_rsc_31_0_cgo_cse,
      ensig_cgo => reg_ensig_cgo_cse,
      mult_12_z_mul_cmp_en => mult_12_z_mul_cmp_en,
      S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg => hybrid_core_wait_dp_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg,
      ensig_cgo_1 => reg_ensig_cgo_1_cse,
      mult_z_mul_cmp_en => mult_z_mul_cmp_en
    );
  hybrid_core_wait_dp_inst_xx_rsc_0_0_cgo_iro <= NOT mux_138_itm;
  hybrid_core_wait_dp_inst_xx_rsc_4_0_cgo_iro <= NOT mux_357_itm;
  hybrid_core_wait_dp_inst_xx_rsc_8_0_cgo_iro <= NOT mux_566_itm;
  hybrid_core_wait_dp_inst_xx_rsc_12_0_cgo_iro <= NOT mux_772_itm;
  hybrid_core_wait_dp_inst_xx_rsc_16_0_cgo_iro <= NOT mux_979_itm;
  hybrid_core_wait_dp_inst_xx_rsc_20_0_cgo_iro <= NOT mux_1196_itm;
  hybrid_core_wait_dp_inst_xx_rsc_24_0_cgo_iro <= NOT mux_1414_itm;
  hybrid_core_wait_dp_inst_xx_rsc_28_0_cgo_iro <= NOT mux_1631_itm;
  hybrid_core_wait_dp_inst_yy_rsc_0_0_cgo_iro <= NOT mux_1843_itm;
  hybrid_core_wait_dp_inst_yy_rsc_1_0_cgo_iro <= NOT mux_1902_itm;
  hybrid_core_wait_dp_inst_yy_rsc_2_0_cgo_iro <= NOT mux_1950_itm;
  hybrid_core_wait_dp_inst_yy_rsc_3_0_cgo_iro <= NOT mux_2010_itm;
  hybrid_core_wait_dp_inst_yy_rsc_4_0_cgo_iro <= NOT mux_2075_itm;
  hybrid_core_wait_dp_inst_yy_rsc_5_0_cgo_iro <= NOT mux_2130_itm;
  hybrid_core_wait_dp_inst_yy_rsc_6_0_cgo_iro <= NOT mux_2175_itm;
  hybrid_core_wait_dp_inst_yy_rsc_7_0_cgo_iro <= NOT mux_2233_itm;
  hybrid_core_wait_dp_inst_yy_rsc_8_0_cgo_iro <= NOT mux_2295_itm;
  hybrid_core_wait_dp_inst_yy_rsc_9_0_cgo_iro <= NOT mux_2350_itm;
  hybrid_core_wait_dp_inst_yy_rsc_10_0_cgo_iro <= NOT mux_2395_itm;
  hybrid_core_wait_dp_inst_yy_rsc_11_0_cgo_iro <= NOT mux_2453_itm;
  hybrid_core_wait_dp_inst_yy_rsc_12_0_cgo_iro <= NOT mux_2515_itm;
  hybrid_core_wait_dp_inst_yy_rsc_13_0_cgo_iro <= NOT mux_2570_itm;
  hybrid_core_wait_dp_inst_yy_rsc_14_0_cgo_iro <= NOT mux_2615_itm;
  hybrid_core_wait_dp_inst_yy_rsc_15_0_cgo_iro <= NOT mux_2673_itm;
  hybrid_core_wait_dp_inst_yy_rsc_16_0_cgo_iro <= NOT mux_2735_itm;
  hybrid_core_wait_dp_inst_yy_rsc_17_0_cgo_iro <= NOT mux_2790_itm;
  hybrid_core_wait_dp_inst_yy_rsc_18_0_cgo_iro <= NOT mux_2835_itm;
  hybrid_core_wait_dp_inst_yy_rsc_19_0_cgo_iro <= NOT mux_2893_itm;
  hybrid_core_wait_dp_inst_yy_rsc_20_0_cgo_iro <= NOT mux_2955_itm;
  hybrid_core_wait_dp_inst_yy_rsc_21_0_cgo_iro <= NOT mux_3010_itm;
  hybrid_core_wait_dp_inst_yy_rsc_22_0_cgo_iro <= NOT mux_3055_itm;
  hybrid_core_wait_dp_inst_yy_rsc_23_0_cgo_iro <= NOT mux_3113_itm;
  hybrid_core_wait_dp_inst_yy_rsc_24_0_cgo_iro <= NOT mux_3175_itm;
  hybrid_core_wait_dp_inst_yy_rsc_25_0_cgo_iro <= NOT mux_3230_itm;
  hybrid_core_wait_dp_inst_yy_rsc_26_0_cgo_iro <= NOT mux_3275_itm;
  hybrid_core_wait_dp_inst_yy_rsc_27_0_cgo_iro <= NOT mux_3333_itm;
  hybrid_core_wait_dp_inst_yy_rsc_28_0_cgo_iro <= NOT mux_3395_itm;
  hybrid_core_wait_dp_inst_yy_rsc_29_0_cgo_iro <= NOT mux_3450_itm;
  hybrid_core_wait_dp_inst_yy_rsc_30_0_cgo_iro <= NOT mux_3495_itm;
  hybrid_core_wait_dp_inst_yy_rsc_31_0_cgo_iro <= NOT mux_3553_itm;
  hybrid_core_wait_dp_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z <= S34_OUTER_LOOP_for_tf_mul_cmp_z;
  hybrid_core_wait_dp_inst_ensig_cgo_iro_1 <= NOT mux_3669_itm;
  S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg <= hybrid_core_wait_dp_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg;

  hybrid_core_twiddle_h_rsci_1_inst : hybrid_core_twiddle_h_rsci_1
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsci_adrb_d => hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_adrb_d,
      twiddle_h_rsci_qb_d => hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_qb_d,
      twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_h_rsci_oswt => reg_twiddle_rsci_oswt_cse,
      twiddle_h_rsci_adrb_d_core => hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_adrb_d_core,
      twiddle_h_rsci_qb_d_mxwt => hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_qb_d_mxwt,
      twiddle_h_rsci_oswt_pff => mux_111_rmff
    );
  twiddle_h_rsci_adrb_d_reg <= hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_adrb_d;
  hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_qb_d <= twiddle_h_rsci_qb_d;
  hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_adrb_d_core <= '0' & S2_INNER_LOOP1_tfh_S2_INNER_LOOP1_tfh_mux_rmff
      & S2_INNER_LOOP1_tfh_mux1h_rmff;
  twiddle_h_rsci_qb_d_mxwt <= hybrid_core_twiddle_h_rsci_1_inst_twiddle_h_rsci_qb_d_mxwt;

  hybrid_core_revArr_rsci_inst : hybrid_core_revArr_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      revArr_rsc_s_tdone => revArr_rsc_s_tdone,
      revArr_rsc_tr_write_done => revArr_rsc_tr_write_done,
      revArr_rsc_RREADY => revArr_rsc_RREADY,
      revArr_rsc_RVALID => revArr_rsc_RVALID,
      revArr_rsc_RUSER => revArr_rsc_RUSER,
      revArr_rsc_RLAST => revArr_rsc_RLAST,
      revArr_rsc_RRESP => hybrid_core_revArr_rsci_inst_revArr_rsc_RRESP,
      revArr_rsc_RDATA => hybrid_core_revArr_rsci_inst_revArr_rsc_RDATA,
      revArr_rsc_RID => revArr_rsc_RID,
      revArr_rsc_ARREADY => revArr_rsc_ARREADY,
      revArr_rsc_ARVALID => revArr_rsc_ARVALID,
      revArr_rsc_ARUSER => revArr_rsc_ARUSER,
      revArr_rsc_ARREGION => hybrid_core_revArr_rsci_inst_revArr_rsc_ARREGION,
      revArr_rsc_ARQOS => hybrid_core_revArr_rsci_inst_revArr_rsc_ARQOS,
      revArr_rsc_ARPROT => hybrid_core_revArr_rsci_inst_revArr_rsc_ARPROT,
      revArr_rsc_ARCACHE => hybrid_core_revArr_rsci_inst_revArr_rsc_ARCACHE,
      revArr_rsc_ARLOCK => revArr_rsc_ARLOCK,
      revArr_rsc_ARBURST => hybrid_core_revArr_rsci_inst_revArr_rsc_ARBURST,
      revArr_rsc_ARSIZE => hybrid_core_revArr_rsci_inst_revArr_rsc_ARSIZE,
      revArr_rsc_ARLEN => hybrid_core_revArr_rsci_inst_revArr_rsc_ARLEN,
      revArr_rsc_ARADDR => hybrid_core_revArr_rsci_inst_revArr_rsc_ARADDR,
      revArr_rsc_ARID => revArr_rsc_ARID,
      revArr_rsc_BREADY => revArr_rsc_BREADY,
      revArr_rsc_BVALID => revArr_rsc_BVALID,
      revArr_rsc_BUSER => revArr_rsc_BUSER,
      revArr_rsc_BRESP => hybrid_core_revArr_rsci_inst_revArr_rsc_BRESP,
      revArr_rsc_BID => revArr_rsc_BID,
      revArr_rsc_WREADY => revArr_rsc_WREADY,
      revArr_rsc_WVALID => revArr_rsc_WVALID,
      revArr_rsc_WUSER => revArr_rsc_WUSER,
      revArr_rsc_WLAST => revArr_rsc_WLAST,
      revArr_rsc_WSTRB => hybrid_core_revArr_rsci_inst_revArr_rsc_WSTRB,
      revArr_rsc_WDATA => hybrid_core_revArr_rsci_inst_revArr_rsc_WDATA,
      revArr_rsc_AWREADY => revArr_rsc_AWREADY,
      revArr_rsc_AWVALID => revArr_rsc_AWVALID,
      revArr_rsc_AWUSER => revArr_rsc_AWUSER,
      revArr_rsc_AWREGION => hybrid_core_revArr_rsci_inst_revArr_rsc_AWREGION,
      revArr_rsc_AWQOS => hybrid_core_revArr_rsci_inst_revArr_rsc_AWQOS,
      revArr_rsc_AWPROT => hybrid_core_revArr_rsci_inst_revArr_rsc_AWPROT,
      revArr_rsc_AWCACHE => hybrid_core_revArr_rsci_inst_revArr_rsc_AWCACHE,
      revArr_rsc_AWLOCK => revArr_rsc_AWLOCK,
      revArr_rsc_AWBURST => hybrid_core_revArr_rsci_inst_revArr_rsc_AWBURST,
      revArr_rsc_AWSIZE => hybrid_core_revArr_rsci_inst_revArr_rsc_AWSIZE,
      revArr_rsc_AWLEN => hybrid_core_revArr_rsci_inst_revArr_rsc_AWLEN,
      revArr_rsc_AWADDR => hybrid_core_revArr_rsci_inst_revArr_rsc_AWADDR,
      revArr_rsc_AWID => revArr_rsc_AWID,
      core_wen => core_wen,
      revArr_rsci_oswt => reg_revArr_rsci_oswt_cse,
      revArr_rsci_wen_comp => revArr_rsci_wen_comp,
      revArr_rsci_s_raddr_core => hybrid_core_revArr_rsci_inst_revArr_rsci_s_raddr_core,
      revArr_rsci_s_din_mxwt => hybrid_core_revArr_rsci_inst_revArr_rsci_s_din_mxwt
    );
  revArr_rsc_RRESP <= hybrid_core_revArr_rsci_inst_revArr_rsc_RRESP;
  revArr_rsc_RDATA <= hybrid_core_revArr_rsci_inst_revArr_rsc_RDATA;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARREGION <= revArr_rsc_ARREGION;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARQOS <= revArr_rsc_ARQOS;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARPROT <= revArr_rsc_ARPROT;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARCACHE <= revArr_rsc_ARCACHE;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARBURST <= revArr_rsc_ARBURST;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARSIZE <= revArr_rsc_ARSIZE;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARLEN <= revArr_rsc_ARLEN;
  hybrid_core_revArr_rsci_inst_revArr_rsc_ARADDR <= revArr_rsc_ARADDR;
  revArr_rsc_BRESP <= hybrid_core_revArr_rsci_inst_revArr_rsc_BRESP;
  hybrid_core_revArr_rsci_inst_revArr_rsc_WSTRB <= revArr_rsc_WSTRB;
  hybrid_core_revArr_rsci_inst_revArr_rsc_WDATA <= revArr_rsc_WDATA;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWREGION <= revArr_rsc_AWREGION;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWQOS <= revArr_rsc_AWQOS;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWPROT <= revArr_rsc_AWPROT;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWCACHE <= revArr_rsc_AWCACHE;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWBURST <= revArr_rsc_AWBURST;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWSIZE <= revArr_rsc_AWSIZE;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWLEN <= revArr_rsc_AWLEN;
  hybrid_core_revArr_rsci_inst_revArr_rsc_AWADDR <= revArr_rsc_AWADDR;
  hybrid_core_revArr_rsci_inst_revArr_rsci_s_raddr_core <= revArr_rsci_s_raddr_core_4
      & revArr_rsci_s_raddr_core_3_0;
  revArr_rsci_s_din_mxwt <= hybrid_core_revArr_rsci_inst_revArr_rsci_s_din_mxwt;

  hybrid_core_tw_rsci_inst : hybrid_core_tw_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      tw_rsc_s_tdone => tw_rsc_s_tdone,
      tw_rsc_tr_write_done => tw_rsc_tr_write_done,
      tw_rsc_RREADY => tw_rsc_RREADY,
      tw_rsc_RVALID => tw_rsc_RVALID,
      tw_rsc_RUSER => tw_rsc_RUSER,
      tw_rsc_RLAST => tw_rsc_RLAST,
      tw_rsc_RRESP => hybrid_core_tw_rsci_inst_tw_rsc_RRESP,
      tw_rsc_RDATA => hybrid_core_tw_rsci_inst_tw_rsc_RDATA,
      tw_rsc_RID => tw_rsc_RID,
      tw_rsc_ARREADY => tw_rsc_ARREADY,
      tw_rsc_ARVALID => tw_rsc_ARVALID,
      tw_rsc_ARUSER => tw_rsc_ARUSER,
      tw_rsc_ARREGION => hybrid_core_tw_rsci_inst_tw_rsc_ARREGION,
      tw_rsc_ARQOS => hybrid_core_tw_rsci_inst_tw_rsc_ARQOS,
      tw_rsc_ARPROT => hybrid_core_tw_rsci_inst_tw_rsc_ARPROT,
      tw_rsc_ARCACHE => hybrid_core_tw_rsci_inst_tw_rsc_ARCACHE,
      tw_rsc_ARLOCK => tw_rsc_ARLOCK,
      tw_rsc_ARBURST => hybrid_core_tw_rsci_inst_tw_rsc_ARBURST,
      tw_rsc_ARSIZE => hybrid_core_tw_rsci_inst_tw_rsc_ARSIZE,
      tw_rsc_ARLEN => hybrid_core_tw_rsci_inst_tw_rsc_ARLEN,
      tw_rsc_ARADDR => hybrid_core_tw_rsci_inst_tw_rsc_ARADDR,
      tw_rsc_ARID => tw_rsc_ARID,
      tw_rsc_BREADY => tw_rsc_BREADY,
      tw_rsc_BVALID => tw_rsc_BVALID,
      tw_rsc_BUSER => tw_rsc_BUSER,
      tw_rsc_BRESP => hybrid_core_tw_rsci_inst_tw_rsc_BRESP,
      tw_rsc_BID => tw_rsc_BID,
      tw_rsc_WREADY => tw_rsc_WREADY,
      tw_rsc_WVALID => tw_rsc_WVALID,
      tw_rsc_WUSER => tw_rsc_WUSER,
      tw_rsc_WLAST => tw_rsc_WLAST,
      tw_rsc_WSTRB => hybrid_core_tw_rsci_inst_tw_rsc_WSTRB,
      tw_rsc_WDATA => hybrid_core_tw_rsci_inst_tw_rsc_WDATA,
      tw_rsc_AWREADY => tw_rsc_AWREADY,
      tw_rsc_AWVALID => tw_rsc_AWVALID,
      tw_rsc_AWUSER => tw_rsc_AWUSER,
      tw_rsc_AWREGION => hybrid_core_tw_rsci_inst_tw_rsc_AWREGION,
      tw_rsc_AWQOS => hybrid_core_tw_rsci_inst_tw_rsc_AWQOS,
      tw_rsc_AWPROT => hybrid_core_tw_rsci_inst_tw_rsc_AWPROT,
      tw_rsc_AWCACHE => hybrid_core_tw_rsci_inst_tw_rsc_AWCACHE,
      tw_rsc_AWLOCK => tw_rsc_AWLOCK,
      tw_rsc_AWBURST => hybrid_core_tw_rsci_inst_tw_rsc_AWBURST,
      tw_rsc_AWSIZE => hybrid_core_tw_rsci_inst_tw_rsc_AWSIZE,
      tw_rsc_AWLEN => hybrid_core_tw_rsci_inst_tw_rsc_AWLEN,
      tw_rsc_AWADDR => hybrid_core_tw_rsci_inst_tw_rsc_AWADDR,
      tw_rsc_AWID => tw_rsc_AWID,
      core_wen => core_wen,
      tw_rsci_oswt => reg_tw_rsci_oswt_cse,
      tw_rsci_wen_comp => tw_rsci_wen_comp,
      tw_rsci_s_raddr_core => hybrid_core_tw_rsci_inst_tw_rsci_s_raddr_core,
      tw_rsci_s_din_mxwt => hybrid_core_tw_rsci_inst_tw_rsci_s_din_mxwt
    );
  tw_rsc_RRESP <= hybrid_core_tw_rsci_inst_tw_rsc_RRESP;
  tw_rsc_RDATA <= hybrid_core_tw_rsci_inst_tw_rsc_RDATA;
  hybrid_core_tw_rsci_inst_tw_rsc_ARREGION <= tw_rsc_ARREGION;
  hybrid_core_tw_rsci_inst_tw_rsc_ARQOS <= tw_rsc_ARQOS;
  hybrid_core_tw_rsci_inst_tw_rsc_ARPROT <= tw_rsc_ARPROT;
  hybrid_core_tw_rsci_inst_tw_rsc_ARCACHE <= tw_rsc_ARCACHE;
  hybrid_core_tw_rsci_inst_tw_rsc_ARBURST <= tw_rsc_ARBURST;
  hybrid_core_tw_rsci_inst_tw_rsc_ARSIZE <= tw_rsc_ARSIZE;
  hybrid_core_tw_rsci_inst_tw_rsc_ARLEN <= tw_rsc_ARLEN;
  hybrid_core_tw_rsci_inst_tw_rsc_ARADDR <= tw_rsc_ARADDR;
  tw_rsc_BRESP <= hybrid_core_tw_rsci_inst_tw_rsc_BRESP;
  hybrid_core_tw_rsci_inst_tw_rsc_WSTRB <= tw_rsc_WSTRB;
  hybrid_core_tw_rsci_inst_tw_rsc_WDATA <= tw_rsc_WDATA;
  hybrid_core_tw_rsci_inst_tw_rsc_AWREGION <= tw_rsc_AWREGION;
  hybrid_core_tw_rsci_inst_tw_rsc_AWQOS <= tw_rsc_AWQOS;
  hybrid_core_tw_rsci_inst_tw_rsc_AWPROT <= tw_rsc_AWPROT;
  hybrid_core_tw_rsci_inst_tw_rsc_AWCACHE <= tw_rsc_AWCACHE;
  hybrid_core_tw_rsci_inst_tw_rsc_AWBURST <= tw_rsc_AWBURST;
  hybrid_core_tw_rsci_inst_tw_rsc_AWSIZE <= tw_rsc_AWSIZE;
  hybrid_core_tw_rsci_inst_tw_rsc_AWLEN <= tw_rsc_AWLEN;
  hybrid_core_tw_rsci_inst_tw_rsc_AWADDR <= tw_rsc_AWADDR;
  hybrid_core_tw_rsci_inst_tw_rsci_s_raddr_core <= reg_tw_rsci_s_raddr_core_cse;
  tw_rsci_s_din_mxwt <= hybrid_core_tw_rsci_inst_tw_rsci_s_din_mxwt;

  hybrid_core_tw_h_rsci_inst : hybrid_core_tw_h_rsci
    PORT MAP(
      clk => clk,
      rst => rst,
      tw_h_rsc_s_tdone => tw_h_rsc_s_tdone,
      tw_h_rsc_tr_write_done => tw_h_rsc_tr_write_done,
      tw_h_rsc_RREADY => tw_h_rsc_RREADY,
      tw_h_rsc_RVALID => tw_h_rsc_RVALID,
      tw_h_rsc_RUSER => tw_h_rsc_RUSER,
      tw_h_rsc_RLAST => tw_h_rsc_RLAST,
      tw_h_rsc_RRESP => hybrid_core_tw_h_rsci_inst_tw_h_rsc_RRESP,
      tw_h_rsc_RDATA => hybrid_core_tw_h_rsci_inst_tw_h_rsc_RDATA,
      tw_h_rsc_RID => tw_h_rsc_RID,
      tw_h_rsc_ARREADY => tw_h_rsc_ARREADY,
      tw_h_rsc_ARVALID => tw_h_rsc_ARVALID,
      tw_h_rsc_ARUSER => tw_h_rsc_ARUSER,
      tw_h_rsc_ARREGION => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARREGION,
      tw_h_rsc_ARQOS => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARQOS,
      tw_h_rsc_ARPROT => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARPROT,
      tw_h_rsc_ARCACHE => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARCACHE,
      tw_h_rsc_ARLOCK => tw_h_rsc_ARLOCK,
      tw_h_rsc_ARBURST => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARBURST,
      tw_h_rsc_ARSIZE => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARSIZE,
      tw_h_rsc_ARLEN => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARLEN,
      tw_h_rsc_ARADDR => hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARADDR,
      tw_h_rsc_ARID => tw_h_rsc_ARID,
      tw_h_rsc_BREADY => tw_h_rsc_BREADY,
      tw_h_rsc_BVALID => tw_h_rsc_BVALID,
      tw_h_rsc_BUSER => tw_h_rsc_BUSER,
      tw_h_rsc_BRESP => hybrid_core_tw_h_rsci_inst_tw_h_rsc_BRESP,
      tw_h_rsc_BID => tw_h_rsc_BID,
      tw_h_rsc_WREADY => tw_h_rsc_WREADY,
      tw_h_rsc_WVALID => tw_h_rsc_WVALID,
      tw_h_rsc_WUSER => tw_h_rsc_WUSER,
      tw_h_rsc_WLAST => tw_h_rsc_WLAST,
      tw_h_rsc_WSTRB => hybrid_core_tw_h_rsci_inst_tw_h_rsc_WSTRB,
      tw_h_rsc_WDATA => hybrid_core_tw_h_rsci_inst_tw_h_rsc_WDATA,
      tw_h_rsc_AWREADY => tw_h_rsc_AWREADY,
      tw_h_rsc_AWVALID => tw_h_rsc_AWVALID,
      tw_h_rsc_AWUSER => tw_h_rsc_AWUSER,
      tw_h_rsc_AWREGION => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWREGION,
      tw_h_rsc_AWQOS => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWQOS,
      tw_h_rsc_AWPROT => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWPROT,
      tw_h_rsc_AWCACHE => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWCACHE,
      tw_h_rsc_AWLOCK => tw_h_rsc_AWLOCK,
      tw_h_rsc_AWBURST => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWBURST,
      tw_h_rsc_AWSIZE => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWSIZE,
      tw_h_rsc_AWLEN => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWLEN,
      tw_h_rsc_AWADDR => hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWADDR,
      tw_h_rsc_AWID => tw_h_rsc_AWID,
      core_wen => core_wen,
      tw_h_rsci_oswt => reg_tw_rsci_oswt_cse,
      tw_h_rsci_wen_comp => tw_h_rsci_wen_comp,
      tw_h_rsci_s_raddr_core => hybrid_core_tw_h_rsci_inst_tw_h_rsci_s_raddr_core,
      tw_h_rsci_s_din_mxwt => hybrid_core_tw_h_rsci_inst_tw_h_rsci_s_din_mxwt
    );
  tw_h_rsc_RRESP <= hybrid_core_tw_h_rsci_inst_tw_h_rsc_RRESP;
  tw_h_rsc_RDATA <= hybrid_core_tw_h_rsci_inst_tw_h_rsc_RDATA;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARREGION <= tw_h_rsc_ARREGION;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARQOS <= tw_h_rsc_ARQOS;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARPROT <= tw_h_rsc_ARPROT;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARCACHE <= tw_h_rsc_ARCACHE;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARBURST <= tw_h_rsc_ARBURST;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARSIZE <= tw_h_rsc_ARSIZE;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARLEN <= tw_h_rsc_ARLEN;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_ARADDR <= tw_h_rsc_ARADDR;
  tw_h_rsc_BRESP <= hybrid_core_tw_h_rsci_inst_tw_h_rsc_BRESP;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_WSTRB <= tw_h_rsc_WSTRB;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_WDATA <= tw_h_rsc_WDATA;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWREGION <= tw_h_rsc_AWREGION;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWQOS <= tw_h_rsc_AWQOS;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWPROT <= tw_h_rsc_AWPROT;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWCACHE <= tw_h_rsc_AWCACHE;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWBURST <= tw_h_rsc_AWBURST;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWSIZE <= tw_h_rsc_AWSIZE;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWLEN <= tw_h_rsc_AWLEN;
  hybrid_core_tw_h_rsci_inst_tw_h_rsc_AWADDR <= tw_h_rsc_AWADDR;
  hybrid_core_tw_h_rsci_inst_tw_h_rsci_s_raddr_core <= reg_tw_rsci_s_raddr_core_cse;
  tw_h_rsci_s_din_mxwt <= hybrid_core_tw_h_rsci_inst_tw_h_rsci_s_din_mxwt;

  hybrid_core_x_rsc_0_0_i_inst : hybrid_core_x_rsc_0_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_0_0_s_tdone => x_rsc_0_0_s_tdone,
      x_rsc_0_0_tr_write_done => x_rsc_0_0_tr_write_done,
      x_rsc_0_0_RREADY => x_rsc_0_0_RREADY,
      x_rsc_0_0_RVALID => x_rsc_0_0_RVALID,
      x_rsc_0_0_RUSER => x_rsc_0_0_RUSER,
      x_rsc_0_0_RLAST => x_rsc_0_0_RLAST,
      x_rsc_0_0_RRESP => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_RRESP,
      x_rsc_0_0_RDATA => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_RDATA,
      x_rsc_0_0_RID => x_rsc_0_0_RID,
      x_rsc_0_0_ARREADY => x_rsc_0_0_ARREADY,
      x_rsc_0_0_ARVALID => x_rsc_0_0_ARVALID,
      x_rsc_0_0_ARUSER => x_rsc_0_0_ARUSER,
      x_rsc_0_0_ARREGION => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARREGION,
      x_rsc_0_0_ARQOS => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARQOS,
      x_rsc_0_0_ARPROT => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARPROT,
      x_rsc_0_0_ARCACHE => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARCACHE,
      x_rsc_0_0_ARLOCK => x_rsc_0_0_ARLOCK,
      x_rsc_0_0_ARBURST => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARBURST,
      x_rsc_0_0_ARSIZE => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARSIZE,
      x_rsc_0_0_ARLEN => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARLEN,
      x_rsc_0_0_ARADDR => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARADDR,
      x_rsc_0_0_ARID => x_rsc_0_0_ARID,
      x_rsc_0_0_BREADY => x_rsc_0_0_BREADY,
      x_rsc_0_0_BVALID => x_rsc_0_0_BVALID,
      x_rsc_0_0_BUSER => x_rsc_0_0_BUSER,
      x_rsc_0_0_BRESP => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_BRESP,
      x_rsc_0_0_BID => x_rsc_0_0_BID,
      x_rsc_0_0_WREADY => x_rsc_0_0_WREADY,
      x_rsc_0_0_WVALID => x_rsc_0_0_WVALID,
      x_rsc_0_0_WUSER => x_rsc_0_0_WUSER,
      x_rsc_0_0_WLAST => x_rsc_0_0_WLAST,
      x_rsc_0_0_WSTRB => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_WSTRB,
      x_rsc_0_0_WDATA => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_WDATA,
      x_rsc_0_0_AWREADY => x_rsc_0_0_AWREADY,
      x_rsc_0_0_AWVALID => x_rsc_0_0_AWVALID,
      x_rsc_0_0_AWUSER => x_rsc_0_0_AWUSER,
      x_rsc_0_0_AWREGION => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWREGION,
      x_rsc_0_0_AWQOS => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWQOS,
      x_rsc_0_0_AWPROT => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWPROT,
      x_rsc_0_0_AWCACHE => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWCACHE,
      x_rsc_0_0_AWLOCK => x_rsc_0_0_AWLOCK,
      x_rsc_0_0_AWBURST => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWBURST,
      x_rsc_0_0_AWSIZE => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWSIZE,
      x_rsc_0_0_AWLEN => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWLEN,
      x_rsc_0_0_AWADDR => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWADDR,
      x_rsc_0_0_AWID => x_rsc_0_0_AWID,
      core_wen => core_wen,
      x_rsc_0_0_i_oswt => reg_x_rsc_0_0_i_oswt_cse,
      x_rsc_0_0_i_wen_comp => x_rsc_0_0_i_wen_comp,
      x_rsc_0_0_i_oswt_1 => reg_x_rsc_0_0_i_oswt_1_cse,
      x_rsc_0_0_i_wen_comp_1 => x_rsc_0_0_i_wen_comp_1,
      x_rsc_0_0_i_s_raddr_core => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_raddr_core,
      x_rsc_0_0_i_s_waddr_core => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_waddr_core,
      x_rsc_0_0_i_s_din_mxwt => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_din_mxwt,
      x_rsc_0_0_i_s_dout_core => hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_dout_core
    );
  x_rsc_0_0_RRESP <= hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_RRESP;
  x_rsc_0_0_RDATA <= hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_RDATA;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARREGION <= x_rsc_0_0_ARREGION;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARQOS <= x_rsc_0_0_ARQOS;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARPROT <= x_rsc_0_0_ARPROT;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARCACHE <= x_rsc_0_0_ARCACHE;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARBURST <= x_rsc_0_0_ARBURST;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARSIZE <= x_rsc_0_0_ARSIZE;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARLEN <= x_rsc_0_0_ARLEN;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_ARADDR <= x_rsc_0_0_ARADDR;
  x_rsc_0_0_BRESP <= hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_BRESP;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_WSTRB <= x_rsc_0_0_WSTRB;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_WDATA <= x_rsc_0_0_WDATA;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWREGION <= x_rsc_0_0_AWREGION;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWQOS <= x_rsc_0_0_AWQOS;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWPROT <= x_rsc_0_0_AWPROT;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWCACHE <= x_rsc_0_0_AWCACHE;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWBURST <= x_rsc_0_0_AWBURST;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWSIZE <= x_rsc_0_0_AWSIZE;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWLEN <= x_rsc_0_0_AWLEN;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_AWADDR <= x_rsc_0_0_AWADDR;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_0_0_i_s_din_mxwt <= hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_din_mxwt;
  hybrid_core_x_rsc_0_0_i_inst_x_rsc_0_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_1_0_i_inst : hybrid_core_x_rsc_1_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_1_0_s_tdone => x_rsc_1_0_s_tdone,
      x_rsc_1_0_tr_write_done => x_rsc_1_0_tr_write_done,
      x_rsc_1_0_RREADY => x_rsc_1_0_RREADY,
      x_rsc_1_0_RVALID => x_rsc_1_0_RVALID,
      x_rsc_1_0_RUSER => x_rsc_1_0_RUSER,
      x_rsc_1_0_RLAST => x_rsc_1_0_RLAST,
      x_rsc_1_0_RRESP => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_RRESP,
      x_rsc_1_0_RDATA => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_RDATA,
      x_rsc_1_0_RID => x_rsc_1_0_RID,
      x_rsc_1_0_ARREADY => x_rsc_1_0_ARREADY,
      x_rsc_1_0_ARVALID => x_rsc_1_0_ARVALID,
      x_rsc_1_0_ARUSER => x_rsc_1_0_ARUSER,
      x_rsc_1_0_ARREGION => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARREGION,
      x_rsc_1_0_ARQOS => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARQOS,
      x_rsc_1_0_ARPROT => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARPROT,
      x_rsc_1_0_ARCACHE => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARCACHE,
      x_rsc_1_0_ARLOCK => x_rsc_1_0_ARLOCK,
      x_rsc_1_0_ARBURST => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARBURST,
      x_rsc_1_0_ARSIZE => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARSIZE,
      x_rsc_1_0_ARLEN => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARLEN,
      x_rsc_1_0_ARADDR => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARADDR,
      x_rsc_1_0_ARID => x_rsc_1_0_ARID,
      x_rsc_1_0_BREADY => x_rsc_1_0_BREADY,
      x_rsc_1_0_BVALID => x_rsc_1_0_BVALID,
      x_rsc_1_0_BUSER => x_rsc_1_0_BUSER,
      x_rsc_1_0_BRESP => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_BRESP,
      x_rsc_1_0_BID => x_rsc_1_0_BID,
      x_rsc_1_0_WREADY => x_rsc_1_0_WREADY,
      x_rsc_1_0_WVALID => x_rsc_1_0_WVALID,
      x_rsc_1_0_WUSER => x_rsc_1_0_WUSER,
      x_rsc_1_0_WLAST => x_rsc_1_0_WLAST,
      x_rsc_1_0_WSTRB => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_WSTRB,
      x_rsc_1_0_WDATA => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_WDATA,
      x_rsc_1_0_AWREADY => x_rsc_1_0_AWREADY,
      x_rsc_1_0_AWVALID => x_rsc_1_0_AWVALID,
      x_rsc_1_0_AWUSER => x_rsc_1_0_AWUSER,
      x_rsc_1_0_AWREGION => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWREGION,
      x_rsc_1_0_AWQOS => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWQOS,
      x_rsc_1_0_AWPROT => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWPROT,
      x_rsc_1_0_AWCACHE => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWCACHE,
      x_rsc_1_0_AWLOCK => x_rsc_1_0_AWLOCK,
      x_rsc_1_0_AWBURST => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWBURST,
      x_rsc_1_0_AWSIZE => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWSIZE,
      x_rsc_1_0_AWLEN => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWLEN,
      x_rsc_1_0_AWADDR => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWADDR,
      x_rsc_1_0_AWID => x_rsc_1_0_AWID,
      core_wen => core_wen,
      x_rsc_1_0_i_oswt => reg_x_rsc_1_0_i_oswt_cse,
      x_rsc_1_0_i_wen_comp => x_rsc_1_0_i_wen_comp,
      x_rsc_1_0_i_oswt_1 => reg_x_rsc_1_0_i_oswt_1_cse,
      x_rsc_1_0_i_wen_comp_1 => x_rsc_1_0_i_wen_comp_1,
      x_rsc_1_0_i_s_raddr_core => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_raddr_core,
      x_rsc_1_0_i_s_waddr_core => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_waddr_core,
      x_rsc_1_0_i_s_din_mxwt => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_din_mxwt,
      x_rsc_1_0_i_s_dout_core => hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_dout_core
    );
  x_rsc_1_0_RRESP <= hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_RRESP;
  x_rsc_1_0_RDATA <= hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_RDATA;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARREGION <= x_rsc_1_0_ARREGION;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARQOS <= x_rsc_1_0_ARQOS;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARPROT <= x_rsc_1_0_ARPROT;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARCACHE <= x_rsc_1_0_ARCACHE;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARBURST <= x_rsc_1_0_ARBURST;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARSIZE <= x_rsc_1_0_ARSIZE;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARLEN <= x_rsc_1_0_ARLEN;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_ARADDR <= x_rsc_1_0_ARADDR;
  x_rsc_1_0_BRESP <= hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_BRESP;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_WSTRB <= x_rsc_1_0_WSTRB;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_WDATA <= x_rsc_1_0_WDATA;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWREGION <= x_rsc_1_0_AWREGION;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWQOS <= x_rsc_1_0_AWQOS;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWPROT <= x_rsc_1_0_AWPROT;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWCACHE <= x_rsc_1_0_AWCACHE;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWBURST <= x_rsc_1_0_AWBURST;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWSIZE <= x_rsc_1_0_AWSIZE;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWLEN <= x_rsc_1_0_AWLEN;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_AWADDR <= x_rsc_1_0_AWADDR;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_1_0_i_s_din_mxwt <= hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_din_mxwt;
  hybrid_core_x_rsc_1_0_i_inst_x_rsc_1_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_2_0_i_inst : hybrid_core_x_rsc_2_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_2_0_s_tdone => x_rsc_2_0_s_tdone,
      x_rsc_2_0_tr_write_done => x_rsc_2_0_tr_write_done,
      x_rsc_2_0_RREADY => x_rsc_2_0_RREADY,
      x_rsc_2_0_RVALID => x_rsc_2_0_RVALID,
      x_rsc_2_0_RUSER => x_rsc_2_0_RUSER,
      x_rsc_2_0_RLAST => x_rsc_2_0_RLAST,
      x_rsc_2_0_RRESP => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_RRESP,
      x_rsc_2_0_RDATA => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_RDATA,
      x_rsc_2_0_RID => x_rsc_2_0_RID,
      x_rsc_2_0_ARREADY => x_rsc_2_0_ARREADY,
      x_rsc_2_0_ARVALID => x_rsc_2_0_ARVALID,
      x_rsc_2_0_ARUSER => x_rsc_2_0_ARUSER,
      x_rsc_2_0_ARREGION => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARREGION,
      x_rsc_2_0_ARQOS => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARQOS,
      x_rsc_2_0_ARPROT => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARPROT,
      x_rsc_2_0_ARCACHE => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARCACHE,
      x_rsc_2_0_ARLOCK => x_rsc_2_0_ARLOCK,
      x_rsc_2_0_ARBURST => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARBURST,
      x_rsc_2_0_ARSIZE => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARSIZE,
      x_rsc_2_0_ARLEN => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARLEN,
      x_rsc_2_0_ARADDR => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARADDR,
      x_rsc_2_0_ARID => x_rsc_2_0_ARID,
      x_rsc_2_0_BREADY => x_rsc_2_0_BREADY,
      x_rsc_2_0_BVALID => x_rsc_2_0_BVALID,
      x_rsc_2_0_BUSER => x_rsc_2_0_BUSER,
      x_rsc_2_0_BRESP => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_BRESP,
      x_rsc_2_0_BID => x_rsc_2_0_BID,
      x_rsc_2_0_WREADY => x_rsc_2_0_WREADY,
      x_rsc_2_0_WVALID => x_rsc_2_0_WVALID,
      x_rsc_2_0_WUSER => x_rsc_2_0_WUSER,
      x_rsc_2_0_WLAST => x_rsc_2_0_WLAST,
      x_rsc_2_0_WSTRB => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_WSTRB,
      x_rsc_2_0_WDATA => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_WDATA,
      x_rsc_2_0_AWREADY => x_rsc_2_0_AWREADY,
      x_rsc_2_0_AWVALID => x_rsc_2_0_AWVALID,
      x_rsc_2_0_AWUSER => x_rsc_2_0_AWUSER,
      x_rsc_2_0_AWREGION => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWREGION,
      x_rsc_2_0_AWQOS => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWQOS,
      x_rsc_2_0_AWPROT => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWPROT,
      x_rsc_2_0_AWCACHE => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWCACHE,
      x_rsc_2_0_AWLOCK => x_rsc_2_0_AWLOCK,
      x_rsc_2_0_AWBURST => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWBURST,
      x_rsc_2_0_AWSIZE => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWSIZE,
      x_rsc_2_0_AWLEN => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWLEN,
      x_rsc_2_0_AWADDR => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWADDR,
      x_rsc_2_0_AWID => x_rsc_2_0_AWID,
      core_wen => core_wen,
      x_rsc_2_0_i_oswt => reg_x_rsc_2_0_i_oswt_cse,
      x_rsc_2_0_i_wen_comp => x_rsc_2_0_i_wen_comp,
      x_rsc_2_0_i_oswt_1 => reg_x_rsc_2_0_i_oswt_1_cse,
      x_rsc_2_0_i_wen_comp_1 => x_rsc_2_0_i_wen_comp_1,
      x_rsc_2_0_i_s_raddr_core => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_raddr_core,
      x_rsc_2_0_i_s_waddr_core => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_waddr_core,
      x_rsc_2_0_i_s_din_mxwt => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_din_mxwt,
      x_rsc_2_0_i_s_dout_core => hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_dout_core
    );
  x_rsc_2_0_RRESP <= hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_RRESP;
  x_rsc_2_0_RDATA <= hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_RDATA;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARREGION <= x_rsc_2_0_ARREGION;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARQOS <= x_rsc_2_0_ARQOS;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARPROT <= x_rsc_2_0_ARPROT;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARCACHE <= x_rsc_2_0_ARCACHE;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARBURST <= x_rsc_2_0_ARBURST;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARSIZE <= x_rsc_2_0_ARSIZE;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARLEN <= x_rsc_2_0_ARLEN;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_ARADDR <= x_rsc_2_0_ARADDR;
  x_rsc_2_0_BRESP <= hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_BRESP;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_WSTRB <= x_rsc_2_0_WSTRB;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_WDATA <= x_rsc_2_0_WDATA;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWREGION <= x_rsc_2_0_AWREGION;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWQOS <= x_rsc_2_0_AWQOS;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWPROT <= x_rsc_2_0_AWPROT;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWCACHE <= x_rsc_2_0_AWCACHE;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWBURST <= x_rsc_2_0_AWBURST;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWSIZE <= x_rsc_2_0_AWSIZE;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWLEN <= x_rsc_2_0_AWLEN;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_AWADDR <= x_rsc_2_0_AWADDR;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_2_0_i_s_din_mxwt <= hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_din_mxwt;
  hybrid_core_x_rsc_2_0_i_inst_x_rsc_2_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_3_0_i_inst : hybrid_core_x_rsc_3_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_3_0_s_tdone => x_rsc_3_0_s_tdone,
      x_rsc_3_0_tr_write_done => x_rsc_3_0_tr_write_done,
      x_rsc_3_0_RREADY => x_rsc_3_0_RREADY,
      x_rsc_3_0_RVALID => x_rsc_3_0_RVALID,
      x_rsc_3_0_RUSER => x_rsc_3_0_RUSER,
      x_rsc_3_0_RLAST => x_rsc_3_0_RLAST,
      x_rsc_3_0_RRESP => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_RRESP,
      x_rsc_3_0_RDATA => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_RDATA,
      x_rsc_3_0_RID => x_rsc_3_0_RID,
      x_rsc_3_0_ARREADY => x_rsc_3_0_ARREADY,
      x_rsc_3_0_ARVALID => x_rsc_3_0_ARVALID,
      x_rsc_3_0_ARUSER => x_rsc_3_0_ARUSER,
      x_rsc_3_0_ARREGION => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARREGION,
      x_rsc_3_0_ARQOS => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARQOS,
      x_rsc_3_0_ARPROT => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARPROT,
      x_rsc_3_0_ARCACHE => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARCACHE,
      x_rsc_3_0_ARLOCK => x_rsc_3_0_ARLOCK,
      x_rsc_3_0_ARBURST => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARBURST,
      x_rsc_3_0_ARSIZE => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARSIZE,
      x_rsc_3_0_ARLEN => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARLEN,
      x_rsc_3_0_ARADDR => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARADDR,
      x_rsc_3_0_ARID => x_rsc_3_0_ARID,
      x_rsc_3_0_BREADY => x_rsc_3_0_BREADY,
      x_rsc_3_0_BVALID => x_rsc_3_0_BVALID,
      x_rsc_3_0_BUSER => x_rsc_3_0_BUSER,
      x_rsc_3_0_BRESP => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_BRESP,
      x_rsc_3_0_BID => x_rsc_3_0_BID,
      x_rsc_3_0_WREADY => x_rsc_3_0_WREADY,
      x_rsc_3_0_WVALID => x_rsc_3_0_WVALID,
      x_rsc_3_0_WUSER => x_rsc_3_0_WUSER,
      x_rsc_3_0_WLAST => x_rsc_3_0_WLAST,
      x_rsc_3_0_WSTRB => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_WSTRB,
      x_rsc_3_0_WDATA => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_WDATA,
      x_rsc_3_0_AWREADY => x_rsc_3_0_AWREADY,
      x_rsc_3_0_AWVALID => x_rsc_3_0_AWVALID,
      x_rsc_3_0_AWUSER => x_rsc_3_0_AWUSER,
      x_rsc_3_0_AWREGION => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWREGION,
      x_rsc_3_0_AWQOS => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWQOS,
      x_rsc_3_0_AWPROT => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWPROT,
      x_rsc_3_0_AWCACHE => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWCACHE,
      x_rsc_3_0_AWLOCK => x_rsc_3_0_AWLOCK,
      x_rsc_3_0_AWBURST => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWBURST,
      x_rsc_3_0_AWSIZE => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWSIZE,
      x_rsc_3_0_AWLEN => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWLEN,
      x_rsc_3_0_AWADDR => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWADDR,
      x_rsc_3_0_AWID => x_rsc_3_0_AWID,
      core_wen => core_wen,
      x_rsc_3_0_i_oswt => reg_x_rsc_3_0_i_oswt_cse,
      x_rsc_3_0_i_wen_comp => x_rsc_3_0_i_wen_comp,
      x_rsc_3_0_i_oswt_1 => reg_x_rsc_3_0_i_oswt_1_cse,
      x_rsc_3_0_i_wen_comp_1 => x_rsc_3_0_i_wen_comp_1,
      x_rsc_3_0_i_s_raddr_core => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_raddr_core,
      x_rsc_3_0_i_s_waddr_core => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_waddr_core,
      x_rsc_3_0_i_s_din_mxwt => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_din_mxwt,
      x_rsc_3_0_i_s_dout_core => hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_dout_core
    );
  x_rsc_3_0_RRESP <= hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_RRESP;
  x_rsc_3_0_RDATA <= hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_RDATA;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARREGION <= x_rsc_3_0_ARREGION;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARQOS <= x_rsc_3_0_ARQOS;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARPROT <= x_rsc_3_0_ARPROT;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARCACHE <= x_rsc_3_0_ARCACHE;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARBURST <= x_rsc_3_0_ARBURST;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARSIZE <= x_rsc_3_0_ARSIZE;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARLEN <= x_rsc_3_0_ARLEN;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_ARADDR <= x_rsc_3_0_ARADDR;
  x_rsc_3_0_BRESP <= hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_BRESP;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_WSTRB <= x_rsc_3_0_WSTRB;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_WDATA <= x_rsc_3_0_WDATA;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWREGION <= x_rsc_3_0_AWREGION;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWQOS <= x_rsc_3_0_AWQOS;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWPROT <= x_rsc_3_0_AWPROT;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWCACHE <= x_rsc_3_0_AWCACHE;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWBURST <= x_rsc_3_0_AWBURST;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWSIZE <= x_rsc_3_0_AWSIZE;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWLEN <= x_rsc_3_0_AWLEN;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_AWADDR <= x_rsc_3_0_AWADDR;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_3_0_i_s_din_mxwt <= hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_din_mxwt;
  hybrid_core_x_rsc_3_0_i_inst_x_rsc_3_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_4_0_i_inst : hybrid_core_x_rsc_4_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_4_0_s_tdone => x_rsc_4_0_s_tdone,
      x_rsc_4_0_tr_write_done => x_rsc_4_0_tr_write_done,
      x_rsc_4_0_RREADY => x_rsc_4_0_RREADY,
      x_rsc_4_0_RVALID => x_rsc_4_0_RVALID,
      x_rsc_4_0_RUSER => x_rsc_4_0_RUSER,
      x_rsc_4_0_RLAST => x_rsc_4_0_RLAST,
      x_rsc_4_0_RRESP => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_RRESP,
      x_rsc_4_0_RDATA => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_RDATA,
      x_rsc_4_0_RID => x_rsc_4_0_RID,
      x_rsc_4_0_ARREADY => x_rsc_4_0_ARREADY,
      x_rsc_4_0_ARVALID => x_rsc_4_0_ARVALID,
      x_rsc_4_0_ARUSER => x_rsc_4_0_ARUSER,
      x_rsc_4_0_ARREGION => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARREGION,
      x_rsc_4_0_ARQOS => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARQOS,
      x_rsc_4_0_ARPROT => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARPROT,
      x_rsc_4_0_ARCACHE => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARCACHE,
      x_rsc_4_0_ARLOCK => x_rsc_4_0_ARLOCK,
      x_rsc_4_0_ARBURST => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARBURST,
      x_rsc_4_0_ARSIZE => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARSIZE,
      x_rsc_4_0_ARLEN => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARLEN,
      x_rsc_4_0_ARADDR => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARADDR,
      x_rsc_4_0_ARID => x_rsc_4_0_ARID,
      x_rsc_4_0_BREADY => x_rsc_4_0_BREADY,
      x_rsc_4_0_BVALID => x_rsc_4_0_BVALID,
      x_rsc_4_0_BUSER => x_rsc_4_0_BUSER,
      x_rsc_4_0_BRESP => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_BRESP,
      x_rsc_4_0_BID => x_rsc_4_0_BID,
      x_rsc_4_0_WREADY => x_rsc_4_0_WREADY,
      x_rsc_4_0_WVALID => x_rsc_4_0_WVALID,
      x_rsc_4_0_WUSER => x_rsc_4_0_WUSER,
      x_rsc_4_0_WLAST => x_rsc_4_0_WLAST,
      x_rsc_4_0_WSTRB => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_WSTRB,
      x_rsc_4_0_WDATA => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_WDATA,
      x_rsc_4_0_AWREADY => x_rsc_4_0_AWREADY,
      x_rsc_4_0_AWVALID => x_rsc_4_0_AWVALID,
      x_rsc_4_0_AWUSER => x_rsc_4_0_AWUSER,
      x_rsc_4_0_AWREGION => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWREGION,
      x_rsc_4_0_AWQOS => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWQOS,
      x_rsc_4_0_AWPROT => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWPROT,
      x_rsc_4_0_AWCACHE => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWCACHE,
      x_rsc_4_0_AWLOCK => x_rsc_4_0_AWLOCK,
      x_rsc_4_0_AWBURST => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWBURST,
      x_rsc_4_0_AWSIZE => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWSIZE,
      x_rsc_4_0_AWLEN => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWLEN,
      x_rsc_4_0_AWADDR => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWADDR,
      x_rsc_4_0_AWID => x_rsc_4_0_AWID,
      core_wen => core_wen,
      x_rsc_4_0_i_oswt => reg_x_rsc_4_0_i_oswt_cse,
      x_rsc_4_0_i_wen_comp => x_rsc_4_0_i_wen_comp,
      x_rsc_4_0_i_oswt_1 => reg_x_rsc_4_0_i_oswt_1_cse,
      x_rsc_4_0_i_wen_comp_1 => x_rsc_4_0_i_wen_comp_1,
      x_rsc_4_0_i_s_raddr_core => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_raddr_core,
      x_rsc_4_0_i_s_waddr_core => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_waddr_core,
      x_rsc_4_0_i_s_din_mxwt => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_din_mxwt,
      x_rsc_4_0_i_s_dout_core => hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_dout_core
    );
  x_rsc_4_0_RRESP <= hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_RRESP;
  x_rsc_4_0_RDATA <= hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_RDATA;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARREGION <= x_rsc_4_0_ARREGION;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARQOS <= x_rsc_4_0_ARQOS;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARPROT <= x_rsc_4_0_ARPROT;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARCACHE <= x_rsc_4_0_ARCACHE;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARBURST <= x_rsc_4_0_ARBURST;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARSIZE <= x_rsc_4_0_ARSIZE;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARLEN <= x_rsc_4_0_ARLEN;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_ARADDR <= x_rsc_4_0_ARADDR;
  x_rsc_4_0_BRESP <= hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_BRESP;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_WSTRB <= x_rsc_4_0_WSTRB;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_WDATA <= x_rsc_4_0_WDATA;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWREGION <= x_rsc_4_0_AWREGION;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWQOS <= x_rsc_4_0_AWQOS;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWPROT <= x_rsc_4_0_AWPROT;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWCACHE <= x_rsc_4_0_AWCACHE;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWBURST <= x_rsc_4_0_AWBURST;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWSIZE <= x_rsc_4_0_AWSIZE;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWLEN <= x_rsc_4_0_AWLEN;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_AWADDR <= x_rsc_4_0_AWADDR;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_4_0_i_s_din_mxwt <= hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_din_mxwt;
  hybrid_core_x_rsc_4_0_i_inst_x_rsc_4_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_5_0_i_inst : hybrid_core_x_rsc_5_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_5_0_s_tdone => x_rsc_5_0_s_tdone,
      x_rsc_5_0_tr_write_done => x_rsc_5_0_tr_write_done,
      x_rsc_5_0_RREADY => x_rsc_5_0_RREADY,
      x_rsc_5_0_RVALID => x_rsc_5_0_RVALID,
      x_rsc_5_0_RUSER => x_rsc_5_0_RUSER,
      x_rsc_5_0_RLAST => x_rsc_5_0_RLAST,
      x_rsc_5_0_RRESP => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_RRESP,
      x_rsc_5_0_RDATA => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_RDATA,
      x_rsc_5_0_RID => x_rsc_5_0_RID,
      x_rsc_5_0_ARREADY => x_rsc_5_0_ARREADY,
      x_rsc_5_0_ARVALID => x_rsc_5_0_ARVALID,
      x_rsc_5_0_ARUSER => x_rsc_5_0_ARUSER,
      x_rsc_5_0_ARREGION => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARREGION,
      x_rsc_5_0_ARQOS => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARQOS,
      x_rsc_5_0_ARPROT => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARPROT,
      x_rsc_5_0_ARCACHE => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARCACHE,
      x_rsc_5_0_ARLOCK => x_rsc_5_0_ARLOCK,
      x_rsc_5_0_ARBURST => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARBURST,
      x_rsc_5_0_ARSIZE => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARSIZE,
      x_rsc_5_0_ARLEN => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARLEN,
      x_rsc_5_0_ARADDR => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARADDR,
      x_rsc_5_0_ARID => x_rsc_5_0_ARID,
      x_rsc_5_0_BREADY => x_rsc_5_0_BREADY,
      x_rsc_5_0_BVALID => x_rsc_5_0_BVALID,
      x_rsc_5_0_BUSER => x_rsc_5_0_BUSER,
      x_rsc_5_0_BRESP => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_BRESP,
      x_rsc_5_0_BID => x_rsc_5_0_BID,
      x_rsc_5_0_WREADY => x_rsc_5_0_WREADY,
      x_rsc_5_0_WVALID => x_rsc_5_0_WVALID,
      x_rsc_5_0_WUSER => x_rsc_5_0_WUSER,
      x_rsc_5_0_WLAST => x_rsc_5_0_WLAST,
      x_rsc_5_0_WSTRB => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_WSTRB,
      x_rsc_5_0_WDATA => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_WDATA,
      x_rsc_5_0_AWREADY => x_rsc_5_0_AWREADY,
      x_rsc_5_0_AWVALID => x_rsc_5_0_AWVALID,
      x_rsc_5_0_AWUSER => x_rsc_5_0_AWUSER,
      x_rsc_5_0_AWREGION => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWREGION,
      x_rsc_5_0_AWQOS => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWQOS,
      x_rsc_5_0_AWPROT => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWPROT,
      x_rsc_5_0_AWCACHE => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWCACHE,
      x_rsc_5_0_AWLOCK => x_rsc_5_0_AWLOCK,
      x_rsc_5_0_AWBURST => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWBURST,
      x_rsc_5_0_AWSIZE => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWSIZE,
      x_rsc_5_0_AWLEN => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWLEN,
      x_rsc_5_0_AWADDR => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWADDR,
      x_rsc_5_0_AWID => x_rsc_5_0_AWID,
      core_wen => core_wen,
      x_rsc_5_0_i_oswt => reg_x_rsc_5_0_i_oswt_cse,
      x_rsc_5_0_i_wen_comp => x_rsc_5_0_i_wen_comp,
      x_rsc_5_0_i_oswt_1 => reg_x_rsc_5_0_i_oswt_1_cse,
      x_rsc_5_0_i_wen_comp_1 => x_rsc_5_0_i_wen_comp_1,
      x_rsc_5_0_i_s_raddr_core => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_raddr_core,
      x_rsc_5_0_i_s_waddr_core => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_waddr_core,
      x_rsc_5_0_i_s_din_mxwt => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_din_mxwt,
      x_rsc_5_0_i_s_dout_core => hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_dout_core
    );
  x_rsc_5_0_RRESP <= hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_RRESP;
  x_rsc_5_0_RDATA <= hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_RDATA;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARREGION <= x_rsc_5_0_ARREGION;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARQOS <= x_rsc_5_0_ARQOS;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARPROT <= x_rsc_5_0_ARPROT;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARCACHE <= x_rsc_5_0_ARCACHE;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARBURST <= x_rsc_5_0_ARBURST;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARSIZE <= x_rsc_5_0_ARSIZE;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARLEN <= x_rsc_5_0_ARLEN;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_ARADDR <= x_rsc_5_0_ARADDR;
  x_rsc_5_0_BRESP <= hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_BRESP;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_WSTRB <= x_rsc_5_0_WSTRB;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_WDATA <= x_rsc_5_0_WDATA;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWREGION <= x_rsc_5_0_AWREGION;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWQOS <= x_rsc_5_0_AWQOS;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWPROT <= x_rsc_5_0_AWPROT;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWCACHE <= x_rsc_5_0_AWCACHE;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWBURST <= x_rsc_5_0_AWBURST;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWSIZE <= x_rsc_5_0_AWSIZE;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWLEN <= x_rsc_5_0_AWLEN;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_AWADDR <= x_rsc_5_0_AWADDR;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_5_0_i_s_din_mxwt <= hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_din_mxwt;
  hybrid_core_x_rsc_5_0_i_inst_x_rsc_5_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_6_0_i_inst : hybrid_core_x_rsc_6_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_6_0_s_tdone => x_rsc_6_0_s_tdone,
      x_rsc_6_0_tr_write_done => x_rsc_6_0_tr_write_done,
      x_rsc_6_0_RREADY => x_rsc_6_0_RREADY,
      x_rsc_6_0_RVALID => x_rsc_6_0_RVALID,
      x_rsc_6_0_RUSER => x_rsc_6_0_RUSER,
      x_rsc_6_0_RLAST => x_rsc_6_0_RLAST,
      x_rsc_6_0_RRESP => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_RRESP,
      x_rsc_6_0_RDATA => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_RDATA,
      x_rsc_6_0_RID => x_rsc_6_0_RID,
      x_rsc_6_0_ARREADY => x_rsc_6_0_ARREADY,
      x_rsc_6_0_ARVALID => x_rsc_6_0_ARVALID,
      x_rsc_6_0_ARUSER => x_rsc_6_0_ARUSER,
      x_rsc_6_0_ARREGION => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARREGION,
      x_rsc_6_0_ARQOS => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARQOS,
      x_rsc_6_0_ARPROT => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARPROT,
      x_rsc_6_0_ARCACHE => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARCACHE,
      x_rsc_6_0_ARLOCK => x_rsc_6_0_ARLOCK,
      x_rsc_6_0_ARBURST => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARBURST,
      x_rsc_6_0_ARSIZE => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARSIZE,
      x_rsc_6_0_ARLEN => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARLEN,
      x_rsc_6_0_ARADDR => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARADDR,
      x_rsc_6_0_ARID => x_rsc_6_0_ARID,
      x_rsc_6_0_BREADY => x_rsc_6_0_BREADY,
      x_rsc_6_0_BVALID => x_rsc_6_0_BVALID,
      x_rsc_6_0_BUSER => x_rsc_6_0_BUSER,
      x_rsc_6_0_BRESP => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_BRESP,
      x_rsc_6_0_BID => x_rsc_6_0_BID,
      x_rsc_6_0_WREADY => x_rsc_6_0_WREADY,
      x_rsc_6_0_WVALID => x_rsc_6_0_WVALID,
      x_rsc_6_0_WUSER => x_rsc_6_0_WUSER,
      x_rsc_6_0_WLAST => x_rsc_6_0_WLAST,
      x_rsc_6_0_WSTRB => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_WSTRB,
      x_rsc_6_0_WDATA => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_WDATA,
      x_rsc_6_0_AWREADY => x_rsc_6_0_AWREADY,
      x_rsc_6_0_AWVALID => x_rsc_6_0_AWVALID,
      x_rsc_6_0_AWUSER => x_rsc_6_0_AWUSER,
      x_rsc_6_0_AWREGION => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWREGION,
      x_rsc_6_0_AWQOS => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWQOS,
      x_rsc_6_0_AWPROT => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWPROT,
      x_rsc_6_0_AWCACHE => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWCACHE,
      x_rsc_6_0_AWLOCK => x_rsc_6_0_AWLOCK,
      x_rsc_6_0_AWBURST => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWBURST,
      x_rsc_6_0_AWSIZE => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWSIZE,
      x_rsc_6_0_AWLEN => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWLEN,
      x_rsc_6_0_AWADDR => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWADDR,
      x_rsc_6_0_AWID => x_rsc_6_0_AWID,
      core_wen => core_wen,
      x_rsc_6_0_i_oswt => reg_x_rsc_6_0_i_oswt_cse,
      x_rsc_6_0_i_wen_comp => x_rsc_6_0_i_wen_comp,
      x_rsc_6_0_i_oswt_1 => reg_x_rsc_6_0_i_oswt_1_cse,
      x_rsc_6_0_i_wen_comp_1 => x_rsc_6_0_i_wen_comp_1,
      x_rsc_6_0_i_s_raddr_core => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_raddr_core,
      x_rsc_6_0_i_s_waddr_core => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_waddr_core,
      x_rsc_6_0_i_s_din_mxwt => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_din_mxwt,
      x_rsc_6_0_i_s_dout_core => hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_dout_core
    );
  x_rsc_6_0_RRESP <= hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_RRESP;
  x_rsc_6_0_RDATA <= hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_RDATA;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARREGION <= x_rsc_6_0_ARREGION;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARQOS <= x_rsc_6_0_ARQOS;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARPROT <= x_rsc_6_0_ARPROT;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARCACHE <= x_rsc_6_0_ARCACHE;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARBURST <= x_rsc_6_0_ARBURST;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARSIZE <= x_rsc_6_0_ARSIZE;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARLEN <= x_rsc_6_0_ARLEN;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_ARADDR <= x_rsc_6_0_ARADDR;
  x_rsc_6_0_BRESP <= hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_BRESP;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_WSTRB <= x_rsc_6_0_WSTRB;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_WDATA <= x_rsc_6_0_WDATA;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWREGION <= x_rsc_6_0_AWREGION;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWQOS <= x_rsc_6_0_AWQOS;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWPROT <= x_rsc_6_0_AWPROT;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWCACHE <= x_rsc_6_0_AWCACHE;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWBURST <= x_rsc_6_0_AWBURST;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWSIZE <= x_rsc_6_0_AWSIZE;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWLEN <= x_rsc_6_0_AWLEN;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_AWADDR <= x_rsc_6_0_AWADDR;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_6_0_i_s_din_mxwt <= hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_din_mxwt;
  hybrid_core_x_rsc_6_0_i_inst_x_rsc_6_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_7_0_i_inst : hybrid_core_x_rsc_7_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_7_0_s_tdone => x_rsc_7_0_s_tdone,
      x_rsc_7_0_tr_write_done => x_rsc_7_0_tr_write_done,
      x_rsc_7_0_RREADY => x_rsc_7_0_RREADY,
      x_rsc_7_0_RVALID => x_rsc_7_0_RVALID,
      x_rsc_7_0_RUSER => x_rsc_7_0_RUSER,
      x_rsc_7_0_RLAST => x_rsc_7_0_RLAST,
      x_rsc_7_0_RRESP => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_RRESP,
      x_rsc_7_0_RDATA => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_RDATA,
      x_rsc_7_0_RID => x_rsc_7_0_RID,
      x_rsc_7_0_ARREADY => x_rsc_7_0_ARREADY,
      x_rsc_7_0_ARVALID => x_rsc_7_0_ARVALID,
      x_rsc_7_0_ARUSER => x_rsc_7_0_ARUSER,
      x_rsc_7_0_ARREGION => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARREGION,
      x_rsc_7_0_ARQOS => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARQOS,
      x_rsc_7_0_ARPROT => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARPROT,
      x_rsc_7_0_ARCACHE => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARCACHE,
      x_rsc_7_0_ARLOCK => x_rsc_7_0_ARLOCK,
      x_rsc_7_0_ARBURST => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARBURST,
      x_rsc_7_0_ARSIZE => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARSIZE,
      x_rsc_7_0_ARLEN => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARLEN,
      x_rsc_7_0_ARADDR => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARADDR,
      x_rsc_7_0_ARID => x_rsc_7_0_ARID,
      x_rsc_7_0_BREADY => x_rsc_7_0_BREADY,
      x_rsc_7_0_BVALID => x_rsc_7_0_BVALID,
      x_rsc_7_0_BUSER => x_rsc_7_0_BUSER,
      x_rsc_7_0_BRESP => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_BRESP,
      x_rsc_7_0_BID => x_rsc_7_0_BID,
      x_rsc_7_0_WREADY => x_rsc_7_0_WREADY,
      x_rsc_7_0_WVALID => x_rsc_7_0_WVALID,
      x_rsc_7_0_WUSER => x_rsc_7_0_WUSER,
      x_rsc_7_0_WLAST => x_rsc_7_0_WLAST,
      x_rsc_7_0_WSTRB => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_WSTRB,
      x_rsc_7_0_WDATA => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_WDATA,
      x_rsc_7_0_AWREADY => x_rsc_7_0_AWREADY,
      x_rsc_7_0_AWVALID => x_rsc_7_0_AWVALID,
      x_rsc_7_0_AWUSER => x_rsc_7_0_AWUSER,
      x_rsc_7_0_AWREGION => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWREGION,
      x_rsc_7_0_AWQOS => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWQOS,
      x_rsc_7_0_AWPROT => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWPROT,
      x_rsc_7_0_AWCACHE => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWCACHE,
      x_rsc_7_0_AWLOCK => x_rsc_7_0_AWLOCK,
      x_rsc_7_0_AWBURST => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWBURST,
      x_rsc_7_0_AWSIZE => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWSIZE,
      x_rsc_7_0_AWLEN => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWLEN,
      x_rsc_7_0_AWADDR => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWADDR,
      x_rsc_7_0_AWID => x_rsc_7_0_AWID,
      core_wen => core_wen,
      x_rsc_7_0_i_oswt => reg_x_rsc_7_0_i_oswt_cse,
      x_rsc_7_0_i_wen_comp => x_rsc_7_0_i_wen_comp,
      x_rsc_7_0_i_oswt_1 => reg_x_rsc_7_0_i_oswt_1_cse,
      x_rsc_7_0_i_wen_comp_1 => x_rsc_7_0_i_wen_comp_1,
      x_rsc_7_0_i_s_raddr_core => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_raddr_core,
      x_rsc_7_0_i_s_waddr_core => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_waddr_core,
      x_rsc_7_0_i_s_din_mxwt => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_din_mxwt,
      x_rsc_7_0_i_s_dout_core => hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_dout_core
    );
  x_rsc_7_0_RRESP <= hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_RRESP;
  x_rsc_7_0_RDATA <= hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_RDATA;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARREGION <= x_rsc_7_0_ARREGION;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARQOS <= x_rsc_7_0_ARQOS;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARPROT <= x_rsc_7_0_ARPROT;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARCACHE <= x_rsc_7_0_ARCACHE;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARBURST <= x_rsc_7_0_ARBURST;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARSIZE <= x_rsc_7_0_ARSIZE;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARLEN <= x_rsc_7_0_ARLEN;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_ARADDR <= x_rsc_7_0_ARADDR;
  x_rsc_7_0_BRESP <= hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_BRESP;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_WSTRB <= x_rsc_7_0_WSTRB;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_WDATA <= x_rsc_7_0_WDATA;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWREGION <= x_rsc_7_0_AWREGION;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWQOS <= x_rsc_7_0_AWQOS;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWPROT <= x_rsc_7_0_AWPROT;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWCACHE <= x_rsc_7_0_AWCACHE;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWBURST <= x_rsc_7_0_AWBURST;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWSIZE <= x_rsc_7_0_AWSIZE;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWLEN <= x_rsc_7_0_AWLEN;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_AWADDR <= x_rsc_7_0_AWADDR;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_7_0_i_s_din_mxwt <= hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_din_mxwt;
  hybrid_core_x_rsc_7_0_i_inst_x_rsc_7_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_8_0_i_inst : hybrid_core_x_rsc_8_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_8_0_s_tdone => x_rsc_8_0_s_tdone,
      x_rsc_8_0_tr_write_done => x_rsc_8_0_tr_write_done,
      x_rsc_8_0_RREADY => x_rsc_8_0_RREADY,
      x_rsc_8_0_RVALID => x_rsc_8_0_RVALID,
      x_rsc_8_0_RUSER => x_rsc_8_0_RUSER,
      x_rsc_8_0_RLAST => x_rsc_8_0_RLAST,
      x_rsc_8_0_RRESP => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_RRESP,
      x_rsc_8_0_RDATA => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_RDATA,
      x_rsc_8_0_RID => x_rsc_8_0_RID,
      x_rsc_8_0_ARREADY => x_rsc_8_0_ARREADY,
      x_rsc_8_0_ARVALID => x_rsc_8_0_ARVALID,
      x_rsc_8_0_ARUSER => x_rsc_8_0_ARUSER,
      x_rsc_8_0_ARREGION => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARREGION,
      x_rsc_8_0_ARQOS => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARQOS,
      x_rsc_8_0_ARPROT => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARPROT,
      x_rsc_8_0_ARCACHE => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARCACHE,
      x_rsc_8_0_ARLOCK => x_rsc_8_0_ARLOCK,
      x_rsc_8_0_ARBURST => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARBURST,
      x_rsc_8_0_ARSIZE => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARSIZE,
      x_rsc_8_0_ARLEN => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARLEN,
      x_rsc_8_0_ARADDR => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARADDR,
      x_rsc_8_0_ARID => x_rsc_8_0_ARID,
      x_rsc_8_0_BREADY => x_rsc_8_0_BREADY,
      x_rsc_8_0_BVALID => x_rsc_8_0_BVALID,
      x_rsc_8_0_BUSER => x_rsc_8_0_BUSER,
      x_rsc_8_0_BRESP => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_BRESP,
      x_rsc_8_0_BID => x_rsc_8_0_BID,
      x_rsc_8_0_WREADY => x_rsc_8_0_WREADY,
      x_rsc_8_0_WVALID => x_rsc_8_0_WVALID,
      x_rsc_8_0_WUSER => x_rsc_8_0_WUSER,
      x_rsc_8_0_WLAST => x_rsc_8_0_WLAST,
      x_rsc_8_0_WSTRB => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_WSTRB,
      x_rsc_8_0_WDATA => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_WDATA,
      x_rsc_8_0_AWREADY => x_rsc_8_0_AWREADY,
      x_rsc_8_0_AWVALID => x_rsc_8_0_AWVALID,
      x_rsc_8_0_AWUSER => x_rsc_8_0_AWUSER,
      x_rsc_8_0_AWREGION => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWREGION,
      x_rsc_8_0_AWQOS => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWQOS,
      x_rsc_8_0_AWPROT => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWPROT,
      x_rsc_8_0_AWCACHE => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWCACHE,
      x_rsc_8_0_AWLOCK => x_rsc_8_0_AWLOCK,
      x_rsc_8_0_AWBURST => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWBURST,
      x_rsc_8_0_AWSIZE => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWSIZE,
      x_rsc_8_0_AWLEN => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWLEN,
      x_rsc_8_0_AWADDR => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWADDR,
      x_rsc_8_0_AWID => x_rsc_8_0_AWID,
      core_wen => core_wen,
      x_rsc_8_0_i_oswt => reg_x_rsc_8_0_i_oswt_cse,
      x_rsc_8_0_i_wen_comp => x_rsc_8_0_i_wen_comp,
      x_rsc_8_0_i_oswt_1 => reg_x_rsc_8_0_i_oswt_1_cse,
      x_rsc_8_0_i_wen_comp_1 => x_rsc_8_0_i_wen_comp_1,
      x_rsc_8_0_i_s_raddr_core => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_raddr_core,
      x_rsc_8_0_i_s_waddr_core => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_waddr_core,
      x_rsc_8_0_i_s_din_mxwt => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_din_mxwt,
      x_rsc_8_0_i_s_dout_core => hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_dout_core
    );
  x_rsc_8_0_RRESP <= hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_RRESP;
  x_rsc_8_0_RDATA <= hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_RDATA;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARREGION <= x_rsc_8_0_ARREGION;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARQOS <= x_rsc_8_0_ARQOS;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARPROT <= x_rsc_8_0_ARPROT;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARCACHE <= x_rsc_8_0_ARCACHE;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARBURST <= x_rsc_8_0_ARBURST;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARSIZE <= x_rsc_8_0_ARSIZE;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARLEN <= x_rsc_8_0_ARLEN;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_ARADDR <= x_rsc_8_0_ARADDR;
  x_rsc_8_0_BRESP <= hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_BRESP;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_WSTRB <= x_rsc_8_0_WSTRB;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_WDATA <= x_rsc_8_0_WDATA;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWREGION <= x_rsc_8_0_AWREGION;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWQOS <= x_rsc_8_0_AWQOS;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWPROT <= x_rsc_8_0_AWPROT;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWCACHE <= x_rsc_8_0_AWCACHE;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWBURST <= x_rsc_8_0_AWBURST;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWSIZE <= x_rsc_8_0_AWSIZE;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWLEN <= x_rsc_8_0_AWLEN;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_AWADDR <= x_rsc_8_0_AWADDR;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_8_0_i_s_din_mxwt <= hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_din_mxwt;
  hybrid_core_x_rsc_8_0_i_inst_x_rsc_8_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_9_0_i_inst : hybrid_core_x_rsc_9_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_9_0_s_tdone => x_rsc_9_0_s_tdone,
      x_rsc_9_0_tr_write_done => x_rsc_9_0_tr_write_done,
      x_rsc_9_0_RREADY => x_rsc_9_0_RREADY,
      x_rsc_9_0_RVALID => x_rsc_9_0_RVALID,
      x_rsc_9_0_RUSER => x_rsc_9_0_RUSER,
      x_rsc_9_0_RLAST => x_rsc_9_0_RLAST,
      x_rsc_9_0_RRESP => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_RRESP,
      x_rsc_9_0_RDATA => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_RDATA,
      x_rsc_9_0_RID => x_rsc_9_0_RID,
      x_rsc_9_0_ARREADY => x_rsc_9_0_ARREADY,
      x_rsc_9_0_ARVALID => x_rsc_9_0_ARVALID,
      x_rsc_9_0_ARUSER => x_rsc_9_0_ARUSER,
      x_rsc_9_0_ARREGION => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARREGION,
      x_rsc_9_0_ARQOS => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARQOS,
      x_rsc_9_0_ARPROT => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARPROT,
      x_rsc_9_0_ARCACHE => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARCACHE,
      x_rsc_9_0_ARLOCK => x_rsc_9_0_ARLOCK,
      x_rsc_9_0_ARBURST => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARBURST,
      x_rsc_9_0_ARSIZE => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARSIZE,
      x_rsc_9_0_ARLEN => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARLEN,
      x_rsc_9_0_ARADDR => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARADDR,
      x_rsc_9_0_ARID => x_rsc_9_0_ARID,
      x_rsc_9_0_BREADY => x_rsc_9_0_BREADY,
      x_rsc_9_0_BVALID => x_rsc_9_0_BVALID,
      x_rsc_9_0_BUSER => x_rsc_9_0_BUSER,
      x_rsc_9_0_BRESP => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_BRESP,
      x_rsc_9_0_BID => x_rsc_9_0_BID,
      x_rsc_9_0_WREADY => x_rsc_9_0_WREADY,
      x_rsc_9_0_WVALID => x_rsc_9_0_WVALID,
      x_rsc_9_0_WUSER => x_rsc_9_0_WUSER,
      x_rsc_9_0_WLAST => x_rsc_9_0_WLAST,
      x_rsc_9_0_WSTRB => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_WSTRB,
      x_rsc_9_0_WDATA => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_WDATA,
      x_rsc_9_0_AWREADY => x_rsc_9_0_AWREADY,
      x_rsc_9_0_AWVALID => x_rsc_9_0_AWVALID,
      x_rsc_9_0_AWUSER => x_rsc_9_0_AWUSER,
      x_rsc_9_0_AWREGION => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWREGION,
      x_rsc_9_0_AWQOS => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWQOS,
      x_rsc_9_0_AWPROT => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWPROT,
      x_rsc_9_0_AWCACHE => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWCACHE,
      x_rsc_9_0_AWLOCK => x_rsc_9_0_AWLOCK,
      x_rsc_9_0_AWBURST => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWBURST,
      x_rsc_9_0_AWSIZE => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWSIZE,
      x_rsc_9_0_AWLEN => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWLEN,
      x_rsc_9_0_AWADDR => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWADDR,
      x_rsc_9_0_AWID => x_rsc_9_0_AWID,
      core_wen => core_wen,
      x_rsc_9_0_i_oswt => reg_x_rsc_9_0_i_oswt_cse,
      x_rsc_9_0_i_wen_comp => x_rsc_9_0_i_wen_comp,
      x_rsc_9_0_i_oswt_1 => reg_x_rsc_9_0_i_oswt_1_cse,
      x_rsc_9_0_i_wen_comp_1 => x_rsc_9_0_i_wen_comp_1,
      x_rsc_9_0_i_s_raddr_core => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_raddr_core,
      x_rsc_9_0_i_s_waddr_core => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_waddr_core,
      x_rsc_9_0_i_s_din_mxwt => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_din_mxwt,
      x_rsc_9_0_i_s_dout_core => hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_dout_core
    );
  x_rsc_9_0_RRESP <= hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_RRESP;
  x_rsc_9_0_RDATA <= hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_RDATA;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARREGION <= x_rsc_9_0_ARREGION;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARQOS <= x_rsc_9_0_ARQOS;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARPROT <= x_rsc_9_0_ARPROT;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARCACHE <= x_rsc_9_0_ARCACHE;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARBURST <= x_rsc_9_0_ARBURST;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARSIZE <= x_rsc_9_0_ARSIZE;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARLEN <= x_rsc_9_0_ARLEN;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_ARADDR <= x_rsc_9_0_ARADDR;
  x_rsc_9_0_BRESP <= hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_BRESP;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_WSTRB <= x_rsc_9_0_WSTRB;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_WDATA <= x_rsc_9_0_WDATA;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWREGION <= x_rsc_9_0_AWREGION;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWQOS <= x_rsc_9_0_AWQOS;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWPROT <= x_rsc_9_0_AWPROT;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWCACHE <= x_rsc_9_0_AWCACHE;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWBURST <= x_rsc_9_0_AWBURST;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWSIZE <= x_rsc_9_0_AWSIZE;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWLEN <= x_rsc_9_0_AWLEN;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_AWADDR <= x_rsc_9_0_AWADDR;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_9_0_i_s_din_mxwt <= hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_din_mxwt;
  hybrid_core_x_rsc_9_0_i_inst_x_rsc_9_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_10_0_i_inst : hybrid_core_x_rsc_10_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_10_0_s_tdone => x_rsc_10_0_s_tdone,
      x_rsc_10_0_tr_write_done => x_rsc_10_0_tr_write_done,
      x_rsc_10_0_RREADY => x_rsc_10_0_RREADY,
      x_rsc_10_0_RVALID => x_rsc_10_0_RVALID,
      x_rsc_10_0_RUSER => x_rsc_10_0_RUSER,
      x_rsc_10_0_RLAST => x_rsc_10_0_RLAST,
      x_rsc_10_0_RRESP => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_RRESP,
      x_rsc_10_0_RDATA => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_RDATA,
      x_rsc_10_0_RID => x_rsc_10_0_RID,
      x_rsc_10_0_ARREADY => x_rsc_10_0_ARREADY,
      x_rsc_10_0_ARVALID => x_rsc_10_0_ARVALID,
      x_rsc_10_0_ARUSER => x_rsc_10_0_ARUSER,
      x_rsc_10_0_ARREGION => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARREGION,
      x_rsc_10_0_ARQOS => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARQOS,
      x_rsc_10_0_ARPROT => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARPROT,
      x_rsc_10_0_ARCACHE => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARCACHE,
      x_rsc_10_0_ARLOCK => x_rsc_10_0_ARLOCK,
      x_rsc_10_0_ARBURST => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARBURST,
      x_rsc_10_0_ARSIZE => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARSIZE,
      x_rsc_10_0_ARLEN => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARLEN,
      x_rsc_10_0_ARADDR => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARADDR,
      x_rsc_10_0_ARID => x_rsc_10_0_ARID,
      x_rsc_10_0_BREADY => x_rsc_10_0_BREADY,
      x_rsc_10_0_BVALID => x_rsc_10_0_BVALID,
      x_rsc_10_0_BUSER => x_rsc_10_0_BUSER,
      x_rsc_10_0_BRESP => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_BRESP,
      x_rsc_10_0_BID => x_rsc_10_0_BID,
      x_rsc_10_0_WREADY => x_rsc_10_0_WREADY,
      x_rsc_10_0_WVALID => x_rsc_10_0_WVALID,
      x_rsc_10_0_WUSER => x_rsc_10_0_WUSER,
      x_rsc_10_0_WLAST => x_rsc_10_0_WLAST,
      x_rsc_10_0_WSTRB => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_WSTRB,
      x_rsc_10_0_WDATA => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_WDATA,
      x_rsc_10_0_AWREADY => x_rsc_10_0_AWREADY,
      x_rsc_10_0_AWVALID => x_rsc_10_0_AWVALID,
      x_rsc_10_0_AWUSER => x_rsc_10_0_AWUSER,
      x_rsc_10_0_AWREGION => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWREGION,
      x_rsc_10_0_AWQOS => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWQOS,
      x_rsc_10_0_AWPROT => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWPROT,
      x_rsc_10_0_AWCACHE => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWCACHE,
      x_rsc_10_0_AWLOCK => x_rsc_10_0_AWLOCK,
      x_rsc_10_0_AWBURST => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWBURST,
      x_rsc_10_0_AWSIZE => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWSIZE,
      x_rsc_10_0_AWLEN => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWLEN,
      x_rsc_10_0_AWADDR => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWADDR,
      x_rsc_10_0_AWID => x_rsc_10_0_AWID,
      core_wen => core_wen,
      x_rsc_10_0_i_oswt => reg_x_rsc_10_0_i_oswt_cse,
      x_rsc_10_0_i_wen_comp => x_rsc_10_0_i_wen_comp,
      x_rsc_10_0_i_oswt_1 => reg_x_rsc_10_0_i_oswt_1_cse,
      x_rsc_10_0_i_wen_comp_1 => x_rsc_10_0_i_wen_comp_1,
      x_rsc_10_0_i_s_raddr_core => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_raddr_core,
      x_rsc_10_0_i_s_waddr_core => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_waddr_core,
      x_rsc_10_0_i_s_din_mxwt => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_din_mxwt,
      x_rsc_10_0_i_s_dout_core => hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_dout_core
    );
  x_rsc_10_0_RRESP <= hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_RRESP;
  x_rsc_10_0_RDATA <= hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_RDATA;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARREGION <= x_rsc_10_0_ARREGION;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARQOS <= x_rsc_10_0_ARQOS;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARPROT <= x_rsc_10_0_ARPROT;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARCACHE <= x_rsc_10_0_ARCACHE;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARBURST <= x_rsc_10_0_ARBURST;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARSIZE <= x_rsc_10_0_ARSIZE;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARLEN <= x_rsc_10_0_ARLEN;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_ARADDR <= x_rsc_10_0_ARADDR;
  x_rsc_10_0_BRESP <= hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_BRESP;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_WSTRB <= x_rsc_10_0_WSTRB;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_WDATA <= x_rsc_10_0_WDATA;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWREGION <= x_rsc_10_0_AWREGION;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWQOS <= x_rsc_10_0_AWQOS;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWPROT <= x_rsc_10_0_AWPROT;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWCACHE <= x_rsc_10_0_AWCACHE;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWBURST <= x_rsc_10_0_AWBURST;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWSIZE <= x_rsc_10_0_AWSIZE;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWLEN <= x_rsc_10_0_AWLEN;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_AWADDR <= x_rsc_10_0_AWADDR;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_10_0_i_s_din_mxwt <= hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_din_mxwt;
  hybrid_core_x_rsc_10_0_i_inst_x_rsc_10_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_11_0_i_inst : hybrid_core_x_rsc_11_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_11_0_s_tdone => x_rsc_11_0_s_tdone,
      x_rsc_11_0_tr_write_done => x_rsc_11_0_tr_write_done,
      x_rsc_11_0_RREADY => x_rsc_11_0_RREADY,
      x_rsc_11_0_RVALID => x_rsc_11_0_RVALID,
      x_rsc_11_0_RUSER => x_rsc_11_0_RUSER,
      x_rsc_11_0_RLAST => x_rsc_11_0_RLAST,
      x_rsc_11_0_RRESP => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_RRESP,
      x_rsc_11_0_RDATA => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_RDATA,
      x_rsc_11_0_RID => x_rsc_11_0_RID,
      x_rsc_11_0_ARREADY => x_rsc_11_0_ARREADY,
      x_rsc_11_0_ARVALID => x_rsc_11_0_ARVALID,
      x_rsc_11_0_ARUSER => x_rsc_11_0_ARUSER,
      x_rsc_11_0_ARREGION => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARREGION,
      x_rsc_11_0_ARQOS => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARQOS,
      x_rsc_11_0_ARPROT => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARPROT,
      x_rsc_11_0_ARCACHE => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARCACHE,
      x_rsc_11_0_ARLOCK => x_rsc_11_0_ARLOCK,
      x_rsc_11_0_ARBURST => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARBURST,
      x_rsc_11_0_ARSIZE => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARSIZE,
      x_rsc_11_0_ARLEN => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARLEN,
      x_rsc_11_0_ARADDR => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARADDR,
      x_rsc_11_0_ARID => x_rsc_11_0_ARID,
      x_rsc_11_0_BREADY => x_rsc_11_0_BREADY,
      x_rsc_11_0_BVALID => x_rsc_11_0_BVALID,
      x_rsc_11_0_BUSER => x_rsc_11_0_BUSER,
      x_rsc_11_0_BRESP => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_BRESP,
      x_rsc_11_0_BID => x_rsc_11_0_BID,
      x_rsc_11_0_WREADY => x_rsc_11_0_WREADY,
      x_rsc_11_0_WVALID => x_rsc_11_0_WVALID,
      x_rsc_11_0_WUSER => x_rsc_11_0_WUSER,
      x_rsc_11_0_WLAST => x_rsc_11_0_WLAST,
      x_rsc_11_0_WSTRB => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_WSTRB,
      x_rsc_11_0_WDATA => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_WDATA,
      x_rsc_11_0_AWREADY => x_rsc_11_0_AWREADY,
      x_rsc_11_0_AWVALID => x_rsc_11_0_AWVALID,
      x_rsc_11_0_AWUSER => x_rsc_11_0_AWUSER,
      x_rsc_11_0_AWREGION => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWREGION,
      x_rsc_11_0_AWQOS => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWQOS,
      x_rsc_11_0_AWPROT => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWPROT,
      x_rsc_11_0_AWCACHE => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWCACHE,
      x_rsc_11_0_AWLOCK => x_rsc_11_0_AWLOCK,
      x_rsc_11_0_AWBURST => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWBURST,
      x_rsc_11_0_AWSIZE => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWSIZE,
      x_rsc_11_0_AWLEN => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWLEN,
      x_rsc_11_0_AWADDR => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWADDR,
      x_rsc_11_0_AWID => x_rsc_11_0_AWID,
      core_wen => core_wen,
      x_rsc_11_0_i_oswt => reg_x_rsc_11_0_i_oswt_cse,
      x_rsc_11_0_i_wen_comp => x_rsc_11_0_i_wen_comp,
      x_rsc_11_0_i_oswt_1 => reg_x_rsc_11_0_i_oswt_1_cse,
      x_rsc_11_0_i_wen_comp_1 => x_rsc_11_0_i_wen_comp_1,
      x_rsc_11_0_i_s_raddr_core => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_raddr_core,
      x_rsc_11_0_i_s_waddr_core => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_waddr_core,
      x_rsc_11_0_i_s_din_mxwt => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_din_mxwt,
      x_rsc_11_0_i_s_dout_core => hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_dout_core
    );
  x_rsc_11_0_RRESP <= hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_RRESP;
  x_rsc_11_0_RDATA <= hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_RDATA;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARREGION <= x_rsc_11_0_ARREGION;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARQOS <= x_rsc_11_0_ARQOS;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARPROT <= x_rsc_11_0_ARPROT;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARCACHE <= x_rsc_11_0_ARCACHE;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARBURST <= x_rsc_11_0_ARBURST;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARSIZE <= x_rsc_11_0_ARSIZE;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARLEN <= x_rsc_11_0_ARLEN;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_ARADDR <= x_rsc_11_0_ARADDR;
  x_rsc_11_0_BRESP <= hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_BRESP;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_WSTRB <= x_rsc_11_0_WSTRB;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_WDATA <= x_rsc_11_0_WDATA;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWREGION <= x_rsc_11_0_AWREGION;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWQOS <= x_rsc_11_0_AWQOS;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWPROT <= x_rsc_11_0_AWPROT;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWCACHE <= x_rsc_11_0_AWCACHE;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWBURST <= x_rsc_11_0_AWBURST;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWSIZE <= x_rsc_11_0_AWSIZE;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWLEN <= x_rsc_11_0_AWLEN;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_AWADDR <= x_rsc_11_0_AWADDR;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_11_0_i_s_din_mxwt <= hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_din_mxwt;
  hybrid_core_x_rsc_11_0_i_inst_x_rsc_11_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_12_0_i_inst : hybrid_core_x_rsc_12_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_12_0_s_tdone => x_rsc_12_0_s_tdone,
      x_rsc_12_0_tr_write_done => x_rsc_12_0_tr_write_done,
      x_rsc_12_0_RREADY => x_rsc_12_0_RREADY,
      x_rsc_12_0_RVALID => x_rsc_12_0_RVALID,
      x_rsc_12_0_RUSER => x_rsc_12_0_RUSER,
      x_rsc_12_0_RLAST => x_rsc_12_0_RLAST,
      x_rsc_12_0_RRESP => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_RRESP,
      x_rsc_12_0_RDATA => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_RDATA,
      x_rsc_12_0_RID => x_rsc_12_0_RID,
      x_rsc_12_0_ARREADY => x_rsc_12_0_ARREADY,
      x_rsc_12_0_ARVALID => x_rsc_12_0_ARVALID,
      x_rsc_12_0_ARUSER => x_rsc_12_0_ARUSER,
      x_rsc_12_0_ARREGION => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARREGION,
      x_rsc_12_0_ARQOS => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARQOS,
      x_rsc_12_0_ARPROT => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARPROT,
      x_rsc_12_0_ARCACHE => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARCACHE,
      x_rsc_12_0_ARLOCK => x_rsc_12_0_ARLOCK,
      x_rsc_12_0_ARBURST => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARBURST,
      x_rsc_12_0_ARSIZE => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARSIZE,
      x_rsc_12_0_ARLEN => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARLEN,
      x_rsc_12_0_ARADDR => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARADDR,
      x_rsc_12_0_ARID => x_rsc_12_0_ARID,
      x_rsc_12_0_BREADY => x_rsc_12_0_BREADY,
      x_rsc_12_0_BVALID => x_rsc_12_0_BVALID,
      x_rsc_12_0_BUSER => x_rsc_12_0_BUSER,
      x_rsc_12_0_BRESP => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_BRESP,
      x_rsc_12_0_BID => x_rsc_12_0_BID,
      x_rsc_12_0_WREADY => x_rsc_12_0_WREADY,
      x_rsc_12_0_WVALID => x_rsc_12_0_WVALID,
      x_rsc_12_0_WUSER => x_rsc_12_0_WUSER,
      x_rsc_12_0_WLAST => x_rsc_12_0_WLAST,
      x_rsc_12_0_WSTRB => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_WSTRB,
      x_rsc_12_0_WDATA => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_WDATA,
      x_rsc_12_0_AWREADY => x_rsc_12_0_AWREADY,
      x_rsc_12_0_AWVALID => x_rsc_12_0_AWVALID,
      x_rsc_12_0_AWUSER => x_rsc_12_0_AWUSER,
      x_rsc_12_0_AWREGION => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWREGION,
      x_rsc_12_0_AWQOS => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWQOS,
      x_rsc_12_0_AWPROT => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWPROT,
      x_rsc_12_0_AWCACHE => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWCACHE,
      x_rsc_12_0_AWLOCK => x_rsc_12_0_AWLOCK,
      x_rsc_12_0_AWBURST => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWBURST,
      x_rsc_12_0_AWSIZE => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWSIZE,
      x_rsc_12_0_AWLEN => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWLEN,
      x_rsc_12_0_AWADDR => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWADDR,
      x_rsc_12_0_AWID => x_rsc_12_0_AWID,
      core_wen => core_wen,
      x_rsc_12_0_i_oswt => reg_x_rsc_12_0_i_oswt_cse,
      x_rsc_12_0_i_wen_comp => x_rsc_12_0_i_wen_comp,
      x_rsc_12_0_i_oswt_1 => reg_x_rsc_12_0_i_oswt_1_cse,
      x_rsc_12_0_i_wen_comp_1 => x_rsc_12_0_i_wen_comp_1,
      x_rsc_12_0_i_s_raddr_core => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_raddr_core,
      x_rsc_12_0_i_s_waddr_core => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_waddr_core,
      x_rsc_12_0_i_s_din_mxwt => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_din_mxwt,
      x_rsc_12_0_i_s_dout_core => hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_dout_core
    );
  x_rsc_12_0_RRESP <= hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_RRESP;
  x_rsc_12_0_RDATA <= hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_RDATA;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARREGION <= x_rsc_12_0_ARREGION;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARQOS <= x_rsc_12_0_ARQOS;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARPROT <= x_rsc_12_0_ARPROT;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARCACHE <= x_rsc_12_0_ARCACHE;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARBURST <= x_rsc_12_0_ARBURST;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARSIZE <= x_rsc_12_0_ARSIZE;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARLEN <= x_rsc_12_0_ARLEN;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_ARADDR <= x_rsc_12_0_ARADDR;
  x_rsc_12_0_BRESP <= hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_BRESP;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_WSTRB <= x_rsc_12_0_WSTRB;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_WDATA <= x_rsc_12_0_WDATA;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWREGION <= x_rsc_12_0_AWREGION;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWQOS <= x_rsc_12_0_AWQOS;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWPROT <= x_rsc_12_0_AWPROT;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWCACHE <= x_rsc_12_0_AWCACHE;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWBURST <= x_rsc_12_0_AWBURST;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWSIZE <= x_rsc_12_0_AWSIZE;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWLEN <= x_rsc_12_0_AWLEN;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_AWADDR <= x_rsc_12_0_AWADDR;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_12_0_i_s_din_mxwt <= hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_din_mxwt;
  hybrid_core_x_rsc_12_0_i_inst_x_rsc_12_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_13_0_i_inst : hybrid_core_x_rsc_13_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_13_0_s_tdone => x_rsc_13_0_s_tdone,
      x_rsc_13_0_tr_write_done => x_rsc_13_0_tr_write_done,
      x_rsc_13_0_RREADY => x_rsc_13_0_RREADY,
      x_rsc_13_0_RVALID => x_rsc_13_0_RVALID,
      x_rsc_13_0_RUSER => x_rsc_13_0_RUSER,
      x_rsc_13_0_RLAST => x_rsc_13_0_RLAST,
      x_rsc_13_0_RRESP => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_RRESP,
      x_rsc_13_0_RDATA => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_RDATA,
      x_rsc_13_0_RID => x_rsc_13_0_RID,
      x_rsc_13_0_ARREADY => x_rsc_13_0_ARREADY,
      x_rsc_13_0_ARVALID => x_rsc_13_0_ARVALID,
      x_rsc_13_0_ARUSER => x_rsc_13_0_ARUSER,
      x_rsc_13_0_ARREGION => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARREGION,
      x_rsc_13_0_ARQOS => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARQOS,
      x_rsc_13_0_ARPROT => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARPROT,
      x_rsc_13_0_ARCACHE => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARCACHE,
      x_rsc_13_0_ARLOCK => x_rsc_13_0_ARLOCK,
      x_rsc_13_0_ARBURST => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARBURST,
      x_rsc_13_0_ARSIZE => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARSIZE,
      x_rsc_13_0_ARLEN => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARLEN,
      x_rsc_13_0_ARADDR => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARADDR,
      x_rsc_13_0_ARID => x_rsc_13_0_ARID,
      x_rsc_13_0_BREADY => x_rsc_13_0_BREADY,
      x_rsc_13_0_BVALID => x_rsc_13_0_BVALID,
      x_rsc_13_0_BUSER => x_rsc_13_0_BUSER,
      x_rsc_13_0_BRESP => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_BRESP,
      x_rsc_13_0_BID => x_rsc_13_0_BID,
      x_rsc_13_0_WREADY => x_rsc_13_0_WREADY,
      x_rsc_13_0_WVALID => x_rsc_13_0_WVALID,
      x_rsc_13_0_WUSER => x_rsc_13_0_WUSER,
      x_rsc_13_0_WLAST => x_rsc_13_0_WLAST,
      x_rsc_13_0_WSTRB => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_WSTRB,
      x_rsc_13_0_WDATA => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_WDATA,
      x_rsc_13_0_AWREADY => x_rsc_13_0_AWREADY,
      x_rsc_13_0_AWVALID => x_rsc_13_0_AWVALID,
      x_rsc_13_0_AWUSER => x_rsc_13_0_AWUSER,
      x_rsc_13_0_AWREGION => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWREGION,
      x_rsc_13_0_AWQOS => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWQOS,
      x_rsc_13_0_AWPROT => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWPROT,
      x_rsc_13_0_AWCACHE => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWCACHE,
      x_rsc_13_0_AWLOCK => x_rsc_13_0_AWLOCK,
      x_rsc_13_0_AWBURST => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWBURST,
      x_rsc_13_0_AWSIZE => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWSIZE,
      x_rsc_13_0_AWLEN => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWLEN,
      x_rsc_13_0_AWADDR => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWADDR,
      x_rsc_13_0_AWID => x_rsc_13_0_AWID,
      core_wen => core_wen,
      x_rsc_13_0_i_oswt => reg_x_rsc_13_0_i_oswt_cse,
      x_rsc_13_0_i_wen_comp => x_rsc_13_0_i_wen_comp,
      x_rsc_13_0_i_oswt_1 => reg_x_rsc_13_0_i_oswt_1_cse,
      x_rsc_13_0_i_wen_comp_1 => x_rsc_13_0_i_wen_comp_1,
      x_rsc_13_0_i_s_raddr_core => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_raddr_core,
      x_rsc_13_0_i_s_waddr_core => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_waddr_core,
      x_rsc_13_0_i_s_din_mxwt => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_din_mxwt,
      x_rsc_13_0_i_s_dout_core => hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_dout_core
    );
  x_rsc_13_0_RRESP <= hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_RRESP;
  x_rsc_13_0_RDATA <= hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_RDATA;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARREGION <= x_rsc_13_0_ARREGION;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARQOS <= x_rsc_13_0_ARQOS;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARPROT <= x_rsc_13_0_ARPROT;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARCACHE <= x_rsc_13_0_ARCACHE;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARBURST <= x_rsc_13_0_ARBURST;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARSIZE <= x_rsc_13_0_ARSIZE;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARLEN <= x_rsc_13_0_ARLEN;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_ARADDR <= x_rsc_13_0_ARADDR;
  x_rsc_13_0_BRESP <= hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_BRESP;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_WSTRB <= x_rsc_13_0_WSTRB;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_WDATA <= x_rsc_13_0_WDATA;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWREGION <= x_rsc_13_0_AWREGION;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWQOS <= x_rsc_13_0_AWQOS;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWPROT <= x_rsc_13_0_AWPROT;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWCACHE <= x_rsc_13_0_AWCACHE;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWBURST <= x_rsc_13_0_AWBURST;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWSIZE <= x_rsc_13_0_AWSIZE;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWLEN <= x_rsc_13_0_AWLEN;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_AWADDR <= x_rsc_13_0_AWADDR;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_13_0_i_s_din_mxwt <= hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_din_mxwt;
  hybrid_core_x_rsc_13_0_i_inst_x_rsc_13_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_14_0_i_inst : hybrid_core_x_rsc_14_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_14_0_s_tdone => x_rsc_14_0_s_tdone,
      x_rsc_14_0_tr_write_done => x_rsc_14_0_tr_write_done,
      x_rsc_14_0_RREADY => x_rsc_14_0_RREADY,
      x_rsc_14_0_RVALID => x_rsc_14_0_RVALID,
      x_rsc_14_0_RUSER => x_rsc_14_0_RUSER,
      x_rsc_14_0_RLAST => x_rsc_14_0_RLAST,
      x_rsc_14_0_RRESP => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_RRESP,
      x_rsc_14_0_RDATA => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_RDATA,
      x_rsc_14_0_RID => x_rsc_14_0_RID,
      x_rsc_14_0_ARREADY => x_rsc_14_0_ARREADY,
      x_rsc_14_0_ARVALID => x_rsc_14_0_ARVALID,
      x_rsc_14_0_ARUSER => x_rsc_14_0_ARUSER,
      x_rsc_14_0_ARREGION => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARREGION,
      x_rsc_14_0_ARQOS => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARQOS,
      x_rsc_14_0_ARPROT => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARPROT,
      x_rsc_14_0_ARCACHE => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARCACHE,
      x_rsc_14_0_ARLOCK => x_rsc_14_0_ARLOCK,
      x_rsc_14_0_ARBURST => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARBURST,
      x_rsc_14_0_ARSIZE => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARSIZE,
      x_rsc_14_0_ARLEN => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARLEN,
      x_rsc_14_0_ARADDR => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARADDR,
      x_rsc_14_0_ARID => x_rsc_14_0_ARID,
      x_rsc_14_0_BREADY => x_rsc_14_0_BREADY,
      x_rsc_14_0_BVALID => x_rsc_14_0_BVALID,
      x_rsc_14_0_BUSER => x_rsc_14_0_BUSER,
      x_rsc_14_0_BRESP => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_BRESP,
      x_rsc_14_0_BID => x_rsc_14_0_BID,
      x_rsc_14_0_WREADY => x_rsc_14_0_WREADY,
      x_rsc_14_0_WVALID => x_rsc_14_0_WVALID,
      x_rsc_14_0_WUSER => x_rsc_14_0_WUSER,
      x_rsc_14_0_WLAST => x_rsc_14_0_WLAST,
      x_rsc_14_0_WSTRB => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_WSTRB,
      x_rsc_14_0_WDATA => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_WDATA,
      x_rsc_14_0_AWREADY => x_rsc_14_0_AWREADY,
      x_rsc_14_0_AWVALID => x_rsc_14_0_AWVALID,
      x_rsc_14_0_AWUSER => x_rsc_14_0_AWUSER,
      x_rsc_14_0_AWREGION => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWREGION,
      x_rsc_14_0_AWQOS => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWQOS,
      x_rsc_14_0_AWPROT => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWPROT,
      x_rsc_14_0_AWCACHE => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWCACHE,
      x_rsc_14_0_AWLOCK => x_rsc_14_0_AWLOCK,
      x_rsc_14_0_AWBURST => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWBURST,
      x_rsc_14_0_AWSIZE => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWSIZE,
      x_rsc_14_0_AWLEN => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWLEN,
      x_rsc_14_0_AWADDR => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWADDR,
      x_rsc_14_0_AWID => x_rsc_14_0_AWID,
      core_wen => core_wen,
      x_rsc_14_0_i_oswt => reg_x_rsc_14_0_i_oswt_cse,
      x_rsc_14_0_i_wen_comp => x_rsc_14_0_i_wen_comp,
      x_rsc_14_0_i_oswt_1 => reg_x_rsc_14_0_i_oswt_1_cse,
      x_rsc_14_0_i_wen_comp_1 => x_rsc_14_0_i_wen_comp_1,
      x_rsc_14_0_i_s_raddr_core => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_raddr_core,
      x_rsc_14_0_i_s_waddr_core => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_waddr_core,
      x_rsc_14_0_i_s_din_mxwt => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_din_mxwt,
      x_rsc_14_0_i_s_dout_core => hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_dout_core
    );
  x_rsc_14_0_RRESP <= hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_RRESP;
  x_rsc_14_0_RDATA <= hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_RDATA;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARREGION <= x_rsc_14_0_ARREGION;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARQOS <= x_rsc_14_0_ARQOS;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARPROT <= x_rsc_14_0_ARPROT;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARCACHE <= x_rsc_14_0_ARCACHE;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARBURST <= x_rsc_14_0_ARBURST;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARSIZE <= x_rsc_14_0_ARSIZE;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARLEN <= x_rsc_14_0_ARLEN;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_ARADDR <= x_rsc_14_0_ARADDR;
  x_rsc_14_0_BRESP <= hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_BRESP;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_WSTRB <= x_rsc_14_0_WSTRB;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_WDATA <= x_rsc_14_0_WDATA;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWREGION <= x_rsc_14_0_AWREGION;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWQOS <= x_rsc_14_0_AWQOS;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWPROT <= x_rsc_14_0_AWPROT;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWCACHE <= x_rsc_14_0_AWCACHE;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWBURST <= x_rsc_14_0_AWBURST;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWSIZE <= x_rsc_14_0_AWSIZE;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWLEN <= x_rsc_14_0_AWLEN;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_AWADDR <= x_rsc_14_0_AWADDR;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_14_0_i_s_din_mxwt <= hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_din_mxwt;
  hybrid_core_x_rsc_14_0_i_inst_x_rsc_14_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_15_0_i_inst : hybrid_core_x_rsc_15_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_15_0_s_tdone => x_rsc_15_0_s_tdone,
      x_rsc_15_0_tr_write_done => x_rsc_15_0_tr_write_done,
      x_rsc_15_0_RREADY => x_rsc_15_0_RREADY,
      x_rsc_15_0_RVALID => x_rsc_15_0_RVALID,
      x_rsc_15_0_RUSER => x_rsc_15_0_RUSER,
      x_rsc_15_0_RLAST => x_rsc_15_0_RLAST,
      x_rsc_15_0_RRESP => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_RRESP,
      x_rsc_15_0_RDATA => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_RDATA,
      x_rsc_15_0_RID => x_rsc_15_0_RID,
      x_rsc_15_0_ARREADY => x_rsc_15_0_ARREADY,
      x_rsc_15_0_ARVALID => x_rsc_15_0_ARVALID,
      x_rsc_15_0_ARUSER => x_rsc_15_0_ARUSER,
      x_rsc_15_0_ARREGION => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARREGION,
      x_rsc_15_0_ARQOS => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARQOS,
      x_rsc_15_0_ARPROT => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARPROT,
      x_rsc_15_0_ARCACHE => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARCACHE,
      x_rsc_15_0_ARLOCK => x_rsc_15_0_ARLOCK,
      x_rsc_15_0_ARBURST => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARBURST,
      x_rsc_15_0_ARSIZE => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARSIZE,
      x_rsc_15_0_ARLEN => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARLEN,
      x_rsc_15_0_ARADDR => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARADDR,
      x_rsc_15_0_ARID => x_rsc_15_0_ARID,
      x_rsc_15_0_BREADY => x_rsc_15_0_BREADY,
      x_rsc_15_0_BVALID => x_rsc_15_0_BVALID,
      x_rsc_15_0_BUSER => x_rsc_15_0_BUSER,
      x_rsc_15_0_BRESP => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_BRESP,
      x_rsc_15_0_BID => x_rsc_15_0_BID,
      x_rsc_15_0_WREADY => x_rsc_15_0_WREADY,
      x_rsc_15_0_WVALID => x_rsc_15_0_WVALID,
      x_rsc_15_0_WUSER => x_rsc_15_0_WUSER,
      x_rsc_15_0_WLAST => x_rsc_15_0_WLAST,
      x_rsc_15_0_WSTRB => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_WSTRB,
      x_rsc_15_0_WDATA => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_WDATA,
      x_rsc_15_0_AWREADY => x_rsc_15_0_AWREADY,
      x_rsc_15_0_AWVALID => x_rsc_15_0_AWVALID,
      x_rsc_15_0_AWUSER => x_rsc_15_0_AWUSER,
      x_rsc_15_0_AWREGION => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWREGION,
      x_rsc_15_0_AWQOS => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWQOS,
      x_rsc_15_0_AWPROT => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWPROT,
      x_rsc_15_0_AWCACHE => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWCACHE,
      x_rsc_15_0_AWLOCK => x_rsc_15_0_AWLOCK,
      x_rsc_15_0_AWBURST => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWBURST,
      x_rsc_15_0_AWSIZE => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWSIZE,
      x_rsc_15_0_AWLEN => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWLEN,
      x_rsc_15_0_AWADDR => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWADDR,
      x_rsc_15_0_AWID => x_rsc_15_0_AWID,
      core_wen => core_wen,
      x_rsc_15_0_i_oswt => reg_x_rsc_15_0_i_oswt_cse,
      x_rsc_15_0_i_wen_comp => x_rsc_15_0_i_wen_comp,
      x_rsc_15_0_i_oswt_1 => reg_x_rsc_15_0_i_oswt_1_cse,
      x_rsc_15_0_i_wen_comp_1 => x_rsc_15_0_i_wen_comp_1,
      x_rsc_15_0_i_s_raddr_core => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_raddr_core,
      x_rsc_15_0_i_s_waddr_core => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_waddr_core,
      x_rsc_15_0_i_s_din_mxwt => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_din_mxwt,
      x_rsc_15_0_i_s_dout_core => hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_dout_core
    );
  x_rsc_15_0_RRESP <= hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_RRESP;
  x_rsc_15_0_RDATA <= hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_RDATA;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARREGION <= x_rsc_15_0_ARREGION;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARQOS <= x_rsc_15_0_ARQOS;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARPROT <= x_rsc_15_0_ARPROT;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARCACHE <= x_rsc_15_0_ARCACHE;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARBURST <= x_rsc_15_0_ARBURST;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARSIZE <= x_rsc_15_0_ARSIZE;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARLEN <= x_rsc_15_0_ARLEN;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_ARADDR <= x_rsc_15_0_ARADDR;
  x_rsc_15_0_BRESP <= hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_BRESP;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_WSTRB <= x_rsc_15_0_WSTRB;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_WDATA <= x_rsc_15_0_WDATA;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWREGION <= x_rsc_15_0_AWREGION;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWQOS <= x_rsc_15_0_AWQOS;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWPROT <= x_rsc_15_0_AWPROT;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWCACHE <= x_rsc_15_0_AWCACHE;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWBURST <= x_rsc_15_0_AWBURST;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWSIZE <= x_rsc_15_0_AWSIZE;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWLEN <= x_rsc_15_0_AWLEN;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_AWADDR <= x_rsc_15_0_AWADDR;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_15_0_i_s_din_mxwt <= hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_din_mxwt;
  hybrid_core_x_rsc_15_0_i_inst_x_rsc_15_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_16_0_i_inst : hybrid_core_x_rsc_16_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_16_0_s_tdone => x_rsc_16_0_s_tdone,
      x_rsc_16_0_tr_write_done => x_rsc_16_0_tr_write_done,
      x_rsc_16_0_RREADY => x_rsc_16_0_RREADY,
      x_rsc_16_0_RVALID => x_rsc_16_0_RVALID,
      x_rsc_16_0_RUSER => x_rsc_16_0_RUSER,
      x_rsc_16_0_RLAST => x_rsc_16_0_RLAST,
      x_rsc_16_0_RRESP => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_RRESP,
      x_rsc_16_0_RDATA => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_RDATA,
      x_rsc_16_0_RID => x_rsc_16_0_RID,
      x_rsc_16_0_ARREADY => x_rsc_16_0_ARREADY,
      x_rsc_16_0_ARVALID => x_rsc_16_0_ARVALID,
      x_rsc_16_0_ARUSER => x_rsc_16_0_ARUSER,
      x_rsc_16_0_ARREGION => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARREGION,
      x_rsc_16_0_ARQOS => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARQOS,
      x_rsc_16_0_ARPROT => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARPROT,
      x_rsc_16_0_ARCACHE => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARCACHE,
      x_rsc_16_0_ARLOCK => x_rsc_16_0_ARLOCK,
      x_rsc_16_0_ARBURST => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARBURST,
      x_rsc_16_0_ARSIZE => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARSIZE,
      x_rsc_16_0_ARLEN => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARLEN,
      x_rsc_16_0_ARADDR => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARADDR,
      x_rsc_16_0_ARID => x_rsc_16_0_ARID,
      x_rsc_16_0_BREADY => x_rsc_16_0_BREADY,
      x_rsc_16_0_BVALID => x_rsc_16_0_BVALID,
      x_rsc_16_0_BUSER => x_rsc_16_0_BUSER,
      x_rsc_16_0_BRESP => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_BRESP,
      x_rsc_16_0_BID => x_rsc_16_0_BID,
      x_rsc_16_0_WREADY => x_rsc_16_0_WREADY,
      x_rsc_16_0_WVALID => x_rsc_16_0_WVALID,
      x_rsc_16_0_WUSER => x_rsc_16_0_WUSER,
      x_rsc_16_0_WLAST => x_rsc_16_0_WLAST,
      x_rsc_16_0_WSTRB => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_WSTRB,
      x_rsc_16_0_WDATA => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_WDATA,
      x_rsc_16_0_AWREADY => x_rsc_16_0_AWREADY,
      x_rsc_16_0_AWVALID => x_rsc_16_0_AWVALID,
      x_rsc_16_0_AWUSER => x_rsc_16_0_AWUSER,
      x_rsc_16_0_AWREGION => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWREGION,
      x_rsc_16_0_AWQOS => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWQOS,
      x_rsc_16_0_AWPROT => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWPROT,
      x_rsc_16_0_AWCACHE => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWCACHE,
      x_rsc_16_0_AWLOCK => x_rsc_16_0_AWLOCK,
      x_rsc_16_0_AWBURST => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWBURST,
      x_rsc_16_0_AWSIZE => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWSIZE,
      x_rsc_16_0_AWLEN => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWLEN,
      x_rsc_16_0_AWADDR => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWADDR,
      x_rsc_16_0_AWID => x_rsc_16_0_AWID,
      core_wen => core_wen,
      x_rsc_16_0_i_oswt => reg_x_rsc_16_0_i_oswt_cse,
      x_rsc_16_0_i_wen_comp => x_rsc_16_0_i_wen_comp,
      x_rsc_16_0_i_oswt_1 => reg_x_rsc_16_0_i_oswt_1_cse,
      x_rsc_16_0_i_wen_comp_1 => x_rsc_16_0_i_wen_comp_1,
      x_rsc_16_0_i_s_raddr_core => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_raddr_core,
      x_rsc_16_0_i_s_waddr_core => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_waddr_core,
      x_rsc_16_0_i_s_din_mxwt => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_din_mxwt,
      x_rsc_16_0_i_s_dout_core => hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_dout_core
    );
  x_rsc_16_0_RRESP <= hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_RRESP;
  x_rsc_16_0_RDATA <= hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_RDATA;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARREGION <= x_rsc_16_0_ARREGION;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARQOS <= x_rsc_16_0_ARQOS;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARPROT <= x_rsc_16_0_ARPROT;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARCACHE <= x_rsc_16_0_ARCACHE;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARBURST <= x_rsc_16_0_ARBURST;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARSIZE <= x_rsc_16_0_ARSIZE;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARLEN <= x_rsc_16_0_ARLEN;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_ARADDR <= x_rsc_16_0_ARADDR;
  x_rsc_16_0_BRESP <= hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_BRESP;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_WSTRB <= x_rsc_16_0_WSTRB;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_WDATA <= x_rsc_16_0_WDATA;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWREGION <= x_rsc_16_0_AWREGION;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWQOS <= x_rsc_16_0_AWQOS;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWPROT <= x_rsc_16_0_AWPROT;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWCACHE <= x_rsc_16_0_AWCACHE;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWBURST <= x_rsc_16_0_AWBURST;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWSIZE <= x_rsc_16_0_AWSIZE;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWLEN <= x_rsc_16_0_AWLEN;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_AWADDR <= x_rsc_16_0_AWADDR;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_16_0_i_s_din_mxwt <= hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_din_mxwt;
  hybrid_core_x_rsc_16_0_i_inst_x_rsc_16_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_17_0_i_inst : hybrid_core_x_rsc_17_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_17_0_s_tdone => x_rsc_17_0_s_tdone,
      x_rsc_17_0_tr_write_done => x_rsc_17_0_tr_write_done,
      x_rsc_17_0_RREADY => x_rsc_17_0_RREADY,
      x_rsc_17_0_RVALID => x_rsc_17_0_RVALID,
      x_rsc_17_0_RUSER => x_rsc_17_0_RUSER,
      x_rsc_17_0_RLAST => x_rsc_17_0_RLAST,
      x_rsc_17_0_RRESP => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_RRESP,
      x_rsc_17_0_RDATA => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_RDATA,
      x_rsc_17_0_RID => x_rsc_17_0_RID,
      x_rsc_17_0_ARREADY => x_rsc_17_0_ARREADY,
      x_rsc_17_0_ARVALID => x_rsc_17_0_ARVALID,
      x_rsc_17_0_ARUSER => x_rsc_17_0_ARUSER,
      x_rsc_17_0_ARREGION => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARREGION,
      x_rsc_17_0_ARQOS => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARQOS,
      x_rsc_17_0_ARPROT => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARPROT,
      x_rsc_17_0_ARCACHE => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARCACHE,
      x_rsc_17_0_ARLOCK => x_rsc_17_0_ARLOCK,
      x_rsc_17_0_ARBURST => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARBURST,
      x_rsc_17_0_ARSIZE => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARSIZE,
      x_rsc_17_0_ARLEN => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARLEN,
      x_rsc_17_0_ARADDR => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARADDR,
      x_rsc_17_0_ARID => x_rsc_17_0_ARID,
      x_rsc_17_0_BREADY => x_rsc_17_0_BREADY,
      x_rsc_17_0_BVALID => x_rsc_17_0_BVALID,
      x_rsc_17_0_BUSER => x_rsc_17_0_BUSER,
      x_rsc_17_0_BRESP => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_BRESP,
      x_rsc_17_0_BID => x_rsc_17_0_BID,
      x_rsc_17_0_WREADY => x_rsc_17_0_WREADY,
      x_rsc_17_0_WVALID => x_rsc_17_0_WVALID,
      x_rsc_17_0_WUSER => x_rsc_17_0_WUSER,
      x_rsc_17_0_WLAST => x_rsc_17_0_WLAST,
      x_rsc_17_0_WSTRB => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_WSTRB,
      x_rsc_17_0_WDATA => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_WDATA,
      x_rsc_17_0_AWREADY => x_rsc_17_0_AWREADY,
      x_rsc_17_0_AWVALID => x_rsc_17_0_AWVALID,
      x_rsc_17_0_AWUSER => x_rsc_17_0_AWUSER,
      x_rsc_17_0_AWREGION => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWREGION,
      x_rsc_17_0_AWQOS => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWQOS,
      x_rsc_17_0_AWPROT => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWPROT,
      x_rsc_17_0_AWCACHE => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWCACHE,
      x_rsc_17_0_AWLOCK => x_rsc_17_0_AWLOCK,
      x_rsc_17_0_AWBURST => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWBURST,
      x_rsc_17_0_AWSIZE => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWSIZE,
      x_rsc_17_0_AWLEN => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWLEN,
      x_rsc_17_0_AWADDR => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWADDR,
      x_rsc_17_0_AWID => x_rsc_17_0_AWID,
      core_wen => core_wen,
      x_rsc_17_0_i_oswt => reg_x_rsc_17_0_i_oswt_cse,
      x_rsc_17_0_i_wen_comp => x_rsc_17_0_i_wen_comp,
      x_rsc_17_0_i_oswt_1 => reg_x_rsc_17_0_i_oswt_1_cse,
      x_rsc_17_0_i_wen_comp_1 => x_rsc_17_0_i_wen_comp_1,
      x_rsc_17_0_i_s_raddr_core => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_raddr_core,
      x_rsc_17_0_i_s_waddr_core => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_waddr_core,
      x_rsc_17_0_i_s_din_mxwt => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_din_mxwt,
      x_rsc_17_0_i_s_dout_core => hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_dout_core
    );
  x_rsc_17_0_RRESP <= hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_RRESP;
  x_rsc_17_0_RDATA <= hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_RDATA;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARREGION <= x_rsc_17_0_ARREGION;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARQOS <= x_rsc_17_0_ARQOS;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARPROT <= x_rsc_17_0_ARPROT;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARCACHE <= x_rsc_17_0_ARCACHE;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARBURST <= x_rsc_17_0_ARBURST;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARSIZE <= x_rsc_17_0_ARSIZE;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARLEN <= x_rsc_17_0_ARLEN;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_ARADDR <= x_rsc_17_0_ARADDR;
  x_rsc_17_0_BRESP <= hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_BRESP;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_WSTRB <= x_rsc_17_0_WSTRB;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_WDATA <= x_rsc_17_0_WDATA;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWREGION <= x_rsc_17_0_AWREGION;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWQOS <= x_rsc_17_0_AWQOS;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWPROT <= x_rsc_17_0_AWPROT;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWCACHE <= x_rsc_17_0_AWCACHE;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWBURST <= x_rsc_17_0_AWBURST;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWSIZE <= x_rsc_17_0_AWSIZE;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWLEN <= x_rsc_17_0_AWLEN;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_AWADDR <= x_rsc_17_0_AWADDR;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_17_0_i_s_din_mxwt <= hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_din_mxwt;
  hybrid_core_x_rsc_17_0_i_inst_x_rsc_17_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_18_0_i_inst : hybrid_core_x_rsc_18_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_18_0_s_tdone => x_rsc_18_0_s_tdone,
      x_rsc_18_0_tr_write_done => x_rsc_18_0_tr_write_done,
      x_rsc_18_0_RREADY => x_rsc_18_0_RREADY,
      x_rsc_18_0_RVALID => x_rsc_18_0_RVALID,
      x_rsc_18_0_RUSER => x_rsc_18_0_RUSER,
      x_rsc_18_0_RLAST => x_rsc_18_0_RLAST,
      x_rsc_18_0_RRESP => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_RRESP,
      x_rsc_18_0_RDATA => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_RDATA,
      x_rsc_18_0_RID => x_rsc_18_0_RID,
      x_rsc_18_0_ARREADY => x_rsc_18_0_ARREADY,
      x_rsc_18_0_ARVALID => x_rsc_18_0_ARVALID,
      x_rsc_18_0_ARUSER => x_rsc_18_0_ARUSER,
      x_rsc_18_0_ARREGION => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARREGION,
      x_rsc_18_0_ARQOS => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARQOS,
      x_rsc_18_0_ARPROT => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARPROT,
      x_rsc_18_0_ARCACHE => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARCACHE,
      x_rsc_18_0_ARLOCK => x_rsc_18_0_ARLOCK,
      x_rsc_18_0_ARBURST => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARBURST,
      x_rsc_18_0_ARSIZE => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARSIZE,
      x_rsc_18_0_ARLEN => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARLEN,
      x_rsc_18_0_ARADDR => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARADDR,
      x_rsc_18_0_ARID => x_rsc_18_0_ARID,
      x_rsc_18_0_BREADY => x_rsc_18_0_BREADY,
      x_rsc_18_0_BVALID => x_rsc_18_0_BVALID,
      x_rsc_18_0_BUSER => x_rsc_18_0_BUSER,
      x_rsc_18_0_BRESP => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_BRESP,
      x_rsc_18_0_BID => x_rsc_18_0_BID,
      x_rsc_18_0_WREADY => x_rsc_18_0_WREADY,
      x_rsc_18_0_WVALID => x_rsc_18_0_WVALID,
      x_rsc_18_0_WUSER => x_rsc_18_0_WUSER,
      x_rsc_18_0_WLAST => x_rsc_18_0_WLAST,
      x_rsc_18_0_WSTRB => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_WSTRB,
      x_rsc_18_0_WDATA => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_WDATA,
      x_rsc_18_0_AWREADY => x_rsc_18_0_AWREADY,
      x_rsc_18_0_AWVALID => x_rsc_18_0_AWVALID,
      x_rsc_18_0_AWUSER => x_rsc_18_0_AWUSER,
      x_rsc_18_0_AWREGION => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWREGION,
      x_rsc_18_0_AWQOS => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWQOS,
      x_rsc_18_0_AWPROT => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWPROT,
      x_rsc_18_0_AWCACHE => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWCACHE,
      x_rsc_18_0_AWLOCK => x_rsc_18_0_AWLOCK,
      x_rsc_18_0_AWBURST => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWBURST,
      x_rsc_18_0_AWSIZE => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWSIZE,
      x_rsc_18_0_AWLEN => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWLEN,
      x_rsc_18_0_AWADDR => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWADDR,
      x_rsc_18_0_AWID => x_rsc_18_0_AWID,
      core_wen => core_wen,
      x_rsc_18_0_i_oswt => reg_x_rsc_18_0_i_oswt_cse,
      x_rsc_18_0_i_wen_comp => x_rsc_18_0_i_wen_comp,
      x_rsc_18_0_i_oswt_1 => reg_x_rsc_18_0_i_oswt_1_cse,
      x_rsc_18_0_i_wen_comp_1 => x_rsc_18_0_i_wen_comp_1,
      x_rsc_18_0_i_s_raddr_core => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_raddr_core,
      x_rsc_18_0_i_s_waddr_core => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_waddr_core,
      x_rsc_18_0_i_s_din_mxwt => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_din_mxwt,
      x_rsc_18_0_i_s_dout_core => hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_dout_core
    );
  x_rsc_18_0_RRESP <= hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_RRESP;
  x_rsc_18_0_RDATA <= hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_RDATA;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARREGION <= x_rsc_18_0_ARREGION;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARQOS <= x_rsc_18_0_ARQOS;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARPROT <= x_rsc_18_0_ARPROT;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARCACHE <= x_rsc_18_0_ARCACHE;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARBURST <= x_rsc_18_0_ARBURST;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARSIZE <= x_rsc_18_0_ARSIZE;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARLEN <= x_rsc_18_0_ARLEN;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_ARADDR <= x_rsc_18_0_ARADDR;
  x_rsc_18_0_BRESP <= hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_BRESP;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_WSTRB <= x_rsc_18_0_WSTRB;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_WDATA <= x_rsc_18_0_WDATA;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWREGION <= x_rsc_18_0_AWREGION;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWQOS <= x_rsc_18_0_AWQOS;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWPROT <= x_rsc_18_0_AWPROT;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWCACHE <= x_rsc_18_0_AWCACHE;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWBURST <= x_rsc_18_0_AWBURST;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWSIZE <= x_rsc_18_0_AWSIZE;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWLEN <= x_rsc_18_0_AWLEN;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_AWADDR <= x_rsc_18_0_AWADDR;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_18_0_i_s_din_mxwt <= hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_din_mxwt;
  hybrid_core_x_rsc_18_0_i_inst_x_rsc_18_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_19_0_i_inst : hybrid_core_x_rsc_19_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_19_0_s_tdone => x_rsc_19_0_s_tdone,
      x_rsc_19_0_tr_write_done => x_rsc_19_0_tr_write_done,
      x_rsc_19_0_RREADY => x_rsc_19_0_RREADY,
      x_rsc_19_0_RVALID => x_rsc_19_0_RVALID,
      x_rsc_19_0_RUSER => x_rsc_19_0_RUSER,
      x_rsc_19_0_RLAST => x_rsc_19_0_RLAST,
      x_rsc_19_0_RRESP => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_RRESP,
      x_rsc_19_0_RDATA => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_RDATA,
      x_rsc_19_0_RID => x_rsc_19_0_RID,
      x_rsc_19_0_ARREADY => x_rsc_19_0_ARREADY,
      x_rsc_19_0_ARVALID => x_rsc_19_0_ARVALID,
      x_rsc_19_0_ARUSER => x_rsc_19_0_ARUSER,
      x_rsc_19_0_ARREGION => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARREGION,
      x_rsc_19_0_ARQOS => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARQOS,
      x_rsc_19_0_ARPROT => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARPROT,
      x_rsc_19_0_ARCACHE => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARCACHE,
      x_rsc_19_0_ARLOCK => x_rsc_19_0_ARLOCK,
      x_rsc_19_0_ARBURST => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARBURST,
      x_rsc_19_0_ARSIZE => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARSIZE,
      x_rsc_19_0_ARLEN => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARLEN,
      x_rsc_19_0_ARADDR => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARADDR,
      x_rsc_19_0_ARID => x_rsc_19_0_ARID,
      x_rsc_19_0_BREADY => x_rsc_19_0_BREADY,
      x_rsc_19_0_BVALID => x_rsc_19_0_BVALID,
      x_rsc_19_0_BUSER => x_rsc_19_0_BUSER,
      x_rsc_19_0_BRESP => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_BRESP,
      x_rsc_19_0_BID => x_rsc_19_0_BID,
      x_rsc_19_0_WREADY => x_rsc_19_0_WREADY,
      x_rsc_19_0_WVALID => x_rsc_19_0_WVALID,
      x_rsc_19_0_WUSER => x_rsc_19_0_WUSER,
      x_rsc_19_0_WLAST => x_rsc_19_0_WLAST,
      x_rsc_19_0_WSTRB => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_WSTRB,
      x_rsc_19_0_WDATA => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_WDATA,
      x_rsc_19_0_AWREADY => x_rsc_19_0_AWREADY,
      x_rsc_19_0_AWVALID => x_rsc_19_0_AWVALID,
      x_rsc_19_0_AWUSER => x_rsc_19_0_AWUSER,
      x_rsc_19_0_AWREGION => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWREGION,
      x_rsc_19_0_AWQOS => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWQOS,
      x_rsc_19_0_AWPROT => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWPROT,
      x_rsc_19_0_AWCACHE => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWCACHE,
      x_rsc_19_0_AWLOCK => x_rsc_19_0_AWLOCK,
      x_rsc_19_0_AWBURST => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWBURST,
      x_rsc_19_0_AWSIZE => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWSIZE,
      x_rsc_19_0_AWLEN => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWLEN,
      x_rsc_19_0_AWADDR => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWADDR,
      x_rsc_19_0_AWID => x_rsc_19_0_AWID,
      core_wen => core_wen,
      x_rsc_19_0_i_oswt => reg_x_rsc_19_0_i_oswt_cse,
      x_rsc_19_0_i_wen_comp => x_rsc_19_0_i_wen_comp,
      x_rsc_19_0_i_oswt_1 => reg_x_rsc_19_0_i_oswt_1_cse,
      x_rsc_19_0_i_wen_comp_1 => x_rsc_19_0_i_wen_comp_1,
      x_rsc_19_0_i_s_raddr_core => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_raddr_core,
      x_rsc_19_0_i_s_waddr_core => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_waddr_core,
      x_rsc_19_0_i_s_din_mxwt => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_din_mxwt,
      x_rsc_19_0_i_s_dout_core => hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_dout_core
    );
  x_rsc_19_0_RRESP <= hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_RRESP;
  x_rsc_19_0_RDATA <= hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_RDATA;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARREGION <= x_rsc_19_0_ARREGION;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARQOS <= x_rsc_19_0_ARQOS;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARPROT <= x_rsc_19_0_ARPROT;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARCACHE <= x_rsc_19_0_ARCACHE;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARBURST <= x_rsc_19_0_ARBURST;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARSIZE <= x_rsc_19_0_ARSIZE;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARLEN <= x_rsc_19_0_ARLEN;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_ARADDR <= x_rsc_19_0_ARADDR;
  x_rsc_19_0_BRESP <= hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_BRESP;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_WSTRB <= x_rsc_19_0_WSTRB;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_WDATA <= x_rsc_19_0_WDATA;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWREGION <= x_rsc_19_0_AWREGION;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWQOS <= x_rsc_19_0_AWQOS;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWPROT <= x_rsc_19_0_AWPROT;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWCACHE <= x_rsc_19_0_AWCACHE;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWBURST <= x_rsc_19_0_AWBURST;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWSIZE <= x_rsc_19_0_AWSIZE;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWLEN <= x_rsc_19_0_AWLEN;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_AWADDR <= x_rsc_19_0_AWADDR;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_19_0_i_s_din_mxwt <= hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_din_mxwt;
  hybrid_core_x_rsc_19_0_i_inst_x_rsc_19_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_20_0_i_inst : hybrid_core_x_rsc_20_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_20_0_s_tdone => x_rsc_20_0_s_tdone,
      x_rsc_20_0_tr_write_done => x_rsc_20_0_tr_write_done,
      x_rsc_20_0_RREADY => x_rsc_20_0_RREADY,
      x_rsc_20_0_RVALID => x_rsc_20_0_RVALID,
      x_rsc_20_0_RUSER => x_rsc_20_0_RUSER,
      x_rsc_20_0_RLAST => x_rsc_20_0_RLAST,
      x_rsc_20_0_RRESP => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_RRESP,
      x_rsc_20_0_RDATA => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_RDATA,
      x_rsc_20_0_RID => x_rsc_20_0_RID,
      x_rsc_20_0_ARREADY => x_rsc_20_0_ARREADY,
      x_rsc_20_0_ARVALID => x_rsc_20_0_ARVALID,
      x_rsc_20_0_ARUSER => x_rsc_20_0_ARUSER,
      x_rsc_20_0_ARREGION => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARREGION,
      x_rsc_20_0_ARQOS => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARQOS,
      x_rsc_20_0_ARPROT => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARPROT,
      x_rsc_20_0_ARCACHE => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARCACHE,
      x_rsc_20_0_ARLOCK => x_rsc_20_0_ARLOCK,
      x_rsc_20_0_ARBURST => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARBURST,
      x_rsc_20_0_ARSIZE => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARSIZE,
      x_rsc_20_0_ARLEN => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARLEN,
      x_rsc_20_0_ARADDR => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARADDR,
      x_rsc_20_0_ARID => x_rsc_20_0_ARID,
      x_rsc_20_0_BREADY => x_rsc_20_0_BREADY,
      x_rsc_20_0_BVALID => x_rsc_20_0_BVALID,
      x_rsc_20_0_BUSER => x_rsc_20_0_BUSER,
      x_rsc_20_0_BRESP => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_BRESP,
      x_rsc_20_0_BID => x_rsc_20_0_BID,
      x_rsc_20_0_WREADY => x_rsc_20_0_WREADY,
      x_rsc_20_0_WVALID => x_rsc_20_0_WVALID,
      x_rsc_20_0_WUSER => x_rsc_20_0_WUSER,
      x_rsc_20_0_WLAST => x_rsc_20_0_WLAST,
      x_rsc_20_0_WSTRB => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_WSTRB,
      x_rsc_20_0_WDATA => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_WDATA,
      x_rsc_20_0_AWREADY => x_rsc_20_0_AWREADY,
      x_rsc_20_0_AWVALID => x_rsc_20_0_AWVALID,
      x_rsc_20_0_AWUSER => x_rsc_20_0_AWUSER,
      x_rsc_20_0_AWREGION => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWREGION,
      x_rsc_20_0_AWQOS => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWQOS,
      x_rsc_20_0_AWPROT => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWPROT,
      x_rsc_20_0_AWCACHE => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWCACHE,
      x_rsc_20_0_AWLOCK => x_rsc_20_0_AWLOCK,
      x_rsc_20_0_AWBURST => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWBURST,
      x_rsc_20_0_AWSIZE => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWSIZE,
      x_rsc_20_0_AWLEN => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWLEN,
      x_rsc_20_0_AWADDR => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWADDR,
      x_rsc_20_0_AWID => x_rsc_20_0_AWID,
      core_wen => core_wen,
      x_rsc_20_0_i_oswt => reg_x_rsc_20_0_i_oswt_cse,
      x_rsc_20_0_i_wen_comp => x_rsc_20_0_i_wen_comp,
      x_rsc_20_0_i_oswt_1 => reg_x_rsc_20_0_i_oswt_1_cse,
      x_rsc_20_0_i_wen_comp_1 => x_rsc_20_0_i_wen_comp_1,
      x_rsc_20_0_i_s_raddr_core => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_raddr_core,
      x_rsc_20_0_i_s_waddr_core => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_waddr_core,
      x_rsc_20_0_i_s_din_mxwt => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_din_mxwt,
      x_rsc_20_0_i_s_dout_core => hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_dout_core
    );
  x_rsc_20_0_RRESP <= hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_RRESP;
  x_rsc_20_0_RDATA <= hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_RDATA;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARREGION <= x_rsc_20_0_ARREGION;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARQOS <= x_rsc_20_0_ARQOS;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARPROT <= x_rsc_20_0_ARPROT;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARCACHE <= x_rsc_20_0_ARCACHE;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARBURST <= x_rsc_20_0_ARBURST;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARSIZE <= x_rsc_20_0_ARSIZE;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARLEN <= x_rsc_20_0_ARLEN;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_ARADDR <= x_rsc_20_0_ARADDR;
  x_rsc_20_0_BRESP <= hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_BRESP;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_WSTRB <= x_rsc_20_0_WSTRB;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_WDATA <= x_rsc_20_0_WDATA;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWREGION <= x_rsc_20_0_AWREGION;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWQOS <= x_rsc_20_0_AWQOS;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWPROT <= x_rsc_20_0_AWPROT;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWCACHE <= x_rsc_20_0_AWCACHE;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWBURST <= x_rsc_20_0_AWBURST;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWSIZE <= x_rsc_20_0_AWSIZE;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWLEN <= x_rsc_20_0_AWLEN;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_AWADDR <= x_rsc_20_0_AWADDR;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_20_0_i_s_din_mxwt <= hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_din_mxwt;
  hybrid_core_x_rsc_20_0_i_inst_x_rsc_20_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_21_0_i_inst : hybrid_core_x_rsc_21_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_21_0_s_tdone => x_rsc_21_0_s_tdone,
      x_rsc_21_0_tr_write_done => x_rsc_21_0_tr_write_done,
      x_rsc_21_0_RREADY => x_rsc_21_0_RREADY,
      x_rsc_21_0_RVALID => x_rsc_21_0_RVALID,
      x_rsc_21_0_RUSER => x_rsc_21_0_RUSER,
      x_rsc_21_0_RLAST => x_rsc_21_0_RLAST,
      x_rsc_21_0_RRESP => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_RRESP,
      x_rsc_21_0_RDATA => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_RDATA,
      x_rsc_21_0_RID => x_rsc_21_0_RID,
      x_rsc_21_0_ARREADY => x_rsc_21_0_ARREADY,
      x_rsc_21_0_ARVALID => x_rsc_21_0_ARVALID,
      x_rsc_21_0_ARUSER => x_rsc_21_0_ARUSER,
      x_rsc_21_0_ARREGION => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARREGION,
      x_rsc_21_0_ARQOS => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARQOS,
      x_rsc_21_0_ARPROT => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARPROT,
      x_rsc_21_0_ARCACHE => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARCACHE,
      x_rsc_21_0_ARLOCK => x_rsc_21_0_ARLOCK,
      x_rsc_21_0_ARBURST => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARBURST,
      x_rsc_21_0_ARSIZE => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARSIZE,
      x_rsc_21_0_ARLEN => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARLEN,
      x_rsc_21_0_ARADDR => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARADDR,
      x_rsc_21_0_ARID => x_rsc_21_0_ARID,
      x_rsc_21_0_BREADY => x_rsc_21_0_BREADY,
      x_rsc_21_0_BVALID => x_rsc_21_0_BVALID,
      x_rsc_21_0_BUSER => x_rsc_21_0_BUSER,
      x_rsc_21_0_BRESP => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_BRESP,
      x_rsc_21_0_BID => x_rsc_21_0_BID,
      x_rsc_21_0_WREADY => x_rsc_21_0_WREADY,
      x_rsc_21_0_WVALID => x_rsc_21_0_WVALID,
      x_rsc_21_0_WUSER => x_rsc_21_0_WUSER,
      x_rsc_21_0_WLAST => x_rsc_21_0_WLAST,
      x_rsc_21_0_WSTRB => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_WSTRB,
      x_rsc_21_0_WDATA => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_WDATA,
      x_rsc_21_0_AWREADY => x_rsc_21_0_AWREADY,
      x_rsc_21_0_AWVALID => x_rsc_21_0_AWVALID,
      x_rsc_21_0_AWUSER => x_rsc_21_0_AWUSER,
      x_rsc_21_0_AWREGION => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWREGION,
      x_rsc_21_0_AWQOS => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWQOS,
      x_rsc_21_0_AWPROT => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWPROT,
      x_rsc_21_0_AWCACHE => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWCACHE,
      x_rsc_21_0_AWLOCK => x_rsc_21_0_AWLOCK,
      x_rsc_21_0_AWBURST => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWBURST,
      x_rsc_21_0_AWSIZE => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWSIZE,
      x_rsc_21_0_AWLEN => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWLEN,
      x_rsc_21_0_AWADDR => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWADDR,
      x_rsc_21_0_AWID => x_rsc_21_0_AWID,
      core_wen => core_wen,
      x_rsc_21_0_i_oswt => reg_x_rsc_21_0_i_oswt_cse,
      x_rsc_21_0_i_wen_comp => x_rsc_21_0_i_wen_comp,
      x_rsc_21_0_i_oswt_1 => reg_x_rsc_21_0_i_oswt_1_cse,
      x_rsc_21_0_i_wen_comp_1 => x_rsc_21_0_i_wen_comp_1,
      x_rsc_21_0_i_s_raddr_core => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_raddr_core,
      x_rsc_21_0_i_s_waddr_core => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_waddr_core,
      x_rsc_21_0_i_s_din_mxwt => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_din_mxwt,
      x_rsc_21_0_i_s_dout_core => hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_dout_core
    );
  x_rsc_21_0_RRESP <= hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_RRESP;
  x_rsc_21_0_RDATA <= hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_RDATA;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARREGION <= x_rsc_21_0_ARREGION;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARQOS <= x_rsc_21_0_ARQOS;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARPROT <= x_rsc_21_0_ARPROT;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARCACHE <= x_rsc_21_0_ARCACHE;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARBURST <= x_rsc_21_0_ARBURST;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARSIZE <= x_rsc_21_0_ARSIZE;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARLEN <= x_rsc_21_0_ARLEN;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_ARADDR <= x_rsc_21_0_ARADDR;
  x_rsc_21_0_BRESP <= hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_BRESP;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_WSTRB <= x_rsc_21_0_WSTRB;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_WDATA <= x_rsc_21_0_WDATA;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWREGION <= x_rsc_21_0_AWREGION;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWQOS <= x_rsc_21_0_AWQOS;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWPROT <= x_rsc_21_0_AWPROT;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWCACHE <= x_rsc_21_0_AWCACHE;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWBURST <= x_rsc_21_0_AWBURST;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWSIZE <= x_rsc_21_0_AWSIZE;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWLEN <= x_rsc_21_0_AWLEN;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_AWADDR <= x_rsc_21_0_AWADDR;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_21_0_i_s_din_mxwt <= hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_din_mxwt;
  hybrid_core_x_rsc_21_0_i_inst_x_rsc_21_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_22_0_i_inst : hybrid_core_x_rsc_22_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_22_0_s_tdone => x_rsc_22_0_s_tdone,
      x_rsc_22_0_tr_write_done => x_rsc_22_0_tr_write_done,
      x_rsc_22_0_RREADY => x_rsc_22_0_RREADY,
      x_rsc_22_0_RVALID => x_rsc_22_0_RVALID,
      x_rsc_22_0_RUSER => x_rsc_22_0_RUSER,
      x_rsc_22_0_RLAST => x_rsc_22_0_RLAST,
      x_rsc_22_0_RRESP => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_RRESP,
      x_rsc_22_0_RDATA => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_RDATA,
      x_rsc_22_0_RID => x_rsc_22_0_RID,
      x_rsc_22_0_ARREADY => x_rsc_22_0_ARREADY,
      x_rsc_22_0_ARVALID => x_rsc_22_0_ARVALID,
      x_rsc_22_0_ARUSER => x_rsc_22_0_ARUSER,
      x_rsc_22_0_ARREGION => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARREGION,
      x_rsc_22_0_ARQOS => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARQOS,
      x_rsc_22_0_ARPROT => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARPROT,
      x_rsc_22_0_ARCACHE => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARCACHE,
      x_rsc_22_0_ARLOCK => x_rsc_22_0_ARLOCK,
      x_rsc_22_0_ARBURST => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARBURST,
      x_rsc_22_0_ARSIZE => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARSIZE,
      x_rsc_22_0_ARLEN => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARLEN,
      x_rsc_22_0_ARADDR => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARADDR,
      x_rsc_22_0_ARID => x_rsc_22_0_ARID,
      x_rsc_22_0_BREADY => x_rsc_22_0_BREADY,
      x_rsc_22_0_BVALID => x_rsc_22_0_BVALID,
      x_rsc_22_0_BUSER => x_rsc_22_0_BUSER,
      x_rsc_22_0_BRESP => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_BRESP,
      x_rsc_22_0_BID => x_rsc_22_0_BID,
      x_rsc_22_0_WREADY => x_rsc_22_0_WREADY,
      x_rsc_22_0_WVALID => x_rsc_22_0_WVALID,
      x_rsc_22_0_WUSER => x_rsc_22_0_WUSER,
      x_rsc_22_0_WLAST => x_rsc_22_0_WLAST,
      x_rsc_22_0_WSTRB => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_WSTRB,
      x_rsc_22_0_WDATA => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_WDATA,
      x_rsc_22_0_AWREADY => x_rsc_22_0_AWREADY,
      x_rsc_22_0_AWVALID => x_rsc_22_0_AWVALID,
      x_rsc_22_0_AWUSER => x_rsc_22_0_AWUSER,
      x_rsc_22_0_AWREGION => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWREGION,
      x_rsc_22_0_AWQOS => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWQOS,
      x_rsc_22_0_AWPROT => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWPROT,
      x_rsc_22_0_AWCACHE => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWCACHE,
      x_rsc_22_0_AWLOCK => x_rsc_22_0_AWLOCK,
      x_rsc_22_0_AWBURST => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWBURST,
      x_rsc_22_0_AWSIZE => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWSIZE,
      x_rsc_22_0_AWLEN => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWLEN,
      x_rsc_22_0_AWADDR => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWADDR,
      x_rsc_22_0_AWID => x_rsc_22_0_AWID,
      core_wen => core_wen,
      x_rsc_22_0_i_oswt => reg_x_rsc_22_0_i_oswt_cse,
      x_rsc_22_0_i_wen_comp => x_rsc_22_0_i_wen_comp,
      x_rsc_22_0_i_oswt_1 => reg_x_rsc_22_0_i_oswt_1_cse,
      x_rsc_22_0_i_wen_comp_1 => x_rsc_22_0_i_wen_comp_1,
      x_rsc_22_0_i_s_raddr_core => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_raddr_core,
      x_rsc_22_0_i_s_waddr_core => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_waddr_core,
      x_rsc_22_0_i_s_din_mxwt => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_din_mxwt,
      x_rsc_22_0_i_s_dout_core => hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_dout_core
    );
  x_rsc_22_0_RRESP <= hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_RRESP;
  x_rsc_22_0_RDATA <= hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_RDATA;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARREGION <= x_rsc_22_0_ARREGION;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARQOS <= x_rsc_22_0_ARQOS;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARPROT <= x_rsc_22_0_ARPROT;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARCACHE <= x_rsc_22_0_ARCACHE;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARBURST <= x_rsc_22_0_ARBURST;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARSIZE <= x_rsc_22_0_ARSIZE;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARLEN <= x_rsc_22_0_ARLEN;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_ARADDR <= x_rsc_22_0_ARADDR;
  x_rsc_22_0_BRESP <= hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_BRESP;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_WSTRB <= x_rsc_22_0_WSTRB;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_WDATA <= x_rsc_22_0_WDATA;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWREGION <= x_rsc_22_0_AWREGION;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWQOS <= x_rsc_22_0_AWQOS;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWPROT <= x_rsc_22_0_AWPROT;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWCACHE <= x_rsc_22_0_AWCACHE;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWBURST <= x_rsc_22_0_AWBURST;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWSIZE <= x_rsc_22_0_AWSIZE;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWLEN <= x_rsc_22_0_AWLEN;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_AWADDR <= x_rsc_22_0_AWADDR;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_22_0_i_s_din_mxwt <= hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_din_mxwt;
  hybrid_core_x_rsc_22_0_i_inst_x_rsc_22_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_23_0_i_inst : hybrid_core_x_rsc_23_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_23_0_s_tdone => x_rsc_23_0_s_tdone,
      x_rsc_23_0_tr_write_done => x_rsc_23_0_tr_write_done,
      x_rsc_23_0_RREADY => x_rsc_23_0_RREADY,
      x_rsc_23_0_RVALID => x_rsc_23_0_RVALID,
      x_rsc_23_0_RUSER => x_rsc_23_0_RUSER,
      x_rsc_23_0_RLAST => x_rsc_23_0_RLAST,
      x_rsc_23_0_RRESP => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_RRESP,
      x_rsc_23_0_RDATA => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_RDATA,
      x_rsc_23_0_RID => x_rsc_23_0_RID,
      x_rsc_23_0_ARREADY => x_rsc_23_0_ARREADY,
      x_rsc_23_0_ARVALID => x_rsc_23_0_ARVALID,
      x_rsc_23_0_ARUSER => x_rsc_23_0_ARUSER,
      x_rsc_23_0_ARREGION => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARREGION,
      x_rsc_23_0_ARQOS => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARQOS,
      x_rsc_23_0_ARPROT => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARPROT,
      x_rsc_23_0_ARCACHE => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARCACHE,
      x_rsc_23_0_ARLOCK => x_rsc_23_0_ARLOCK,
      x_rsc_23_0_ARBURST => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARBURST,
      x_rsc_23_0_ARSIZE => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARSIZE,
      x_rsc_23_0_ARLEN => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARLEN,
      x_rsc_23_0_ARADDR => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARADDR,
      x_rsc_23_0_ARID => x_rsc_23_0_ARID,
      x_rsc_23_0_BREADY => x_rsc_23_0_BREADY,
      x_rsc_23_0_BVALID => x_rsc_23_0_BVALID,
      x_rsc_23_0_BUSER => x_rsc_23_0_BUSER,
      x_rsc_23_0_BRESP => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_BRESP,
      x_rsc_23_0_BID => x_rsc_23_0_BID,
      x_rsc_23_0_WREADY => x_rsc_23_0_WREADY,
      x_rsc_23_0_WVALID => x_rsc_23_0_WVALID,
      x_rsc_23_0_WUSER => x_rsc_23_0_WUSER,
      x_rsc_23_0_WLAST => x_rsc_23_0_WLAST,
      x_rsc_23_0_WSTRB => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_WSTRB,
      x_rsc_23_0_WDATA => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_WDATA,
      x_rsc_23_0_AWREADY => x_rsc_23_0_AWREADY,
      x_rsc_23_0_AWVALID => x_rsc_23_0_AWVALID,
      x_rsc_23_0_AWUSER => x_rsc_23_0_AWUSER,
      x_rsc_23_0_AWREGION => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWREGION,
      x_rsc_23_0_AWQOS => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWQOS,
      x_rsc_23_0_AWPROT => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWPROT,
      x_rsc_23_0_AWCACHE => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWCACHE,
      x_rsc_23_0_AWLOCK => x_rsc_23_0_AWLOCK,
      x_rsc_23_0_AWBURST => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWBURST,
      x_rsc_23_0_AWSIZE => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWSIZE,
      x_rsc_23_0_AWLEN => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWLEN,
      x_rsc_23_0_AWADDR => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWADDR,
      x_rsc_23_0_AWID => x_rsc_23_0_AWID,
      core_wen => core_wen,
      x_rsc_23_0_i_oswt => reg_x_rsc_23_0_i_oswt_cse,
      x_rsc_23_0_i_wen_comp => x_rsc_23_0_i_wen_comp,
      x_rsc_23_0_i_oswt_1 => reg_x_rsc_23_0_i_oswt_1_cse,
      x_rsc_23_0_i_wen_comp_1 => x_rsc_23_0_i_wen_comp_1,
      x_rsc_23_0_i_s_raddr_core => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_raddr_core,
      x_rsc_23_0_i_s_waddr_core => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_waddr_core,
      x_rsc_23_0_i_s_din_mxwt => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_din_mxwt,
      x_rsc_23_0_i_s_dout_core => hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_dout_core
    );
  x_rsc_23_0_RRESP <= hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_RRESP;
  x_rsc_23_0_RDATA <= hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_RDATA;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARREGION <= x_rsc_23_0_ARREGION;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARQOS <= x_rsc_23_0_ARQOS;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARPROT <= x_rsc_23_0_ARPROT;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARCACHE <= x_rsc_23_0_ARCACHE;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARBURST <= x_rsc_23_0_ARBURST;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARSIZE <= x_rsc_23_0_ARSIZE;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARLEN <= x_rsc_23_0_ARLEN;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_ARADDR <= x_rsc_23_0_ARADDR;
  x_rsc_23_0_BRESP <= hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_BRESP;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_WSTRB <= x_rsc_23_0_WSTRB;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_WDATA <= x_rsc_23_0_WDATA;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWREGION <= x_rsc_23_0_AWREGION;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWQOS <= x_rsc_23_0_AWQOS;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWPROT <= x_rsc_23_0_AWPROT;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWCACHE <= x_rsc_23_0_AWCACHE;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWBURST <= x_rsc_23_0_AWBURST;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWSIZE <= x_rsc_23_0_AWSIZE;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWLEN <= x_rsc_23_0_AWLEN;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_AWADDR <= x_rsc_23_0_AWADDR;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_23_0_i_s_din_mxwt <= hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_din_mxwt;
  hybrid_core_x_rsc_23_0_i_inst_x_rsc_23_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_24_0_i_inst : hybrid_core_x_rsc_24_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_24_0_s_tdone => x_rsc_24_0_s_tdone,
      x_rsc_24_0_tr_write_done => x_rsc_24_0_tr_write_done,
      x_rsc_24_0_RREADY => x_rsc_24_0_RREADY,
      x_rsc_24_0_RVALID => x_rsc_24_0_RVALID,
      x_rsc_24_0_RUSER => x_rsc_24_0_RUSER,
      x_rsc_24_0_RLAST => x_rsc_24_0_RLAST,
      x_rsc_24_0_RRESP => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_RRESP,
      x_rsc_24_0_RDATA => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_RDATA,
      x_rsc_24_0_RID => x_rsc_24_0_RID,
      x_rsc_24_0_ARREADY => x_rsc_24_0_ARREADY,
      x_rsc_24_0_ARVALID => x_rsc_24_0_ARVALID,
      x_rsc_24_0_ARUSER => x_rsc_24_0_ARUSER,
      x_rsc_24_0_ARREGION => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARREGION,
      x_rsc_24_0_ARQOS => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARQOS,
      x_rsc_24_0_ARPROT => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARPROT,
      x_rsc_24_0_ARCACHE => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARCACHE,
      x_rsc_24_0_ARLOCK => x_rsc_24_0_ARLOCK,
      x_rsc_24_0_ARBURST => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARBURST,
      x_rsc_24_0_ARSIZE => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARSIZE,
      x_rsc_24_0_ARLEN => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARLEN,
      x_rsc_24_0_ARADDR => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARADDR,
      x_rsc_24_0_ARID => x_rsc_24_0_ARID,
      x_rsc_24_0_BREADY => x_rsc_24_0_BREADY,
      x_rsc_24_0_BVALID => x_rsc_24_0_BVALID,
      x_rsc_24_0_BUSER => x_rsc_24_0_BUSER,
      x_rsc_24_0_BRESP => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_BRESP,
      x_rsc_24_0_BID => x_rsc_24_0_BID,
      x_rsc_24_0_WREADY => x_rsc_24_0_WREADY,
      x_rsc_24_0_WVALID => x_rsc_24_0_WVALID,
      x_rsc_24_0_WUSER => x_rsc_24_0_WUSER,
      x_rsc_24_0_WLAST => x_rsc_24_0_WLAST,
      x_rsc_24_0_WSTRB => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_WSTRB,
      x_rsc_24_0_WDATA => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_WDATA,
      x_rsc_24_0_AWREADY => x_rsc_24_0_AWREADY,
      x_rsc_24_0_AWVALID => x_rsc_24_0_AWVALID,
      x_rsc_24_0_AWUSER => x_rsc_24_0_AWUSER,
      x_rsc_24_0_AWREGION => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWREGION,
      x_rsc_24_0_AWQOS => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWQOS,
      x_rsc_24_0_AWPROT => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWPROT,
      x_rsc_24_0_AWCACHE => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWCACHE,
      x_rsc_24_0_AWLOCK => x_rsc_24_0_AWLOCK,
      x_rsc_24_0_AWBURST => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWBURST,
      x_rsc_24_0_AWSIZE => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWSIZE,
      x_rsc_24_0_AWLEN => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWLEN,
      x_rsc_24_0_AWADDR => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWADDR,
      x_rsc_24_0_AWID => x_rsc_24_0_AWID,
      core_wen => core_wen,
      x_rsc_24_0_i_oswt => reg_x_rsc_24_0_i_oswt_cse,
      x_rsc_24_0_i_wen_comp => x_rsc_24_0_i_wen_comp,
      x_rsc_24_0_i_oswt_1 => reg_x_rsc_24_0_i_oswt_1_cse,
      x_rsc_24_0_i_wen_comp_1 => x_rsc_24_0_i_wen_comp_1,
      x_rsc_24_0_i_s_raddr_core => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_raddr_core,
      x_rsc_24_0_i_s_waddr_core => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_waddr_core,
      x_rsc_24_0_i_s_din_mxwt => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_din_mxwt,
      x_rsc_24_0_i_s_dout_core => hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_dout_core
    );
  x_rsc_24_0_RRESP <= hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_RRESP;
  x_rsc_24_0_RDATA <= hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_RDATA;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARREGION <= x_rsc_24_0_ARREGION;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARQOS <= x_rsc_24_0_ARQOS;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARPROT <= x_rsc_24_0_ARPROT;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARCACHE <= x_rsc_24_0_ARCACHE;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARBURST <= x_rsc_24_0_ARBURST;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARSIZE <= x_rsc_24_0_ARSIZE;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARLEN <= x_rsc_24_0_ARLEN;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_ARADDR <= x_rsc_24_0_ARADDR;
  x_rsc_24_0_BRESP <= hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_BRESP;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_WSTRB <= x_rsc_24_0_WSTRB;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_WDATA <= x_rsc_24_0_WDATA;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWREGION <= x_rsc_24_0_AWREGION;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWQOS <= x_rsc_24_0_AWQOS;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWPROT <= x_rsc_24_0_AWPROT;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWCACHE <= x_rsc_24_0_AWCACHE;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWBURST <= x_rsc_24_0_AWBURST;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWSIZE <= x_rsc_24_0_AWSIZE;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWLEN <= x_rsc_24_0_AWLEN;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_AWADDR <= x_rsc_24_0_AWADDR;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_24_0_i_s_din_mxwt <= hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_din_mxwt;
  hybrid_core_x_rsc_24_0_i_inst_x_rsc_24_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_25_0_i_inst : hybrid_core_x_rsc_25_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_25_0_s_tdone => x_rsc_25_0_s_tdone,
      x_rsc_25_0_tr_write_done => x_rsc_25_0_tr_write_done,
      x_rsc_25_0_RREADY => x_rsc_25_0_RREADY,
      x_rsc_25_0_RVALID => x_rsc_25_0_RVALID,
      x_rsc_25_0_RUSER => x_rsc_25_0_RUSER,
      x_rsc_25_0_RLAST => x_rsc_25_0_RLAST,
      x_rsc_25_0_RRESP => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_RRESP,
      x_rsc_25_0_RDATA => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_RDATA,
      x_rsc_25_0_RID => x_rsc_25_0_RID,
      x_rsc_25_0_ARREADY => x_rsc_25_0_ARREADY,
      x_rsc_25_0_ARVALID => x_rsc_25_0_ARVALID,
      x_rsc_25_0_ARUSER => x_rsc_25_0_ARUSER,
      x_rsc_25_0_ARREGION => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARREGION,
      x_rsc_25_0_ARQOS => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARQOS,
      x_rsc_25_0_ARPROT => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARPROT,
      x_rsc_25_0_ARCACHE => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARCACHE,
      x_rsc_25_0_ARLOCK => x_rsc_25_0_ARLOCK,
      x_rsc_25_0_ARBURST => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARBURST,
      x_rsc_25_0_ARSIZE => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARSIZE,
      x_rsc_25_0_ARLEN => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARLEN,
      x_rsc_25_0_ARADDR => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARADDR,
      x_rsc_25_0_ARID => x_rsc_25_0_ARID,
      x_rsc_25_0_BREADY => x_rsc_25_0_BREADY,
      x_rsc_25_0_BVALID => x_rsc_25_0_BVALID,
      x_rsc_25_0_BUSER => x_rsc_25_0_BUSER,
      x_rsc_25_0_BRESP => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_BRESP,
      x_rsc_25_0_BID => x_rsc_25_0_BID,
      x_rsc_25_0_WREADY => x_rsc_25_0_WREADY,
      x_rsc_25_0_WVALID => x_rsc_25_0_WVALID,
      x_rsc_25_0_WUSER => x_rsc_25_0_WUSER,
      x_rsc_25_0_WLAST => x_rsc_25_0_WLAST,
      x_rsc_25_0_WSTRB => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_WSTRB,
      x_rsc_25_0_WDATA => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_WDATA,
      x_rsc_25_0_AWREADY => x_rsc_25_0_AWREADY,
      x_rsc_25_0_AWVALID => x_rsc_25_0_AWVALID,
      x_rsc_25_0_AWUSER => x_rsc_25_0_AWUSER,
      x_rsc_25_0_AWREGION => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWREGION,
      x_rsc_25_0_AWQOS => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWQOS,
      x_rsc_25_0_AWPROT => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWPROT,
      x_rsc_25_0_AWCACHE => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWCACHE,
      x_rsc_25_0_AWLOCK => x_rsc_25_0_AWLOCK,
      x_rsc_25_0_AWBURST => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWBURST,
      x_rsc_25_0_AWSIZE => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWSIZE,
      x_rsc_25_0_AWLEN => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWLEN,
      x_rsc_25_0_AWADDR => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWADDR,
      x_rsc_25_0_AWID => x_rsc_25_0_AWID,
      core_wen => core_wen,
      x_rsc_25_0_i_oswt => reg_x_rsc_25_0_i_oswt_cse,
      x_rsc_25_0_i_wen_comp => x_rsc_25_0_i_wen_comp,
      x_rsc_25_0_i_oswt_1 => reg_x_rsc_25_0_i_oswt_1_cse,
      x_rsc_25_0_i_wen_comp_1 => x_rsc_25_0_i_wen_comp_1,
      x_rsc_25_0_i_s_raddr_core => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_raddr_core,
      x_rsc_25_0_i_s_waddr_core => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_waddr_core,
      x_rsc_25_0_i_s_din_mxwt => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_din_mxwt,
      x_rsc_25_0_i_s_dout_core => hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_dout_core
    );
  x_rsc_25_0_RRESP <= hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_RRESP;
  x_rsc_25_0_RDATA <= hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_RDATA;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARREGION <= x_rsc_25_0_ARREGION;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARQOS <= x_rsc_25_0_ARQOS;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARPROT <= x_rsc_25_0_ARPROT;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARCACHE <= x_rsc_25_0_ARCACHE;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARBURST <= x_rsc_25_0_ARBURST;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARSIZE <= x_rsc_25_0_ARSIZE;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARLEN <= x_rsc_25_0_ARLEN;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_ARADDR <= x_rsc_25_0_ARADDR;
  x_rsc_25_0_BRESP <= hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_BRESP;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_WSTRB <= x_rsc_25_0_WSTRB;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_WDATA <= x_rsc_25_0_WDATA;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWREGION <= x_rsc_25_0_AWREGION;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWQOS <= x_rsc_25_0_AWQOS;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWPROT <= x_rsc_25_0_AWPROT;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWCACHE <= x_rsc_25_0_AWCACHE;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWBURST <= x_rsc_25_0_AWBURST;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWSIZE <= x_rsc_25_0_AWSIZE;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWLEN <= x_rsc_25_0_AWLEN;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_AWADDR <= x_rsc_25_0_AWADDR;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_25_0_i_s_din_mxwt <= hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_din_mxwt;
  hybrid_core_x_rsc_25_0_i_inst_x_rsc_25_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_26_0_i_inst : hybrid_core_x_rsc_26_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_26_0_s_tdone => x_rsc_26_0_s_tdone,
      x_rsc_26_0_tr_write_done => x_rsc_26_0_tr_write_done,
      x_rsc_26_0_RREADY => x_rsc_26_0_RREADY,
      x_rsc_26_0_RVALID => x_rsc_26_0_RVALID,
      x_rsc_26_0_RUSER => x_rsc_26_0_RUSER,
      x_rsc_26_0_RLAST => x_rsc_26_0_RLAST,
      x_rsc_26_0_RRESP => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_RRESP,
      x_rsc_26_0_RDATA => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_RDATA,
      x_rsc_26_0_RID => x_rsc_26_0_RID,
      x_rsc_26_0_ARREADY => x_rsc_26_0_ARREADY,
      x_rsc_26_0_ARVALID => x_rsc_26_0_ARVALID,
      x_rsc_26_0_ARUSER => x_rsc_26_0_ARUSER,
      x_rsc_26_0_ARREGION => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARREGION,
      x_rsc_26_0_ARQOS => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARQOS,
      x_rsc_26_0_ARPROT => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARPROT,
      x_rsc_26_0_ARCACHE => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARCACHE,
      x_rsc_26_0_ARLOCK => x_rsc_26_0_ARLOCK,
      x_rsc_26_0_ARBURST => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARBURST,
      x_rsc_26_0_ARSIZE => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARSIZE,
      x_rsc_26_0_ARLEN => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARLEN,
      x_rsc_26_0_ARADDR => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARADDR,
      x_rsc_26_0_ARID => x_rsc_26_0_ARID,
      x_rsc_26_0_BREADY => x_rsc_26_0_BREADY,
      x_rsc_26_0_BVALID => x_rsc_26_0_BVALID,
      x_rsc_26_0_BUSER => x_rsc_26_0_BUSER,
      x_rsc_26_0_BRESP => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_BRESP,
      x_rsc_26_0_BID => x_rsc_26_0_BID,
      x_rsc_26_0_WREADY => x_rsc_26_0_WREADY,
      x_rsc_26_0_WVALID => x_rsc_26_0_WVALID,
      x_rsc_26_0_WUSER => x_rsc_26_0_WUSER,
      x_rsc_26_0_WLAST => x_rsc_26_0_WLAST,
      x_rsc_26_0_WSTRB => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_WSTRB,
      x_rsc_26_0_WDATA => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_WDATA,
      x_rsc_26_0_AWREADY => x_rsc_26_0_AWREADY,
      x_rsc_26_0_AWVALID => x_rsc_26_0_AWVALID,
      x_rsc_26_0_AWUSER => x_rsc_26_0_AWUSER,
      x_rsc_26_0_AWREGION => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWREGION,
      x_rsc_26_0_AWQOS => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWQOS,
      x_rsc_26_0_AWPROT => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWPROT,
      x_rsc_26_0_AWCACHE => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWCACHE,
      x_rsc_26_0_AWLOCK => x_rsc_26_0_AWLOCK,
      x_rsc_26_0_AWBURST => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWBURST,
      x_rsc_26_0_AWSIZE => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWSIZE,
      x_rsc_26_0_AWLEN => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWLEN,
      x_rsc_26_0_AWADDR => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWADDR,
      x_rsc_26_0_AWID => x_rsc_26_0_AWID,
      core_wen => core_wen,
      x_rsc_26_0_i_oswt => reg_x_rsc_26_0_i_oswt_cse,
      x_rsc_26_0_i_wen_comp => x_rsc_26_0_i_wen_comp,
      x_rsc_26_0_i_oswt_1 => reg_x_rsc_26_0_i_oswt_1_cse,
      x_rsc_26_0_i_wen_comp_1 => x_rsc_26_0_i_wen_comp_1,
      x_rsc_26_0_i_s_raddr_core => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_raddr_core,
      x_rsc_26_0_i_s_waddr_core => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_waddr_core,
      x_rsc_26_0_i_s_din_mxwt => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_din_mxwt,
      x_rsc_26_0_i_s_dout_core => hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_dout_core
    );
  x_rsc_26_0_RRESP <= hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_RRESP;
  x_rsc_26_0_RDATA <= hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_RDATA;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARREGION <= x_rsc_26_0_ARREGION;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARQOS <= x_rsc_26_0_ARQOS;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARPROT <= x_rsc_26_0_ARPROT;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARCACHE <= x_rsc_26_0_ARCACHE;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARBURST <= x_rsc_26_0_ARBURST;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARSIZE <= x_rsc_26_0_ARSIZE;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARLEN <= x_rsc_26_0_ARLEN;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_ARADDR <= x_rsc_26_0_ARADDR;
  x_rsc_26_0_BRESP <= hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_BRESP;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_WSTRB <= x_rsc_26_0_WSTRB;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_WDATA <= x_rsc_26_0_WDATA;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWREGION <= x_rsc_26_0_AWREGION;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWQOS <= x_rsc_26_0_AWQOS;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWPROT <= x_rsc_26_0_AWPROT;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWCACHE <= x_rsc_26_0_AWCACHE;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWBURST <= x_rsc_26_0_AWBURST;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWSIZE <= x_rsc_26_0_AWSIZE;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWLEN <= x_rsc_26_0_AWLEN;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_AWADDR <= x_rsc_26_0_AWADDR;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_26_0_i_s_din_mxwt <= hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_din_mxwt;
  hybrid_core_x_rsc_26_0_i_inst_x_rsc_26_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_27_0_i_inst : hybrid_core_x_rsc_27_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_27_0_s_tdone => x_rsc_27_0_s_tdone,
      x_rsc_27_0_tr_write_done => x_rsc_27_0_tr_write_done,
      x_rsc_27_0_RREADY => x_rsc_27_0_RREADY,
      x_rsc_27_0_RVALID => x_rsc_27_0_RVALID,
      x_rsc_27_0_RUSER => x_rsc_27_0_RUSER,
      x_rsc_27_0_RLAST => x_rsc_27_0_RLAST,
      x_rsc_27_0_RRESP => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_RRESP,
      x_rsc_27_0_RDATA => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_RDATA,
      x_rsc_27_0_RID => x_rsc_27_0_RID,
      x_rsc_27_0_ARREADY => x_rsc_27_0_ARREADY,
      x_rsc_27_0_ARVALID => x_rsc_27_0_ARVALID,
      x_rsc_27_0_ARUSER => x_rsc_27_0_ARUSER,
      x_rsc_27_0_ARREGION => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARREGION,
      x_rsc_27_0_ARQOS => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARQOS,
      x_rsc_27_0_ARPROT => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARPROT,
      x_rsc_27_0_ARCACHE => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARCACHE,
      x_rsc_27_0_ARLOCK => x_rsc_27_0_ARLOCK,
      x_rsc_27_0_ARBURST => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARBURST,
      x_rsc_27_0_ARSIZE => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARSIZE,
      x_rsc_27_0_ARLEN => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARLEN,
      x_rsc_27_0_ARADDR => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARADDR,
      x_rsc_27_0_ARID => x_rsc_27_0_ARID,
      x_rsc_27_0_BREADY => x_rsc_27_0_BREADY,
      x_rsc_27_0_BVALID => x_rsc_27_0_BVALID,
      x_rsc_27_0_BUSER => x_rsc_27_0_BUSER,
      x_rsc_27_0_BRESP => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_BRESP,
      x_rsc_27_0_BID => x_rsc_27_0_BID,
      x_rsc_27_0_WREADY => x_rsc_27_0_WREADY,
      x_rsc_27_0_WVALID => x_rsc_27_0_WVALID,
      x_rsc_27_0_WUSER => x_rsc_27_0_WUSER,
      x_rsc_27_0_WLAST => x_rsc_27_0_WLAST,
      x_rsc_27_0_WSTRB => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_WSTRB,
      x_rsc_27_0_WDATA => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_WDATA,
      x_rsc_27_0_AWREADY => x_rsc_27_0_AWREADY,
      x_rsc_27_0_AWVALID => x_rsc_27_0_AWVALID,
      x_rsc_27_0_AWUSER => x_rsc_27_0_AWUSER,
      x_rsc_27_0_AWREGION => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWREGION,
      x_rsc_27_0_AWQOS => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWQOS,
      x_rsc_27_0_AWPROT => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWPROT,
      x_rsc_27_0_AWCACHE => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWCACHE,
      x_rsc_27_0_AWLOCK => x_rsc_27_0_AWLOCK,
      x_rsc_27_0_AWBURST => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWBURST,
      x_rsc_27_0_AWSIZE => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWSIZE,
      x_rsc_27_0_AWLEN => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWLEN,
      x_rsc_27_0_AWADDR => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWADDR,
      x_rsc_27_0_AWID => x_rsc_27_0_AWID,
      core_wen => core_wen,
      x_rsc_27_0_i_oswt => reg_x_rsc_27_0_i_oswt_cse,
      x_rsc_27_0_i_wen_comp => x_rsc_27_0_i_wen_comp,
      x_rsc_27_0_i_oswt_1 => reg_x_rsc_27_0_i_oswt_1_cse,
      x_rsc_27_0_i_wen_comp_1 => x_rsc_27_0_i_wen_comp_1,
      x_rsc_27_0_i_s_raddr_core => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_raddr_core,
      x_rsc_27_0_i_s_waddr_core => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_waddr_core,
      x_rsc_27_0_i_s_din_mxwt => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_din_mxwt,
      x_rsc_27_0_i_s_dout_core => hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_dout_core
    );
  x_rsc_27_0_RRESP <= hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_RRESP;
  x_rsc_27_0_RDATA <= hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_RDATA;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARREGION <= x_rsc_27_0_ARREGION;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARQOS <= x_rsc_27_0_ARQOS;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARPROT <= x_rsc_27_0_ARPROT;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARCACHE <= x_rsc_27_0_ARCACHE;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARBURST <= x_rsc_27_0_ARBURST;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARSIZE <= x_rsc_27_0_ARSIZE;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARLEN <= x_rsc_27_0_ARLEN;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_ARADDR <= x_rsc_27_0_ARADDR;
  x_rsc_27_0_BRESP <= hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_BRESP;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_WSTRB <= x_rsc_27_0_WSTRB;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_WDATA <= x_rsc_27_0_WDATA;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWREGION <= x_rsc_27_0_AWREGION;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWQOS <= x_rsc_27_0_AWQOS;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWPROT <= x_rsc_27_0_AWPROT;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWCACHE <= x_rsc_27_0_AWCACHE;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWBURST <= x_rsc_27_0_AWBURST;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWSIZE <= x_rsc_27_0_AWSIZE;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWLEN <= x_rsc_27_0_AWLEN;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_AWADDR <= x_rsc_27_0_AWADDR;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_27_0_i_s_din_mxwt <= hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_din_mxwt;
  hybrid_core_x_rsc_27_0_i_inst_x_rsc_27_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_28_0_i_inst : hybrid_core_x_rsc_28_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_28_0_s_tdone => x_rsc_28_0_s_tdone,
      x_rsc_28_0_tr_write_done => x_rsc_28_0_tr_write_done,
      x_rsc_28_0_RREADY => x_rsc_28_0_RREADY,
      x_rsc_28_0_RVALID => x_rsc_28_0_RVALID,
      x_rsc_28_0_RUSER => x_rsc_28_0_RUSER,
      x_rsc_28_0_RLAST => x_rsc_28_0_RLAST,
      x_rsc_28_0_RRESP => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_RRESP,
      x_rsc_28_0_RDATA => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_RDATA,
      x_rsc_28_0_RID => x_rsc_28_0_RID,
      x_rsc_28_0_ARREADY => x_rsc_28_0_ARREADY,
      x_rsc_28_0_ARVALID => x_rsc_28_0_ARVALID,
      x_rsc_28_0_ARUSER => x_rsc_28_0_ARUSER,
      x_rsc_28_0_ARREGION => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARREGION,
      x_rsc_28_0_ARQOS => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARQOS,
      x_rsc_28_0_ARPROT => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARPROT,
      x_rsc_28_0_ARCACHE => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARCACHE,
      x_rsc_28_0_ARLOCK => x_rsc_28_0_ARLOCK,
      x_rsc_28_0_ARBURST => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARBURST,
      x_rsc_28_0_ARSIZE => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARSIZE,
      x_rsc_28_0_ARLEN => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARLEN,
      x_rsc_28_0_ARADDR => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARADDR,
      x_rsc_28_0_ARID => x_rsc_28_0_ARID,
      x_rsc_28_0_BREADY => x_rsc_28_0_BREADY,
      x_rsc_28_0_BVALID => x_rsc_28_0_BVALID,
      x_rsc_28_0_BUSER => x_rsc_28_0_BUSER,
      x_rsc_28_0_BRESP => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_BRESP,
      x_rsc_28_0_BID => x_rsc_28_0_BID,
      x_rsc_28_0_WREADY => x_rsc_28_0_WREADY,
      x_rsc_28_0_WVALID => x_rsc_28_0_WVALID,
      x_rsc_28_0_WUSER => x_rsc_28_0_WUSER,
      x_rsc_28_0_WLAST => x_rsc_28_0_WLAST,
      x_rsc_28_0_WSTRB => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_WSTRB,
      x_rsc_28_0_WDATA => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_WDATA,
      x_rsc_28_0_AWREADY => x_rsc_28_0_AWREADY,
      x_rsc_28_0_AWVALID => x_rsc_28_0_AWVALID,
      x_rsc_28_0_AWUSER => x_rsc_28_0_AWUSER,
      x_rsc_28_0_AWREGION => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWREGION,
      x_rsc_28_0_AWQOS => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWQOS,
      x_rsc_28_0_AWPROT => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWPROT,
      x_rsc_28_0_AWCACHE => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWCACHE,
      x_rsc_28_0_AWLOCK => x_rsc_28_0_AWLOCK,
      x_rsc_28_0_AWBURST => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWBURST,
      x_rsc_28_0_AWSIZE => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWSIZE,
      x_rsc_28_0_AWLEN => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWLEN,
      x_rsc_28_0_AWADDR => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWADDR,
      x_rsc_28_0_AWID => x_rsc_28_0_AWID,
      core_wen => core_wen,
      x_rsc_28_0_i_oswt => reg_x_rsc_28_0_i_oswt_cse,
      x_rsc_28_0_i_wen_comp => x_rsc_28_0_i_wen_comp,
      x_rsc_28_0_i_oswt_1 => reg_x_rsc_28_0_i_oswt_1_cse,
      x_rsc_28_0_i_wen_comp_1 => x_rsc_28_0_i_wen_comp_1,
      x_rsc_28_0_i_s_raddr_core => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_raddr_core,
      x_rsc_28_0_i_s_waddr_core => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_waddr_core,
      x_rsc_28_0_i_s_din_mxwt => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_din_mxwt,
      x_rsc_28_0_i_s_dout_core => hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_dout_core
    );
  x_rsc_28_0_RRESP <= hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_RRESP;
  x_rsc_28_0_RDATA <= hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_RDATA;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARREGION <= x_rsc_28_0_ARREGION;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARQOS <= x_rsc_28_0_ARQOS;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARPROT <= x_rsc_28_0_ARPROT;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARCACHE <= x_rsc_28_0_ARCACHE;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARBURST <= x_rsc_28_0_ARBURST;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARSIZE <= x_rsc_28_0_ARSIZE;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARLEN <= x_rsc_28_0_ARLEN;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_ARADDR <= x_rsc_28_0_ARADDR;
  x_rsc_28_0_BRESP <= hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_BRESP;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_WSTRB <= x_rsc_28_0_WSTRB;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_WDATA <= x_rsc_28_0_WDATA;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWREGION <= x_rsc_28_0_AWREGION;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWQOS <= x_rsc_28_0_AWQOS;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWPROT <= x_rsc_28_0_AWPROT;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWCACHE <= x_rsc_28_0_AWCACHE;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWBURST <= x_rsc_28_0_AWBURST;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWSIZE <= x_rsc_28_0_AWSIZE;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWLEN <= x_rsc_28_0_AWLEN;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_AWADDR <= x_rsc_28_0_AWADDR;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_28_0_i_s_din_mxwt <= hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_din_mxwt;
  hybrid_core_x_rsc_28_0_i_inst_x_rsc_28_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_29_0_i_inst : hybrid_core_x_rsc_29_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_29_0_s_tdone => x_rsc_29_0_s_tdone,
      x_rsc_29_0_tr_write_done => x_rsc_29_0_tr_write_done,
      x_rsc_29_0_RREADY => x_rsc_29_0_RREADY,
      x_rsc_29_0_RVALID => x_rsc_29_0_RVALID,
      x_rsc_29_0_RUSER => x_rsc_29_0_RUSER,
      x_rsc_29_0_RLAST => x_rsc_29_0_RLAST,
      x_rsc_29_0_RRESP => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_RRESP,
      x_rsc_29_0_RDATA => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_RDATA,
      x_rsc_29_0_RID => x_rsc_29_0_RID,
      x_rsc_29_0_ARREADY => x_rsc_29_0_ARREADY,
      x_rsc_29_0_ARVALID => x_rsc_29_0_ARVALID,
      x_rsc_29_0_ARUSER => x_rsc_29_0_ARUSER,
      x_rsc_29_0_ARREGION => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARREGION,
      x_rsc_29_0_ARQOS => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARQOS,
      x_rsc_29_0_ARPROT => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARPROT,
      x_rsc_29_0_ARCACHE => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARCACHE,
      x_rsc_29_0_ARLOCK => x_rsc_29_0_ARLOCK,
      x_rsc_29_0_ARBURST => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARBURST,
      x_rsc_29_0_ARSIZE => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARSIZE,
      x_rsc_29_0_ARLEN => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARLEN,
      x_rsc_29_0_ARADDR => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARADDR,
      x_rsc_29_0_ARID => x_rsc_29_0_ARID,
      x_rsc_29_0_BREADY => x_rsc_29_0_BREADY,
      x_rsc_29_0_BVALID => x_rsc_29_0_BVALID,
      x_rsc_29_0_BUSER => x_rsc_29_0_BUSER,
      x_rsc_29_0_BRESP => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_BRESP,
      x_rsc_29_0_BID => x_rsc_29_0_BID,
      x_rsc_29_0_WREADY => x_rsc_29_0_WREADY,
      x_rsc_29_0_WVALID => x_rsc_29_0_WVALID,
      x_rsc_29_0_WUSER => x_rsc_29_0_WUSER,
      x_rsc_29_0_WLAST => x_rsc_29_0_WLAST,
      x_rsc_29_0_WSTRB => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_WSTRB,
      x_rsc_29_0_WDATA => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_WDATA,
      x_rsc_29_0_AWREADY => x_rsc_29_0_AWREADY,
      x_rsc_29_0_AWVALID => x_rsc_29_0_AWVALID,
      x_rsc_29_0_AWUSER => x_rsc_29_0_AWUSER,
      x_rsc_29_0_AWREGION => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWREGION,
      x_rsc_29_0_AWQOS => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWQOS,
      x_rsc_29_0_AWPROT => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWPROT,
      x_rsc_29_0_AWCACHE => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWCACHE,
      x_rsc_29_0_AWLOCK => x_rsc_29_0_AWLOCK,
      x_rsc_29_0_AWBURST => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWBURST,
      x_rsc_29_0_AWSIZE => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWSIZE,
      x_rsc_29_0_AWLEN => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWLEN,
      x_rsc_29_0_AWADDR => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWADDR,
      x_rsc_29_0_AWID => x_rsc_29_0_AWID,
      core_wen => core_wen,
      x_rsc_29_0_i_oswt => reg_x_rsc_29_0_i_oswt_cse,
      x_rsc_29_0_i_wen_comp => x_rsc_29_0_i_wen_comp,
      x_rsc_29_0_i_oswt_1 => reg_x_rsc_29_0_i_oswt_1_cse,
      x_rsc_29_0_i_wen_comp_1 => x_rsc_29_0_i_wen_comp_1,
      x_rsc_29_0_i_s_raddr_core => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_raddr_core,
      x_rsc_29_0_i_s_waddr_core => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_waddr_core,
      x_rsc_29_0_i_s_din_mxwt => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_din_mxwt,
      x_rsc_29_0_i_s_dout_core => hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_dout_core
    );
  x_rsc_29_0_RRESP <= hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_RRESP;
  x_rsc_29_0_RDATA <= hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_RDATA;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARREGION <= x_rsc_29_0_ARREGION;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARQOS <= x_rsc_29_0_ARQOS;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARPROT <= x_rsc_29_0_ARPROT;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARCACHE <= x_rsc_29_0_ARCACHE;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARBURST <= x_rsc_29_0_ARBURST;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARSIZE <= x_rsc_29_0_ARSIZE;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARLEN <= x_rsc_29_0_ARLEN;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_ARADDR <= x_rsc_29_0_ARADDR;
  x_rsc_29_0_BRESP <= hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_BRESP;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_WSTRB <= x_rsc_29_0_WSTRB;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_WDATA <= x_rsc_29_0_WDATA;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWREGION <= x_rsc_29_0_AWREGION;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWQOS <= x_rsc_29_0_AWQOS;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWPROT <= x_rsc_29_0_AWPROT;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWCACHE <= x_rsc_29_0_AWCACHE;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWBURST <= x_rsc_29_0_AWBURST;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWSIZE <= x_rsc_29_0_AWSIZE;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWLEN <= x_rsc_29_0_AWLEN;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_AWADDR <= x_rsc_29_0_AWADDR;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_29_0_i_s_din_mxwt <= hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_din_mxwt;
  hybrid_core_x_rsc_29_0_i_inst_x_rsc_29_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_30_0_i_inst : hybrid_core_x_rsc_30_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_30_0_s_tdone => x_rsc_30_0_s_tdone,
      x_rsc_30_0_tr_write_done => x_rsc_30_0_tr_write_done,
      x_rsc_30_0_RREADY => x_rsc_30_0_RREADY,
      x_rsc_30_0_RVALID => x_rsc_30_0_RVALID,
      x_rsc_30_0_RUSER => x_rsc_30_0_RUSER,
      x_rsc_30_0_RLAST => x_rsc_30_0_RLAST,
      x_rsc_30_0_RRESP => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_RRESP,
      x_rsc_30_0_RDATA => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_RDATA,
      x_rsc_30_0_RID => x_rsc_30_0_RID,
      x_rsc_30_0_ARREADY => x_rsc_30_0_ARREADY,
      x_rsc_30_0_ARVALID => x_rsc_30_0_ARVALID,
      x_rsc_30_0_ARUSER => x_rsc_30_0_ARUSER,
      x_rsc_30_0_ARREGION => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARREGION,
      x_rsc_30_0_ARQOS => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARQOS,
      x_rsc_30_0_ARPROT => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARPROT,
      x_rsc_30_0_ARCACHE => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARCACHE,
      x_rsc_30_0_ARLOCK => x_rsc_30_0_ARLOCK,
      x_rsc_30_0_ARBURST => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARBURST,
      x_rsc_30_0_ARSIZE => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARSIZE,
      x_rsc_30_0_ARLEN => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARLEN,
      x_rsc_30_0_ARADDR => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARADDR,
      x_rsc_30_0_ARID => x_rsc_30_0_ARID,
      x_rsc_30_0_BREADY => x_rsc_30_0_BREADY,
      x_rsc_30_0_BVALID => x_rsc_30_0_BVALID,
      x_rsc_30_0_BUSER => x_rsc_30_0_BUSER,
      x_rsc_30_0_BRESP => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_BRESP,
      x_rsc_30_0_BID => x_rsc_30_0_BID,
      x_rsc_30_0_WREADY => x_rsc_30_0_WREADY,
      x_rsc_30_0_WVALID => x_rsc_30_0_WVALID,
      x_rsc_30_0_WUSER => x_rsc_30_0_WUSER,
      x_rsc_30_0_WLAST => x_rsc_30_0_WLAST,
      x_rsc_30_0_WSTRB => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_WSTRB,
      x_rsc_30_0_WDATA => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_WDATA,
      x_rsc_30_0_AWREADY => x_rsc_30_0_AWREADY,
      x_rsc_30_0_AWVALID => x_rsc_30_0_AWVALID,
      x_rsc_30_0_AWUSER => x_rsc_30_0_AWUSER,
      x_rsc_30_0_AWREGION => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWREGION,
      x_rsc_30_0_AWQOS => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWQOS,
      x_rsc_30_0_AWPROT => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWPROT,
      x_rsc_30_0_AWCACHE => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWCACHE,
      x_rsc_30_0_AWLOCK => x_rsc_30_0_AWLOCK,
      x_rsc_30_0_AWBURST => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWBURST,
      x_rsc_30_0_AWSIZE => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWSIZE,
      x_rsc_30_0_AWLEN => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWLEN,
      x_rsc_30_0_AWADDR => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWADDR,
      x_rsc_30_0_AWID => x_rsc_30_0_AWID,
      core_wen => core_wen,
      x_rsc_30_0_i_oswt => reg_x_rsc_30_0_i_oswt_cse,
      x_rsc_30_0_i_wen_comp => x_rsc_30_0_i_wen_comp,
      x_rsc_30_0_i_oswt_1 => reg_x_rsc_30_0_i_oswt_1_cse,
      x_rsc_30_0_i_wen_comp_1 => x_rsc_30_0_i_wen_comp_1,
      x_rsc_30_0_i_s_raddr_core => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_raddr_core,
      x_rsc_30_0_i_s_waddr_core => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_waddr_core,
      x_rsc_30_0_i_s_din_mxwt => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_din_mxwt,
      x_rsc_30_0_i_s_dout_core => hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_dout_core
    );
  x_rsc_30_0_RRESP <= hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_RRESP;
  x_rsc_30_0_RDATA <= hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_RDATA;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARREGION <= x_rsc_30_0_ARREGION;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARQOS <= x_rsc_30_0_ARQOS;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARPROT <= x_rsc_30_0_ARPROT;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARCACHE <= x_rsc_30_0_ARCACHE;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARBURST <= x_rsc_30_0_ARBURST;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARSIZE <= x_rsc_30_0_ARSIZE;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARLEN <= x_rsc_30_0_ARLEN;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_ARADDR <= x_rsc_30_0_ARADDR;
  x_rsc_30_0_BRESP <= hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_BRESP;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_WSTRB <= x_rsc_30_0_WSTRB;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_WDATA <= x_rsc_30_0_WDATA;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWREGION <= x_rsc_30_0_AWREGION;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWQOS <= x_rsc_30_0_AWQOS;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWPROT <= x_rsc_30_0_AWPROT;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWCACHE <= x_rsc_30_0_AWCACHE;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWBURST <= x_rsc_30_0_AWBURST;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWSIZE <= x_rsc_30_0_AWSIZE;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWLEN <= x_rsc_30_0_AWLEN;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_AWADDR <= x_rsc_30_0_AWADDR;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_30_0_i_s_din_mxwt <= hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_din_mxwt;
  hybrid_core_x_rsc_30_0_i_inst_x_rsc_30_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_31_0_i_inst : hybrid_core_x_rsc_31_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_31_0_s_tdone => x_rsc_31_0_s_tdone,
      x_rsc_31_0_tr_write_done => x_rsc_31_0_tr_write_done,
      x_rsc_31_0_RREADY => x_rsc_31_0_RREADY,
      x_rsc_31_0_RVALID => x_rsc_31_0_RVALID,
      x_rsc_31_0_RUSER => x_rsc_31_0_RUSER,
      x_rsc_31_0_RLAST => x_rsc_31_0_RLAST,
      x_rsc_31_0_RRESP => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_RRESP,
      x_rsc_31_0_RDATA => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_RDATA,
      x_rsc_31_0_RID => x_rsc_31_0_RID,
      x_rsc_31_0_ARREADY => x_rsc_31_0_ARREADY,
      x_rsc_31_0_ARVALID => x_rsc_31_0_ARVALID,
      x_rsc_31_0_ARUSER => x_rsc_31_0_ARUSER,
      x_rsc_31_0_ARREGION => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARREGION,
      x_rsc_31_0_ARQOS => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARQOS,
      x_rsc_31_0_ARPROT => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARPROT,
      x_rsc_31_0_ARCACHE => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARCACHE,
      x_rsc_31_0_ARLOCK => x_rsc_31_0_ARLOCK,
      x_rsc_31_0_ARBURST => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARBURST,
      x_rsc_31_0_ARSIZE => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARSIZE,
      x_rsc_31_0_ARLEN => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARLEN,
      x_rsc_31_0_ARADDR => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARADDR,
      x_rsc_31_0_ARID => x_rsc_31_0_ARID,
      x_rsc_31_0_BREADY => x_rsc_31_0_BREADY,
      x_rsc_31_0_BVALID => x_rsc_31_0_BVALID,
      x_rsc_31_0_BUSER => x_rsc_31_0_BUSER,
      x_rsc_31_0_BRESP => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_BRESP,
      x_rsc_31_0_BID => x_rsc_31_0_BID,
      x_rsc_31_0_WREADY => x_rsc_31_0_WREADY,
      x_rsc_31_0_WVALID => x_rsc_31_0_WVALID,
      x_rsc_31_0_WUSER => x_rsc_31_0_WUSER,
      x_rsc_31_0_WLAST => x_rsc_31_0_WLAST,
      x_rsc_31_0_WSTRB => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_WSTRB,
      x_rsc_31_0_WDATA => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_WDATA,
      x_rsc_31_0_AWREADY => x_rsc_31_0_AWREADY,
      x_rsc_31_0_AWVALID => x_rsc_31_0_AWVALID,
      x_rsc_31_0_AWUSER => x_rsc_31_0_AWUSER,
      x_rsc_31_0_AWREGION => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWREGION,
      x_rsc_31_0_AWQOS => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWQOS,
      x_rsc_31_0_AWPROT => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWPROT,
      x_rsc_31_0_AWCACHE => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWCACHE,
      x_rsc_31_0_AWLOCK => x_rsc_31_0_AWLOCK,
      x_rsc_31_0_AWBURST => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWBURST,
      x_rsc_31_0_AWSIZE => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWSIZE,
      x_rsc_31_0_AWLEN => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWLEN,
      x_rsc_31_0_AWADDR => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWADDR,
      x_rsc_31_0_AWID => x_rsc_31_0_AWID,
      core_wen => core_wen,
      x_rsc_31_0_i_oswt => reg_x_rsc_31_0_i_oswt_cse,
      x_rsc_31_0_i_wen_comp => x_rsc_31_0_i_wen_comp,
      x_rsc_31_0_i_oswt_1 => reg_x_rsc_31_0_i_oswt_1_cse,
      x_rsc_31_0_i_wen_comp_1 => x_rsc_31_0_i_wen_comp_1,
      x_rsc_31_0_i_s_raddr_core => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_raddr_core,
      x_rsc_31_0_i_s_waddr_core => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_waddr_core,
      x_rsc_31_0_i_s_din_mxwt => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_din_mxwt,
      x_rsc_31_0_i_s_dout_core => hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_dout_core
    );
  x_rsc_31_0_RRESP <= hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_RRESP;
  x_rsc_31_0_RDATA <= hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_RDATA;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARREGION <= x_rsc_31_0_ARREGION;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARQOS <= x_rsc_31_0_ARQOS;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARPROT <= x_rsc_31_0_ARPROT;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARCACHE <= x_rsc_31_0_ARCACHE;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARBURST <= x_rsc_31_0_ARBURST;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARSIZE <= x_rsc_31_0_ARSIZE;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARLEN <= x_rsc_31_0_ARLEN;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_ARADDR <= x_rsc_31_0_ARADDR;
  x_rsc_31_0_BRESP <= hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_BRESP;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_WSTRB <= x_rsc_31_0_WSTRB;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_WDATA <= x_rsc_31_0_WDATA;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWREGION <= x_rsc_31_0_AWREGION;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWQOS <= x_rsc_31_0_AWQOS;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWPROT <= x_rsc_31_0_AWPROT;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWCACHE <= x_rsc_31_0_AWCACHE;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWBURST <= x_rsc_31_0_AWBURST;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWSIZE <= x_rsc_31_0_AWSIZE;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWLEN <= x_rsc_31_0_AWLEN;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_AWADDR <= x_rsc_31_0_AWADDR;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_raddr_core <= reg_x_rsc_0_0_i_s_raddr_core_cse;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_waddr_core <= reg_x_rsc_0_0_i_s_waddr_core_cse;
  x_rsc_31_0_i_s_din_mxwt <= hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_din_mxwt;
  hybrid_core_x_rsc_31_0_i_inst_x_rsc_31_0_i_s_dout_core <= reg_x_rsc_0_0_i_s_dout_core_cse;

  hybrid_core_x_rsc_triosy_31_0_obj_inst : hybrid_core_x_rsc_triosy_31_0_obj
    PORT MAP(
      x_rsc_triosy_31_0_lz => x_rsc_triosy_31_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_31_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_30_0_obj_inst : hybrid_core_x_rsc_triosy_30_0_obj
    PORT MAP(
      x_rsc_triosy_30_0_lz => x_rsc_triosy_30_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_30_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_29_0_obj_inst : hybrid_core_x_rsc_triosy_29_0_obj
    PORT MAP(
      x_rsc_triosy_29_0_lz => x_rsc_triosy_29_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_29_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_28_0_obj_inst : hybrid_core_x_rsc_triosy_28_0_obj
    PORT MAP(
      x_rsc_triosy_28_0_lz => x_rsc_triosy_28_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_28_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_27_0_obj_inst : hybrid_core_x_rsc_triosy_27_0_obj
    PORT MAP(
      x_rsc_triosy_27_0_lz => x_rsc_triosy_27_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_27_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_26_0_obj_inst : hybrid_core_x_rsc_triosy_26_0_obj
    PORT MAP(
      x_rsc_triosy_26_0_lz => x_rsc_triosy_26_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_26_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_25_0_obj_inst : hybrid_core_x_rsc_triosy_25_0_obj
    PORT MAP(
      x_rsc_triosy_25_0_lz => x_rsc_triosy_25_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_25_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_24_0_obj_inst : hybrid_core_x_rsc_triosy_24_0_obj
    PORT MAP(
      x_rsc_triosy_24_0_lz => x_rsc_triosy_24_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_24_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_23_0_obj_inst : hybrid_core_x_rsc_triosy_23_0_obj
    PORT MAP(
      x_rsc_triosy_23_0_lz => x_rsc_triosy_23_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_23_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_22_0_obj_inst : hybrid_core_x_rsc_triosy_22_0_obj
    PORT MAP(
      x_rsc_triosy_22_0_lz => x_rsc_triosy_22_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_22_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_21_0_obj_inst : hybrid_core_x_rsc_triosy_21_0_obj
    PORT MAP(
      x_rsc_triosy_21_0_lz => x_rsc_triosy_21_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_21_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_20_0_obj_inst : hybrid_core_x_rsc_triosy_20_0_obj
    PORT MAP(
      x_rsc_triosy_20_0_lz => x_rsc_triosy_20_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_20_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_19_0_obj_inst : hybrid_core_x_rsc_triosy_19_0_obj
    PORT MAP(
      x_rsc_triosy_19_0_lz => x_rsc_triosy_19_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_19_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_18_0_obj_inst : hybrid_core_x_rsc_triosy_18_0_obj
    PORT MAP(
      x_rsc_triosy_18_0_lz => x_rsc_triosy_18_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_18_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_17_0_obj_inst : hybrid_core_x_rsc_triosy_17_0_obj
    PORT MAP(
      x_rsc_triosy_17_0_lz => x_rsc_triosy_17_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_17_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_16_0_obj_inst : hybrid_core_x_rsc_triosy_16_0_obj
    PORT MAP(
      x_rsc_triosy_16_0_lz => x_rsc_triosy_16_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_16_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_15_0_obj_inst : hybrid_core_x_rsc_triosy_15_0_obj
    PORT MAP(
      x_rsc_triosy_15_0_lz => x_rsc_triosy_15_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_15_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_14_0_obj_inst : hybrid_core_x_rsc_triosy_14_0_obj
    PORT MAP(
      x_rsc_triosy_14_0_lz => x_rsc_triosy_14_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_14_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_13_0_obj_inst : hybrid_core_x_rsc_triosy_13_0_obj
    PORT MAP(
      x_rsc_triosy_13_0_lz => x_rsc_triosy_13_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_13_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_12_0_obj_inst : hybrid_core_x_rsc_triosy_12_0_obj
    PORT MAP(
      x_rsc_triosy_12_0_lz => x_rsc_triosy_12_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_12_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_11_0_obj_inst : hybrid_core_x_rsc_triosy_11_0_obj
    PORT MAP(
      x_rsc_triosy_11_0_lz => x_rsc_triosy_11_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_11_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_10_0_obj_inst : hybrid_core_x_rsc_triosy_10_0_obj
    PORT MAP(
      x_rsc_triosy_10_0_lz => x_rsc_triosy_10_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_10_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_9_0_obj_inst : hybrid_core_x_rsc_triosy_9_0_obj
    PORT MAP(
      x_rsc_triosy_9_0_lz => x_rsc_triosy_9_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_9_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_8_0_obj_inst : hybrid_core_x_rsc_triosy_8_0_obj
    PORT MAP(
      x_rsc_triosy_8_0_lz => x_rsc_triosy_8_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_8_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_7_0_obj_inst : hybrid_core_x_rsc_triosy_7_0_obj
    PORT MAP(
      x_rsc_triosy_7_0_lz => x_rsc_triosy_7_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_7_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_6_0_obj_inst : hybrid_core_x_rsc_triosy_6_0_obj
    PORT MAP(
      x_rsc_triosy_6_0_lz => x_rsc_triosy_6_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_6_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_5_0_obj_inst : hybrid_core_x_rsc_triosy_5_0_obj
    PORT MAP(
      x_rsc_triosy_5_0_lz => x_rsc_triosy_5_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_5_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_4_0_obj_inst : hybrid_core_x_rsc_triosy_4_0_obj
    PORT MAP(
      x_rsc_triosy_4_0_lz => x_rsc_triosy_4_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_4_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_3_0_obj_inst : hybrid_core_x_rsc_triosy_3_0_obj
    PORT MAP(
      x_rsc_triosy_3_0_lz => x_rsc_triosy_3_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_3_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_2_0_obj_inst : hybrid_core_x_rsc_triosy_2_0_obj
    PORT MAP(
      x_rsc_triosy_2_0_lz => x_rsc_triosy_2_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_2_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_1_0_obj_inst : hybrid_core_x_rsc_triosy_1_0_obj
    PORT MAP(
      x_rsc_triosy_1_0_lz => x_rsc_triosy_1_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_1_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_x_rsc_triosy_0_0_obj_inst : hybrid_core_x_rsc_triosy_0_0_obj
    PORT MAP(
      x_rsc_triosy_0_0_lz => x_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      x_rsc_triosy_0_0_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_m_rsc_triosy_obj_inst : hybrid_core_m_rsc_triosy_obj
    PORT MAP(
      m_rsc_triosy_lz => m_rsc_triosy_lz,
      core_wten => core_wten,
      m_rsc_triosy_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_twiddle_rsc_triosy_obj_inst : hybrid_core_twiddle_rsc_triosy_obj
    PORT MAP(
      twiddle_rsc_triosy_lz => twiddle_rsc_triosy_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_twiddle_h_rsc_triosy_obj_inst : hybrid_core_twiddle_h_rsc_triosy_obj
    PORT MAP(
      twiddle_h_rsc_triosy_lz => twiddle_h_rsc_triosy_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_revArr_rsc_triosy_obj_inst : hybrid_core_revArr_rsc_triosy_obj
    PORT MAP(
      revArr_rsc_triosy_lz => revArr_rsc_triosy_lz,
      core_wten => core_wten,
      revArr_rsc_triosy_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_tw_rsc_triosy_obj_inst : hybrid_core_tw_rsc_triosy_obj
    PORT MAP(
      tw_rsc_triosy_lz => tw_rsc_triosy_lz,
      core_wten => core_wten,
      tw_rsc_triosy_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_tw_h_rsc_triosy_obj_inst : hybrid_core_tw_h_rsc_triosy_obj
    PORT MAP(
      tw_h_rsc_triosy_lz => tw_h_rsc_triosy_lz,
      core_wten => core_wten,
      tw_h_rsc_triosy_obj_iswt0 => reg_x_rsc_triosy_31_0_obj_iswt0_cse
    );
  hybrid_core_staller_inst : hybrid_core_staller
    PORT MAP(
      clk => clk,
      rst => rst,
      core_wen => core_wen,
      core_wten => core_wten,
      revArr_rsci_wen_comp => revArr_rsci_wen_comp,
      tw_rsci_wen_comp => tw_rsci_wen_comp,
      tw_h_rsci_wen_comp => tw_h_rsci_wen_comp,
      x_rsc_0_0_i_wen_comp => x_rsc_0_0_i_wen_comp,
      x_rsc_0_0_i_wen_comp_1 => x_rsc_0_0_i_wen_comp_1,
      x_rsc_1_0_i_wen_comp => x_rsc_1_0_i_wen_comp,
      x_rsc_1_0_i_wen_comp_1 => x_rsc_1_0_i_wen_comp_1,
      x_rsc_2_0_i_wen_comp => x_rsc_2_0_i_wen_comp,
      x_rsc_2_0_i_wen_comp_1 => x_rsc_2_0_i_wen_comp_1,
      x_rsc_3_0_i_wen_comp => x_rsc_3_0_i_wen_comp,
      x_rsc_3_0_i_wen_comp_1 => x_rsc_3_0_i_wen_comp_1,
      x_rsc_4_0_i_wen_comp => x_rsc_4_0_i_wen_comp,
      x_rsc_4_0_i_wen_comp_1 => x_rsc_4_0_i_wen_comp_1,
      x_rsc_5_0_i_wen_comp => x_rsc_5_0_i_wen_comp,
      x_rsc_5_0_i_wen_comp_1 => x_rsc_5_0_i_wen_comp_1,
      x_rsc_6_0_i_wen_comp => x_rsc_6_0_i_wen_comp,
      x_rsc_6_0_i_wen_comp_1 => x_rsc_6_0_i_wen_comp_1,
      x_rsc_7_0_i_wen_comp => x_rsc_7_0_i_wen_comp,
      x_rsc_7_0_i_wen_comp_1 => x_rsc_7_0_i_wen_comp_1,
      x_rsc_8_0_i_wen_comp => x_rsc_8_0_i_wen_comp,
      x_rsc_8_0_i_wen_comp_1 => x_rsc_8_0_i_wen_comp_1,
      x_rsc_9_0_i_wen_comp => x_rsc_9_0_i_wen_comp,
      x_rsc_9_0_i_wen_comp_1 => x_rsc_9_0_i_wen_comp_1,
      x_rsc_10_0_i_wen_comp => x_rsc_10_0_i_wen_comp,
      x_rsc_10_0_i_wen_comp_1 => x_rsc_10_0_i_wen_comp_1,
      x_rsc_11_0_i_wen_comp => x_rsc_11_0_i_wen_comp,
      x_rsc_11_0_i_wen_comp_1 => x_rsc_11_0_i_wen_comp_1,
      x_rsc_12_0_i_wen_comp => x_rsc_12_0_i_wen_comp,
      x_rsc_12_0_i_wen_comp_1 => x_rsc_12_0_i_wen_comp_1,
      x_rsc_13_0_i_wen_comp => x_rsc_13_0_i_wen_comp,
      x_rsc_13_0_i_wen_comp_1 => x_rsc_13_0_i_wen_comp_1,
      x_rsc_14_0_i_wen_comp => x_rsc_14_0_i_wen_comp,
      x_rsc_14_0_i_wen_comp_1 => x_rsc_14_0_i_wen_comp_1,
      x_rsc_15_0_i_wen_comp => x_rsc_15_0_i_wen_comp,
      x_rsc_15_0_i_wen_comp_1 => x_rsc_15_0_i_wen_comp_1,
      x_rsc_16_0_i_wen_comp => x_rsc_16_0_i_wen_comp,
      x_rsc_16_0_i_wen_comp_1 => x_rsc_16_0_i_wen_comp_1,
      x_rsc_17_0_i_wen_comp => x_rsc_17_0_i_wen_comp,
      x_rsc_17_0_i_wen_comp_1 => x_rsc_17_0_i_wen_comp_1,
      x_rsc_18_0_i_wen_comp => x_rsc_18_0_i_wen_comp,
      x_rsc_18_0_i_wen_comp_1 => x_rsc_18_0_i_wen_comp_1,
      x_rsc_19_0_i_wen_comp => x_rsc_19_0_i_wen_comp,
      x_rsc_19_0_i_wen_comp_1 => x_rsc_19_0_i_wen_comp_1,
      x_rsc_20_0_i_wen_comp => x_rsc_20_0_i_wen_comp,
      x_rsc_20_0_i_wen_comp_1 => x_rsc_20_0_i_wen_comp_1,
      x_rsc_21_0_i_wen_comp => x_rsc_21_0_i_wen_comp,
      x_rsc_21_0_i_wen_comp_1 => x_rsc_21_0_i_wen_comp_1,
      x_rsc_22_0_i_wen_comp => x_rsc_22_0_i_wen_comp,
      x_rsc_22_0_i_wen_comp_1 => x_rsc_22_0_i_wen_comp_1,
      x_rsc_23_0_i_wen_comp => x_rsc_23_0_i_wen_comp,
      x_rsc_23_0_i_wen_comp_1 => x_rsc_23_0_i_wen_comp_1,
      x_rsc_24_0_i_wen_comp => x_rsc_24_0_i_wen_comp,
      x_rsc_24_0_i_wen_comp_1 => x_rsc_24_0_i_wen_comp_1,
      x_rsc_25_0_i_wen_comp => x_rsc_25_0_i_wen_comp,
      x_rsc_25_0_i_wen_comp_1 => x_rsc_25_0_i_wen_comp_1,
      x_rsc_26_0_i_wen_comp => x_rsc_26_0_i_wen_comp,
      x_rsc_26_0_i_wen_comp_1 => x_rsc_26_0_i_wen_comp_1,
      x_rsc_27_0_i_wen_comp => x_rsc_27_0_i_wen_comp,
      x_rsc_27_0_i_wen_comp_1 => x_rsc_27_0_i_wen_comp_1,
      x_rsc_28_0_i_wen_comp => x_rsc_28_0_i_wen_comp,
      x_rsc_28_0_i_wen_comp_1 => x_rsc_28_0_i_wen_comp_1,
      x_rsc_29_0_i_wen_comp => x_rsc_29_0_i_wen_comp,
      x_rsc_29_0_i_wen_comp_1 => x_rsc_29_0_i_wen_comp_1,
      x_rsc_30_0_i_wen_comp => x_rsc_30_0_i_wen_comp,
      x_rsc_30_0_i_wen_comp_1 => x_rsc_30_0_i_wen_comp_1,
      x_rsc_31_0_i_wen_comp => x_rsc_31_0_i_wen_comp,
      x_rsc_31_0_i_wen_comp_1 => x_rsc_31_0_i_wen_comp_1
    );
  hybrid_core_core_fsm_inst : hybrid_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      core_wen => core_wen,
      fsm_output => hybrid_core_core_fsm_inst_fsm_output,
      S1_OUTER_LOOP_for_C_5_tr0 => hybrid_core_core_fsm_inst_S1_OUTER_LOOP_for_C_5_tr0,
      S1_OUTER_LOOP_C_0_tr0 => hybrid_core_core_fsm_inst_S1_OUTER_LOOP_C_0_tr0,
      S2_COPY_LOOP_for_C_4_tr0 => hybrid_core_core_fsm_inst_S2_COPY_LOOP_for_C_4_tr0,
      S2_COPY_LOOP_C_0_tr0 => hybrid_core_core_fsm_inst_S2_COPY_LOOP_C_0_tr0,
      S2_INNER_LOOP1_for_C_20_tr0 => hybrid_core_core_fsm_inst_S2_INNER_LOOP1_for_C_20_tr0,
      S2_INNER_LOOP1_C_2_tr0 => hybrid_core_core_fsm_inst_S2_INNER_LOOP1_C_2_tr0,
      S2_INNER_LOOP2_for_C_20_tr0 => hybrid_core_core_fsm_inst_S2_INNER_LOOP2_for_C_20_tr0,
      S2_INNER_LOOP2_C_2_tr0 => hybrid_core_core_fsm_inst_S2_INNER_LOOP2_C_2_tr0,
      S2_INNER_LOOP2_C_2_tr1 => hybrid_core_core_fsm_inst_S2_INNER_LOOP2_C_2_tr1,
      S2_INNER_LOOP3_for_C_20_tr0 => hybrid_core_core_fsm_inst_S2_INNER_LOOP3_for_C_20_tr0,
      S2_INNER_LOOP3_C_2_tr0 => hybrid_core_core_fsm_inst_S2_INNER_LOOP3_C_2_tr0,
      S34_OUTER_LOOP_for_C_12_tr0 => hybrid_core_core_fsm_inst_S34_OUTER_LOOP_for_C_12_tr0,
      S34_OUTER_LOOP_C_0_tr0 => hybrid_core_core_fsm_inst_S34_OUTER_LOOP_C_0_tr0,
      S5_COPY_LOOP_for_C_4_tr0 => hybrid_core_core_fsm_inst_S5_COPY_LOOP_for_C_4_tr0,
      S5_COPY_LOOP_C_0_tr0 => hybrid_core_core_fsm_inst_S5_COPY_LOOP_C_0_tr0,
      S5_INNER_LOOP1_for_C_20_tr0 => hybrid_core_core_fsm_inst_S5_INNER_LOOP1_for_C_20_tr0,
      S5_INNER_LOOP1_C_2_tr0 => hybrid_core_core_fsm_inst_S5_INNER_LOOP1_C_2_tr0,
      S5_INNER_LOOP2_for_C_20_tr0 => hybrid_core_core_fsm_inst_S5_INNER_LOOP2_for_C_20_tr0,
      S5_INNER_LOOP2_C_2_tr0 => hybrid_core_core_fsm_inst_S5_INNER_LOOP2_C_2_tr0,
      S5_INNER_LOOP2_C_2_tr1 => hybrid_core_core_fsm_inst_S5_INNER_LOOP2_C_2_tr1,
      S5_INNER_LOOP3_for_C_20_tr0 => hybrid_core_core_fsm_inst_S5_INNER_LOOP3_for_C_20_tr0,
      S5_INNER_LOOP3_C_2_tr0 => hybrid_core_core_fsm_inst_S5_INNER_LOOP3_C_2_tr0,
      S6_OUTER_LOOP_for_C_4_tr0 => hybrid_core_core_fsm_inst_S6_OUTER_LOOP_for_C_4_tr0,
      S6_OUTER_LOOP_C_0_tr0 => hybrid_core_core_fsm_inst_S6_OUTER_LOOP_C_0_tr0
    );
  fsm_output <= hybrid_core_core_fsm_inst_fsm_output;
  hybrid_core_core_fsm_inst_S1_OUTER_LOOP_for_C_5_tr0 <= NOT operator_20_true_1_slc_operator_20_true_1_acc_14_itm;
  hybrid_core_core_fsm_inst_S1_OUTER_LOOP_C_0_tr0 <= S1_OUTER_LOOP_k_5_0_sva_2(5);
  hybrid_core_core_fsm_inst_S2_COPY_LOOP_for_C_4_tr0 <= S2_COPY_LOOP_for_i_5_0_sva_1_5;
  hybrid_core_core_fsm_inst_S2_COPY_LOOP_C_0_tr0 <= z_out(5);
  hybrid_core_core_fsm_inst_S2_INNER_LOOP1_for_C_20_tr0 <= S1_OUTER_LOOP_for_acc_svs_3_0(3);
  hybrid_core_core_fsm_inst_S2_INNER_LOOP1_C_2_tr0 <= S2_INNER_LOOP1_r_4_0_sva_2(4);
  hybrid_core_core_fsm_inst_S2_INNER_LOOP2_for_C_20_tr0 <= S1_OUTER_LOOP_for_acc_svs_3_0(3);
  hybrid_core_core_fsm_inst_S2_INNER_LOOP2_C_2_tr0 <= and_dcpl_53;
  hybrid_core_core_fsm_inst_S2_INNER_LOOP2_C_2_tr1 <= NOT (S2_INNER_LOOP1_r_4_0_sva_2(4));
  hybrid_core_core_fsm_inst_S2_INNER_LOOP3_for_C_20_tr0 <= S1_OUTER_LOOP_for_acc_svs_3_0(3);
  hybrid_core_core_fsm_inst_S2_INNER_LOOP3_C_2_tr0 <= S2_INNER_LOOP1_r_4_0_sva_2(4);
  hybrid_core_core_fsm_inst_S34_OUTER_LOOP_for_C_12_tr0 <= NOT operator_20_true_8_slc_operator_20_true_8_acc_14_itm;
  hybrid_core_core_fsm_inst_S34_OUTER_LOOP_C_0_tr0 <= S1_OUTER_LOOP_k_5_0_sva_2(5);
  hybrid_core_core_fsm_inst_S5_COPY_LOOP_for_C_4_tr0 <= S2_COPY_LOOP_for_i_5_0_sva_1_5;
  hybrid_core_core_fsm_inst_S5_COPY_LOOP_C_0_tr0 <= z_out(5);
  hybrid_core_core_fsm_inst_S5_INNER_LOOP1_for_C_20_tr0 <= S1_OUTER_LOOP_for_acc_svs_3_0(3);
  hybrid_core_core_fsm_inst_S5_INNER_LOOP1_C_2_tr0 <= S2_INNER_LOOP1_r_4_0_sva_2(4);
  hybrid_core_core_fsm_inst_S5_INNER_LOOP2_for_C_20_tr0 <= S1_OUTER_LOOP_for_acc_svs_3_0(3);
  hybrid_core_core_fsm_inst_S5_INNER_LOOP2_C_2_tr0 <= and_dcpl_53;
  hybrid_core_core_fsm_inst_S5_INNER_LOOP2_C_2_tr1 <= NOT (S2_INNER_LOOP1_r_4_0_sva_2(4));
  hybrid_core_core_fsm_inst_S5_INNER_LOOP3_for_C_20_tr0 <= S1_OUTER_LOOP_for_acc_svs_3_0(3);
  hybrid_core_core_fsm_inst_S5_INNER_LOOP3_C_2_tr0 <= S2_INNER_LOOP1_r_4_0_sva_2(4);
  hybrid_core_core_fsm_inst_S6_OUTER_LOOP_for_C_4_tr0 <= NOT operator_20_true_15_slc_operator_20_true_15_acc_14_itm;
  hybrid_core_core_fsm_inst_S6_OUTER_LOOP_C_0_tr0 <= z_out(5);

  S34_OUTER_LOOP_for_tf_mul_cmp_b <= S34_OUTER_LOOP_for_k_slc_S34_OUTER_LOOP_for_k_sva_19_5_4_0_1
      & S34_OUTER_LOOP_for_k_sva_4_0;
  or_299_nl <= (NOT (fsm_output(6))) OR (fsm_output(1)) OR (fsm_output(5));
  or_298_nl <= (fsm_output(6)) OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  mux_109_nl <= MUX_s_1_2_2(or_299_nl, or_298_nl, fsm_output(3));
  nor_2167_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR mux_109_nl);
  and_2097_nl <= (NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("011"))))
      AND mux_108_cse;
  mux_110_nl <= MUX_s_1_2_2(nor_2167_nl, and_2097_nl, fsm_output(0));
  nor_2170_nl <= NOT((fsm_output(3)) OR (fsm_output(6)) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)));
  nor_2171_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)));
  mux_107_nl <= MUX_s_1_2_2(nor_2170_nl, nor_2171_nl, fsm_output(4));
  and_2098_nl <= (NOT((fsm_output(0)) OR (NOT (fsm_output(2))))) AND mux_107_nl;
  mux_111_rmff <= MUX_s_1_2_2(mux_110_nl, and_2098_nl, fsm_output(7));
  S2_INNER_LOOP2_tf_and_nl <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0))
      AND operator_33_true_return_2_3_0_sva_2_0;
  and_90_nl <= and_dcpl_57 AND and_2893_cse AND and_dcpl_79;
  S2_INNER_LOOP1_tfh_mux1h_rmff <= MUX1HOT_v_3_3_2((S2_INNER_LOOP1_tf_and_psp_sva_1(2
      DOWNTO 0)), S2_INNER_LOOP2_tf_and_nl, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), STD_LOGIC_VECTOR'( and_90_nl & and_dcpl_84 & and_dcpl_86));
  S2_INNER_LOOP1_tfh_or_nl <= and_dcpl_84 OR and_dcpl_86;
  S2_INNER_LOOP1_tfh_S2_INNER_LOOP1_tfh_mux_rmff <= MUX_s_1_2_2((S2_INNER_LOOP1_tf_and_psp_sva_1(3)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), S2_INNER_LOOP1_tfh_or_nl);
  or_340_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_132_nl <= MUX_s_1_2_2(or_340_nl, or_338_cse, fsm_output(3));
  mux_133_nl <= MUX_s_1_2_2(mux_132_nl, or_337_cse, fsm_output(1));
  mux_134_nl <= MUX_s_1_2_2(mux_133_nl, or_tmp_156, fsm_output(4));
  mux_131_nl <= MUX_s_1_2_2(mux_tmp_128, or_336_cse, fsm_output(4));
  mux_135_nl <= MUX_s_1_2_2(mux_134_nl, mux_131_nl, fsm_output(0));
  or_335_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_129_nl <= MUX_s_1_2_2(or_335_nl, or_tmp_156, fsm_output(4));
  or_332_nl <= (fsm_output(4)) OR mux_tmp_128;
  mux_130_nl <= MUX_s_1_2_2(mux_129_nl, or_332_nl, fsm_output(0));
  mux_136_nl <= MUX_s_1_2_2(mux_135_nl, mux_130_nl, or_2186_cse);
  or_327_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_137_nl <= MUX_s_1_2_2(mux_136_nl, or_327_nl, fsm_output(2));
  or_326_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_124_nl <= MUX_s_1_2_2(or_326_nl, mux_tmp_121, fsm_output(4));
  or_323_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_122_nl <= MUX_s_1_2_2(or_324_cse, or_323_nl, or_2189_cse);
  or_325_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_122_nl;
  mux_123_nl <= MUX_s_1_2_2(or_325_nl, mux_tmp_121, fsm_output(4));
  mux_125_nl <= MUX_s_1_2_2(mux_124_nl, mux_123_nl, fsm_output(0));
  or_317_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_118_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_134, or_315_cse);
  or_316_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_118_nl;
  mux_119_nl <= MUX_s_1_2_2(or_317_nl, or_316_nl, fsm_output(4));
  or_313_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_115_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_134, or_309_cse);
  or_312_nl <= (fsm_output(6)) OR mux_115_nl;
  mux_116_nl <= MUX_s_1_2_2(or_312_nl, or_tmp_131, fsm_output(3));
  nand_8_nl <= NOT((fsm_output(1)) AND (NOT mux_116_nl));
  mux_117_nl <= MUX_s_1_2_2(or_313_nl, nand_8_nl, fsm_output(4));
  mux_120_nl <= MUX_s_1_2_2(mux_119_nl, mux_117_nl, fsm_output(0));
  mux_126_nl <= MUX_s_1_2_2(mux_125_nl, mux_120_nl, fsm_output(2));
  mux_138_itm <= MUX_s_1_2_2(mux_137_nl, mux_126_nl, fsm_output(5));
  mux_167_cse <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(7));
  or_4679_cse <= (NOT (fsm_output(3))) OR (fsm_output(7));
  nor_2152_cse <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00000")));
  mux_162_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), fsm_output(1));
  and_2086_nl <= or_4679_cse AND (fsm_output(6));
  mux_169_nl <= MUX_s_1_2_2(mux_213_cse, and_2086_nl, fsm_output(1));
  mux_170_nl <= MUX_s_1_2_2(mux_169_nl, nor_tmp_35, fsm_output(0));
  or_374_nl <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(3));
  mux_168_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_374_nl);
  mux_171_cse <= MUX_s_1_2_2(mux_170_nl, mux_168_nl, fsm_output(4));
  mux_163_cse <= MUX_s_1_2_2(mux_162_cse, mux_213_cse, fsm_output(0));
  nor_2139_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2140_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_187_nl <= MUX_s_1_2_2(nor_2139_nl, nor_2140_nl, fsm_output(2));
  and_2084_nl <= (fsm_output(3)) AND mux_187_nl;
  nor_2141_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_186);
  mux_188_nl <= MUX_s_1_2_2(and_2084_nl, nor_2141_nl, fsm_output(4));
  and_2085_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_186);
  mux_189_nl <= MUX_s_1_2_2(mux_188_nl, and_2085_nl, fsm_output(5));
  mux_182_nl <= MUX_s_1_2_2(nor_2144_cse, (fsm_output(1)), fsm_output(0));
  mux_183_nl <= MUX_s_1_2_2(mux_182_nl, or_401_cse, fsm_output(2));
  or_400_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_184_nl <= MUX_s_1_2_2((NOT mux_183_nl), or_400_nl, or_2245_cse);
  nor_2143_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_184_nl);
  mux_185_nl <= MUX_s_1_2_2(nor_2142_cse, nor_2143_nl, fsm_output(5));
  mux_190_nl <= MUX_s_1_2_2(mux_189_nl, mux_185_nl, fsm_output(6));
  mux_180_nl <= MUX_s_1_2_2(or_395_cse, or_394_cse, fsm_output(3));
  or_396_nl <= (fsm_output(4)) OR mux_180_nl;
  or_392_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  nor_2146_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT or_tmp_207));
  or_389_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0000"));
  mux_176_nl <= MUX_s_1_2_2(nor_2146_nl, or_tmp_207, or_389_nl);
  mux_177_nl <= MUX_s_1_2_2(or_2242_cse, mux_176_nl, fsm_output(1));
  nand_10_nl <= NOT((fsm_output(1)) AND (NOT(or_387_cse AND or_tmp_207)));
  mux_178_nl <= MUX_s_1_2_2(mux_177_nl, nand_10_nl, fsm_output(0));
  mux_179_nl <= MUX_s_1_2_2(or_392_nl, mux_178_nl, fsm_output(2));
  or_393_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_179_nl;
  mux_181_nl <= MUX_s_1_2_2(or_396_nl, or_393_nl, fsm_output(5));
  nor_2145_nl <= NOT((fsm_output(6)) OR mux_181_nl);
  mux_191_rmff <= MUX_s_1_2_2(mux_190_nl, nor_2145_nl, fsm_output(7));
  or_435_cse <= (fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  and_2074_nl <= ((fsm_output(1)) OR (fsm_output(7))) AND (fsm_output(6));
  mux_222_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, fsm_output(1));
  mux_223_cse <= MUX_s_1_2_2(and_2074_nl, mux_222_nl, fsm_output(3));
  mux_224_nl <= MUX_s_1_2_2(mux_223_cse, nor_tmp_35, or_435_cse);
  or_434_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_221_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_434_nl);
  mux_225_nl <= MUX_s_1_2_2(mux_224_nl, mux_221_nl, fsm_output(4));
  mux_226_cse <= MUX_s_1_2_2(mux_225_nl, nor_tmp_35, fsm_output(5));
  mux_213_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), fsm_output(3));
  nor_2124_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_231);
  nor_2122_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2123_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_237_nl <= MUX_s_1_2_2(nor_2122_nl, nor_2123_nl, fsm_output(2));
  and_2073_nl <= (fsm_output(3)) AND mux_237_nl;
  mux_238_nl <= MUX_s_1_2_2(and_2073_nl, nor_2124_cse, fsm_output(4));
  nor_2125_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  mux_239_nl <= MUX_s_1_2_2(mux_238_nl, nor_2125_nl, fsm_output(5));
  nand_494_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_234_nl <= MUX_s_1_2_2(nand_494_nl, nor_2186_cse, fsm_output(2));
  or_458_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_235_nl <= MUX_s_1_2_2(mux_234_nl, or_458_nl, or_2294_cse);
  nor_2127_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_235_nl);
  mux_236_nl <= MUX_s_1_2_2(nor_2142_cse, nor_2127_nl, fsm_output(5));
  mux_240_nl <= MUX_s_1_2_2(mux_239_nl, mux_236_nl, fsm_output(6));
  or_453_nl <= (fsm_output(2)) OR mux_tmp_231;
  mux_232_nl <= MUX_s_1_2_2(or_453_nl, or_394_cse, fsm_output(3));
  or_454_nl <= (fsm_output(4)) OR mux_232_nl;
  nand_495_nl <= NOT(or_447_cse AND or_tmp_263);
  nand_496_nl <= NOT(or_445_cse AND or_tmp_263);
  mux_229_nl <= MUX_s_1_2_2(nand_495_nl, nand_496_nl, fsm_output(0));
  nand_14_nl <= NOT((fsm_output(1)) AND mux_229_nl);
  mux_230_nl <= MUX_s_1_2_2(or_448_cse, nand_14_nl, fsm_output(2));
  or_449_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_230_nl;
  mux_233_nl <= MUX_s_1_2_2(or_454_nl, or_449_nl, fsm_output(5));
  nor_2130_nl <= NOT((fsm_output(6)) OR mux_233_nl);
  mux_241_rmff <= MUX_s_1_2_2(mux_240_nl, nor_2130_nl, fsm_output(7));
  nor_2103_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2104_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_289_nl <= MUX_s_1_2_2(nor_2103_nl, nor_2104_nl, fsm_output(2));
  and_2062_nl <= (fsm_output(3)) AND mux_289_nl;
  mux_290_nl <= MUX_s_1_2_2(and_2062_nl, nor_2124_cse, fsm_output(4));
  nor_2106_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  nor_2107_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  mux_288_nl <= MUX_s_1_2_2(nor_2106_nl, nor_2107_nl, fsm_output(2));
  and_2063_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_288_nl;
  mux_291_nl <= MUX_s_1_2_2(mux_290_nl, and_2063_nl, fsm_output(5));
  nand_491_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_285_nl <= MUX_s_1_2_2(nand_491_nl, nor_2186_cse, fsm_output(2));
  or_512_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_286_nl <= MUX_s_1_2_2(mux_285_nl, or_512_nl, or_2338_cse);
  nor_2109_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_286_nl);
  mux_287_nl <= MUX_s_1_2_2(nor_2142_cse, nor_2109_nl, fsm_output(5));
  mux_292_nl <= MUX_s_1_2_2(mux_291_nl, mux_287_nl, fsm_output(6));
  or_508_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  and_2064_nl <= nand_492_cse AND or_tmp_317;
  or_503_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"));
  mux_280_nl <= MUX_s_1_2_2(and_2064_nl, or_tmp_317, or_503_nl);
  and_203_nl <= or_501_cse AND or_tmp_317;
  mux_281_nl <= MUX_s_1_2_2(mux_280_nl, and_203_nl, fsm_output(0));
  nand_17_nl <= NOT((fsm_output(1)) AND (NOT mux_281_nl));
  mux_283_nl <= MUX_s_1_2_2(mux_tmp_231, nand_17_nl, fsm_output(2));
  or_507_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_283_nl;
  mux_284_nl <= MUX_s_1_2_2(or_508_nl, or_507_nl, fsm_output(5));
  nor_2112_nl <= NOT((fsm_output(6)) OR mux_284_nl);
  mux_293_rmff <= MUX_s_1_2_2(mux_292_nl, nor_2112_nl, fsm_output(7));
  or_579_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_353_nl <= MUX_s_1_2_2(or_579_nl, or_tmp_386, fsm_output(4));
  or_577_nl <= (fsm_output(4)) OR mux_tmp_347;
  mux_354_nl <= MUX_s_1_2_2(mux_353_nl, or_577_nl, fsm_output(0));
  or_576_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_349_nl <= MUX_s_1_2_2(or_576_nl, or_338_cse, fsm_output(3));
  mux_350_nl <= MUX_s_1_2_2(mux_349_nl, or_337_cse, fsm_output(1));
  mux_351_nl <= MUX_s_1_2_2(mux_350_nl, or_tmp_386, fsm_output(4));
  mux_348_nl <= MUX_s_1_2_2(mux_tmp_347, or_336_cse, fsm_output(4));
  mux_352_nl <= MUX_s_1_2_2(mux_351_nl, mux_348_nl, fsm_output(0));
  mux_355_nl <= MUX_s_1_2_2(mux_354_nl, mux_352_nl, nor_690_cse);
  or_567_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_356_nl <= MUX_s_1_2_2(mux_355_nl, or_567_nl, fsm_output(2));
  or_566_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_343_nl <= MUX_s_1_2_2(or_566_nl, mux_tmp_340, fsm_output(4));
  or_563_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_341_nl <= MUX_s_1_2_2(or_324_cse, or_563_nl, or_2386_cse);
  or_565_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_341_nl;
  mux_342_nl <= MUX_s_1_2_2(or_565_nl, mux_tmp_340, fsm_output(4));
  mux_344_nl <= MUX_s_1_2_2(mux_343_nl, mux_342_nl, fsm_output(0));
  or_557_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_337_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_365, or_555_cse);
  or_556_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_337_nl;
  mux_338_nl <= MUX_s_1_2_2(or_557_nl, or_556_nl, fsm_output(4));
  or_553_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_334_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_365, or_549_cse);
  or_552_nl <= (fsm_output(6)) OR mux_334_nl;
  mux_335_nl <= MUX_s_1_2_2(or_552_nl, or_tmp_362, fsm_output(3));
  nand_21_nl <= NOT((fsm_output(1)) AND (NOT mux_335_nl));
  mux_336_nl <= MUX_s_1_2_2(or_553_nl, nand_21_nl, fsm_output(4));
  mux_339_nl <= MUX_s_1_2_2(mux_338_nl, mux_336_nl, fsm_output(0));
  mux_345_nl <= MUX_s_1_2_2(mux_344_nl, mux_339_nl, fsm_output(2));
  mux_357_itm <= MUX_s_1_2_2(mux_356_nl, mux_345_nl, fsm_output(5));
  nor_2078_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(1))));
  nor_2079_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(1)));
  mux_404_nl <= MUX_s_1_2_2(nor_2078_nl, nor_2079_nl, fsm_output(2));
  and_2041_nl <= (fsm_output(3)) AND mux_404_nl;
  nor_2080_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_403);
  mux_405_nl <= MUX_s_1_2_2(and_2041_nl, nor_2080_nl, fsm_output(4));
  and_2042_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_403);
  mux_406_nl <= MUX_s_1_2_2(mux_405_nl, and_2042_nl, fsm_output(5));
  nor_2083_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(1))));
  mux_399_nl <= MUX_s_1_2_2(nor_2083_nl, (fsm_output(1)), fsm_output(0));
  mux_400_nl <= MUX_s_1_2_2(mux_399_nl, or_401_cse, fsm_output(2));
  or_640_nl <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(1)));
  mux_401_nl <= MUX_s_1_2_2((NOT mux_400_nl), or_640_nl, or_2440_cse);
  nor_2082_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_401_nl);
  mux_402_nl <= MUX_s_1_2_2(nor_2081_cse, nor_2082_nl, fsm_output(5));
  mux_407_nl <= MUX_s_1_2_2(mux_406_nl, mux_402_nl, fsm_output(6));
  mux_397_nl <= MUX_s_1_2_2(or_634_cse, or_632_cse, fsm_output(3));
  or_635_nl <= (fsm_output(4)) OR mux_397_nl;
  or_629_nl <= (NOT (fsm_output(0))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR
      (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01"));
  or_627_nl <= (fsm_output(1)) OR (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))));
  mux_392_nl <= MUX_s_1_2_2(or_627_nl, (fsm_output(1)), reg_S2_COPY_LOOP_for_i_5_0_2_reg(2));
  mux_393_nl <= MUX_s_1_2_2(mux_tmp_391, (NOT mux_392_nl), S6_OUTER_LOOP_for_acc_tmp(0));
  or_621_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010"));
  mux_394_nl <= MUX_s_1_2_2(mux_393_nl, mux_tmp_391, or_621_nl);
  or_620_nl <= (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  mux_390_nl <= MUX_s_1_2_2((NOT (fsm_output(1))), or_620_nl, or_618_cse);
  mux_395_nl <= MUX_s_1_2_2(mux_394_nl, mux_390_nl, fsm_output(0));
  mux_396_nl <= MUX_s_1_2_2(or_629_nl, mux_395_nl, fsm_output(2));
  or_630_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_396_nl;
  mux_398_nl <= MUX_s_1_2_2(or_635_nl, or_630_nl, fsm_output(5));
  nor_2084_nl <= NOT((fsm_output(6)) OR mux_398_nl);
  mux_408_rmff <= MUX_s_1_2_2(mux_407_nl, nor_2084_nl, fsm_output(7));
  or_673_cse <= (fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_672_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_435_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_672_nl);
  mux_438_nl <= MUX_s_1_2_2(mux_223_cse, nor_tmp_35, or_673_cse);
  mux_439_nl <= MUX_s_1_2_2(mux_438_nl, mux_435_cse, fsm_output(4));
  mux_440_cse <= MUX_s_1_2_2(mux_439_nl, nor_tmp_35, fsm_output(5));
  nor_2066_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_445);
  nor_2064_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2065_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_451_nl <= MUX_s_1_2_2(nor_2064_nl, nor_2065_nl, fsm_output(2));
  and_2031_nl <= (fsm_output(3)) AND mux_451_nl;
  mux_452_nl <= MUX_s_1_2_2(and_2031_nl, nor_2066_cse, fsm_output(4));
  nor_2067_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_453_nl <= MUX_s_1_2_2(mux_452_nl, nor_2067_nl, fsm_output(5));
  nand_482_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_448_nl <= MUX_s_1_2_2(nand_482_nl, nor_2186_cse, fsm_output(2));
  or_699_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_449_nl <= MUX_s_1_2_2(mux_448_nl, or_699_nl, or_2487_cse);
  nor_2069_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_449_nl);
  mux_450_nl <= MUX_s_1_2_2(nor_2081_cse, nor_2069_nl, fsm_output(5));
  mux_454_nl <= MUX_s_1_2_2(mux_453_nl, mux_450_nl, fsm_output(6));
  or_694_nl <= (fsm_output(2)) OR mux_tmp_445;
  mux_446_nl <= MUX_s_1_2_2(or_694_nl, or_632_cse, fsm_output(3));
  or_695_nl <= (fsm_output(4)) OR mux_446_nl;
  nand_483_nl <= NOT(or_684_cse AND or_tmp_493);
  nand_484_nl <= NOT(or_682_cse AND or_tmp_493);
  mux_443_nl <= MUX_s_1_2_2(nand_483_nl, nand_484_nl, fsm_output(0));
  nand_26_nl <= NOT((fsm_output(1)) AND mux_443_nl);
  mux_444_nl <= MUX_s_1_2_2(or_686_cse, nand_26_nl, fsm_output(2));
  or_687_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_444_nl;
  mux_447_nl <= MUX_s_1_2_2(or_695_nl, or_687_nl, fsm_output(5));
  nor_2072_nl <= NOT((fsm_output(6)) OR mux_447_nl);
  mux_455_rmff <= MUX_s_1_2_2(mux_454_nl, nor_2072_nl, fsm_output(7));
  nor_132_cse <= NOT((fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  and_2020_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111")) AND (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2050_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_500_nl <= MUX_s_1_2_2(and_2020_nl, nor_2050_nl, fsm_output(2));
  and_2019_nl <= (fsm_output(3)) AND mux_500_nl;
  mux_501_nl <= MUX_s_1_2_2(and_2019_nl, nor_2066_cse, fsm_output(4));
  nor_2052_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  nor_2053_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_499_nl <= MUX_s_1_2_2(nor_2052_nl, nor_2053_nl, fsm_output(2));
  and_2021_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_499_nl;
  mux_502_nl <= MUX_s_1_2_2(mux_501_nl, and_2021_nl, fsm_output(5));
  nand_478_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_496_nl <= MUX_s_1_2_2(nand_478_nl, nor_2186_cse, fsm_output(2));
  or_750_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_497_nl <= MUX_s_1_2_2(mux_496_nl, or_750_nl, or_2528_cse);
  nor_2055_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_497_nl);
  mux_498_nl <= MUX_s_1_2_2(nor_2081_cse, nor_2055_nl, fsm_output(5));
  mux_503_nl <= MUX_s_1_2_2(mux_502_nl, mux_498_nl, fsm_output(6));
  or_746_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  and_2022_nl <= nand_479_cse AND or_tmp_545;
  or_738_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  mux_491_nl <= MUX_s_1_2_2(and_2022_nl, or_tmp_545, or_738_nl);
  and_259_nl <= or_735_cse AND or_tmp_545;
  mux_492_nl <= MUX_s_1_2_2(mux_491_nl, and_259_nl, fsm_output(0));
  nand_29_nl <= NOT((fsm_output(1)) AND (NOT mux_492_nl));
  mux_494_nl <= MUX_s_1_2_2(mux_tmp_445, nand_29_nl, fsm_output(2));
  or_744_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_494_nl;
  mux_495_nl <= MUX_s_1_2_2(or_746_nl, or_744_nl, fsm_output(5));
  nor_2058_nl <= NOT((fsm_output(6)) OR mux_495_nl);
  mux_504_rmff <= MUX_s_1_2_2(mux_503_nl, nor_2058_nl, fsm_output(7));
  or_820_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_560_nl <= MUX_s_1_2_2(or_820_nl, or_338_cse, fsm_output(3));
  mux_561_nl <= MUX_s_1_2_2(mux_560_nl, or_337_cse, fsm_output(1));
  mux_562_nl <= MUX_s_1_2_2(mux_561_nl, or_tmp_620, fsm_output(4));
  mux_559_nl <= MUX_s_1_2_2(mux_tmp_556, or_336_cse, fsm_output(4));
  mux_563_nl <= MUX_s_1_2_2(mux_562_nl, mux_559_nl, fsm_output(0));
  or_815_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_557_nl <= MUX_s_1_2_2(or_815_nl, or_tmp_620, fsm_output(4));
  or_812_nl <= (fsm_output(4)) OR mux_tmp_556;
  mux_558_nl <= MUX_s_1_2_2(mux_557_nl, or_812_nl, fsm_output(0));
  mux_564_nl <= MUX_s_1_2_2(mux_563_nl, mux_558_nl, or_2574_cse);
  or_807_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_565_nl <= MUX_s_1_2_2(mux_564_nl, or_807_nl, fsm_output(2));
  or_806_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_552_nl <= MUX_s_1_2_2(or_806_nl, mux_tmp_549, fsm_output(4));
  or_803_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_550_nl <= MUX_s_1_2_2(or_324_cse, or_803_nl, or_2577_cse);
  or_805_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_550_nl;
  mux_551_nl <= MUX_s_1_2_2(or_805_nl, mux_tmp_549, fsm_output(4));
  mux_553_nl <= MUX_s_1_2_2(mux_552_nl, mux_551_nl, fsm_output(0));
  or_797_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_546_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_598, or_795_cse);
  or_796_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_546_nl;
  mux_547_nl <= MUX_s_1_2_2(or_797_nl, or_796_nl, fsm_output(4));
  or_793_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_543_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_598, or_789_cse);
  or_792_nl <= (fsm_output(6)) OR mux_543_nl;
  mux_544_nl <= MUX_s_1_2_2(or_792_nl, or_tmp_595, fsm_output(3));
  nand_33_nl <= NOT((fsm_output(1)) AND (NOT mux_544_nl));
  mux_545_nl <= MUX_s_1_2_2(or_793_nl, nand_33_nl, fsm_output(4));
  mux_548_nl <= MUX_s_1_2_2(mux_547_nl, mux_545_nl, fsm_output(0));
  mux_554_nl <= MUX_s_1_2_2(mux_553_nl, mux_548_nl, fsm_output(2));
  mux_566_itm <= MUX_s_1_2_2(mux_565_nl, mux_554_nl, fsm_output(5));
  nor_2027_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2028_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_610_nl <= MUX_s_1_2_2(nor_2027_nl, nor_2028_nl, fsm_output(2));
  and_1999_nl <= (fsm_output(3)) AND mux_610_nl;
  nor_2029_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_609);
  mux_611_nl <= MUX_s_1_2_2(and_1999_nl, nor_2029_nl, fsm_output(4));
  and_2000_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_609);
  mux_612_nl <= MUX_s_1_2_2(mux_611_nl, and_2000_nl, fsm_output(5));
  mux_605_nl <= MUX_s_1_2_2(nor_2032_cse, (fsm_output(1)), fsm_output(0));
  mux_606_nl <= MUX_s_1_2_2(mux_605_nl, or_401_cse, fsm_output(2));
  or_869_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_607_nl <= MUX_s_1_2_2((NOT mux_606_nl), or_869_nl, or_2622_cse);
  nor_2031_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_607_nl);
  mux_608_nl <= MUX_s_1_2_2(nor_2030_cse, nor_2031_nl, fsm_output(5));
  mux_613_nl <= MUX_s_1_2_2(mux_612_nl, mux_608_nl, fsm_output(6));
  mux_603_nl <= MUX_s_1_2_2(or_864_cse, or_863_cse, fsm_output(3));
  or_865_nl <= (fsm_output(4)) OR mux_603_nl;
  or_861_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  nor_2034_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT or_233_cse));
  or_858_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0100"));
  mux_599_nl <= MUX_s_1_2_2(nor_2034_nl, or_233_cse, or_858_nl);
  mux_600_nl <= MUX_s_1_2_2(or_2619_cse, mux_599_nl, fsm_output(1));
  nand_35_nl <= NOT((fsm_output(1)) AND (NOT(or_856_cse AND or_233_cse)));
  mux_601_nl <= MUX_s_1_2_2(mux_600_nl, nand_35_nl, fsm_output(0));
  mux_602_nl <= MUX_s_1_2_2(or_861_nl, mux_601_nl, fsm_output(2));
  or_862_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_602_nl;
  mux_604_nl <= MUX_s_1_2_2(or_865_nl, or_862_nl, fsm_output(5));
  nor_2033_nl <= NOT((fsm_output(6)) OR mux_604_nl);
  mux_614_rmff <= MUX_s_1_2_2(mux_613_nl, nor_2033_nl, fsm_output(7));
  or_898_cse <= (fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_897_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_641_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_897_nl);
  mux_644_nl <= MUX_s_1_2_2(mux_223_cse, nor_tmp_35, or_898_cse);
  mux_645_nl <= MUX_s_1_2_2(mux_644_nl, mux_641_cse, fsm_output(4));
  mux_646_cse <= MUX_s_1_2_2(mux_645_nl, nor_tmp_35, fsm_output(5));
  nor_2014_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_651);
  nor_2012_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_2013_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_657_nl <= MUX_s_1_2_2(nor_2012_nl, nor_2013_nl, fsm_output(2));
  and_1989_nl <= (fsm_output(3)) AND mux_657_nl;
  mux_658_nl <= MUX_s_1_2_2(and_1989_nl, nor_2014_cse, fsm_output(4));
  nor_2015_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  mux_659_nl <= MUX_s_1_2_2(mux_658_nl, nor_2015_nl, fsm_output(5));
  nand_468_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_654_nl <= MUX_s_1_2_2(nand_468_nl, nor_2186_cse, fsm_output(2));
  or_921_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_655_nl <= MUX_s_1_2_2(mux_654_nl, or_921_nl, or_2664_cse);
  nor_2017_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_655_nl);
  mux_656_nl <= MUX_s_1_2_2(nor_2030_cse, nor_2017_nl, fsm_output(5));
  mux_660_nl <= MUX_s_1_2_2(mux_659_nl, mux_656_nl, fsm_output(6));
  or_916_nl <= (fsm_output(2)) OR mux_tmp_651;
  mux_652_nl <= MUX_s_1_2_2(or_916_nl, or_863_cse, fsm_output(3));
  or_917_nl <= (fsm_output(4)) OR mux_652_nl;
  nand_469_nl <= NOT(or_910_cse AND or_261_cse);
  nand_470_nl <= NOT(or_908_cse AND or_261_cse);
  mux_649_nl <= MUX_s_1_2_2(nand_469_nl, nand_470_nl, fsm_output(0));
  nand_39_nl <= NOT((fsm_output(1)) AND mux_649_nl);
  mux_650_nl <= MUX_s_1_2_2(or_911_cse, nand_39_nl, fsm_output(2));
  or_912_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_650_nl;
  mux_653_nl <= MUX_s_1_2_2(or_917_nl, or_912_nl, fsm_output(5));
  nor_2020_nl <= NOT((fsm_output(6)) OR mux_653_nl);
  mux_661_rmff <= MUX_s_1_2_2(mux_660_nl, nor_2020_nl, fsm_output(7));
  and_1978_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1011")) AND (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_1998_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_706_nl <= MUX_s_1_2_2(and_1978_nl, nor_1998_nl, fsm_output(2));
  and_1977_nl <= (fsm_output(3)) AND mux_706_nl;
  mux_707_nl <= MUX_s_1_2_2(and_1977_nl, nor_2014_cse, fsm_output(4));
  nor_2000_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  nor_2001_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  mux_705_nl <= MUX_s_1_2_2(nor_2000_nl, nor_2001_nl, fsm_output(2));
  and_1979_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_705_nl;
  mux_708_nl <= MUX_s_1_2_2(mux_707_nl, and_1979_nl, fsm_output(5));
  nand_465_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_702_nl <= MUX_s_1_2_2(nand_465_nl, nor_2186_cse, fsm_output(2));
  or_970_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_703_nl <= MUX_s_1_2_2(mux_702_nl, or_970_nl, or_2700_cse);
  nor_2003_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_703_nl);
  mux_704_nl <= MUX_s_1_2_2(nor_2030_cse, nor_2003_nl, fsm_output(5));
  mux_709_nl <= MUX_s_1_2_2(mux_708_nl, mux_704_nl, fsm_output(6));
  or_966_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  and_1980_nl <= nand_492_cse AND or_tmp_759;
  or_958_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("010"));
  mux_697_nl <= MUX_s_1_2_2(and_1980_nl, or_tmp_759, or_958_nl);
  and_313_nl <= or_955_cse AND or_tmp_759;
  mux_698_nl <= MUX_s_1_2_2(mux_697_nl, and_313_nl, fsm_output(0));
  nand_42_nl <= NOT((fsm_output(1)) AND (NOT mux_698_nl));
  mux_700_nl <= MUX_s_1_2_2(mux_tmp_651, nand_42_nl, fsm_output(2));
  or_964_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_700_nl;
  mux_701_nl <= MUX_s_1_2_2(or_966_nl, or_964_nl, fsm_output(5));
  nor_2006_nl <= NOT((fsm_output(6)) OR mux_701_nl);
  mux_710_rmff <= MUX_s_1_2_2(mux_709_nl, nor_2006_nl, fsm_output(7));
  or_1036_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_768_nl <= MUX_s_1_2_2(or_1036_nl, or_tmp_830, fsm_output(4));
  or_1034_nl <= (fsm_output(4)) OR mux_tmp_762;
  mux_769_nl <= MUX_s_1_2_2(mux_768_nl, or_1034_nl, fsm_output(0));
  or_1033_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_764_nl <= MUX_s_1_2_2(or_1033_nl, or_338_cse, fsm_output(3));
  mux_765_nl <= MUX_s_1_2_2(mux_764_nl, or_337_cse, fsm_output(1));
  mux_766_nl <= MUX_s_1_2_2(mux_765_nl, or_tmp_830, fsm_output(4));
  mux_763_nl <= MUX_s_1_2_2(mux_tmp_762, or_336_cse, fsm_output(4));
  mux_767_nl <= MUX_s_1_2_2(mux_766_nl, mux_763_nl, fsm_output(0));
  mux_770_nl <= MUX_s_1_2_2(mux_769_nl, mux_767_nl, nor_805_cse);
  or_1024_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_771_nl <= MUX_s_1_2_2(mux_770_nl, or_1024_nl, fsm_output(2));
  or_1023_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_758_nl <= MUX_s_1_2_2(or_1023_nl, mux_tmp_755, fsm_output(4));
  or_1020_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_756_nl <= MUX_s_1_2_2(or_324_cse, or_1020_nl, or_2747_cse);
  or_1022_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_756_nl;
  mux_757_nl <= MUX_s_1_2_2(or_1022_nl, mux_tmp_755, fsm_output(4));
  mux_759_nl <= MUX_s_1_2_2(mux_758_nl, mux_757_nl, fsm_output(0));
  or_1014_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_752_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_809, or_1012_cse);
  or_1013_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_752_nl;
  mux_753_nl <= MUX_s_1_2_2(or_1014_nl, or_1013_nl, fsm_output(4));
  or_1010_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  mux_749_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_809, or_1006_cse);
  or_1009_nl <= (fsm_output(6)) OR mux_749_nl;
  mux_750_nl <= MUX_s_1_2_2(or_1009_nl, or_tmp_806, fsm_output(3));
  nand_46_nl <= NOT((fsm_output(1)) AND (NOT mux_750_nl));
  mux_751_nl <= MUX_s_1_2_2(or_1010_nl, nand_46_nl, fsm_output(4));
  mux_754_nl <= MUX_s_1_2_2(mux_753_nl, mux_751_nl, fsm_output(0));
  mux_760_nl <= MUX_s_1_2_2(mux_759_nl, mux_754_nl, fsm_output(2));
  mux_772_itm <= MUX_s_1_2_2(mux_771_nl, mux_760_nl, fsm_output(5));
  nor_1978_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389);
  or_1083_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  or_1085_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  and_1957_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1101")) AND (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_1976_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_816_nl <= MUX_s_1_2_2(and_1957_nl, nor_1976_nl, fsm_output(2));
  and_1956_nl <= (fsm_output(3)) AND mux_816_nl;
  nor_1977_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_815);
  mux_817_nl <= MUX_s_1_2_2(and_1956_nl, nor_1977_nl, fsm_output(4));
  and_1958_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_815);
  mux_818_nl <= MUX_s_1_2_2(mux_817_nl, and_1958_nl, fsm_output(5));
  nor_1980_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_811_nl <= MUX_s_1_2_2(nor_1980_nl, (fsm_output(1)), fsm_output(0));
  mux_812_nl <= MUX_s_1_2_2(mux_811_nl, or_401_cse, fsm_output(2));
  or_1090_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_813_nl <= MUX_s_1_2_2((NOT mux_812_nl), or_1090_nl, or_2800_cse);
  nor_1979_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_813_nl);
  mux_814_nl <= MUX_s_1_2_2(nor_1978_cse, nor_1979_nl, fsm_output(5));
  mux_819_nl <= MUX_s_1_2_2(mux_818_nl, mux_814_nl, fsm_output(6));
  mux_809_nl <= MUX_s_1_2_2(or_1085_cse, or_1083_cse, fsm_output(3));
  or_1086_nl <= (fsm_output(4)) OR mux_809_nl;
  or_1080_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  or_1078_nl <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  nor_1982_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT or_tmp_875));
  or_1076_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0110"));
  mux_805_nl <= MUX_s_1_2_2(nor_1982_nl, or_tmp_875, or_1076_nl);
  mux_806_nl <= MUX_s_1_2_2(or_1078_nl, mux_805_nl, fsm_output(1));
  nand_48_nl <= NOT((fsm_output(1)) AND (NOT(or_1073_cse AND or_tmp_875)));
  mux_807_nl <= MUX_s_1_2_2(mux_806_nl, nand_48_nl, fsm_output(0));
  mux_808_nl <= MUX_s_1_2_2(or_1080_nl, mux_807_nl, fsm_output(2));
  or_1081_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_808_nl;
  mux_810_nl <= MUX_s_1_2_2(or_1086_nl, or_1081_nl, fsm_output(5));
  nor_1981_nl <= NOT((fsm_output(6)) OR mux_810_nl);
  mux_820_rmff <= MUX_s_1_2_2(mux_819_nl, nor_1981_nl, fsm_output(7));
  nor_245_cse <= NOT((fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011")));
  or_1121_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_847_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1121_nl);
  mux_850_nl <= MUX_s_1_2_2(nor_tmp_35, mux_223_cse, nor_245_cse);
  mux_851_nl <= MUX_s_1_2_2(mux_850_nl, mux_847_cse, fsm_output(4));
  mux_852_cse <= MUX_s_1_2_2(mux_851_nl, nor_tmp_35, fsm_output(5));
  or_1135_cse <= (NOT (fsm_output(1))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR
      not_tmp_389;
  nor_1963_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_857);
  and_1945_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1110")) AND (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_1962_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_863_nl <= MUX_s_1_2_2(and_1945_nl, nor_1962_nl, fsm_output(2));
  and_1944_nl <= (fsm_output(3)) AND mux_863_nl;
  mux_864_nl <= MUX_s_1_2_2(and_1944_nl, nor_1963_cse, fsm_output(4));
  nor_1964_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389);
  mux_865_nl <= MUX_s_1_2_2(mux_864_nl, nor_1964_nl, fsm_output(5));
  nand_453_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4))));
  mux_860_nl <= MUX_s_1_2_2(nand_453_nl, nor_2186_cse, fsm_output(2));
  or_1148_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_861_nl <= MUX_s_1_2_2(mux_860_nl, or_1148_nl, or_2847_cse);
  nor_1966_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_861_nl);
  mux_862_nl <= MUX_s_1_2_2(nor_1978_cse, nor_1966_nl, fsm_output(5));
  mux_866_nl <= MUX_s_1_2_2(mux_865_nl, mux_862_nl, fsm_output(6));
  or_1143_nl <= (fsm_output(2)) OR mux_tmp_857;
  mux_858_nl <= MUX_s_1_2_2(or_1143_nl, or_1083_cse, fsm_output(3));
  or_1144_nl <= (fsm_output(4)) OR mux_858_nl;
  nand_454_nl <= NOT(or_1133_cse AND or_tmp_931);
  nand_455_nl <= NOT(or_1130_cse AND or_tmp_931);
  mux_855_nl <= MUX_s_1_2_2(nand_454_nl, nand_455_nl, fsm_output(0));
  nand_52_nl <= NOT((fsm_output(1)) AND mux_855_nl);
  mux_856_nl <= MUX_s_1_2_2(or_1135_cse, nand_52_nl, fsm_output(2));
  or_1136_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_856_nl;
  mux_859_nl <= MUX_s_1_2_2(or_1144_nl, or_1136_nl, fsm_output(5));
  nor_1969_nl <= NOT((fsm_output(6)) OR mux_859_nl);
  mux_867_rmff <= MUX_s_1_2_2(mux_866_nl, nor_1969_nl, fsm_output(7));
  and_1931_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111")) AND (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  nor_1949_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1111")) OR
      S1_OUTER_LOOP_for_acc_svs_4);
  mux_912_nl <= MUX_s_1_2_2(and_1931_nl, nor_1949_nl, fsm_output(2));
  and_1930_nl <= (fsm_output(3)) AND mux_912_nl;
  mux_913_nl <= MUX_s_1_2_2(and_1930_nl, nor_1963_cse, fsm_output(4));
  nor_1951_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389);
  nor_1952_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389);
  mux_911_nl <= MUX_s_1_2_2(nor_1951_nl, nor_1952_nl, fsm_output(2));
  and_1932_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_911_nl;
  mux_914_nl <= MUX_s_1_2_2(mux_913_nl, and_1932_nl, fsm_output(5));
  nand_445_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4))));
  mux_908_nl <= MUX_s_1_2_2(nand_445_nl, nor_2186_cse, fsm_output(2));
  nand_446_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111")) AND
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_909_nl <= MUX_s_1_2_2(mux_908_nl, nand_446_nl, nand_317_cse);
  nor_1954_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_909_nl);
  mux_910_nl <= MUX_s_1_2_2(nor_1978_cse, nor_1954_nl, fsm_output(5));
  mux_915_nl <= MUX_s_1_2_2(mux_914_nl, mux_910_nl, fsm_output(6));
  or_1192_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  and_1934_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1111"))))
      AND or_tmp_982;
  mux_903_nl <= MUX_s_1_2_2(and_1934_nl, or_tmp_982, S6_OUTER_LOOP_for_acc_tmp(4));
  and_360_nl <= nand_449_cse AND or_tmp_982;
  mux_904_nl <= MUX_s_1_2_2(mux_903_nl, and_360_nl, fsm_output(0));
  nand_55_nl <= NOT((fsm_output(1)) AND (NOT mux_904_nl));
  mux_906_nl <= MUX_s_1_2_2(mux_tmp_857, nand_55_nl, fsm_output(2));
  or_1190_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_906_nl;
  mux_907_nl <= MUX_s_1_2_2(or_1192_nl, or_1190_nl, fsm_output(5));
  nor_1956_nl <= NOT((fsm_output(6)) OR mux_907_nl);
  mux_916_rmff <= MUX_s_1_2_2(mux_915_nl, nor_1956_nl, fsm_output(7));
  and_1919_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  or_1264_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_973_nl <= MUX_s_1_2_2(or_1264_nl, or_338_cse, fsm_output(3));
  mux_974_nl <= MUX_s_1_2_2(mux_973_nl, or_337_cse, fsm_output(1));
  mux_975_nl <= MUX_s_1_2_2(mux_974_nl, or_tmp_1054, fsm_output(4));
  mux_972_nl <= MUX_s_1_2_2(mux_tmp_969, or_336_cse, fsm_output(4));
  mux_976_nl <= MUX_s_1_2_2(mux_975_nl, mux_972_nl, fsm_output(0));
  or_1259_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_970_nl <= MUX_s_1_2_2(or_1259_nl, or_tmp_1054, fsm_output(4));
  or_1256_nl <= (fsm_output(4)) OR mux_tmp_969;
  mux_971_nl <= MUX_s_1_2_2(mux_970_nl, or_1256_nl, fsm_output(0));
  mux_977_nl <= MUX_s_1_2_2(mux_976_nl, mux_971_nl, or_2947_cse);
  or_1251_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_978_nl <= MUX_s_1_2_2(mux_977_nl, or_1251_nl, fsm_output(2));
  or_1250_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_965_nl <= MUX_s_1_2_2(or_1250_nl, mux_tmp_962, fsm_output(4));
  or_1248_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_963_nl <= MUX_s_1_2_2(or_1248_nl, or_324_cse, nor_873_cse);
  or_1249_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_963_nl;
  mux_964_nl <= MUX_s_1_2_2(or_1249_nl, mux_tmp_962, fsm_output(4));
  mux_966_nl <= MUX_s_1_2_2(mux_965_nl, mux_964_nl, fsm_output(0));
  or_1242_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  or_1240_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10000"));
  mux_959_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_1033, or_1240_nl);
  or_1241_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_959_nl;
  mux_960_nl <= MUX_s_1_2_2(or_1242_nl, or_1241_nl, fsm_output(4));
  or_1238_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_955_nl <= MUX_s_1_2_2(or_tmp_1033, (NOT (fsm_output(7))), S1_OUTER_LOOP_for_acc_svs_4);
  or_1234_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"));
  mux_956_nl <= MUX_s_1_2_2(mux_955_nl, or_tmp_1033, or_1234_nl);
  or_1237_nl <= (fsm_output(6)) OR mux_956_nl;
  mux_957_nl <= MUX_s_1_2_2(or_1237_nl, or_tmp_1030, fsm_output(3));
  nand_59_nl <= NOT((fsm_output(1)) AND (NOT mux_957_nl));
  mux_958_nl <= MUX_s_1_2_2(or_1238_nl, nand_59_nl, fsm_output(4));
  mux_961_nl <= MUX_s_1_2_2(mux_960_nl, mux_958_nl, fsm_output(0));
  mux_967_nl <= MUX_s_1_2_2(mux_966_nl, mux_961_nl, fsm_output(2));
  mux_979_itm <= MUX_s_1_2_2(mux_978_nl, mux_967_nl, fsm_output(5));
  nor_1925_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  nor_1926_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1026_nl <= MUX_s_1_2_2(nor_1925_nl, nor_1926_nl, fsm_output(2));
  and_1905_nl <= (fsm_output(3)) AND mux_1026_nl;
  nor_1927_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1025);
  mux_1027_nl <= MUX_s_1_2_2(and_1905_nl, nor_1927_nl, fsm_output(4));
  and_1906_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_1025);
  mux_1028_nl <= MUX_s_1_2_2(mux_1027_nl, and_1906_nl, fsm_output(5));
  mux_1020_nl <= MUX_s_1_2_2(nor_1930_cse, (fsm_output(1)), fsm_output(0));
  mux_1021_nl <= MUX_s_1_2_2(mux_1020_nl, or_401_cse, fsm_output(2));
  mux_1022_nl <= MUX_s_1_2_2(or_tmp_1110, (NOT mux_1021_nl), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  or_1314_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"));
  mux_1023_nl <= MUX_s_1_2_2(mux_1022_nl, or_tmp_1110, or_1314_nl);
  nor_1929_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1023_nl);
  mux_1024_nl <= MUX_s_1_2_2(nor_1928_cse, nor_1929_nl, fsm_output(5));
  mux_1029_nl <= MUX_s_1_2_2(mux_1028_nl, mux_1024_nl, fsm_output(6));
  mux_1018_nl <= MUX_s_1_2_2(or_1310_cse, or_1309_cse, fsm_output(3));
  or_1311_nl <= (fsm_output(4)) OR mux_1018_nl;
  or_1307_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  nor_1932_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT or_tmp_77));
  or_1304_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1000"));
  mux_1014_nl <= MUX_s_1_2_2(nor_1932_nl, or_tmp_77, or_1304_nl);
  mux_1015_nl <= MUX_s_1_2_2(or_2999_cse, mux_1014_nl, fsm_output(1));
  nor_1933_nl <= NOT(S1_OUTER_LOOP_for_acc_svs_4 OR (NOT or_tmp_77));
  or_1301_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"));
  mux_1013_nl <= MUX_s_1_2_2(nor_1933_nl, or_tmp_77, or_1301_nl);
  nand_61_nl <= NOT((fsm_output(1)) AND (NOT mux_1013_nl));
  mux_1016_nl <= MUX_s_1_2_2(mux_1015_nl, nand_61_nl, fsm_output(0));
  mux_1017_nl <= MUX_s_1_2_2(or_1307_nl, mux_1016_nl, fsm_output(2));
  or_1308_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1017_nl;
  mux_1019_nl <= MUX_s_1_2_2(or_1311_nl, or_1308_nl, fsm_output(5));
  nor_1931_nl <= NOT((fsm_output(6)) OR mux_1019_nl);
  mux_1030_rmff <= MUX_s_1_2_2(mux_1029_nl, nor_1931_nl, fsm_output(7));
  or_1344_cse <= (fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1061_nl <= MUX_s_1_2_2(mux_223_cse, nor_tmp_35, or_1344_cse);
  or_1343_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_1058_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1343_nl);
  mux_1062_nl <= MUX_s_1_2_2(mux_1061_nl, mux_1058_nl, fsm_output(4));
  mux_1063_cse <= MUX_s_1_2_2(mux_1062_nl, nor_tmp_35, fsm_output(5));
  nor_1914_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1069);
  nor_1912_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  nor_1913_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1076_nl <= MUX_s_1_2_2(nor_1912_nl, nor_1913_nl, fsm_output(2));
  and_1895_nl <= (fsm_output(3)) AND mux_1076_nl;
  mux_1077_nl <= MUX_s_1_2_2(and_1895_nl, nor_1914_cse, fsm_output(4));
  nor_1915_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  mux_1078_nl <= MUX_s_1_2_2(mux_1077_nl, nor_1915_nl, fsm_output(5));
  nand_434_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4)))));
  mux_1072_nl <= MUX_s_1_2_2(nand_434_nl, nor_2186_cse, fsm_output(2));
  mux_1073_nl <= MUX_s_1_2_2(or_tmp_1162, mux_1072_nl, reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  or_1367_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"));
  mux_1074_nl <= MUX_s_1_2_2(mux_1073_nl, or_tmp_1162, or_1367_nl);
  nor_1917_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1074_nl);
  mux_1075_nl <= MUX_s_1_2_2(nor_1928_cse, nor_1917_nl, fsm_output(5));
  mux_1079_nl <= MUX_s_1_2_2(mux_1078_nl, mux_1075_nl, fsm_output(6));
  or_1363_nl <= (fsm_output(2)) OR mux_tmp_1069;
  mux_1070_nl <= MUX_s_1_2_2(or_1363_nl, or_1309_cse, fsm_output(3));
  or_1364_nl <= (fsm_output(4)) OR mux_1070_nl;
  and_399_nl <= (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10010")))
      AND or_tmp_59;
  nor_1921_nl <= NOT(S1_OUTER_LOOP_for_acc_svs_4 OR (NOT or_tmp_59));
  or_1354_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"));
  mux_1066_nl <= MUX_s_1_2_2(nor_1921_nl, or_tmp_59, or_1354_nl);
  mux_1067_nl <= MUX_s_1_2_2(and_399_nl, mux_1066_nl, fsm_output(0));
  nand_65_nl <= NOT((fsm_output(1)) AND (NOT mux_1067_nl));
  mux_1068_nl <= MUX_s_1_2_2(or_1358_cse, nand_65_nl, fsm_output(2));
  or_1359_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1068_nl;
  mux_1071_nl <= MUX_s_1_2_2(or_1364_nl, or_1359_nl, fsm_output(5));
  nor_1920_nl <= NOT((fsm_output(6)) OR mux_1071_nl);
  mux_1080_rmff <= MUX_s_1_2_2(mux_1079_nl, nor_1920_nl, fsm_output(7));
  and_2140_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0011")) AND S1_OUTER_LOOP_for_acc_svs_4;
  nor_1898_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1128_nl <= MUX_s_1_2_2(and_2140_nl, nor_1898_nl, fsm_output(2));
  and_1884_nl <= (fsm_output(3)) AND mux_1128_nl;
  mux_1129_nl <= MUX_s_1_2_2(and_1884_nl, nor_1914_cse, fsm_output(4));
  nor_1900_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  nor_1901_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  mux_1127_nl <= MUX_s_1_2_2(nor_1900_nl, nor_1901_nl, fsm_output(2));
  and_1885_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_1127_nl;
  mux_1130_nl <= MUX_s_1_2_2(mux_1129_nl, and_1885_nl, fsm_output(5));
  nand_430_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4)))));
  mux_1123_nl <= MUX_s_1_2_2(nand_430_nl, nor_2186_cse, fsm_output(2));
  mux_1124_nl <= MUX_s_1_2_2(or_tmp_1212, mux_1123_nl, reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  or_1419_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"));
  mux_1125_nl <= MUX_s_1_2_2(mux_1124_nl, or_tmp_1212, or_1419_nl);
  nor_1903_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1125_nl);
  mux_1126_nl <= MUX_s_1_2_2(nor_1928_cse, nor_1903_nl, fsm_output(5));
  mux_1131_nl <= MUX_s_1_2_2(mux_1130_nl, mux_1126_nl, fsm_output(6));
  or_1416_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  and_1886_nl <= nand_492_cse AND or_tmp_1200;
  or_1411_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("100"));
  mux_1118_nl <= MUX_s_1_2_2(and_1886_nl, or_tmp_1200, or_1411_nl);
  nor_1907_nl <= NOT(S1_OUTER_LOOP_for_acc_svs_4 OR (NOT or_tmp_1200));
  or_1407_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"));
  mux_1117_nl <= MUX_s_1_2_2(nor_1907_nl, or_tmp_1200, or_1407_nl);
  mux_1119_nl <= MUX_s_1_2_2(mux_1118_nl, mux_1117_nl, fsm_output(0));
  nand_68_nl <= NOT((fsm_output(1)) AND (NOT mux_1119_nl));
  mux_1121_nl <= MUX_s_1_2_2(mux_tmp_1069, nand_68_nl, fsm_output(2));
  or_1415_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1121_nl;
  mux_1122_nl <= MUX_s_1_2_2(or_1416_nl, or_1415_nl, fsm_output(5));
  nor_1906_nl <= NOT((fsm_output(6)) OR mux_1122_nl);
  mux_1132_rmff <= MUX_s_1_2_2(mux_1131_nl, nor_1906_nl, fsm_output(7));
  or_1488_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_1192_nl <= MUX_s_1_2_2(or_1488_nl, or_tmp_1271, fsm_output(4));
  or_1486_nl <= (fsm_output(4)) OR mux_tmp_1186;
  mux_1193_nl <= MUX_s_1_2_2(mux_1192_nl, or_1486_nl, fsm_output(0));
  or_1485_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_1188_nl <= MUX_s_1_2_2(or_1485_nl, or_338_cse, fsm_output(3));
  mux_1189_nl <= MUX_s_1_2_2(mux_1188_nl, or_337_cse, fsm_output(1));
  mux_1190_nl <= MUX_s_1_2_2(mux_1189_nl, or_tmp_1271, fsm_output(4));
  mux_1187_nl <= MUX_s_1_2_2(mux_tmp_1186, or_336_cse, fsm_output(4));
  mux_1191_nl <= MUX_s_1_2_2(mux_1190_nl, mux_1187_nl, fsm_output(0));
  mux_1194_nl <= MUX_s_1_2_2(mux_1193_nl, mux_1191_nl, nor_934_cse);
  or_1476_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1195_nl <= MUX_s_1_2_2(mux_1194_nl, or_1476_nl, fsm_output(2));
  or_1475_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1182_nl <= MUX_s_1_2_2(or_1475_nl, mux_tmp_1179, fsm_output(4));
  or_1473_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1180_nl <= MUX_s_1_2_2(or_1473_nl, or_324_cse, nor_938_cse);
  or_1474_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_1180_nl;
  mux_1181_nl <= MUX_s_1_2_2(or_1474_nl, mux_tmp_1179, fsm_output(4));
  mux_1183_nl <= MUX_s_1_2_2(mux_1182_nl, mux_1181_nl, fsm_output(0));
  or_1467_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  or_1465_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10100"));
  mux_1176_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_1251, or_1465_nl);
  or_1466_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_1176_nl;
  mux_1177_nl <= MUX_s_1_2_2(or_1467_nl, or_1466_nl, fsm_output(4));
  or_1463_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  mux_1172_nl <= MUX_s_1_2_2(or_tmp_1251, (NOT (fsm_output(7))), S1_OUTER_LOOP_for_acc_svs_4);
  or_1459_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"));
  mux_1173_nl <= MUX_s_1_2_2(mux_1172_nl, or_tmp_1251, or_1459_nl);
  or_1462_nl <= (fsm_output(6)) OR mux_1173_nl;
  mux_1174_nl <= MUX_s_1_2_2(or_1462_nl, or_tmp_1248, fsm_output(3));
  nand_72_nl <= NOT((fsm_output(1)) AND (NOT mux_1174_nl));
  mux_1175_nl <= MUX_s_1_2_2(or_1463_nl, nand_72_nl, fsm_output(4));
  mux_1178_nl <= MUX_s_1_2_2(mux_1177_nl, mux_1175_nl, fsm_output(0));
  mux_1184_nl <= MUX_s_1_2_2(mux_1183_nl, mux_1178_nl, fsm_output(2));
  mux_1196_itm <= MUX_s_1_2_2(mux_1195_nl, mux_1184_nl, fsm_output(5));
  and_2132_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0101")) AND S1_OUTER_LOOP_for_acc_svs_4;
  nor_1872_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1244_nl <= MUX_s_1_2_2(and_2132_nl, nor_1872_nl, fsm_output(2));
  and_1862_nl <= (fsm_output(3)) AND mux_1244_nl;
  nor_1873_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1243);
  mux_1245_nl <= MUX_s_1_2_2(and_1862_nl, nor_1873_nl, fsm_output(4));
  and_1863_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_1243);
  mux_1246_nl <= MUX_s_1_2_2(mux_1245_nl, and_1863_nl, fsm_output(5));
  nor_1874_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  mux_1238_nl <= MUX_s_1_2_2(or_tmp_1316, (NOT (fsm_output(1))), fsm_output(0));
  mux_1239_nl <= MUX_s_1_2_2(mux_1238_nl, nor_2186_cse, fsm_output(2));
  mux_1240_nl <= MUX_s_1_2_2(or_tmp_1340, mux_1239_nl, reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  or_1551_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"));
  mux_1241_nl <= MUX_s_1_2_2(mux_1240_nl, or_tmp_1340, or_1551_nl);
  nor_1875_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1241_nl);
  mux_1242_nl <= MUX_s_1_2_2(nor_1874_nl, nor_1875_nl, fsm_output(5));
  mux_1247_nl <= MUX_s_1_2_2(mux_1246_nl, mux_1242_nl, fsm_output(6));
  or_1545_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_1236_nl <= MUX_s_1_2_2(or_1547_cse, or_1545_nl, fsm_output(3));
  or_1548_nl <= (fsm_output(4)) OR mux_1236_nl;
  nand_547_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101")));
  nor_1878_nl <= NOT((fsm_output(1)) OR nor_947_cse);
  mux_1232_nl <= MUX_s_1_2_2(or_tmp_1324, nor_1878_nl, S6_OUTER_LOOP_for_acc_tmp(0));
  or_1534_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1010"));
  mux_1233_nl <= MUX_s_1_2_2(mux_1232_nl, or_tmp_1324, or_1534_nl);
  nor_1880_nl <= NOT((reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) OR (NOT or_tmp_1319));
  or_1530_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"));
  mux_1230_nl <= MUX_s_1_2_2(nor_1880_nl, or_tmp_1319, or_1530_nl);
  nand_74_nl <= NOT((fsm_output(1)) AND (NOT mux_1230_nl));
  mux_1231_nl <= MUX_s_1_2_2(nand_74_nl, or_tmp_1316, or_1527_cse);
  mux_1234_nl <= MUX_s_1_2_2(mux_1233_nl, mux_1231_nl, fsm_output(0));
  mux_1235_nl <= MUX_s_1_2_2(nand_547_nl, mux_1234_nl, fsm_output(2));
  or_1543_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1235_nl;
  mux_1237_nl <= MUX_s_1_2_2(or_1548_nl, or_1543_nl, fsm_output(5));
  nor_1877_nl <= NOT((fsm_output(6)) OR mux_1237_nl);
  mux_1248_rmff <= MUX_s_1_2_2(mux_1247_nl, nor_1877_nl, fsm_output(7));
  nor_389_cse <= NOT((fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  mux_1279_nl <= MUX_s_1_2_2(nor_tmp_35, mux_223_cse, nor_389_cse);
  or_1581_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_1276_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1581_nl);
  mux_1280_nl <= MUX_s_1_2_2(mux_1279_nl, mux_1276_nl, fsm_output(4));
  mux_1281_cse <= MUX_s_1_2_2(mux_1280_nl, nor_tmp_35, fsm_output(5));
  nor_1862_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR not_tmp_590);
  nor_1860_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1287);
  and_2131_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0110")) AND S1_OUTER_LOOP_for_acc_svs_4;
  nor_1859_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1294_nl <= MUX_s_1_2_2(and_2131_nl, nor_1859_nl, fsm_output(2));
  and_1851_nl <= (fsm_output(3)) AND mux_1294_nl;
  mux_1295_nl <= MUX_s_1_2_2(and_1851_nl, nor_1860_cse, fsm_output(4));
  nor_1861_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1110"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR not_tmp_590);
  mux_1296_nl <= MUX_s_1_2_2(mux_1295_nl, nor_1861_nl, fsm_output(5));
  nand_419_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4)))));
  mux_1290_nl <= MUX_s_1_2_2(nand_419_nl, nor_2186_cse, fsm_output(2));
  mux_1291_nl <= MUX_s_1_2_2(or_tmp_1397, mux_1290_nl, reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  or_1609_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"));
  mux_1292_nl <= MUX_s_1_2_2(mux_1291_nl, or_tmp_1397, or_1609_nl);
  nor_1863_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1292_nl);
  mux_1293_nl <= MUX_s_1_2_2(nor_1862_cse, nor_1863_nl, fsm_output(5));
  mux_1297_nl <= MUX_s_1_2_2(mux_1296_nl, mux_1293_nl, fsm_output(6));
  or_1605_nl <= (fsm_output(2)) OR mux_tmp_1287;
  or_1600_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1))
      OR not_tmp_590;
  mux_1288_nl <= MUX_s_1_2_2(or_1605_nl, or_1600_nl, fsm_output(3));
  or_1606_nl <= (fsm_output(4)) OR mux_1288_nl;
  or_1597_nl <= (NOT (fsm_output(1))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR
      not_tmp_590;
  and_444_nl <= (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10110")))
      AND or_tmp_1379;
  nor_1867_nl <= NOT(S1_OUTER_LOOP_for_acc_svs_4 OR (NOT or_tmp_1379));
  or_1591_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"));
  mux_1284_nl <= MUX_s_1_2_2(nor_1867_nl, or_tmp_1379, or_1591_nl);
  mux_1285_nl <= MUX_s_1_2_2(and_444_nl, mux_1284_nl, fsm_output(0));
  nand_78_nl <= NOT((fsm_output(1)) AND (NOT mux_1285_nl));
  mux_1286_nl <= MUX_s_1_2_2(or_1597_nl, nand_78_nl, fsm_output(2));
  or_1598_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1286_nl;
  mux_1289_nl <= MUX_s_1_2_2(or_1606_nl, or_1598_nl, fsm_output(5));
  nor_1866_nl <= NOT((fsm_output(6)) OR mux_1289_nl);
  mux_1298_rmff <= MUX_s_1_2_2(mux_1297_nl, nor_1866_nl, fsm_output(7));
  and_2139_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111")) AND S1_OUTER_LOOP_for_acc_svs_4;
  nor_1843_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1346_nl <= MUX_s_1_2_2(and_2139_nl, nor_1843_nl, fsm_output(2));
  and_1838_nl <= (fsm_output(3)) AND mux_1346_nl;
  mux_1347_nl <= MUX_s_1_2_2(and_1838_nl, nor_1860_cse, fsm_output(4));
  nor_1845_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR not_tmp_590);
  nor_1846_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR not_tmp_590);
  mux_1345_nl <= MUX_s_1_2_2(nor_1845_nl, nor_1846_nl, fsm_output(2));
  and_1839_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_1345_nl;
  mux_1348_nl <= MUX_s_1_2_2(mux_1347_nl, and_1839_nl, fsm_output(5));
  nand_411_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND S1_OUTER_LOOP_for_acc_svs_4)));
  mux_1341_nl <= MUX_s_1_2_2(nand_411_nl, nor_2186_cse, fsm_output(2));
  mux_1342_nl <= MUX_s_1_2_2(or_tmp_1452, mux_1341_nl, reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  nand_413_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0111")));
  mux_1343_nl <= MUX_s_1_2_2(mux_1342_nl, or_tmp_1452, nand_413_nl);
  nor_1848_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1343_nl);
  mux_1344_nl <= MUX_s_1_2_2(nor_1862_cse, nor_1848_nl, fsm_output(5));
  mux_1349_nl <= MUX_s_1_2_2(mux_1348_nl, mux_1344_nl, fsm_output(6));
  or_1663_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1))
      OR not_tmp_590;
  and_1840_nl <= nand_479_cse AND or_tmp_1437;
  or_1655_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10"));
  mux_1336_nl <= MUX_s_1_2_2(and_1840_nl, or_tmp_1437, or_1655_nl);
  nor_1852_nl <= NOT(S1_OUTER_LOOP_for_acc_svs_4 OR (NOT or_tmp_1437));
  nand_415_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111")));
  mux_1335_nl <= MUX_s_1_2_2(nor_1852_nl, or_tmp_1437, nand_415_nl);
  mux_1337_nl <= MUX_s_1_2_2(mux_1336_nl, mux_1335_nl, fsm_output(0));
  nand_81_nl <= NOT((fsm_output(1)) AND (NOT mux_1337_nl));
  mux_1339_nl <= MUX_s_1_2_2(mux_tmp_1287, nand_81_nl, fsm_output(2));
  or_1661_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1339_nl;
  mux_1340_nl <= MUX_s_1_2_2(or_1663_nl, or_1661_nl, fsm_output(5));
  nor_1851_nl <= NOT((fsm_output(6)) OR mux_1340_nl);
  mux_1350_rmff <= MUX_s_1_2_2(mux_1349_nl, nor_1851_nl, fsm_output(7));
  and_1827_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("10"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  or_1740_nl <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_1408_nl <= MUX_s_1_2_2(or_1740_nl, or_338_cse, fsm_output(3));
  mux_1409_nl <= MUX_s_1_2_2(mux_1408_nl, or_337_cse, fsm_output(1));
  mux_1410_nl <= MUX_s_1_2_2(mux_1409_nl, or_tmp_1516, fsm_output(4));
  mux_1407_nl <= MUX_s_1_2_2(mux_tmp_1404, or_336_cse, fsm_output(4));
  mux_1411_nl <= MUX_s_1_2_2(mux_1410_nl, mux_1407_nl, fsm_output(0));
  or_1735_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_1405_nl <= MUX_s_1_2_2(or_1735_nl, or_tmp_1516, fsm_output(4));
  or_1732_nl <= (fsm_output(4)) OR mux_tmp_1404;
  mux_1406_nl <= MUX_s_1_2_2(mux_1405_nl, or_1732_nl, fsm_output(0));
  mux_1412_nl <= MUX_s_1_2_2(mux_1411_nl, mux_1406_nl, or_3367_cse);
  or_1727_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1413_nl <= MUX_s_1_2_2(mux_1412_nl, or_1727_nl, fsm_output(2));
  or_1726_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1400_nl <= MUX_s_1_2_2(or_1726_nl, mux_tmp_1397, fsm_output(4));
  or_1724_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1398_nl <= MUX_s_1_2_2(or_1724_nl, or_324_cse, nor_1010_cse);
  or_1725_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_1398_nl;
  mux_1399_nl <= MUX_s_1_2_2(or_1725_nl, mux_tmp_1397, fsm_output(4));
  mux_1401_nl <= MUX_s_1_2_2(mux_1400_nl, mux_1399_nl, fsm_output(0));
  or_1718_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  or_1716_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11000"));
  mux_1394_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_1495, or_1716_nl);
  or_1717_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_1394_nl;
  mux_1395_nl <= MUX_s_1_2_2(or_1718_nl, or_1717_nl, fsm_output(4));
  or_1714_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  and_1822_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4;
  mux_1390_nl <= MUX_s_1_2_2(or_tmp_1495, (NOT (fsm_output(7))), and_1822_nl);
  or_1710_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_1391_nl <= MUX_s_1_2_2(mux_1390_nl, or_tmp_1495, or_1710_nl);
  or_1713_nl <= (fsm_output(6)) OR mux_1391_nl;
  mux_1392_nl <= MUX_s_1_2_2(or_1713_nl, or_tmp_1492, fsm_output(3));
  nand_85_nl <= NOT((fsm_output(1)) AND (NOT mux_1392_nl));
  mux_1393_nl <= MUX_s_1_2_2(or_1714_nl, nand_85_nl, fsm_output(4));
  mux_1396_nl <= MUX_s_1_2_2(mux_1395_nl, mux_1393_nl, fsm_output(0));
  mux_1402_nl <= MUX_s_1_2_2(mux_1401_nl, mux_1396_nl, fsm_output(2));
  mux_1414_itm <= MUX_s_1_2_2(mux_1413_nl, mux_1402_nl, fsm_output(5));
  nor_1819_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_520_cse);
  nor_1820_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_520_cse);
  mux_1461_nl <= MUX_s_1_2_2(nor_1819_nl, nor_1820_nl, fsm_output(2));
  and_1810_nl <= (fsm_output(3)) AND mux_1461_nl;
  nor_1821_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1460);
  mux_1462_nl <= MUX_s_1_2_2(and_1810_nl, nor_1821_nl, fsm_output(4));
  and_1811_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_1460);
  mux_1463_nl <= MUX_s_1_2_2(mux_1462_nl, and_1811_nl, fsm_output(5));
  nor_1824_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR nand_520_cse);
  mux_1455_nl <= MUX_s_1_2_2(nor_1824_nl, (fsm_output(1)), fsm_output(0));
  mux_1456_nl <= MUX_s_1_2_2(mux_1455_nl, or_401_cse, fsm_output(2));
  mux_1457_nl <= MUX_s_1_2_2(or_tmp_1572, (NOT mux_1456_nl), and_1812_cse);
  or_1788_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_1458_nl <= MUX_s_1_2_2(mux_1457_nl, or_tmp_1572, or_1788_nl);
  nor_1823_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1458_nl);
  mux_1459_nl <= MUX_s_1_2_2(nor_1822_cse, nor_1823_nl, fsm_output(5));
  mux_1464_nl <= MUX_s_1_2_2(mux_1463_nl, mux_1459_nl, fsm_output(6));
  mux_1453_nl <= MUX_s_1_2_2(or_1784_cse, or_1783_cse, fsm_output(3));
  or_1785_nl <= (fsm_output(4)) OR mux_1453_nl;
  nand_401_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  nor_1826_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT or_tmp_1558));
  or_1778_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("1100"));
  mux_1449_nl <= MUX_s_1_2_2(nor_1826_nl, or_tmp_1558, or_1778_nl);
  mux_1450_nl <= MUX_s_1_2_2(or_3418_cse, mux_1449_nl, fsm_output(1));
  and_2130_nl <= nand_520_cse AND or_tmp_1558;
  or_1774_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"));
  mux_1448_nl <= MUX_s_1_2_2(and_2130_nl, or_tmp_1558, or_1774_nl);
  nand_87_nl <= NOT((fsm_output(1)) AND (NOT mux_1448_nl));
  mux_1451_nl <= MUX_s_1_2_2(mux_1450_nl, nand_87_nl, fsm_output(0));
  mux_1452_nl <= MUX_s_1_2_2(nand_401_nl, mux_1451_nl, fsm_output(2));
  or_1782_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1452_nl;
  mux_1454_nl <= MUX_s_1_2_2(or_1785_nl, or_1782_nl, fsm_output(5));
  nor_1825_nl <= NOT((fsm_output(6)) OR mux_1454_nl);
  mux_1465_rmff <= MUX_s_1_2_2(mux_1464_nl, nor_1825_nl, fsm_output(7));
  or_1818_cse <= (fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_1817_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_1493_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1817_nl);
  mux_1496_nl <= MUX_s_1_2_2(mux_223_cse, nor_tmp_35, or_1818_cse);
  mux_1497_nl <= MUX_s_1_2_2(mux_1496_nl, mux_1493_cse, fsm_output(4));
  mux_1498_cse <= MUX_s_1_2_2(mux_1497_nl, nor_tmp_35, fsm_output(5));
  nor_1810_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1504);
  nor_1808_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_520_cse);
  nor_1809_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_520_cse);
  mux_1511_nl <= MUX_s_1_2_2(nor_1808_nl, nor_1809_nl, fsm_output(2));
  and_1797_nl <= (fsm_output(3)) AND mux_1511_nl;
  mux_1512_nl <= MUX_s_1_2_2(and_1797_nl, nor_1810_cse, fsm_output(4));
  and_1798_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110")) AND
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110"));
  mux_1513_nl <= MUX_s_1_2_2(mux_1512_nl, and_1798_nl, fsm_output(5));
  nand_392_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR nand_520_cse))));
  mux_1507_nl <= MUX_s_1_2_2(nand_392_nl, nor_2186_cse, fsm_output(2));
  mux_1508_nl <= MUX_s_1_2_2(or_tmp_1624, mux_1507_nl, and_1812_cse);
  or_1841_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_1509_nl <= MUX_s_1_2_2(mux_1508_nl, or_tmp_1624, or_1841_nl);
  nor_1812_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1509_nl);
  mux_1510_nl <= MUX_s_1_2_2(nor_1822_cse, nor_1812_nl, fsm_output(5));
  mux_1514_nl <= MUX_s_1_2_2(mux_1513_nl, mux_1510_nl, fsm_output(6));
  or_1837_nl <= (fsm_output(2)) OR mux_tmp_1504;
  mux_1505_nl <= MUX_s_1_2_2(or_1837_nl, or_1783_cse, fsm_output(3));
  or_1838_nl <= (fsm_output(4)) OR mux_1505_nl;
  and_487_nl <= (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11010")))
      AND or_tmp_1610;
  and_1800_nl <= nand_520_cse AND or_tmp_1610;
  or_1828_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"));
  mux_1501_nl <= MUX_s_1_2_2(and_1800_nl, or_tmp_1610, or_1828_nl);
  mux_1502_nl <= MUX_s_1_2_2(and_487_nl, mux_1501_nl, fsm_output(0));
  nand_91_nl <= NOT((fsm_output(1)) AND (NOT mux_1502_nl));
  mux_1503_nl <= MUX_s_1_2_2(nand_393_cse, nand_91_nl, fsm_output(2));
  or_1833_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1503_nl;
  mux_1506_nl <= MUX_s_1_2_2(or_1838_nl, or_1833_nl, fsm_output(5));
  nor_1815_nl <= NOT((fsm_output(6)) OR mux_1506_nl);
  mux_1515_rmff <= MUX_s_1_2_2(mux_1514_nl, nor_1815_nl, fsm_output(7));
  nor_1792_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)=STD_LOGIC_VECTOR'("011"))))
      OR nand_520_cse);
  nor_1793_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_520_cse);
  mux_1563_nl <= MUX_s_1_2_2(nor_1792_nl, nor_1793_nl, fsm_output(2));
  and_1784_nl <= (fsm_output(3)) AND mux_1563_nl;
  mux_1564_nl <= MUX_s_1_2_2(and_1784_nl, nor_1810_cse, fsm_output(4));
  and_2144_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110"));
  nor_1796_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110")));
  mux_1562_nl <= MUX_s_1_2_2(and_2144_nl, nor_1796_nl, fsm_output(2));
  and_1785_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_1562_nl;
  mux_1565_nl <= MUX_s_1_2_2(mux_1564_nl, and_1785_nl, fsm_output(5));
  nand_385_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR nand_520_cse))));
  mux_1558_nl <= MUX_s_1_2_2(nand_385_nl, nor_2186_cse, fsm_output(2));
  mux_1559_nl <= MUX_s_1_2_2(or_tmp_1677, mux_1558_nl, and_1812_cse);
  or_1895_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"));
  mux_1560_nl <= MUX_s_1_2_2(mux_1559_nl, or_tmp_1677, or_1895_nl);
  nor_1798_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1560_nl);
  mux_1561_nl <= MUX_s_1_2_2(nor_1822_cse, nor_1798_nl, fsm_output(5));
  mux_1566_nl <= MUX_s_1_2_2(mux_1565_nl, mux_1561_nl, fsm_output(6));
  or_1892_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  and_1787_nl <= nand_492_cse AND or_tmp_1662;
  or_1884_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("110"));
  mux_1553_nl <= MUX_s_1_2_2(and_1787_nl, or_tmp_1662, or_1884_nl);
  and_2129_nl <= nand_520_cse AND or_tmp_1662;
  or_1880_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"));
  mux_1552_nl <= MUX_s_1_2_2(and_2129_nl, or_tmp_1662, or_1880_nl);
  mux_1554_nl <= MUX_s_1_2_2(mux_1553_nl, mux_1552_nl, fsm_output(0));
  nand_94_nl <= NOT((fsm_output(1)) AND (NOT mux_1554_nl));
  mux_1556_nl <= MUX_s_1_2_2(mux_tmp_1504, nand_94_nl, fsm_output(2));
  or_1890_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1556_nl;
  mux_1557_nl <= MUX_s_1_2_2(or_1892_nl, or_1890_nl, fsm_output(5));
  nor_1801_nl <= NOT((fsm_output(6)) OR mux_1557_nl);
  mux_1567_rmff <= MUX_s_1_2_2(mux_1566_nl, nor_1801_nl, fsm_output(7));
  and_1773_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("011"));
  or_1967_nl <= (fsm_output(1)) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  mux_1627_nl <= MUX_s_1_2_2(or_1967_nl, or_tmp_1739, fsm_output(4));
  or_1965_nl <= (fsm_output(4)) OR mux_tmp_1621;
  mux_1628_nl <= MUX_s_1_2_2(mux_1627_nl, or_1965_nl, fsm_output(0));
  nand_550_nl <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  mux_1623_nl <= MUX_s_1_2_2(nand_550_nl, or_338_cse, fsm_output(3));
  mux_1624_nl <= MUX_s_1_2_2(mux_1623_nl, or_337_cse, fsm_output(1));
  mux_1625_nl <= MUX_s_1_2_2(mux_1624_nl, or_tmp_1739, fsm_output(4));
  mux_1622_nl <= MUX_s_1_2_2(mux_tmp_1621, or_336_cse, fsm_output(4));
  mux_1626_nl <= MUX_s_1_2_2(mux_1625_nl, mux_1622_nl, fsm_output(0));
  mux_1629_nl <= MUX_s_1_2_2(mux_1628_nl, mux_1626_nl, and_1380_cse);
  or_1955_nl <= (fsm_output(0)) OR (fsm_output(4)) OR (fsm_output(1)) OR (NOT (fsm_output(3)))
      OR (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1630_nl <= MUX_s_1_2_2(mux_1629_nl, or_1955_nl, fsm_output(2));
  or_1954_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (NOT (fsm_output(6)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1617_nl <= MUX_s_1_2_2(or_1954_nl, mux_tmp_1614, fsm_output(4));
  or_1952_nl <= (NOT (fsm_output(6))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1615_nl <= MUX_s_1_2_2(or_1952_nl, or_324_cse, nor_1089_cse);
  or_1953_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR mux_1615_nl;
  mux_1616_nl <= MUX_s_1_2_2(or_1953_nl, mux_tmp_1614, fsm_output(4));
  mux_1618_nl <= MUX_s_1_2_2(mux_1617_nl, mux_1616_nl, fsm_output(0));
  or_1946_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  or_1944_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11100"));
  mux_1611_nl <= MUX_s_1_2_2((NOT (fsm_output(7))), or_tmp_1719, or_1944_nl);
  or_1945_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(6)) OR mux_1611_nl;
  mux_1612_nl <= MUX_s_1_2_2(or_1946_nl, or_1945_nl, fsm_output(4));
  or_1942_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR CONV_SL_1_1(fsm_output(7 DOWNTO
      6)/=STD_LOGIC_VECTOR'("01"));
  and_1769_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND S1_OUTER_LOOP_for_acc_svs_4;
  mux_1607_nl <= MUX_s_1_2_2(or_tmp_1719, (NOT (fsm_output(7))), and_1769_nl);
  or_1938_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  mux_1608_nl <= MUX_s_1_2_2(mux_1607_nl, or_tmp_1719, or_1938_nl);
  or_1941_nl <= (fsm_output(6)) OR mux_1608_nl;
  mux_1609_nl <= MUX_s_1_2_2(or_1941_nl, or_tmp_1716, fsm_output(3));
  nand_98_nl <= NOT((fsm_output(1)) AND (NOT mux_1609_nl));
  mux_1610_nl <= MUX_s_1_2_2(or_1942_nl, nand_98_nl, fsm_output(4));
  mux_1613_nl <= MUX_s_1_2_2(mux_1612_nl, mux_1610_nl, fsm_output(0));
  mux_1619_nl <= MUX_s_1_2_2(mux_1618_nl, mux_1613_nl, fsm_output(2));
  mux_1631_itm <= MUX_s_1_2_2(mux_1630_nl, mux_1619_nl, fsm_output(5));
  nor_1771_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR nand_336_cse);
  or_2011_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR
      nand_480_cse;
  nor_1768_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"))))
      OR nand_517_cse);
  nor_1769_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_517_cse);
  mux_1678_nl <= MUX_s_1_2_2(nor_1768_nl, nor_1769_nl, fsm_output(2));
  and_1754_nl <= (fsm_output(3)) AND mux_1678_nl;
  nor_1770_nl <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1677);
  mux_1679_nl <= MUX_s_1_2_2(and_1754_nl, nor_1770_nl, fsm_output(4));
  and_1755_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("111")) AND
      (NOT mux_tmp_1677);
  mux_1680_nl <= MUX_s_1_2_2(mux_1679_nl, and_1755_nl, fsm_output(5));
  nor_1773_nl <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR nand_517_cse);
  mux_1672_nl <= MUX_s_1_2_2(nor_1773_nl, (fsm_output(1)), fsm_output(0));
  mux_1673_nl <= MUX_s_1_2_2(mux_1672_nl, or_401_cse, fsm_output(2));
  and_1756_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  mux_1674_nl <= MUX_s_1_2_2(or_tmp_1796, (NOT mux_1673_nl), and_1756_nl);
  or_2016_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  mux_1675_nl <= MUX_s_1_2_2(mux_1674_nl, or_tmp_1796, or_2016_nl);
  nor_1772_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1675_nl);
  mux_1676_nl <= MUX_s_1_2_2(nor_1771_cse, nor_1772_nl, fsm_output(5));
  mux_1681_nl <= MUX_s_1_2_2(mux_1680_nl, mux_1676_nl, fsm_output(6));
  or_2012_nl <= (fsm_output(2)) OR nand_336_cse;
  mux_1670_nl <= MUX_s_1_2_2(or_2012_nl, or_2011_cse, fsm_output(3));
  or_2013_nl <= (fsm_output(4)) OR mux_1670_nl;
  nand_362_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  nor_1775_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT or_tmp_1783));
  nand_363_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110")));
  mux_1666_nl <= MUX_s_1_2_2(nor_1775_nl, or_tmp_1783, nand_363_nl);
  mux_1667_nl <= MUX_s_1_2_2(nand_480_cse, mux_1666_nl, fsm_output(1));
  and_2128_nl <= nand_517_cse AND or_tmp_1783;
  or_2003_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  mux_1665_nl <= MUX_s_1_2_2(and_2128_nl, or_tmp_1783, or_2003_nl);
  nand_100_nl <= NOT((fsm_output(1)) AND (NOT mux_1665_nl));
  mux_1668_nl <= MUX_s_1_2_2(mux_1667_nl, nand_100_nl, fsm_output(0));
  mux_1669_nl <= MUX_s_1_2_2(nand_362_nl, mux_1668_nl, fsm_output(2));
  or_2009_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1669_nl;
  mux_1671_nl <= MUX_s_1_2_2(or_2013_nl, or_2009_nl, fsm_output(5));
  nor_1774_nl <= NOT((fsm_output(6)) OR mux_1671_nl);
  mux_1682_rmff <= MUX_s_1_2_2(mux_1681_nl, nor_1774_nl, fsm_output(7));
  and_1737_cse <= (NOT (fsm_output(0))) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  and_1740_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101"));
  mux_1713_nl <= MUX_s_1_2_2(nor_tmp_35, mux_223_cse, and_1737_cse);
  or_2045_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(3)) OR (fsm_output(1));
  mux_1710_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2045_nl);
  mux_1714_nl <= MUX_s_1_2_2(mux_1713_nl, mux_1710_nl, fsm_output(4));
  mux_1715_cse <= MUX_s_1_2_2(mux_1714_nl, nor_tmp_35, fsm_output(5));
  nor_1758_cse <= NOT(CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))
      OR mux_tmp_1721);
  nor_1756_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("11"))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR nand_351_cse);
  nor_1757_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR nand_351_cse);
  mux_1728_nl <= MUX_s_1_2_2(nor_1756_nl, nor_1757_nl, fsm_output(2));
  and_1733_nl <= (fsm_output(3)) AND mux_1728_nl;
  mux_1729_nl <= MUX_s_1_2_2(and_1733_nl, nor_1758_cse, fsm_output(4));
  nor_1759_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1110"))))
      OR nand_480_cse);
  mux_1730_nl <= MUX_s_1_2_2(mux_1729_nl, nor_1759_nl, fsm_output(5));
  nand_349_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR (NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0))
      OR nand_351_cse))));
  mux_1724_nl <= MUX_s_1_2_2(nand_349_nl, nor_2186_cse, fsm_output(2));
  and_1734_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  mux_1725_nl <= MUX_s_1_2_2(or_tmp_1845, mux_1724_nl, and_1734_nl);
  mux_1726_nl <= MUX_s_1_2_2(mux_1725_nl, or_tmp_1845, reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0));
  nor_1761_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1726_nl);
  mux_1727_nl <= MUX_s_1_2_2(nor_1771_cse, nor_1761_nl, fsm_output(5));
  mux_1731_nl <= MUX_s_1_2_2(mux_1730_nl, mux_1727_nl, fsm_output(6));
  or_2063_nl <= (fsm_output(2)) OR mux_tmp_1721;
  mux_1722_nl <= MUX_s_1_2_2(or_2063_nl, or_2011_cse, fsm_output(3));
  or_2064_nl <= (fsm_output(4)) OR mux_1722_nl;
  and_529_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11110"))))
      AND or_tmp_1833;
  and_1735_nl <= nand_351_cse AND or_tmp_1833;
  mux_1718_nl <= MUX_s_1_2_2(and_1735_nl, or_tmp_1833, S1_OUTER_LOOP_for_acc_svs_3_0(0));
  mux_1719_nl <= MUX_s_1_2_2(and_529_nl, mux_1718_nl, fsm_output(0));
  nand_104_nl <= NOT((fsm_output(1)) AND (NOT mux_1719_nl));
  mux_1720_nl <= MUX_s_1_2_2(nand_336_cse, nand_104_nl, fsm_output(2));
  or_2059_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1720_nl;
  mux_1723_nl <= MUX_s_1_2_2(or_2064_nl, or_2059_nl, fsm_output(5));
  nor_1764_nl <= NOT((fsm_output(6)) OR mux_1723_nl);
  mux_1732_rmff <= MUX_s_1_2_2(mux_1731_nl, nor_1764_nl, fsm_output(7));
  and_1721_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110"));
  and_1708_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111")) AND S1_OUTER_LOOP_for_acc_svs_4;
  nor_1745_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT and_1713_cse));
  mux_1777_nl <= MUX_s_1_2_2(and_1708_nl, nor_1745_nl, fsm_output(2));
  and_1707_nl <= (fsm_output(3)) AND mux_1777_nl;
  mux_1778_nl <= MUX_s_1_2_2(and_1707_nl, nor_1758_cse, fsm_output(4));
  and_1710_nl <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  nor_1747_nl <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_480_cse);
  mux_1776_nl <= MUX_s_1_2_2(and_1710_nl, nor_1747_nl, fsm_output(2));
  and_1709_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11")) AND
      mux_1776_nl;
  mux_1779_nl <= MUX_s_1_2_2(mux_1778_nl, and_1709_nl, fsm_output(5));
  or_4557_nl <= (fsm_output(2)) OR (NOT((fsm_output(1)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4));
  nand_338_nl <= NOT((fsm_output(1)) AND ((fsm_output(0)) OR and_1713_cse));
  mux_1773_nl <= MUX_s_1_2_2(nand_338_nl, nor_2186_cse, fsm_output(2));
  mux_1774_nl <= MUX_s_1_2_2(or_4557_nl, mux_1773_nl, and_1329_cse);
  nor_1749_nl <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"))
      OR mux_1774_nl);
  mux_1775_nl <= MUX_s_1_2_2(nor_1771_cse, nor_1749_nl, fsm_output(5));
  mux_1780_nl <= MUX_s_1_2_2(mux_1779_nl, mux_1775_nl, fsm_output(6));
  or_2108_nl <= (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR nand_480_cse;
  or_2104_nl <= S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_61_cse OR and_1692_cse;
  or_2103_nl <= and_1713_cse OR and_1692_cse;
  mux_1769_nl <= MUX_s_1_2_2(or_2104_nl, or_2103_nl, fsm_output(0));
  nand_339_nl <= NOT((fsm_output(1)) AND mux_1769_nl);
  mux_1771_nl <= MUX_s_1_2_2(mux_tmp_1721, nand_339_nl, fsm_output(2));
  or_2106_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("10")) OR mux_1771_nl;
  mux_1772_nl <= MUX_s_1_2_2(or_2108_nl, or_2106_nl, fsm_output(5));
  nor_1751_nl <= NOT((fsm_output(6)) OR mux_1772_nl);
  mux_1781_rmff <= MUX_s_1_2_2(mux_1780_nl, nor_1751_nl, fsm_output(7));
  and_1692_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  or_2159_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1838_nl <= MUX_s_1_2_2(or_2159_nl, or_2158_cse, fsm_output(1));
  mux_1839_nl <= MUX_s_1_2_2(mux_1838_nl, or_2157_cse, fsm_output(0));
  or_2160_nl <= (fsm_output(6)) OR mux_1839_nl;
  mux_1840_nl <= MUX_s_1_2_2(or_2161_cse, or_2160_nl, fsm_output(2));
  mux_1837_nl <= MUX_s_1_2_2(or_tmp_1928, mux_tmp_1832, fsm_output(6));
  or_2156_nl <= (fsm_output(2)) OR mux_1837_nl;
  mux_1841_nl <= MUX_s_1_2_2(mux_1840_nl, or_2156_nl, fsm_output(4));
  or_2155_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2151_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00000"));
  mux_1833_nl <= MUX_s_1_2_2(mux_tmp_1832, or_tmp_1918, or_2151_nl);
  or_2150_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1831_nl <= MUX_s_1_2_2(or_2150_nl, or_tmp_1924, fsm_output(1));
  mux_1834_nl <= MUX_s_1_2_2(mux_1833_nl, mux_1831_nl, fsm_output(0));
  mux_1835_nl <= MUX_s_1_2_2(or_tmp_1928, mux_1834_nl, fsm_output(6));
  or_2154_nl <= (fsm_output(2)) OR mux_1835_nl;
  mux_1836_nl <= MUX_s_1_2_2(or_2155_nl, or_2154_nl, fsm_output(4));
  mux_1842_nl <= MUX_s_1_2_2(mux_1841_nl, mux_1836_nl, or_2189_cse);
  or_2146_nl <= (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1824_nl <= MUX_s_1_2_2(or_2146_nl, (fsm_output(7)), fsm_output(3));
  mux_1825_nl <= MUX_s_1_2_2(or_2147_cse, mux_1824_nl, fsm_output(1));
  mux_1826_nl <= MUX_s_1_2_2(mux_1825_nl, mux_tmp_1821, fsm_output(0));
  mux_1827_nl <= MUX_s_1_2_2(mux_1826_nl, mux_tmp_1820, fsm_output(6));
  mux_1828_nl <= MUX_s_1_2_2(mux_1827_nl, nand_331_cse, fsm_output(2));
  mux_1822_nl <= MUX_s_1_2_2(or_tmp_1918, mux_tmp_1821, fsm_output(0));
  mux_1823_nl <= MUX_s_1_2_2(mux_1822_nl, mux_tmp_1820, fsm_output(6));
  or_2144_nl <= (fsm_output(2)) OR mux_1823_nl;
  mux_1829_nl <= MUX_s_1_2_2(mux_1828_nl, or_2144_nl, or_2186_cse);
  or_2137_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1830_nl <= MUX_s_1_2_2(mux_1829_nl, or_2137_nl, fsm_output(4));
  mux_1843_itm <= MUX_s_1_2_2(mux_1842_nl, mux_1830_nl, fsm_output(5));
  nor_1730_cse <= NOT((fsm_output(0)) OR (fsm_output(2)));
  nor_636_cse <= NOT((fsm_output(1)) OR (NOT (fsm_output(3))));
  or_2186_cse <= CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("000"));
  or_2189_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_2194_cse <= (fsm_output(0)) OR (fsm_output(2));
  mux_1876_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2194_cse);
  and_1675_nl <= (nor_1730_cse OR (fsm_output(7))) AND (fsm_output(6));
  mux_1877_cse <= MUX_s_1_2_2(mux_1876_nl, and_1675_nl, fsm_output(4));
  and_1677_nl <= (fsm_output(4)) AND (fsm_output(0)) AND (fsm_output(2));
  mux_1872_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1677_nl);
  mux_1867_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, fsm_output(2));
  and_1678_nl <= ((fsm_output(2)) OR (fsm_output(7))) AND (fsm_output(6));
  mux_1868_cse <= MUX_s_1_2_2(mux_1867_nl, and_1678_nl, fsm_output(0));
  mux_1865_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), fsm_output(2));
  and_1676_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00000"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1878_nl <= MUX_s_1_2_2(mux_1877_cse, and_1676_nl, or_2189_cse);
  mux_1879_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1878_nl, nor_636_cse);
  or_2188_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_1873_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2188_nl);
  mux_1874_nl <= MUX_s_1_2_2(mux_1873_nl, mux_1872_cse, fsm_output(3));
  mux_1869_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_2186_cse);
  mux_1870_nl <= MUX_s_1_2_2(mux_1869_nl, mux_1865_cse, fsm_output(4));
  mux_1871_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1870_nl, fsm_output(3));
  mux_1875_nl <= MUX_s_1_2_2(mux_1874_nl, mux_1871_nl, fsm_output(1));
  mux_1880_seb <= MUX_s_1_2_2(mux_1879_nl, mux_1875_nl, fsm_output(5));
  nor_1727_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_1896_nl <= MUX_s_1_2_2(nor_1727_nl, (fsm_output(2)), fsm_output(0));
  mux_1897_nl <= MUX_s_1_2_2((NOT mux_1896_nl), (fsm_output(2)), fsm_output(3));
  mux_1898_nl <= MUX_s_1_2_2(mux_1897_nl, or_2215_cse, fsm_output(1));
  or_2217_nl <= (fsm_output(4)) OR mux_1898_nl;
  mux_1894_nl <= MUX_s_1_2_2(or_tmp_1983, (fsm_output(2)), fsm_output(3));
  mux_1895_nl <= MUX_s_1_2_2(mux_1894_nl, or_tmp_1981, fsm_output(1));
  nand_114_nl <= NOT((fsm_output(4)) AND (NOT mux_1895_nl));
  mux_1899_nl <= MUX_s_1_2_2(or_2217_nl, nand_114_nl, fsm_output(6));
  mux_1900_nl <= MUX_s_1_2_2(mux_1899_nl, mux_tmp_1887, fsm_output(5));
  or_2213_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2211_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1888_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_1976, fsm_output(0));
  nor_640_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00001")));
  mux_1889_nl <= MUX_s_1_2_2(or_2211_nl, mux_1888_nl, nor_640_nl);
  mux_1890_nl <= MUX_s_1_2_2(or_tmp_1983, mux_1889_nl, fsm_output(3));
  mux_1891_nl <= MUX_s_1_2_2(mux_1890_nl, or_tmp_1981, fsm_output(1));
  nand_113_nl <= NOT((fsm_output(4)) AND (NOT mux_1891_nl));
  mux_1892_nl <= MUX_s_1_2_2(or_2213_nl, nand_113_nl, fsm_output(6));
  mux_1893_nl <= MUX_s_1_2_2(mux_1892_nl, mux_tmp_1887, fsm_output(5));
  mux_1901_nl <= MUX_s_1_2_2(mux_1900_nl, mux_1893_nl, or_2245_cse);
  nor_1728_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  nor_1729_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  mux_1881_nl <= MUX_s_1_2_2(nor_1728_nl, nor_1729_nl, fsm_output(1));
  nand_111_nl <= NOT(nor_2197_cse AND mux_1881_nl);
  mux_1882_nl <= MUX_s_1_2_2(nand_111_nl, or_2199_cse, fsm_output(5));
  mux_1902_itm <= MUX_s_1_2_2(mux_1901_nl, mux_1882_nl, fsm_output(7));
  or_2242_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_2245_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_2244_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_1925_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2244_nl);
  mux_1926_nl <= MUX_s_1_2_2(mux_1925_nl, mux_1872_cse, fsm_output(3));
  mux_1921_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_2242_cse);
  mux_1922_nl <= MUX_s_1_2_2(mux_1921_nl, mux_1865_cse, fsm_output(4));
  mux_1923_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1922_nl, fsm_output(3));
  mux_1927_cse <= MUX_s_1_2_2(mux_1926_nl, mux_1923_nl, fsm_output(1));
  and_1670_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1930_nl <= MUX_s_1_2_2(mux_1877_cse, and_1670_nl, or_2245_cse);
  mux_1931_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1930_nl, nor_636_cse);
  mux_1932_seb <= MUX_s_1_2_2(mux_1931_nl, mux_1927_cse, fsm_output(5));
  or_2274_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1944_nl <= MUX_s_1_2_2(or_2274_nl, or_2273_cse, fsm_output(0));
  mux_1945_nl <= MUX_s_1_2_2(mux_1944_nl, or_2272_cse, fsm_output(3));
  mux_1946_nl <= MUX_s_1_2_2(mux_1945_nl, or_2271_cse, fsm_output(1));
  mux_1943_nl <= MUX_s_1_2_2(or_tmp_2035, or_119_cse, fsm_output(3));
  or_2270_nl <= (fsm_output(1)) OR mux_1943_nl;
  mux_1947_nl <= MUX_s_1_2_2(mux_1946_nl, or_2270_nl, fsm_output(6));
  mux_1948_nl <= MUX_s_1_2_2(mux_1947_nl, mux_tmp_1938, fsm_output(5));
  or_2268_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2265_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_2263_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1939_nl <= MUX_s_1_2_2(or_2265_nl, or_2263_nl, fsm_output(0));
  mux_1940_nl <= MUX_s_1_2_2(or_tmp_2035, mux_1939_nl, fsm_output(3));
  or_2267_nl <= (fsm_output(1)) OR mux_1940_nl;
  mux_1941_nl <= MUX_s_1_2_2(or_2268_nl, or_2267_nl, fsm_output(6));
  mux_1942_nl <= MUX_s_1_2_2(mux_1941_nl, mux_tmp_1938, fsm_output(5));
  mux_1949_nl <= MUX_s_1_2_2(mux_1948_nl, mux_1942_nl, or_2294_cse);
  or_2254_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1933_nl <= MUX_s_1_2_2(or_2254_nl, or_2199_cse, fsm_output(5));
  mux_1950_itm <= MUX_s_1_2_2(mux_1949_nl, mux_1933_nl, fsm_output(7));
  or_2294_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1659_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1988_nl <= MUX_s_1_2_2(mux_1877_cse, and_1659_nl, or_2294_cse);
  mux_1989_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1988_nl, nor_636_cse);
  mux_1990_seb <= MUX_s_1_2_2(mux_1989_nl, mux_1927_cse, fsm_output(5));
  nor_1703_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_2004_nl <= MUX_s_1_2_2(nor_1703_nl, (fsm_output(2)), fsm_output(0));
  mux_2005_nl <= MUX_s_1_2_2((NOT mux_2004_nl), or_4378_cse, fsm_output(1));
  mux_2006_nl <= MUX_s_1_2_2(mux_2005_nl, or_4699_cse, fsm_output(3));
  or_2317_nl <= (fsm_output(6)) OR mux_2006_nl;
  mux_2003_nl <= MUX_s_1_2_2(mux_tmp_1999, or_4699_cse, fsm_output(3));
  nand_119_nl <= NOT((fsm_output(6)) AND (NOT mux_2003_nl));
  mux_2007_nl <= MUX_s_1_2_2(or_2317_nl, nand_119_nl, fsm_output(4));
  mux_2008_nl <= MUX_s_1_2_2(mux_2007_nl, mux_tmp_1996, fsm_output(5));
  or_2313_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_1997_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2075, fsm_output(0));
  nor_664_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00011")));
  mux_1998_nl <= MUX_s_1_2_2(or_tmp_2076, mux_1997_nl, nor_664_nl);
  or_2311_nl <= (fsm_output(1)) OR mux_1998_nl;
  mux_2000_nl <= MUX_s_1_2_2(mux_tmp_1999, or_2311_nl, fsm_output(3));
  nand_118_nl <= NOT((fsm_output(6)) AND (NOT mux_2000_nl));
  mux_2001_nl <= MUX_s_1_2_2(or_2313_nl, nand_118_nl, fsm_output(4));
  mux_2002_nl <= MUX_s_1_2_2(mux_2001_nl, mux_tmp_1996, fsm_output(5));
  mux_2009_nl <= MUX_s_1_2_2(mux_2008_nl, mux_2002_nl, or_2338_cse);
  or_2303_nl <= (fsm_output(0)) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1991_nl <= MUX_s_1_2_2(or_tmp_2071, or_2303_nl, fsm_output(1));
  or_4537_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_1991_nl;
  mux_1992_nl <= MUX_s_1_2_2(or_4537_nl, or_2199_cse, fsm_output(5));
  mux_2010_itm <= MUX_s_1_2_2(mux_2009_nl, mux_1992_nl, fsm_output(7));
  or_2338_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1646_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2049_nl <= MUX_s_1_2_2(mux_1877_cse, and_1646_nl, or_2338_cse);
  mux_2050_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2049_nl, nor_636_cse);
  mux_2051_seb <= MUX_s_1_2_2(mux_2050_nl, mux_1927_cse, fsm_output(5));
  or_2367_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2070_nl <= MUX_s_1_2_2(or_2367_nl, or_2158_cse, fsm_output(1));
  mux_2071_nl <= MUX_s_1_2_2(mux_2070_nl, or_2157_cse, fsm_output(0));
  or_2368_nl <= (fsm_output(6)) OR mux_2071_nl;
  mux_2072_nl <= MUX_s_1_2_2(or_2161_cse, or_2368_nl, fsm_output(2));
  mux_2069_nl <= MUX_s_1_2_2(or_tmp_2126, mux_tmp_2064, fsm_output(6));
  or_2364_nl <= (fsm_output(2)) OR mux_2069_nl;
  mux_2073_nl <= MUX_s_1_2_2(mux_2072_nl, or_2364_nl, fsm_output(4));
  or_2363_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2359_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00100"));
  mux_2065_nl <= MUX_s_1_2_2(mux_tmp_2064, or_tmp_2119, or_2359_nl);
  or_2358_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2063_nl <= MUX_s_1_2_2(or_2358_nl, or_tmp_2122, fsm_output(1));
  mux_2066_nl <= MUX_s_1_2_2(mux_2065_nl, mux_2063_nl, fsm_output(0));
  mux_2067_nl <= MUX_s_1_2_2(or_tmp_2126, mux_2066_nl, fsm_output(6));
  or_2362_nl <= (fsm_output(2)) OR mux_2067_nl;
  mux_2068_nl <= MUX_s_1_2_2(or_2363_nl, or_2362_nl, fsm_output(4));
  mux_2074_nl <= MUX_s_1_2_2(mux_2073_nl, mux_2068_nl, or_2386_cse);
  mux_2059_nl <= MUX_s_1_2_2(or_tmp_2119, mux_tmp_2053, fsm_output(0));
  mux_2060_nl <= MUX_s_1_2_2(mux_2059_nl, mux_tmp_2052, fsm_output(6));
  or_2355_nl <= (fsm_output(2)) OR mux_2060_nl;
  or_2352_nl <= (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2054_nl <= MUX_s_1_2_2(or_2352_nl, (fsm_output(7)), fsm_output(3));
  mux_2055_nl <= MUX_s_1_2_2(or_2147_cse, mux_2054_nl, fsm_output(1));
  mux_2056_nl <= MUX_s_1_2_2(mux_2055_nl, mux_tmp_2053, fsm_output(0));
  mux_2057_nl <= MUX_s_1_2_2(mux_2056_nl, mux_tmp_2052, fsm_output(6));
  mux_2058_nl <= MUX_s_1_2_2(mux_2057_nl, nand_331_cse, fsm_output(2));
  mux_2061_nl <= MUX_s_1_2_2(or_2355_nl, mux_2058_nl, nor_690_cse);
  or_2346_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2062_nl <= MUX_s_1_2_2(mux_2061_nl, or_2346_nl, fsm_output(4));
  mux_2075_itm <= MUX_s_1_2_2(mux_2074_nl, mux_2062_nl, fsm_output(5));
  nor_690_cse <= NOT(CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("001")));
  or_2386_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1636_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00100"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2106_nl <= MUX_s_1_2_2(mux_1877_cse, and_1636_nl, or_2386_cse);
  mux_2107_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2106_nl, nor_636_cse);
  or_2385_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2101_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2385_nl);
  mux_2102_nl <= MUX_s_1_2_2(mux_2101_nl, mux_1872_cse, fsm_output(3));
  mux_2097_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, nor_690_cse);
  mux_2098_nl <= MUX_s_1_2_2(mux_2097_nl, mux_1865_cse, fsm_output(4));
  mux_2099_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2098_nl, fsm_output(3));
  mux_2103_nl <= MUX_s_1_2_2(mux_2102_nl, mux_2099_nl, fsm_output(1));
  mux_2108_seb <= MUX_s_1_2_2(mux_2107_nl, mux_2103_nl, fsm_output(5));
  nor_1683_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_2124_nl <= MUX_s_1_2_2(nor_1683_nl, (fsm_output(2)), fsm_output(0));
  mux_2125_nl <= MUX_s_1_2_2((NOT mux_2124_nl), (fsm_output(2)), fsm_output(3));
  mux_2126_nl <= MUX_s_1_2_2(mux_2125_nl, or_2215_cse, fsm_output(1));
  or_2422_nl <= (fsm_output(4)) OR mux_2126_nl;
  mux_2122_nl <= MUX_s_1_2_2(or_tmp_2179, (fsm_output(2)), fsm_output(3));
  mux_2123_nl <= MUX_s_1_2_2(mux_2122_nl, or_tmp_2176, fsm_output(1));
  nand_123_nl <= NOT((fsm_output(4)) AND (NOT mux_2123_nl));
  mux_2127_nl <= MUX_s_1_2_2(or_2422_nl, nand_123_nl, fsm_output(6));
  mux_2128_nl <= MUX_s_1_2_2(mux_2127_nl, mux_tmp_2115, fsm_output(5));
  or_2418_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2415_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2116_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2168, fsm_output(0));
  nor_697_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00101")));
  mux_2117_nl <= MUX_s_1_2_2(or_2415_nl, mux_2116_nl, nor_697_nl);
  mux_2118_nl <= MUX_s_1_2_2(or_tmp_2179, mux_2117_nl, fsm_output(3));
  mux_2119_nl <= MUX_s_1_2_2(mux_2118_nl, or_tmp_2176, fsm_output(1));
  nand_122_nl <= NOT((fsm_output(4)) AND (NOT mux_2119_nl));
  mux_2120_nl <= MUX_s_1_2_2(or_2418_nl, nand_122_nl, fsm_output(6));
  mux_2121_nl <= MUX_s_1_2_2(mux_2120_nl, mux_tmp_2115, fsm_output(5));
  mux_2129_nl <= MUX_s_1_2_2(mux_2128_nl, mux_2121_nl, or_2440_cse);
  nor_1684_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  nor_1685_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_2109_nl <= MUX_s_1_2_2(nor_1684_nl, nor_1685_nl, fsm_output(1));
  nand_120_nl <= NOT(nor_2197_cse AND mux_2109_nl);
  mux_2110_nl <= MUX_s_1_2_2(nand_120_nl, or_2396_cse, fsm_output(5));
  mux_2130_itm <= MUX_s_1_2_2(mux_2129_nl, mux_2110_nl, fsm_output(7));
  nor_701_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  or_2440_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_2439_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2150_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2439_nl);
  mux_2151_nl <= MUX_s_1_2_2(mux_2150_nl, mux_1872_cse, fsm_output(3));
  mux_2146_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, nor_701_cse);
  mux_2147_nl <= MUX_s_1_2_2(mux_2146_nl, mux_1865_cse, fsm_output(4));
  mux_2148_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2147_nl, fsm_output(3));
  mux_2152_cse <= MUX_s_1_2_2(mux_2151_nl, mux_2148_nl, fsm_output(1));
  and_1630_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2155_nl <= MUX_s_1_2_2(mux_1877_cse, and_1630_nl, or_2440_cse);
  mux_2156_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2155_nl, nor_636_cse);
  mux_2157_seb <= MUX_s_1_2_2(mux_2156_nl, mux_2152_cse, fsm_output(5));
  or_2475_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2169_nl <= MUX_s_1_2_2(or_2475_nl, or_2273_cse, fsm_output(0));
  mux_2170_nl <= MUX_s_1_2_2(mux_2169_nl, or_2272_cse, fsm_output(3));
  mux_2171_nl <= MUX_s_1_2_2(mux_2170_nl, or_2271_cse, fsm_output(1));
  mux_2168_nl <= MUX_s_1_2_2(or_tmp_2228, or_119_cse, fsm_output(3));
  or_2471_nl <= (fsm_output(1)) OR mux_2168_nl;
  mux_2172_nl <= MUX_s_1_2_2(mux_2171_nl, or_2471_nl, fsm_output(6));
  mux_2173_nl <= MUX_s_1_2_2(mux_2172_nl, mux_tmp_2163, fsm_output(5));
  or_2469_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2465_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_2463_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2164_nl <= MUX_s_1_2_2(or_2465_nl, or_2463_nl, fsm_output(0));
  mux_2165_nl <= MUX_s_1_2_2(or_tmp_2228, mux_2164_nl, fsm_output(3));
  or_2468_nl <= (fsm_output(1)) OR mux_2165_nl;
  mux_2166_nl <= MUX_s_1_2_2(or_2469_nl, or_2468_nl, fsm_output(6));
  mux_2167_nl <= MUX_s_1_2_2(mux_2166_nl, mux_tmp_2163, fsm_output(5));
  mux_2174_nl <= MUX_s_1_2_2(mux_2173_nl, mux_2167_nl, or_2487_cse);
  or_2450_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2158_nl <= MUX_s_1_2_2(or_2450_nl, or_2396_cse, fsm_output(5));
  mux_2175_itm <= MUX_s_1_2_2(mux_2174_nl, mux_2158_nl, fsm_output(7));
  or_2487_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1619_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2211_nl <= MUX_s_1_2_2(mux_1877_cse, and_1619_nl, or_2487_cse);
  mux_2212_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2211_nl, nor_636_cse);
  mux_2213_seb <= MUX_s_1_2_2(mux_2212_nl, mux_2152_cse, fsm_output(5));
  nor_1665_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_2227_nl <= MUX_s_1_2_2(nor_1665_nl, (fsm_output(2)), fsm_output(0));
  mux_2228_nl <= MUX_s_1_2_2((NOT mux_2227_nl), or_4378_cse, fsm_output(1));
  mux_2229_nl <= MUX_s_1_2_2(mux_2228_nl, or_4699_cse, fsm_output(3));
  or_2516_nl <= (fsm_output(6)) OR mux_2229_nl;
  mux_2226_nl <= MUX_s_1_2_2(mux_tmp_2222, or_4699_cse, fsm_output(3));
  nand_128_nl <= NOT((fsm_output(6)) AND (NOT mux_2226_nl));
  mux_2230_nl <= MUX_s_1_2_2(or_2516_nl, nand_128_nl, fsm_output(4));
  mux_2231_nl <= MUX_s_1_2_2(mux_2230_nl, mux_tmp_2219, fsm_output(5));
  or_2512_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_2220_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2265, fsm_output(0));
  nor_724_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00111")));
  mux_2221_nl <= MUX_s_1_2_2(or_tmp_2266, mux_2220_nl, nor_724_nl);
  or_2509_nl <= (fsm_output(1)) OR mux_2221_nl;
  mux_2223_nl <= MUX_s_1_2_2(mux_tmp_2222, or_2509_nl, fsm_output(3));
  nand_127_nl <= NOT((fsm_output(6)) AND (NOT mux_2223_nl));
  mux_2224_nl <= MUX_s_1_2_2(or_2512_nl, nand_127_nl, fsm_output(4));
  mux_2225_nl <= MUX_s_1_2_2(mux_2224_nl, mux_tmp_2219, fsm_output(5));
  mux_2232_nl <= MUX_s_1_2_2(mux_2231_nl, mux_2225_nl, or_2528_cse);
  or_2497_nl <= (fsm_output(0)) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2214_nl <= MUX_s_1_2_2(or_tmp_2259, or_2497_nl, fsm_output(1));
  or_4516_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_2214_nl;
  mux_2215_nl <= MUX_s_1_2_2(or_4516_nl, or_2396_cse, fsm_output(5));
  mux_2233_itm <= MUX_s_1_2_2(mux_2232_nl, mux_2215_nl, fsm_output(7));
  or_2528_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0111"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1605_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2269_nl <= MUX_s_1_2_2(mux_1877_cse, and_1605_nl, or_2528_cse);
  mux_2270_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2269_nl, nor_636_cse);
  mux_2271_seb <= MUX_s_1_2_2(mux_2270_nl, mux_2152_cse, fsm_output(5));
  or_2557_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2290_nl <= MUX_s_1_2_2(or_2557_nl, or_2158_cse, fsm_output(1));
  mux_2291_nl <= MUX_s_1_2_2(mux_2290_nl, or_2157_cse, fsm_output(0));
  or_2558_nl <= (fsm_output(6)) OR mux_2291_nl;
  mux_2292_nl <= MUX_s_1_2_2(or_2161_cse, or_2558_nl, fsm_output(2));
  mux_2289_nl <= MUX_s_1_2_2(or_tmp_2310, mux_tmp_2284, fsm_output(6));
  or_2554_nl <= (fsm_output(2)) OR mux_2289_nl;
  mux_2293_nl <= MUX_s_1_2_2(mux_2292_nl, or_2554_nl, fsm_output(4));
  or_2553_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2549_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01000"));
  mux_2285_nl <= MUX_s_1_2_2(mux_tmp_2284, or_tmp_2300, or_2549_nl);
  or_2548_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2283_nl <= MUX_s_1_2_2(or_2548_nl, or_tmp_2306, fsm_output(1));
  mux_2286_nl <= MUX_s_1_2_2(mux_2285_nl, mux_2283_nl, fsm_output(0));
  mux_2287_nl <= MUX_s_1_2_2(or_tmp_2310, mux_2286_nl, fsm_output(6));
  or_2552_nl <= (fsm_output(2)) OR mux_2287_nl;
  mux_2288_nl <= MUX_s_1_2_2(or_2553_nl, or_2552_nl, fsm_output(4));
  mux_2294_nl <= MUX_s_1_2_2(mux_2293_nl, mux_2288_nl, or_2577_cse);
  or_2544_nl <= (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2276_nl <= MUX_s_1_2_2(or_2544_nl, (fsm_output(7)), fsm_output(3));
  mux_2277_nl <= MUX_s_1_2_2(or_2147_cse, mux_2276_nl, fsm_output(1));
  mux_2278_nl <= MUX_s_1_2_2(mux_2277_nl, mux_tmp_2273, fsm_output(0));
  mux_2279_nl <= MUX_s_1_2_2(mux_2278_nl, mux_tmp_2272, fsm_output(6));
  mux_2280_nl <= MUX_s_1_2_2(mux_2279_nl, nand_331_cse, fsm_output(2));
  mux_2274_nl <= MUX_s_1_2_2(or_tmp_2300, mux_tmp_2273, fsm_output(0));
  mux_2275_nl <= MUX_s_1_2_2(mux_2274_nl, mux_tmp_2272, fsm_output(6));
  or_2542_nl <= (fsm_output(2)) OR mux_2275_nl;
  mux_2281_nl <= MUX_s_1_2_2(mux_2280_nl, or_2542_nl, or_2574_cse);
  or_2535_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2282_nl <= MUX_s_1_2_2(mux_2281_nl, or_2535_nl, fsm_output(4));
  mux_2295_itm <= MUX_s_1_2_2(mux_2294_nl, mux_2282_nl, fsm_output(5));
  or_2574_cse <= CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("010"));
  or_2577_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1595_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01000"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2326_nl <= MUX_s_1_2_2(mux_1877_cse, and_1595_nl, or_2577_cse);
  mux_2327_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2326_nl, nor_636_cse);
  or_2576_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2321_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2576_nl);
  mux_2322_nl <= MUX_s_1_2_2(mux_2321_nl, mux_1872_cse, fsm_output(3));
  mux_2317_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_2574_cse);
  mux_2318_nl <= MUX_s_1_2_2(mux_2317_nl, mux_1865_cse, fsm_output(4));
  mux_2319_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2318_nl, fsm_output(3));
  mux_2323_nl <= MUX_s_1_2_2(mux_2322_nl, mux_2319_nl, fsm_output(1));
  mux_2328_seb <= MUX_s_1_2_2(mux_2327_nl, mux_2323_nl, fsm_output(5));
  nor_1650_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_2344_nl <= MUX_s_1_2_2(nor_1650_nl, (fsm_output(2)), fsm_output(0));
  mux_2345_nl <= MUX_s_1_2_2((NOT mux_2344_nl), (fsm_output(2)), fsm_output(3));
  mux_2346_nl <= MUX_s_1_2_2(mux_2345_nl, or_2215_cse, fsm_output(1));
  or_2603_nl <= (fsm_output(4)) OR mux_2346_nl;
  mux_2342_nl <= MUX_s_1_2_2(or_tmp_2355, (fsm_output(2)), fsm_output(3));
  mux_2343_nl <= MUX_s_1_2_2(mux_2342_nl, or_tmp_2353, fsm_output(1));
  nand_132_nl <= NOT((fsm_output(4)) AND (NOT mux_2343_nl));
  mux_2347_nl <= MUX_s_1_2_2(or_2603_nl, nand_132_nl, fsm_output(6));
  mux_2348_nl <= MUX_s_1_2_2(mux_2347_nl, mux_tmp_2335, fsm_output(5));
  or_2599_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2597_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2336_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2348, fsm_output(0));
  nor_756_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01001")));
  mux_2337_nl <= MUX_s_1_2_2(or_2597_nl, mux_2336_nl, nor_756_nl);
  mux_2338_nl <= MUX_s_1_2_2(or_tmp_2355, mux_2337_nl, fsm_output(3));
  mux_2339_nl <= MUX_s_1_2_2(mux_2338_nl, or_tmp_2353, fsm_output(1));
  nand_131_nl <= NOT((fsm_output(4)) AND (NOT mux_2339_nl));
  mux_2340_nl <= MUX_s_1_2_2(or_2599_nl, nand_131_nl, fsm_output(6));
  mux_2341_nl <= MUX_s_1_2_2(mux_2340_nl, mux_tmp_2335, fsm_output(5));
  mux_2349_nl <= MUX_s_1_2_2(mux_2348_nl, mux_2341_nl, or_2622_cse);
  nor_1651_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  nor_1652_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  mux_2329_nl <= MUX_s_1_2_2(nor_1651_nl, nor_1652_nl, fsm_output(1));
  nand_129_nl <= NOT(nor_2197_cse AND mux_2329_nl);
  mux_2330_nl <= MUX_s_1_2_2(nand_129_nl, or_2585_cse, fsm_output(5));
  mux_2350_itm <= MUX_s_1_2_2(mux_2349_nl, mux_2330_nl, fsm_output(7));
  or_2619_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_2622_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_2621_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2370_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2621_nl);
  mux_2371_nl <= MUX_s_1_2_2(mux_2370_nl, mux_1872_cse, fsm_output(3));
  mux_2366_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_2619_cse);
  mux_2367_nl <= MUX_s_1_2_2(mux_2366_nl, mux_1865_cse, fsm_output(4));
  mux_2368_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2367_nl, fsm_output(3));
  mux_2372_cse <= MUX_s_1_2_2(mux_2371_nl, mux_2368_nl, fsm_output(1));
  and_1589_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2375_nl <= MUX_s_1_2_2(mux_1877_cse, and_1589_nl, or_2622_cse);
  mux_2376_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2375_nl, nor_636_cse);
  mux_2377_seb <= MUX_s_1_2_2(mux_2376_nl, mux_2372_cse, fsm_output(5));
  or_2650_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2389_nl <= MUX_s_1_2_2(or_2650_nl, or_2273_cse, fsm_output(0));
  mux_2390_nl <= MUX_s_1_2_2(mux_2389_nl, or_2272_cse, fsm_output(3));
  mux_2391_nl <= MUX_s_1_2_2(mux_2390_nl, or_2271_cse, fsm_output(1));
  mux_2388_nl <= MUX_s_1_2_2(or_tmp_2398, or_119_cse, fsm_output(3));
  or_2646_nl <= (fsm_output(1)) OR mux_2388_nl;
  mux_2392_nl <= MUX_s_1_2_2(mux_2391_nl, or_2646_nl, fsm_output(6));
  mux_2393_nl <= MUX_s_1_2_2(mux_2392_nl, mux_tmp_2383, fsm_output(5));
  or_2644_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2641_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_2639_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2384_nl <= MUX_s_1_2_2(or_2641_nl, or_2639_nl, fsm_output(0));
  mux_2385_nl <= MUX_s_1_2_2(or_tmp_2398, mux_2384_nl, fsm_output(3));
  or_2643_nl <= (fsm_output(1)) OR mux_2385_nl;
  mux_2386_nl <= MUX_s_1_2_2(or_2644_nl, or_2643_nl, fsm_output(6));
  mux_2387_nl <= MUX_s_1_2_2(mux_2386_nl, mux_tmp_2383, fsm_output(5));
  mux_2394_nl <= MUX_s_1_2_2(mux_2393_nl, mux_2387_nl, or_2664_cse);
  or_2630_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2378_nl <= MUX_s_1_2_2(or_2630_nl, or_2585_cse, fsm_output(5));
  mux_2395_itm <= MUX_s_1_2_2(mux_2394_nl, mux_2378_nl, fsm_output(7));
  or_2664_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1578_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2431_nl <= MUX_s_1_2_2(mux_1877_cse, and_1578_nl, or_2664_cse);
  mux_2432_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2431_nl, nor_636_cse);
  mux_2433_seb <= MUX_s_1_2_2(mux_2432_nl, mux_2372_cse, fsm_output(5));
  nor_1632_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_2447_nl <= MUX_s_1_2_2(nor_1632_nl, (fsm_output(2)), fsm_output(0));
  mux_2448_nl <= MUX_s_1_2_2((NOT mux_2447_nl), or_4378_cse, fsm_output(1));
  mux_2449_nl <= MUX_s_1_2_2(mux_2448_nl, or_4699_cse, fsm_output(3));
  or_2686_nl <= (fsm_output(6)) OR mux_2449_nl;
  mux_2446_nl <= MUX_s_1_2_2(mux_tmp_2442, or_4699_cse, fsm_output(3));
  nand_137_nl <= NOT((fsm_output(6)) AND (NOT mux_2446_nl));
  mux_2450_nl <= MUX_s_1_2_2(or_2686_nl, nand_137_nl, fsm_output(4));
  mux_2451_nl <= MUX_s_1_2_2(mux_2450_nl, mux_tmp_2439, fsm_output(5));
  or_2682_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_2440_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2432, fsm_output(0));
  nor_780_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01011")));
  mux_2441_nl <= MUX_s_1_2_2(or_tmp_2433, mux_2440_nl, nor_780_nl);
  or_2680_nl <= (fsm_output(1)) OR mux_2441_nl;
  mux_2443_nl <= MUX_s_1_2_2(mux_tmp_2442, or_2680_nl, fsm_output(3));
  nand_136_nl <= NOT((fsm_output(6)) AND (NOT mux_2443_nl));
  mux_2444_nl <= MUX_s_1_2_2(or_2682_nl, nand_136_nl, fsm_output(4));
  mux_2445_nl <= MUX_s_1_2_2(mux_2444_nl, mux_tmp_2439, fsm_output(5));
  mux_2452_nl <= MUX_s_1_2_2(mux_2451_nl, mux_2445_nl, or_2700_cse);
  or_2672_nl <= (fsm_output(0)) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2434_nl <= MUX_s_1_2_2(or_tmp_2428, or_2672_nl, fsm_output(1));
  or_4495_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_2434_nl;
  mux_2435_nl <= MUX_s_1_2_2(or_4495_nl, or_2585_cse, fsm_output(5));
  mux_2453_itm <= MUX_s_1_2_2(mux_2452_nl, mux_2435_nl, fsm_output(7));
  or_2700_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1564_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2489_nl <= MUX_s_1_2_2(mux_1877_cse, and_1564_nl, or_2700_cse);
  mux_2490_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2489_nl, nor_636_cse);
  mux_2491_seb <= MUX_s_1_2_2(mux_2490_nl, mux_2372_cse, fsm_output(5));
  or_2728_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2510_nl <= MUX_s_1_2_2(or_2728_nl, or_2158_cse, fsm_output(1));
  mux_2511_nl <= MUX_s_1_2_2(mux_2510_nl, or_2157_cse, fsm_output(0));
  or_2729_nl <= (fsm_output(6)) OR mux_2511_nl;
  mux_2512_nl <= MUX_s_1_2_2(or_2161_cse, or_2729_nl, fsm_output(2));
  mux_2509_nl <= MUX_s_1_2_2(or_tmp_2476, mux_tmp_2504, fsm_output(6));
  or_2725_nl <= (fsm_output(2)) OR mux_2509_nl;
  mux_2513_nl <= MUX_s_1_2_2(mux_2512_nl, or_2725_nl, fsm_output(4));
  or_2724_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2720_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01100"));
  mux_2505_nl <= MUX_s_1_2_2(mux_tmp_2504, or_tmp_2469, or_2720_nl);
  or_2719_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2503_nl <= MUX_s_1_2_2(or_2719_nl, or_tmp_2472, fsm_output(1));
  mux_2506_nl <= MUX_s_1_2_2(mux_2505_nl, mux_2503_nl, fsm_output(0));
  mux_2507_nl <= MUX_s_1_2_2(or_tmp_2476, mux_2506_nl, fsm_output(6));
  or_2723_nl <= (fsm_output(2)) OR mux_2507_nl;
  mux_2508_nl <= MUX_s_1_2_2(or_2724_nl, or_2723_nl, fsm_output(4));
  mux_2514_nl <= MUX_s_1_2_2(mux_2513_nl, mux_2508_nl, or_2747_cse);
  mux_2499_nl <= MUX_s_1_2_2(or_tmp_2469, mux_tmp_2493, fsm_output(0));
  mux_2500_nl <= MUX_s_1_2_2(mux_2499_nl, mux_tmp_2492, fsm_output(6));
  or_2716_nl <= (fsm_output(2)) OR mux_2500_nl;
  or_2713_nl <= (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  mux_2494_nl <= MUX_s_1_2_2(or_2713_nl, (fsm_output(7)), fsm_output(3));
  mux_2495_nl <= MUX_s_1_2_2(or_2147_cse, mux_2494_nl, fsm_output(1));
  mux_2496_nl <= MUX_s_1_2_2(mux_2495_nl, mux_tmp_2493, fsm_output(0));
  mux_2497_nl <= MUX_s_1_2_2(mux_2496_nl, mux_tmp_2492, fsm_output(6));
  mux_2498_nl <= MUX_s_1_2_2(mux_2497_nl, nand_331_cse, fsm_output(2));
  mux_2501_nl <= MUX_s_1_2_2(or_2716_nl, mux_2498_nl, nor_805_cse);
  or_2707_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  mux_2502_nl <= MUX_s_1_2_2(mux_2501_nl, or_2707_nl, fsm_output(4));
  mux_2515_itm <= MUX_s_1_2_2(mux_2514_nl, mux_2502_nl, fsm_output(5));
  nor_805_cse <= NOT(CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("011")));
  or_2747_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1554_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01100"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2546_nl <= MUX_s_1_2_2(mux_1877_cse, and_1554_nl, or_2747_cse);
  mux_2547_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2546_nl, nor_636_cse);
  or_2746_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2541_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2746_nl);
  mux_2542_nl <= MUX_s_1_2_2(mux_2541_nl, mux_1872_cse, fsm_output(3));
  mux_2537_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, nor_805_cse);
  mux_2538_nl <= MUX_s_1_2_2(mux_2537_nl, mux_1865_cse, fsm_output(4));
  mux_2539_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2538_nl, fsm_output(3));
  mux_2543_nl <= MUX_s_1_2_2(mux_2542_nl, mux_2539_nl, fsm_output(1));
  mux_2548_seb <= MUX_s_1_2_2(mux_2547_nl, mux_2543_nl, fsm_output(5));
  or_2756_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  nor_1617_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  mux_2564_nl <= MUX_s_1_2_2(nor_1617_nl, (fsm_output(2)), fsm_output(0));
  mux_2565_nl <= MUX_s_1_2_2((NOT mux_2564_nl), (fsm_output(2)), fsm_output(3));
  mux_2566_nl <= MUX_s_1_2_2(mux_2565_nl, or_2215_cse, fsm_output(1));
  or_2782_nl <= (fsm_output(4)) OR mux_2566_nl;
  mux_2562_nl <= MUX_s_1_2_2(or_tmp_2529, (fsm_output(2)), fsm_output(3));
  mux_2563_nl <= MUX_s_1_2_2(mux_2562_nl, or_tmp_2526, fsm_output(1));
  nand_141_nl <= NOT((fsm_output(4)) AND (NOT mux_2563_nl));
  mux_2567_nl <= MUX_s_1_2_2(or_2782_nl, nand_141_nl, fsm_output(6));
  mux_2568_nl <= MUX_s_1_2_2(mux_2567_nl, mux_tmp_2555, fsm_output(5));
  or_2778_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2775_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2556_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2518, fsm_output(0));
  nor_813_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01101")));
  mux_2557_nl <= MUX_s_1_2_2(or_2775_nl, mux_2556_nl, nor_813_nl);
  mux_2558_nl <= MUX_s_1_2_2(or_tmp_2529, mux_2557_nl, fsm_output(3));
  mux_2559_nl <= MUX_s_1_2_2(mux_2558_nl, or_tmp_2526, fsm_output(1));
  nand_140_nl <= NOT((fsm_output(4)) AND (NOT mux_2559_nl));
  mux_2560_nl <= MUX_s_1_2_2(or_2778_nl, nand_140_nl, fsm_output(6));
  mux_2561_nl <= MUX_s_1_2_2(mux_2560_nl, mux_tmp_2555, fsm_output(5));
  mux_2569_nl <= MUX_s_1_2_2(mux_2568_nl, mux_2561_nl, or_2800_cse);
  nor_1618_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389);
  nor_1619_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389);
  mux_2549_nl <= MUX_s_1_2_2(nor_1618_nl, nor_1619_nl, fsm_output(1));
  nand_138_nl <= NOT(nor_2197_cse AND mux_2549_nl);
  mux_2550_nl <= MUX_s_1_2_2(nand_138_nl, or_2756_cse, fsm_output(5));
  mux_2570_itm <= MUX_s_1_2_2(mux_2569_nl, mux_2550_nl, fsm_output(7));
  nor_817_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011")));
  or_2800_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_2799_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2590_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2799_nl);
  mux_2591_nl <= MUX_s_1_2_2(mux_2590_nl, mux_1872_cse, fsm_output(3));
  mux_2586_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, nor_817_cse);
  mux_2587_nl <= MUX_s_1_2_2(mux_2586_nl, mux_1865_cse, fsm_output(4));
  mux_2588_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2587_nl, fsm_output(3));
  mux_2592_cse <= MUX_s_1_2_2(mux_2591_nl, mux_2588_nl, fsm_output(1));
  and_1547_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2595_nl <= MUX_s_1_2_2(mux_1877_cse, and_1547_nl, or_2800_cse);
  mux_2596_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2595_nl, nor_636_cse);
  mux_2597_seb <= MUX_s_1_2_2(mux_2596_nl, mux_2592_cse, fsm_output(5));
  or_2835_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2609_nl <= MUX_s_1_2_2(or_2835_nl, or_2273_cse, fsm_output(0));
  mux_2610_nl <= MUX_s_1_2_2(mux_2609_nl, or_2272_cse, fsm_output(3));
  mux_2611_nl <= MUX_s_1_2_2(mux_2610_nl, or_2271_cse, fsm_output(1));
  mux_2608_nl <= MUX_s_1_2_2(or_tmp_2578, or_119_cse, fsm_output(3));
  or_2831_nl <= (fsm_output(1)) OR mux_2608_nl;
  mux_2612_nl <= MUX_s_1_2_2(mux_2611_nl, or_2831_nl, fsm_output(6));
  mux_2613_nl <= MUX_s_1_2_2(mux_2612_nl, mux_tmp_2603, fsm_output(5));
  or_2829_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110")) OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2825_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_2823_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2604_nl <= MUX_s_1_2_2(or_2825_nl, or_2823_nl, fsm_output(0));
  mux_2605_nl <= MUX_s_1_2_2(or_tmp_2578, mux_2604_nl, fsm_output(3));
  or_2828_nl <= (fsm_output(1)) OR mux_2605_nl;
  mux_2606_nl <= MUX_s_1_2_2(or_2829_nl, or_2828_nl, fsm_output(6));
  mux_2607_nl <= MUX_s_1_2_2(mux_2606_nl, mux_tmp_2603, fsm_output(5));
  mux_2614_nl <= MUX_s_1_2_2(mux_2613_nl, mux_2607_nl, or_2847_cse);
  or_2810_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  mux_2598_nl <= MUX_s_1_2_2(or_2810_nl, or_2756_cse, fsm_output(5));
  mux_2615_itm <= MUX_s_1_2_2(mux_2614_nl, mux_2598_nl, fsm_output(7));
  or_2847_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1534_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2651_nl <= MUX_s_1_2_2(mux_1877_cse, and_1534_nl, or_2847_cse);
  mux_2652_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2651_nl, nor_636_cse);
  mux_2653_seb <= MUX_s_1_2_2(mux_2652_nl, mux_2592_cse, fsm_output(5));
  and_1531_nl <= (fsm_output(2)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2667_nl <= MUX_s_1_2_2(and_1531_nl, (fsm_output(2)), fsm_output(0));
  mux_2668_nl <= MUX_s_1_2_2((NOT mux_2667_nl), or_4378_cse, fsm_output(1));
  mux_2669_nl <= MUX_s_1_2_2(mux_2668_nl, or_4699_cse, fsm_output(3));
  or_2876_nl <= (fsm_output(6)) OR mux_2669_nl;
  mux_2666_nl <= MUX_s_1_2_2(mux_tmp_2662, or_4699_cse, fsm_output(3));
  nand_146_nl <= NOT((fsm_output(6)) AND (NOT mux_2666_nl));
  mux_2670_nl <= MUX_s_1_2_2(or_2876_nl, nand_146_nl, fsm_output(4));
  mux_2671_nl <= MUX_s_1_2_2(mux_2670_nl, mux_tmp_2659, fsm_output(5));
  or_2872_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1111")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_2660_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2615, fsm_output(0));
  mux_2661_nl <= MUX_s_1_2_2(or_tmp_2616, mux_2660_nl, and_1532_cse);
  or_2869_nl <= (fsm_output(1)) OR mux_2661_nl;
  mux_2663_nl <= MUX_s_1_2_2(mux_tmp_2662, or_2869_nl, fsm_output(3));
  nand_145_nl <= NOT((fsm_output(6)) AND (NOT mux_2663_nl));
  mux_2664_nl <= MUX_s_1_2_2(or_2872_nl, nand_145_nl, fsm_output(4));
  mux_2665_nl <= MUX_s_1_2_2(mux_2664_nl, mux_tmp_2659, fsm_output(5));
  mux_2672_nl <= MUX_s_1_2_2(mux_2671_nl, mux_2665_nl, nand_317_cse);
  or_2857_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  mux_2654_nl <= MUX_s_1_2_2(or_tmp_2609, or_2857_nl, fsm_output(1));
  or_4474_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_2654_nl;
  mux_2655_nl <= MUX_s_1_2_2(or_4474_nl, or_2756_cse, fsm_output(5));
  mux_2673_itm <= MUX_s_1_2_2(mux_2672_nl, mux_2655_nl, fsm_output(7));
  nand_317_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1518_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("01111"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2709_nl <= MUX_s_1_2_2(mux_1877_cse, and_1518_nl, nand_317_cse);
  mux_2710_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2709_nl, nor_636_cse);
  mux_2711_seb <= MUX_s_1_2_2(mux_2710_nl, mux_2592_cse, fsm_output(5));
  or_2930_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_2927_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10000"));
  mux_2730_nl <= MUX_s_1_2_2(mux_tmp_2723, or_tmp_2656, or_2927_nl);
  or_2926_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2729_nl <= MUX_s_1_2_2(or_2926_nl, or_tmp_2663, fsm_output(1));
  mux_2731_nl <= MUX_s_1_2_2(mux_2730_nl, mux_2729_nl, fsm_output(0));
  mux_2732_nl <= MUX_s_1_2_2(or_tmp_2666, mux_2731_nl, fsm_output(6));
  or_2928_nl <= (fsm_output(2)) OR mux_2732_nl;
  mux_2733_nl <= MUX_s_1_2_2(or_2930_nl, or_2928_nl, fsm_output(4));
  or_2922_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2725_nl <= MUX_s_1_2_2(or_2922_nl, or_2158_cse, fsm_output(1));
  mux_2726_nl <= MUX_s_1_2_2(mux_2725_nl, or_2157_cse, fsm_output(0));
  or_2923_nl <= (fsm_output(6)) OR mux_2726_nl;
  mux_2727_nl <= MUX_s_1_2_2(or_2161_cse, or_2923_nl, fsm_output(2));
  mux_2724_nl <= MUX_s_1_2_2(or_tmp_2666, mux_tmp_2723, fsm_output(6));
  or_2918_nl <= (fsm_output(2)) OR mux_2724_nl;
  mux_2728_nl <= MUX_s_1_2_2(mux_2727_nl, or_2918_nl, fsm_output(4));
  mux_2734_nl <= MUX_s_1_2_2(mux_2733_nl, mux_2728_nl, nor_873_cse);
  or_2911_nl <= (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2716_nl <= MUX_s_1_2_2(or_2911_nl, (fsm_output(7)), fsm_output(3));
  mux_2717_nl <= MUX_s_1_2_2(or_2147_cse, mux_2716_nl, fsm_output(1));
  mux_2718_nl <= MUX_s_1_2_2(mux_2717_nl, mux_tmp_2713, fsm_output(0));
  mux_2719_nl <= MUX_s_1_2_2(mux_2718_nl, mux_tmp_2712, fsm_output(6));
  mux_2720_nl <= MUX_s_1_2_2(mux_2719_nl, nand_331_cse, fsm_output(2));
  mux_2714_nl <= MUX_s_1_2_2(or_tmp_2656, mux_tmp_2713, fsm_output(0));
  mux_2715_nl <= MUX_s_1_2_2(mux_2714_nl, mux_tmp_2712, fsm_output(6));
  or_2908_nl <= (fsm_output(2)) OR mux_2715_nl;
  mux_2721_nl <= MUX_s_1_2_2(mux_2720_nl, or_2908_nl, or_2947_cse);
  or_2896_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2722_nl <= MUX_s_1_2_2(mux_2721_nl, or_2896_nl, fsm_output(4));
  mux_2735_itm <= MUX_s_1_2_2(mux_2734_nl, mux_2722_nl, fsm_output(5));
  or_2947_cse <= CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("100"));
  nor_873_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1507_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10000"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2766_nl <= MUX_s_1_2_2(and_1507_nl, mux_1877_cse, nor_873_cse);
  mux_2767_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2766_nl, nor_636_cse);
  or_2949_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2761_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_2949_nl);
  mux_2762_nl <= MUX_s_1_2_2(mux_2761_nl, mux_1872_cse, fsm_output(3));
  mux_2757_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_2947_cse);
  mux_2758_nl <= MUX_s_1_2_2(mux_2757_nl, mux_1865_cse, fsm_output(4));
  mux_2759_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2758_nl, fsm_output(3));
  mux_2763_nl <= MUX_s_1_2_2(mux_2762_nl, mux_2759_nl, fsm_output(1));
  mux_2768_seb <= MUX_s_1_2_2(mux_2767_nl, mux_2763_nl, fsm_output(5));
  or_2980_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  or_2978_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2783_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2710, fsm_output(0));
  nor_878_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10001")));
  mux_2784_nl <= MUX_s_1_2_2(or_2978_nl, mux_2783_nl, nor_878_nl);
  mux_2785_nl <= MUX_s_1_2_2(or_tmp_2717, mux_2784_nl, fsm_output(3));
  mux_2786_nl <= MUX_s_1_2_2(mux_2785_nl, or_tmp_2716, fsm_output(1));
  nand_150_nl <= NOT((fsm_output(4)) AND (NOT mux_2786_nl));
  mux_2787_nl <= MUX_s_1_2_2(or_2980_nl, nand_150_nl, fsm_output(6));
  mux_2788_nl <= MUX_s_1_2_2(mux_2787_nl, mux_tmp_2775, fsm_output(5));
  nor_1587_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_2778_nl <= MUX_s_1_2_2(nor_1587_nl, (fsm_output(2)), fsm_output(0));
  mux_2779_nl <= MUX_s_1_2_2((NOT mux_2778_nl), (fsm_output(2)), fsm_output(3));
  mux_2780_nl <= MUX_s_1_2_2(mux_2779_nl, or_2215_cse, fsm_output(1));
  or_2976_nl <= (fsm_output(4)) OR mux_2780_nl;
  mux_2776_nl <= MUX_s_1_2_2(or_tmp_2717, (fsm_output(2)), fsm_output(3));
  mux_2777_nl <= MUX_s_1_2_2(mux_2776_nl, or_tmp_2716, fsm_output(1));
  nand_149_nl <= NOT((fsm_output(4)) AND (NOT mux_2777_nl));
  mux_2781_nl <= MUX_s_1_2_2(or_2976_nl, nand_149_nl, fsm_output(6));
  mux_2782_nl <= MUX_s_1_2_2(mux_2781_nl, mux_tmp_2775, fsm_output(5));
  mux_2789_nl <= MUX_s_1_2_2(mux_2788_nl, mux_2782_nl, nor_885_cse);
  nor_1588_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  nor_1589_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  mux_2769_nl <= MUX_s_1_2_2(nor_1588_nl, nor_1589_nl, fsm_output(1));
  nand_147_nl <= NOT(nor_2197_cse AND mux_2769_nl);
  mux_2770_nl <= MUX_s_1_2_2(nand_147_nl, or_2958_cse, fsm_output(5));
  mux_2790_itm <= MUX_s_1_2_2(mux_2789_nl, mux_2770_nl, fsm_output(7));
  or_2999_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  nor_885_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  or_3001_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2810_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3001_nl);
  mux_2811_nl <= MUX_s_1_2_2(mux_2810_nl, mux_1872_cse, fsm_output(3));
  mux_2806_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_2999_cse);
  mux_2807_nl <= MUX_s_1_2_2(mux_2806_nl, mux_1865_cse, fsm_output(4));
  mux_2808_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2807_nl, fsm_output(3));
  mux_2812_cse <= MUX_s_1_2_2(mux_2811_nl, mux_2808_nl, fsm_output(1));
  and_1501_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2815_nl <= MUX_s_1_2_2(and_1501_nl, mux_1877_cse, nor_885_cse);
  mux_2816_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2815_nl, nor_636_cse);
  mux_2817_seb <= MUX_s_1_2_2(mux_2816_nl, mux_2812_cse, fsm_output(5));
  or_3033_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  or_3030_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_3028_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2830_nl <= MUX_s_1_2_2(or_3030_nl, or_3028_nl, fsm_output(0));
  mux_2831_nl <= MUX_s_1_2_2(or_tmp_2765, mux_2830_nl, fsm_output(3));
  or_3031_nl <= (fsm_output(1)) OR mux_2831_nl;
  mux_2832_nl <= MUX_s_1_2_2(or_3033_nl, or_3031_nl, fsm_output(6));
  mux_2833_nl <= MUX_s_1_2_2(mux_2832_nl, mux_tmp_2823, fsm_output(5));
  or_3026_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2825_nl <= MUX_s_1_2_2(or_3026_nl, or_2273_cse, fsm_output(0));
  mux_2826_nl <= MUX_s_1_2_2(mux_2825_nl, or_2272_cse, fsm_output(3));
  mux_2827_nl <= MUX_s_1_2_2(mux_2826_nl, or_2271_cse, fsm_output(1));
  mux_2824_nl <= MUX_s_1_2_2(or_tmp_2765, or_119_cse, fsm_output(3));
  or_3021_nl <= (fsm_output(1)) OR mux_2824_nl;
  mux_2828_nl <= MUX_s_1_2_2(mux_2827_nl, or_3021_nl, fsm_output(6));
  mux_2829_nl <= MUX_s_1_2_2(mux_2828_nl, mux_tmp_2823, fsm_output(5));
  mux_2834_nl <= MUX_s_1_2_2(mux_2833_nl, mux_2829_nl, nor_901_cse);
  or_3009_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2818_nl <= MUX_s_1_2_2(or_3009_nl, or_2958_cse, fsm_output(5));
  mux_2835_itm <= MUX_s_1_2_2(mux_2834_nl, mux_2818_nl, fsm_output(7));
  nor_901_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1490_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2871_nl <= MUX_s_1_2_2(and_1490_nl, mux_1877_cse, nor_901_cse);
  mux_2872_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2871_nl, nor_636_cse);
  mux_2873_seb <= MUX_s_1_2_2(mux_2872_nl, mux_2812_cse, fsm_output(5));
  or_3074_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2887_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2806, fsm_output(0));
  nor_906_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10011")));
  mux_2888_nl <= MUX_s_1_2_2(or_tmp_2808, mux_2887_nl, nor_906_nl);
  or_3072_nl <= (fsm_output(1)) OR mux_2888_nl;
  mux_2889_nl <= MUX_s_1_2_2(mux_tmp_2880, or_3072_nl, fsm_output(3));
  nand_155_nl <= NOT((fsm_output(6)) AND (NOT mux_2889_nl));
  mux_2890_nl <= MUX_s_1_2_2(or_3074_nl, nand_155_nl, fsm_output(4));
  mux_2891_nl <= MUX_s_1_2_2(mux_2890_nl, mux_tmp_2879, fsm_output(5));
  nor_1569_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_2882_nl <= MUX_s_1_2_2(nor_1569_nl, (fsm_output(2)), fsm_output(0));
  mux_2883_nl <= MUX_s_1_2_2((NOT mux_2882_nl), or_4378_cse, fsm_output(1));
  mux_2884_nl <= MUX_s_1_2_2(mux_2883_nl, or_4699_cse, fsm_output(3));
  or_3071_nl <= (fsm_output(6)) OR mux_2884_nl;
  mux_2881_nl <= MUX_s_1_2_2(mux_tmp_2880, or_4699_cse, fsm_output(3));
  nand_154_nl <= NOT((fsm_output(6)) AND (NOT mux_2881_nl));
  mux_2885_nl <= MUX_s_1_2_2(or_3071_nl, nand_154_nl, fsm_output(4));
  mux_2886_nl <= MUX_s_1_2_2(mux_2885_nl, mux_tmp_2879, fsm_output(5));
  mux_2892_nl <= MUX_s_1_2_2(mux_2891_nl, mux_2886_nl, nor_920_cse);
  or_3057_nl <= (fsm_output(0)) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2874_nl <= MUX_s_1_2_2(or_tmp_2802, or_3057_nl, fsm_output(1));
  or_4453_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_2874_nl;
  mux_2875_nl <= MUX_s_1_2_2(or_4453_nl, or_2958_cse, fsm_output(5));
  mux_2893_itm <= MUX_s_1_2_2(mux_2892_nl, mux_2875_nl, fsm_output(7));
  nor_920_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1477_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2929_nl <= MUX_s_1_2_2(and_1477_nl, mux_1877_cse, nor_920_cse);
  mux_2930_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2929_nl, nor_636_cse);
  mux_2931_seb <= MUX_s_1_2_2(mux_2930_nl, mux_2812_cse, fsm_output(5));
  or_3131_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_3128_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10100"));
  mux_2950_nl <= MUX_s_1_2_2(mux_tmp_2943, or_tmp_2855, or_3128_nl);
  or_3127_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2949_nl <= MUX_s_1_2_2(or_3127_nl, or_tmp_2858, fsm_output(1));
  mux_2951_nl <= MUX_s_1_2_2(mux_2950_nl, mux_2949_nl, fsm_output(0));
  mux_2952_nl <= MUX_s_1_2_2(or_tmp_2861, mux_2951_nl, fsm_output(6));
  or_3129_nl <= (fsm_output(2)) OR mux_2952_nl;
  mux_2953_nl <= MUX_s_1_2_2(or_3131_nl, or_3129_nl, fsm_output(4));
  or_3123_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2945_nl <= MUX_s_1_2_2(or_3123_nl, or_2158_cse, fsm_output(1));
  mux_2946_nl <= MUX_s_1_2_2(mux_2945_nl, or_2157_cse, fsm_output(0));
  or_3124_nl <= (fsm_output(6)) OR mux_2946_nl;
  mux_2947_nl <= MUX_s_1_2_2(or_2161_cse, or_3124_nl, fsm_output(2));
  mux_2944_nl <= MUX_s_1_2_2(or_tmp_2861, mux_tmp_2943, fsm_output(6));
  or_3119_nl <= (fsm_output(2)) OR mux_2944_nl;
  mux_2948_nl <= MUX_s_1_2_2(mux_2947_nl, or_3119_nl, fsm_output(4));
  mux_2954_nl <= MUX_s_1_2_2(mux_2953_nl, mux_2948_nl, nor_938_cse);
  mux_2939_nl <= MUX_s_1_2_2(or_tmp_2855, mux_tmp_2933, fsm_output(0));
  mux_2940_nl <= MUX_s_1_2_2(mux_2939_nl, mux_tmp_2932, fsm_output(6));
  or_3113_nl <= (fsm_output(2)) OR mux_2940_nl;
  or_3109_nl <= (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  mux_2934_nl <= MUX_s_1_2_2(or_3109_nl, (fsm_output(7)), fsm_output(3));
  mux_2935_nl <= MUX_s_1_2_2(or_2147_cse, mux_2934_nl, fsm_output(1));
  mux_2936_nl <= MUX_s_1_2_2(mux_2935_nl, mux_tmp_2933, fsm_output(0));
  mux_2937_nl <= MUX_s_1_2_2(mux_2936_nl, mux_tmp_2932, fsm_output(6));
  mux_2938_nl <= MUX_s_1_2_2(mux_2937_nl, nand_331_cse, fsm_output(2));
  mux_2941_nl <= MUX_s_1_2_2(or_3113_nl, mux_2938_nl, nor_934_cse);
  or_3098_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  mux_2942_nl <= MUX_s_1_2_2(mux_2941_nl, or_3098_nl, fsm_output(4));
  mux_2955_itm <= MUX_s_1_2_2(mux_2954_nl, mux_2942_nl, fsm_output(5));
  nor_934_cse <= NOT(CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("101")));
  nor_938_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1467_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10100"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2986_nl <= MUX_s_1_2_2(and_1467_nl, mux_1877_cse, nor_938_cse);
  mux_2987_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2986_nl, nor_636_cse);
  or_3149_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_2981_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3149_nl);
  mux_2982_nl <= MUX_s_1_2_2(mux_2981_nl, mux_1872_cse, fsm_output(3));
  mux_2977_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, nor_934_cse);
  mux_2978_nl <= MUX_s_1_2_2(mux_2977_nl, mux_1865_cse, fsm_output(4));
  mux_2979_nl <= MUX_s_1_2_2(nor_tmp_35, mux_2978_nl, fsm_output(3));
  mux_2983_nl <= MUX_s_1_2_2(mux_2982_nl, mux_2979_nl, fsm_output(1));
  mux_2988_seb <= MUX_s_1_2_2(mux_2987_nl, mux_2983_nl, fsm_output(5));
  or_3189_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  or_3187_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_3003_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_2909, fsm_output(0));
  nor_943_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10101")));
  mux_3004_nl <= MUX_s_1_2_2(or_3187_nl, mux_3003_nl, nor_943_nl);
  mux_3005_nl <= MUX_s_1_2_2(or_tmp_2920, mux_3004_nl, fsm_output(3));
  mux_3006_nl <= MUX_s_1_2_2(mux_3005_nl, or_tmp_2918, fsm_output(1));
  nand_159_nl <= NOT((fsm_output(4)) AND (NOT mux_3006_nl));
  mux_3007_nl <= MUX_s_1_2_2(or_3189_nl, nand_159_nl, fsm_output(6));
  mux_3008_nl <= MUX_s_1_2_2(mux_3007_nl, mux_tmp_2995, fsm_output(5));
  nor_1553_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_2998_nl <= MUX_s_1_2_2(nor_1553_nl, (fsm_output(2)), fsm_output(0));
  mux_2999_nl <= MUX_s_1_2_2((NOT mux_2998_nl), (fsm_output(2)), fsm_output(3));
  mux_3000_nl <= MUX_s_1_2_2(mux_2999_nl, or_2215_cse, fsm_output(1));
  or_3185_nl <= (fsm_output(4)) OR mux_3000_nl;
  mux_2996_nl <= MUX_s_1_2_2(or_tmp_2920, (fsm_output(2)), fsm_output(3));
  mux_2997_nl <= MUX_s_1_2_2(mux_2996_nl, or_tmp_2918, fsm_output(1));
  nand_158_nl <= NOT((fsm_output(4)) AND (NOT mux_2997_nl));
  mux_3001_nl <= MUX_s_1_2_2(or_3185_nl, nand_158_nl, fsm_output(6));
  mux_3002_nl <= MUX_s_1_2_2(mux_3001_nl, mux_tmp_2995, fsm_output(5));
  mux_3009_nl <= MUX_s_1_2_2(mux_3008_nl, mux_3002_nl, nor_951_cse);
  nor_1554_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  nor_1555_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  mux_2989_nl <= MUX_s_1_2_2(nor_1554_nl, nor_1555_nl, fsm_output(1));
  nand_156_nl <= NOT(nor_2197_cse AND mux_2989_nl);
  mux_2990_nl <= MUX_s_1_2_2(nand_156_nl, or_3159_cse, fsm_output(5));
  mux_3010_itm <= MUX_s_1_2_2(mux_3009_nl, mux_2990_nl, fsm_output(7));
  nor_947_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  nor_951_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  or_3209_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_3030_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3209_nl);
  mux_3031_nl <= MUX_s_1_2_2(mux_3030_nl, mux_1872_cse, fsm_output(3));
  mux_3026_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, nor_947_cse);
  mux_3027_nl <= MUX_s_1_2_2(mux_3026_nl, mux_1865_cse, fsm_output(4));
  mux_3028_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3027_nl, fsm_output(3));
  mux_3032_cse <= MUX_s_1_2_2(mux_3031_nl, mux_3028_nl, fsm_output(1));
  and_1461_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3035_nl <= MUX_s_1_2_2(and_1461_nl, mux_1877_cse, nor_951_cse);
  mux_3036_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3035_nl, nor_636_cse);
  mux_3037_seb <= MUX_s_1_2_2(mux_3036_nl, mux_3032_cse, fsm_output(5));
  or_3248_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  or_3245_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10110"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_3243_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_3050_nl <= MUX_s_1_2_2(or_3245_nl, or_3243_nl, fsm_output(0));
  mux_3051_nl <= MUX_s_1_2_2(or_tmp_2974, mux_3050_nl, fsm_output(3));
  or_3246_nl <= (fsm_output(1)) OR mux_3051_nl;
  mux_3052_nl <= MUX_s_1_2_2(or_3248_nl, or_3246_nl, fsm_output(6));
  mux_3053_nl <= MUX_s_1_2_2(mux_3052_nl, mux_tmp_3043, fsm_output(5));
  or_3241_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_3045_nl <= MUX_s_1_2_2(or_3241_nl, or_2273_cse, fsm_output(0));
  mux_3046_nl <= MUX_s_1_2_2(mux_3045_nl, or_2272_cse, fsm_output(3));
  mux_3047_nl <= MUX_s_1_2_2(mux_3046_nl, or_2271_cse, fsm_output(1));
  mux_3044_nl <= MUX_s_1_2_2(or_tmp_2974, or_119_cse, fsm_output(3));
  or_3236_nl <= (fsm_output(1)) OR mux_3044_nl;
  mux_3048_nl <= MUX_s_1_2_2(mux_3047_nl, or_3236_nl, fsm_output(6));
  mux_3049_nl <= MUX_s_1_2_2(mux_3048_nl, mux_tmp_3043, fsm_output(5));
  mux_3054_nl <= MUX_s_1_2_2(mux_3053_nl, mux_3049_nl, nor_969_cse);
  or_3219_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_3038_nl <= MUX_s_1_2_2(or_3219_nl, or_3159_cse, fsm_output(5));
  mux_3055_itm <= MUX_s_1_2_2(mux_3054_nl, mux_3038_nl, fsm_output(7));
  nor_969_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1449_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3091_nl <= MUX_s_1_2_2(and_1449_nl, mux_1877_cse, nor_969_cse);
  mux_3092_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3091_nl, nor_636_cse);
  mux_3093_seb <= MUX_s_1_2_2(mux_3092_nl, mux_3032_cse, fsm_output(5));
  or_3294_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_3107_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_3018, fsm_output(0));
  mux_3108_nl <= MUX_s_1_2_2(or_tmp_3020, mux_3107_nl, and_1447_cse);
  or_3292_nl <= (fsm_output(1)) OR mux_3108_nl;
  mux_3109_nl <= MUX_s_1_2_2(mux_tmp_3100, or_3292_nl, fsm_output(3));
  nand_164_nl <= NOT((fsm_output(6)) AND (NOT mux_3109_nl));
  mux_3110_nl <= MUX_s_1_2_2(or_3294_nl, nand_164_nl, fsm_output(4));
  mux_3111_nl <= MUX_s_1_2_2(mux_3110_nl, mux_tmp_3099, fsm_output(5));
  and_2143_nl <= (fsm_output(2)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND S1_OUTER_LOOP_for_acc_svs_4;
  mux_3102_nl <= MUX_s_1_2_2(and_2143_nl, (fsm_output(2)), fsm_output(0));
  mux_3103_nl <= MUX_s_1_2_2((NOT mux_3102_nl), or_4378_cse, fsm_output(1));
  mux_3104_nl <= MUX_s_1_2_2(mux_3103_nl, or_4699_cse, fsm_output(3));
  or_3291_nl <= (fsm_output(6)) OR mux_3104_nl;
  mux_3101_nl <= MUX_s_1_2_2(mux_tmp_3100, or_4699_cse, fsm_output(3));
  nand_163_nl <= NOT((fsm_output(6)) AND (NOT mux_3101_nl));
  mux_3105_nl <= MUX_s_1_2_2(or_3291_nl, nand_163_nl, fsm_output(4));
  mux_3106_nl <= MUX_s_1_2_2(mux_3105_nl, mux_tmp_3099, fsm_output(5));
  mux_3112_nl <= MUX_s_1_2_2(mux_3111_nl, mux_3106_nl, and_1435_cse);
  or_3272_nl <= (fsm_output(0)) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_3094_nl <= MUX_s_1_2_2(or_tmp_3012, or_3272_nl, fsm_output(1));
  or_4432_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_3094_nl;
  mux_3095_nl <= MUX_s_1_2_2(or_4432_nl, or_3159_cse, fsm_output(5));
  mux_3113_itm <= MUX_s_1_2_2(mux_3112_nl, mux_3095_nl, fsm_output(7));
  and_1435_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1433_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("10111"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3149_nl <= MUX_s_1_2_2(and_1433_nl, mux_1877_cse, and_1435_cse);
  mux_3150_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3149_nl, nor_636_cse);
  mux_3151_seb <= MUX_s_1_2_2(mux_3150_nl, mux_3032_cse, fsm_output(5));
  or_3350_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_520_cse;
  or_3347_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11000"));
  mux_3170_nl <= MUX_s_1_2_2(mux_tmp_3163, or_tmp_3064, or_3347_nl);
  or_3346_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR nand_520_cse;
  mux_3169_nl <= MUX_s_1_2_2(or_3346_nl, or_tmp_3071, fsm_output(1));
  mux_3171_nl <= MUX_s_1_2_2(mux_3170_nl, mux_3169_nl, fsm_output(0));
  mux_3172_nl <= MUX_s_1_2_2(or_tmp_3074, mux_3171_nl, fsm_output(6));
  or_3348_nl <= (fsm_output(2)) OR mux_3172_nl;
  mux_3173_nl <= MUX_s_1_2_2(or_3350_nl, or_3348_nl, fsm_output(4));
  or_3342_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR nand_520_cse;
  mux_3165_nl <= MUX_s_1_2_2(or_3342_nl, or_2158_cse, fsm_output(1));
  mux_3166_nl <= MUX_s_1_2_2(mux_3165_nl, or_2157_cse, fsm_output(0));
  or_3343_nl <= (fsm_output(6)) OR mux_3166_nl;
  mux_3167_nl <= MUX_s_1_2_2(or_2161_cse, or_3343_nl, fsm_output(2));
  mux_3164_nl <= MUX_s_1_2_2(or_tmp_3074, mux_tmp_3163, fsm_output(6));
  or_3338_nl <= (fsm_output(2)) OR mux_3164_nl;
  mux_3168_nl <= MUX_s_1_2_2(mux_3167_nl, or_3338_nl, fsm_output(4));
  mux_3174_nl <= MUX_s_1_2_2(mux_3173_nl, mux_3168_nl, nor_1010_cse);
  or_3331_nl <= (fsm_output(7)) OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)) OR not_tmp_1143;
  mux_3156_nl <= MUX_s_1_2_2(or_3331_nl, (fsm_output(7)), fsm_output(3));
  mux_3157_nl <= MUX_s_1_2_2(or_2147_cse, mux_3156_nl, fsm_output(1));
  mux_3158_nl <= MUX_s_1_2_2(mux_3157_nl, mux_tmp_3153, fsm_output(0));
  mux_3159_nl <= MUX_s_1_2_2(mux_3158_nl, mux_tmp_3152, fsm_output(6));
  mux_3160_nl <= MUX_s_1_2_2(mux_3159_nl, nand_331_cse, fsm_output(2));
  mux_3154_nl <= MUX_s_1_2_2(or_tmp_3064, mux_tmp_3153, fsm_output(0));
  mux_3155_nl <= MUX_s_1_2_2(mux_3154_nl, mux_tmp_3152, fsm_output(6));
  or_3328_nl <= (fsm_output(2)) OR mux_3155_nl;
  mux_3161_nl <= MUX_s_1_2_2(mux_3160_nl, or_3328_nl, or_3367_cse);
  or_3316_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0))
      OR not_tmp_1143;
  mux_3162_nl <= MUX_s_1_2_2(mux_3161_nl, or_3316_nl, fsm_output(4));
  mux_3175_itm <= MUX_s_1_2_2(mux_3174_nl, mux_3162_nl, fsm_output(5));
  or_3367_cse <= CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("110"));
  nor_1010_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1423_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11000"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3206_nl <= MUX_s_1_2_2(and_1423_nl, mux_1877_cse, nor_1010_cse);
  mux_3207_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3206_nl, nor_636_cse);
  or_3369_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_3201_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3369_nl);
  mux_3202_nl <= MUX_s_1_2_2(mux_3201_nl, mux_1872_cse, fsm_output(3));
  mux_3197_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_3367_cse);
  mux_3198_nl <= MUX_s_1_2_2(mux_3197_nl, mux_1865_cse, fsm_output(4));
  mux_3199_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3198_nl, fsm_output(3));
  mux_3203_nl <= MUX_s_1_2_2(mux_3202_nl, mux_3199_nl, fsm_output(1));
  mux_3208_seb <= MUX_s_1_2_2(mux_3207_nl, mux_3203_nl, fsm_output(5));
  or_3399_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_520_cse;
  or_3397_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR nand_520_cse;
  mux_3223_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_3118, fsm_output(0));
  nor_1016_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11001")));
  mux_3224_nl <= MUX_s_1_2_2(or_3397_nl, mux_3223_nl, nor_1016_nl);
  mux_3225_nl <= MUX_s_1_2_2(or_tmp_3125, mux_3224_nl, fsm_output(3));
  mux_3226_nl <= MUX_s_1_2_2(mux_3225_nl, or_tmp_3124, fsm_output(1));
  nand_168_nl <= NOT((fsm_output(4)) AND (NOT mux_3226_nl));
  mux_3227_nl <= MUX_s_1_2_2(or_3399_nl, nand_168_nl, fsm_output(6));
  mux_3228_nl <= MUX_s_1_2_2(mux_3227_nl, mux_tmp_3215, fsm_output(5));
  nor_1519_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("001")) OR nand_520_cse);
  mux_3218_nl <= MUX_s_1_2_2(nor_1519_nl, (fsm_output(2)), fsm_output(0));
  mux_3219_nl <= MUX_s_1_2_2((NOT mux_3218_nl), (fsm_output(2)), fsm_output(3));
  mux_3220_nl <= MUX_s_1_2_2(mux_3219_nl, or_2215_cse, fsm_output(1));
  or_3395_nl <= (fsm_output(4)) OR mux_3220_nl;
  mux_3216_nl <= MUX_s_1_2_2(or_tmp_3125, (fsm_output(2)), fsm_output(3));
  mux_3217_nl <= MUX_s_1_2_2(mux_3216_nl, or_tmp_3124, fsm_output(1));
  nand_167_nl <= NOT((fsm_output(4)) AND (NOT mux_3217_nl));
  mux_3221_nl <= MUX_s_1_2_2(or_3395_nl, nand_167_nl, fsm_output(6));
  mux_3222_nl <= MUX_s_1_2_2(mux_3221_nl, mux_tmp_3215, fsm_output(5));
  mux_3229_nl <= MUX_s_1_2_2(mux_3228_nl, mux_3222_nl, nor_1025_cse);
  nor_1520_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110")));
  nor_1521_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110")));
  mux_3209_nl <= MUX_s_1_2_2(nor_1520_nl, nor_1521_nl, fsm_output(1));
  nand_165_nl <= NOT(nor_2197_cse AND mux_3209_nl);
  mux_3210_nl <= MUX_s_1_2_2(nand_165_nl, or_3377_cse, fsm_output(5));
  mux_3230_itm <= MUX_s_1_2_2(mux_3229_nl, mux_3210_nl, fsm_output(7));
  or_3418_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  nor_1025_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  or_3420_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_3250_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3420_nl);
  mux_3251_nl <= MUX_s_1_2_2(mux_3250_nl, mux_1872_cse, fsm_output(3));
  mux_3246_nl <= MUX_s_1_2_2(mux_1868_cse, nor_tmp_35, or_3418_cse);
  mux_3247_nl <= MUX_s_1_2_2(mux_3246_nl, mux_1865_cse, fsm_output(4));
  mux_3248_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3247_nl, fsm_output(3));
  mux_3252_cse <= MUX_s_1_2_2(mux_3251_nl, mux_3248_nl, fsm_output(1));
  and_1417_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3255_nl <= MUX_s_1_2_2(and_1417_nl, mux_1877_cse, nor_1025_cse);
  mux_3256_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3255_nl, nor_636_cse);
  mux_3257_seb <= MUX_s_1_2_2(mux_3256_nl, mux_3252_cse, fsm_output(5));
  or_3452_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_520_cse;
  or_3449_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11010"))
      OR (fsm_output(2)) OR (NOT (fsm_output(4)));
  or_3447_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR nand_520_cse;
  mux_3270_nl <= MUX_s_1_2_2(or_3449_nl, or_3447_nl, fsm_output(0));
  mux_3271_nl <= MUX_s_1_2_2(or_tmp_3173, mux_3270_nl, fsm_output(3));
  or_3450_nl <= (fsm_output(1)) OR mux_3271_nl;
  mux_3272_nl <= MUX_s_1_2_2(or_3452_nl, or_3450_nl, fsm_output(6));
  mux_3273_nl <= MUX_s_1_2_2(mux_3272_nl, mux_tmp_3263, fsm_output(5));
  or_3445_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR nand_520_cse;
  mux_3265_nl <= MUX_s_1_2_2(or_3445_nl, or_2273_cse, fsm_output(0));
  mux_3266_nl <= MUX_s_1_2_2(mux_3265_nl, or_2272_cse, fsm_output(3));
  mux_3267_nl <= MUX_s_1_2_2(mux_3266_nl, or_2271_cse, fsm_output(1));
  mux_3264_nl <= MUX_s_1_2_2(or_tmp_3173, or_119_cse, fsm_output(3));
  or_3440_nl <= (fsm_output(1)) OR mux_3264_nl;
  mux_3268_nl <= MUX_s_1_2_2(mux_3267_nl, or_3440_nl, fsm_output(6));
  mux_3269_nl <= MUX_s_1_2_2(mux_3268_nl, mux_tmp_3263, fsm_output(5));
  mux_3274_nl <= MUX_s_1_2_2(mux_3273_nl, mux_3269_nl, nor_1044_cse);
  or_3428_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_3258_nl <= MUX_s_1_2_2(or_3428_nl, or_3377_cse, fsm_output(5));
  mux_3275_itm <= MUX_s_1_2_2(mux_3274_nl, mux_3258_nl, fsm_output(7));
  nor_1044_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1405_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3311_nl <= MUX_s_1_2_2(and_1405_nl, mux_1877_cse, nor_1044_cse);
  mux_3312_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3311_nl, nor_636_cse);
  mux_3313_seb <= MUX_s_1_2_2(mux_3312_nl, mux_3252_cse, fsm_output(5));
  or_3493_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT (fsm_output(2)))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_520_cse;
  mux_3327_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_3214, fsm_output(0));
  mux_3328_nl <= MUX_s_1_2_2(or_tmp_3216, mux_3327_nl, and_1403_cse);
  or_3491_nl <= (fsm_output(1)) OR mux_3328_nl;
  mux_3329_nl <= MUX_s_1_2_2(mux_tmp_3320, or_3491_nl, fsm_output(3));
  nand_173_nl <= NOT((fsm_output(6)) AND (NOT mux_3329_nl));
  mux_3330_nl <= MUX_s_1_2_2(or_3493_nl, nand_173_nl, fsm_output(4));
  mux_3331_nl <= MUX_s_1_2_2(mux_3330_nl, mux_tmp_3319, fsm_output(5));
  nor_1501_nl <= NOT((NOT((fsm_output(2)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("011")))) OR nand_520_cse);
  mux_3322_nl <= MUX_s_1_2_2(nor_1501_nl, (fsm_output(2)), fsm_output(0));
  mux_3323_nl <= MUX_s_1_2_2((NOT mux_3322_nl), or_4378_cse, fsm_output(1));
  mux_3324_nl <= MUX_s_1_2_2(mux_3323_nl, or_4699_cse, fsm_output(3));
  or_3490_nl <= (fsm_output(6)) OR mux_3324_nl;
  mux_3321_nl <= MUX_s_1_2_2(mux_tmp_3320, or_4699_cse, fsm_output(3));
  nand_172_nl <= NOT((fsm_output(6)) AND (NOT mux_3321_nl));
  mux_3325_nl <= MUX_s_1_2_2(or_3490_nl, nand_172_nl, fsm_output(4));
  mux_3326_nl <= MUX_s_1_2_2(mux_3325_nl, mux_tmp_3319, fsm_output(5));
  mux_3332_nl <= MUX_s_1_2_2(mux_3331_nl, mux_3326_nl, and_1391_cse);
  or_3476_nl <= (fsm_output(0)) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_3314_nl <= MUX_s_1_2_2(or_tmp_3210, or_3476_nl, fsm_output(1));
  or_4411_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_3314_nl;
  mux_3315_nl <= MUX_s_1_2_2(or_4411_nl, or_3377_cse, fsm_output(5));
  mux_3333_itm <= MUX_s_1_2_2(mux_3332_nl, mux_3315_nl, fsm_output(7));
  and_1391_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1011"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1389_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11011"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3369_nl <= MUX_s_1_2_2(and_1389_nl, mux_1877_cse, and_1391_cse);
  mux_3370_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3369_nl, nor_636_cse);
  mux_3371_seb <= MUX_s_1_2_2(mux_3370_nl, mux_3252_cse, fsm_output(5));
  or_3547_nl <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_517_cse;
  or_3544_nl <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11100"));
  mux_3390_nl <= MUX_s_1_2_2(mux_tmp_3383, or_tmp_3261, or_3544_nl);
  or_3543_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR nand_517_cse;
  mux_3389_nl <= MUX_s_1_2_2(or_3543_nl, or_tmp_3264, fsm_output(1));
  mux_3391_nl <= MUX_s_1_2_2(mux_3390_nl, mux_3389_nl, fsm_output(0));
  mux_3392_nl <= MUX_s_1_2_2(or_tmp_3266, mux_3391_nl, fsm_output(6));
  or_3545_nl <= (fsm_output(2)) OR mux_3392_nl;
  mux_3393_nl <= MUX_s_1_2_2(or_3547_nl, or_3545_nl, fsm_output(4));
  or_3539_nl <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR nand_517_cse;
  mux_3385_nl <= MUX_s_1_2_2(or_3539_nl, or_2158_cse, fsm_output(1));
  mux_3386_nl <= MUX_s_1_2_2(mux_3385_nl, or_2157_cse, fsm_output(0));
  or_3540_nl <= (fsm_output(6)) OR mux_3386_nl;
  mux_3387_nl <= MUX_s_1_2_2(or_2161_cse, or_3540_nl, fsm_output(2));
  mux_3384_nl <= MUX_s_1_2_2(or_tmp_3266, mux_tmp_3383, fsm_output(6));
  or_3535_nl <= (fsm_output(2)) OR mux_3384_nl;
  mux_3388_nl <= MUX_s_1_2_2(mux_3387_nl, or_3535_nl, fsm_output(4));
  mux_3394_nl <= MUX_s_1_2_2(mux_3393_nl, mux_3388_nl, nor_1089_cse);
  mux_3379_nl <= MUX_s_1_2_2(or_tmp_3261, mux_tmp_3373, fsm_output(0));
  mux_3380_nl <= MUX_s_1_2_2(mux_3379_nl, mux_tmp_3372, fsm_output(6));
  or_3530_nl <= (fsm_output(2)) OR mux_3380_nl;
  or_3526_nl <= (fsm_output(7)) OR not_tmp_1199;
  mux_3374_nl <= MUX_s_1_2_2(or_3526_nl, (fsm_output(7)), fsm_output(3));
  mux_3375_nl <= MUX_s_1_2_2(or_2147_cse, mux_3374_nl, fsm_output(1));
  mux_3376_nl <= MUX_s_1_2_2(mux_3375_nl, mux_tmp_3373, fsm_output(0));
  mux_3377_nl <= MUX_s_1_2_2(mux_3376_nl, mux_tmp_3372, fsm_output(6));
  mux_3378_nl <= MUX_s_1_2_2(mux_3377_nl, nand_331_cse, fsm_output(2));
  mux_3381_nl <= MUX_s_1_2_2(or_3530_nl, mux_3378_nl, and_1380_cse);
  or_3517_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(0)) OR (fsm_output(1))
      OR (fsm_output(3)) OR (fsm_output(7)) OR not_tmp_1199;
  mux_3382_nl <= MUX_s_1_2_2(mux_3381_nl, or_3517_nl, fsm_output(4));
  mux_3395_itm <= MUX_s_1_2_2(mux_3394_nl, mux_3382_nl, fsm_output(5));
  and_1380_cse <= CONV_SL_1_1(operator_20_true_28_acc_tmp=STD_LOGIC_VECTOR'("111"));
  nor_1089_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg));
  and_1376_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11100"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3426_nl <= MUX_s_1_2_2(and_1376_nl, mux_1877_cse, nor_1089_cse);
  mux_3427_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3426_nl, nor_636_cse);
  or_3565_nl <= (fsm_output(4)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_3421_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3565_nl);
  mux_3422_nl <= MUX_s_1_2_2(mux_3421_nl, mux_1872_cse, fsm_output(3));
  mux_3417_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, and_1380_cse);
  mux_3418_nl <= MUX_s_1_2_2(mux_3417_nl, mux_1865_cse, fsm_output(4));
  mux_3419_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3418_nl, fsm_output(3));
  mux_3423_nl <= MUX_s_1_2_2(mux_3422_nl, mux_3419_nl, fsm_output(1));
  mux_3428_seb <= MUX_s_1_2_2(mux_3427_nl, mux_3423_nl, fsm_output(5));
  or_3574_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR nand_480_cse;
  or_3599_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_517_cse;
  or_3597_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR nand_517_cse;
  mux_3443_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_3312, fsm_output(0));
  mux_3444_nl <= MUX_s_1_2_2(or_3597_nl, mux_3443_nl, and_1373_cse);
  mux_3445_nl <= MUX_s_1_2_2(not_tmp_1218, mux_3444_nl, fsm_output(3));
  mux_3446_nl <= MUX_s_1_2_2(mux_3445_nl, or_tmp_3320, fsm_output(1));
  nand_176_nl <= NOT((fsm_output(4)) AND (NOT mux_3446_nl));
  mux_3447_nl <= MUX_s_1_2_2(or_3599_nl, nand_176_nl, fsm_output(6));
  mux_3448_nl <= MUX_s_1_2_2(mux_3447_nl, mux_tmp_3435, fsm_output(5));
  nor_1485_nl <= NOT((NOT (fsm_output(2))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")) OR nand_517_cse);
  mux_3438_nl <= MUX_s_1_2_2(nor_1485_nl, (fsm_output(2)), fsm_output(0));
  mux_3439_nl <= MUX_s_1_2_2((NOT mux_3438_nl), (fsm_output(2)), fsm_output(3));
  mux_3440_nl <= MUX_s_1_2_2(mux_3439_nl, or_2215_cse, fsm_output(1));
  or_3595_nl <= (fsm_output(4)) OR mux_3440_nl;
  mux_3436_nl <= MUX_s_1_2_2(not_tmp_1218, (fsm_output(2)), fsm_output(3));
  mux_3437_nl <= MUX_s_1_2_2(mux_3436_nl, or_tmp_3320, fsm_output(1));
  nand_175_nl <= NOT((fsm_output(4)) AND (NOT mux_3437_nl));
  mux_3441_nl <= MUX_s_1_2_2(or_3595_nl, nand_175_nl, fsm_output(6));
  mux_3442_nl <= MUX_s_1_2_2(mux_3441_nl, mux_tmp_3435, fsm_output(5));
  mux_3449_nl <= MUX_s_1_2_2(mux_3448_nl, mux_3442_nl, and_1366_cse);
  nor_1486_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(0)) OR (NOT nor_tmp_1094));
  nor_1487_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR nand_480_cse);
  mux_3429_nl <= MUX_s_1_2_2(nor_1486_nl, nor_1487_nl, fsm_output(1));
  nand_174_nl <= NOT(nor_2197_cse AND mux_3429_nl);
  mux_3430_nl <= MUX_s_1_2_2(nand_174_nl, or_3574_cse, fsm_output(5));
  mux_3450_itm <= MUX_s_1_2_2(mux_3449_nl, mux_3430_nl, fsm_output(7));
  and_1369_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  and_1366_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1101"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_3619_nl <= (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(0)) OR (fsm_output(2));
  mux_3470_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_3619_nl);
  mux_3471_nl <= MUX_s_1_2_2(mux_3470_nl, mux_1872_cse, fsm_output(3));
  mux_3466_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1868_cse, and_1369_cse);
  mux_3467_nl <= MUX_s_1_2_2(mux_3466_nl, mux_1865_cse, fsm_output(4));
  mux_3468_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3467_nl, fsm_output(3));
  mux_3472_cse <= MUX_s_1_2_2(mux_3471_nl, mux_3468_nl, fsm_output(1));
  and_1364_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11101"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3475_nl <= MUX_s_1_2_2(and_1364_nl, mux_1877_cse, and_1366_cse);
  mux_3476_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3475_nl, nor_636_cse);
  mux_3477_seb <= MUX_s_1_2_2(mux_3476_nl, mux_3472_cse, fsm_output(5));
  or_3656_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0010")) OR
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR nand_351_cse;
  nand_513_nl <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11110"))
      AND (NOT (fsm_output(2))) AND (fsm_output(4)));
  or_3651_nl <= (fsm_output(2)) OR (NOT (fsm_output(4))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(0))
      OR nand_351_cse;
  mux_3490_nl <= MUX_s_1_2_2(nand_513_nl, or_3651_nl, fsm_output(0));
  mux_3491_nl <= MUX_s_1_2_2(not_tmp_1239, mux_3490_nl, fsm_output(3));
  or_3654_nl <= (fsm_output(1)) OR mux_3491_nl;
  mux_3492_nl <= MUX_s_1_2_2(or_3656_nl, or_3654_nl, fsm_output(6));
  mux_3493_nl <= MUX_s_1_2_2(mux_3492_nl, mux_tmp_3483, fsm_output(5));
  or_3649_nl <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(0))
      OR nand_351_cse;
  mux_3485_nl <= MUX_s_1_2_2(or_3649_nl, or_2273_cse, fsm_output(0));
  mux_3486_nl <= MUX_s_1_2_2(mux_3485_nl, or_2272_cse, fsm_output(3));
  mux_3487_nl <= MUX_s_1_2_2(mux_3486_nl, or_2271_cse, fsm_output(1));
  mux_3484_nl <= MUX_s_1_2_2(not_tmp_1239, or_119_cse, fsm_output(3));
  or_3644_nl <= (fsm_output(1)) OR mux_3484_nl;
  mux_3488_nl <= MUX_s_1_2_2(mux_3487_nl, or_3644_nl, fsm_output(6));
  mux_3489_nl <= MUX_s_1_2_2(mux_3488_nl, mux_tmp_3483, fsm_output(5));
  mux_3494_nl <= MUX_s_1_2_2(mux_3493_nl, mux_3489_nl, and_1350_cse);
  or_3629_nl <= (fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(3)))
      OR (fsm_output(2)) OR not_tmp_1235;
  mux_3478_nl <= MUX_s_1_2_2(or_3629_nl, or_3574_cse, fsm_output(5));
  mux_3495_itm <= MUX_s_1_2_2(mux_3494_nl, mux_3478_nl, fsm_output(7));
  and_1350_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1110"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1348_nl <= ((NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("11110"))
      OR (NOT (fsm_output(4))) OR (fsm_output(0)) OR (fsm_output(2)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3531_nl <= MUX_s_1_2_2(and_1348_nl, mux_1877_cse, and_1350_cse);
  mux_3532_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3531_nl, nor_636_cse);
  mux_3533_seb <= MUX_s_1_2_2(mux_3532_nl, mux_3472_cse, fsm_output(5));
  or_3696_nl <= (fsm_output(6)) OR (fsm_output(3)) OR (fsm_output(1)) OR (NOT nor_tmp_1140);
  mux_3547_nl <= MUX_s_1_2_2((fsm_output(2)), or_tmp_3413, fsm_output(0));
  mux_3548_nl <= MUX_s_1_2_2(or_tmp_3415, mux_3547_nl, and_1344_cse);
  or_3694_nl <= (fsm_output(1)) OR mux_3548_nl;
  mux_3549_nl <= MUX_s_1_2_2(mux_tmp_3540, or_3694_nl, fsm_output(3));
  nand_180_nl <= NOT((fsm_output(6)) AND (NOT mux_3549_nl));
  mux_3550_nl <= MUX_s_1_2_2(or_3696_nl, nand_180_nl, fsm_output(4));
  mux_3551_nl <= MUX_s_1_2_2(mux_3550_nl, mux_tmp_3539, fsm_output(5));
  mux_3542_nl <= MUX_s_1_2_2(nor_tmp_1140, (fsm_output(2)), fsm_output(0));
  mux_3543_nl <= MUX_s_1_2_2((NOT mux_3542_nl), or_4378_cse, fsm_output(1));
  mux_3544_nl <= MUX_s_1_2_2(mux_3543_nl, or_4699_cse, fsm_output(3));
  or_3693_nl <= (fsm_output(6)) OR mux_3544_nl;
  mux_3541_nl <= MUX_s_1_2_2(mux_tmp_3540, or_4699_cse, fsm_output(3));
  nand_179_nl <= NOT((fsm_output(6)) AND (NOT mux_3541_nl));
  mux_3545_nl <= MUX_s_1_2_2(or_3693_nl, nand_179_nl, fsm_output(4));
  mux_3546_nl <= MUX_s_1_2_2(mux_3545_nl, mux_tmp_3539, fsm_output(5));
  mux_3552_nl <= MUX_s_1_2_2(mux_3551_nl, mux_3546_nl, and_1329_cse);
  or_3680_nl <= (fsm_output(0)) OR (fsm_output(2)) OR nand_480_cse;
  mux_3534_nl <= MUX_s_1_2_2(or_tmp_3410, or_3680_nl, fsm_output(1));
  or_4388_nl <= (NOT (fsm_output(4))) OR (fsm_output(6)) OR (NOT (fsm_output(3)))
      OR mux_3534_nl;
  mux_3535_nl <= MUX_s_1_2_2(or_4388_nl, or_3574_cse, fsm_output(5));
  mux_3553_itm <= MUX_s_1_2_2(mux_3552_nl, mux_3535_nl, fsm_output(7));
  and_1329_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  and_1326_nl <= ((CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(4)) AND (NOT (fsm_output(0))) AND (NOT (fsm_output(2)))) OR
      (fsm_output(7))) AND (fsm_output(6));
  mux_3589_nl <= MUX_s_1_2_2(and_1326_nl, mux_1877_cse, and_1329_cse);
  mux_3590_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3589_nl, nor_636_cse);
  mux_3591_seb <= MUX_s_1_2_2(mux_3590_nl, mux_3472_cse, fsm_output(5));
  and_1109_rmff <= ((fsm_output(1)) XOR (fsm_output(2))) AND (fsm_output(4)) AND
      (fsm_output(6)) AND and_dcpl_461;
  nand_531_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")));
  and_1322_nl <= or_4699_cse AND (fsm_output(4));
  mux_3665_nl <= MUX_s_1_2_2(nor_tmp_4, and_1322_nl, fsm_output(0));
  mux_3666_nl <= MUX_s_1_2_2(mux_3665_nl, (NOT mux_tmp_3659), fsm_output(6));
  or_3820_nl <= nor_2183_cse OR (fsm_output(4));
  mux_3663_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), or_4342_cse);
  mux_3664_nl <= MUX_s_1_2_2(or_3820_nl, mux_3663_nl, fsm_output(6));
  mux_3667_nl <= MUX_s_1_2_2(mux_3666_nl, mux_3664_nl, fsm_output(5));
  or_3817_nl <= (fsm_output(2)) OR (fsm_output(1)) OR (NOT (fsm_output(4)));
  mux_3661_nl <= MUX_s_1_2_2((fsm_output(4)), or_3817_nl, fsm_output(6));
  nand_530_nl <= NOT(nand_531_cse AND (fsm_output(4)));
  mux_3660_nl <= MUX_s_1_2_2(mux_tmp_3659, nand_530_nl, fsm_output(6));
  mux_3662_nl <= MUX_s_1_2_2((NOT mux_3661_nl), mux_3660_nl, fsm_output(5));
  mux_3668_nl <= MUX_s_1_2_2((NOT mux_3667_nl), mux_3662_nl, fsm_output(3));
  mux_3657_nl <= MUX_s_1_2_2(or_tmp_3538, or_tmp_3537, fsm_output(5));
  mux_3656_nl <= MUX_s_1_2_2(or_tmp_3537, or_4376_cse, fsm_output(5));
  mux_3658_nl <= MUX_s_1_2_2(mux_3657_nl, mux_3656_nl, fsm_output(3));
  mux_3669_itm <= MUX_s_1_2_2(mux_3668_nl, mux_3658_nl, fsm_output(7));
  or_3852_cse <= (fsm_output(4)) OR (NOT (fsm_output(3))) OR (fsm_output(1));
  nor_1395_cse <= NOT((fsm_output(3)) OR (fsm_output(6)));
  nor_1393_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 2)/=STD_LOGIC_VECTOR'("001101")));
  nor_1394_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(6)));
  mux_3675_nl <= MUX_s_1_2_2(nor_1394_nl, nor_1395_cse, fsm_output(7));
  and_1319_nl <= (fsm_output(4)) AND mux_3675_nl;
  nor_1396_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR not_tmp_1345);
  mux_3676_nl <= MUX_s_1_2_2(and_1319_nl, nor_1396_nl, fsm_output(2));
  nor_1397_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR (NOT (fsm_output(7)))
      OR (NOT (fsm_output(3))) OR (fsm_output(6)));
  mux_3677_nl <= MUX_s_1_2_2(mux_3676_nl, nor_1397_nl, fsm_output(5));
  mux_3678_cse <= MUX_s_1_2_2(nor_1393_nl, mux_3677_nl, fsm_output(1));
  and_1317_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  or_3894_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  and_2141_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  nor_1368_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01")));
  nor_1375_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  nor_2247_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10")));
  or_3918_cse <= (fsm_output(2)) OR (fsm_output(6));
  and_1306_cse <= (fsm_output(4)) AND (fsm_output(1)) AND (fsm_output(2));
  and_2112_cse <= (fsm_output(5)) AND (fsm_output(7));
  and_1272_cse <= (S2_INNER_LOOP1_r_4_0_sva_2(4)) AND (fsm_output(0));
  nor_1262_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(5)));
  mux_4106_nl <= MUX_s_1_2_2((NOT or_tmp_48), and_2112_cse, fsm_output(4));
  mux_4107_nl <= MUX_s_1_2_2(nor_1262_nl, mux_4106_nl, fsm_output(3));
  mux_4102_nl <= MUX_s_1_2_2((fsm_output(5)), (fsm_output(7)), fsm_output(1));
  mux_4103_nl <= MUX_s_1_2_2(or_tmp_48, mux_4102_nl, fsm_output(0));
  and_1270_nl <= (fsm_output(1)) AND (fsm_output(7)) AND (fsm_output(5));
  mux_4104_nl <= MUX_s_1_2_2((NOT mux_4103_nl), and_1270_nl, fsm_output(4));
  nor_1263_nl <= NOT(and_1317_cse OR (fsm_output(7)) OR (fsm_output(5)));
  mux_4099_nl <= MUX_s_1_2_2((fsm_output(7)), (fsm_output(5)), fsm_output(1));
  mux_4100_nl <= MUX_s_1_2_2(and_2112_cse, mux_4099_nl, and_1272_cse);
  mux_4101_nl <= MUX_s_1_2_2(nor_1263_nl, mux_4100_nl, fsm_output(4));
  mux_4105_nl <= MUX_s_1_2_2(mux_4104_nl, mux_4101_nl, fsm_output(3));
  mux_4108_nl <= MUX_s_1_2_2(mux_4107_nl, mux_4105_nl, fsm_output(2));
  mux_4096_nl <= MUX_s_1_2_2(or_tmp_48, or_4162_cse, fsm_output(4));
  mux_4097_nl <= MUX_s_1_2_2(mux_tmp_4094, mux_4096_nl, fsm_output(3));
  mux_4092_nl <= MUX_s_1_2_2(or_tmp_48, (fsm_output(7)), or_3894_cse);
  mux_4093_nl <= MUX_s_1_2_2(mux_4092_nl, or_4162_cse, fsm_output(4));
  mux_4095_nl <= MUX_s_1_2_2(mux_tmp_4094, mux_4093_nl, fsm_output(3));
  mux_4098_nl <= MUX_s_1_2_2(mux_4097_nl, mux_4095_nl, fsm_output(2));
  mux_4109_nl <= MUX_s_1_2_2(mux_4108_nl, mux_4098_nl, fsm_output(6));
  not_9789_nl <= NOT mux_4109_nl;
  S2_INNER_LOOP1_r_S2_INNER_LOOP1_r_and_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"),
      (S2_INNER_LOOP1_r_4_0_sva_2(3 DOWNTO 0)), not_9789_nl);
  and_1172_nl <= and_dcpl_57 AND and_dcpl_110 AND and_dcpl_54;
  S1_OUTER_LOOP_k_or_nl <= (and_dcpl_95 AND (fsm_output(2)) AND and_dcpl_1000 AND
      nor_1711_cse AND and_dcpl_1070) OR (and_dcpl_71 AND (fsm_output(2)) AND and_dcpl_1031
      AND and_dcpl_103 AND and_dcpl_1070);
  nor_2306_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(2))) OR (fsm_output(1))
      OR (fsm_output(4)));
  mux_3728_nl <= MUX_s_1_2_2(nor_2306_nl, nor_2307_cse, fsm_output(5));
  nor_2308_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(2))
      OR (NOT nor_tmp_3));
  mux_3729_nl <= MUX_s_1_2_2(mux_3728_nl, nor_2308_nl, fsm_output(7));
  and_1179_nl <= mux_3729_nl AND (fsm_output(0)) AND (fsm_output(3));
  mux_3739_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), or_tmp_48);
  or_3906_nl <= (fsm_output(1)) OR (fsm_output(5));
  mux_3738_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3906_nl);
  and_1307_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"));
  mux_3740_nl <= MUX_s_1_2_2(mux_3739_nl, mux_3738_nl, and_1307_nl);
  mux_3733_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1274_cse);
  mux_3732_nl <= MUX_s_1_2_2(mux_3731_cse, mux_tmp_3730, fsm_output(1));
  mux_3734_nl <= MUX_s_1_2_2(mux_3733_nl, mux_3732_nl, and_1272_cse);
  mux_3735_nl <= MUX_s_1_2_2(nor_tmp_35, mux_3734_nl, fsm_output(2));
  mux_3736_nl <= MUX_s_1_2_2(mux_3735_nl, mux_tmp_3730, fsm_output(3));
  mux_3741_nl <= MUX_s_1_2_2(mux_3740_nl, mux_3736_nl, fsm_output(4));
  S1_OUTER_LOOP_k_mux1h_1_nl <= MUX1HOT_v_5_4_2((S1_OUTER_LOOP_for_p_sva_1(4 DOWNTO
      0)), (S1_OUTER_LOOP_k_5_0_sva_2(4 DOWNTO 0)), (z_out(4 DOWNTO 0)), ('0' & S2_INNER_LOOP1_r_S2_INNER_LOOP1_r_and_nl),
      STD_LOGIC_VECTOR'( and_1172_nl & S1_OUTER_LOOP_k_or_nl & and_1179_nl & (NOT
      mux_3741_nl)));
  or_4690_nl <= (fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(6))
      OR (fsm_output(1)) OR (fsm_output(5));
  and_1312_nl <= (NOT((fsm_output(7)) OR (NOT (S1_OUTER_LOOP_k_5_0_sva_2(5))))) AND
      mux_108_cse;
  nor_1362_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(1))) OR (fsm_output(5)));
  nor_1363_nl <= NOT((fsm_output(6)) OR (fsm_output(1)) OR (NOT (fsm_output(5))));
  mux_3724_nl <= MUX_s_1_2_2(nor_1362_nl, nor_1363_nl, fsm_output(7));
  and_1313_nl <= (S2_INNER_LOOP1_r_4_0_sva_2(4)) AND mux_3724_nl;
  mux_3726_nl <= MUX_s_1_2_2(and_1312_nl, and_1313_nl, fsm_output(4));
  nand_534_nl <= NOT((fsm_output(2)) AND mux_3726_nl);
  mux_3727_nl <= MUX_s_1_2_2(or_4690_nl, nand_534_nl, fsm_output(0));
  S2_COPY_LOOP_p_or_nl <= mux_3727_nl OR (fsm_output(3));
  S2_COPY_LOOP_p_asn_S2_COPY_LOOP_p_5_0_sva_4_0_S1_OUTER_LOOP_k_and_rgt <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      S1_OUTER_LOOP_k_mux1h_1_nl, S2_COPY_LOOP_p_or_nl);
  and_2893_cse <= (fsm_output(0)) AND (fsm_output(2));
  or_4854_cse <= (fsm_output(3)) OR (fsm_output(6));
  nor_2186_cse <= NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01")));
  nor_2183_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  and_2120_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111"));
  nor_2178_cse_1 <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  mux_45_cse <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(6));
  or_129_cse <= (NOT (fsm_output(2))) OR (fsm_output(4)) OR (NOT (fsm_output(1)));
  or_115_nl <= (fsm_output(4)) OR (NOT (fsm_output(1)));
  mux_37_cse <= MUX_s_1_2_2(or_115_nl, or_tmp_35, fsm_output(2));
  or_124_cse <= (fsm_output(6)) OR nor_tmp_4;
  nand_536_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11")));
  and_67_nl <= and_dcpl_57 AND and_2893_cse AND and_dcpl_54;
  and_74_nl <= and_dcpl_64 AND and_dcpl_61;
  and_77_nl <= and_dcpl_67 AND and_dcpl_61;
  S1_OUTER_LOOP_k_mux1h_nl <= MUX1HOT_v_5_3_2((S1_OUTER_LOOP_k_5_0_sva_2(4 DOWNTO
      0)), (S1_OUTER_LOOP_for_p_sva_1(4 DOWNTO 0)), (z_out(4 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_67_nl & and_74_nl & and_77_nl));
  or_271_nl <= nor_2183_cse OR (fsm_output(6));
  nand_535_nl <= NOT(nand_536_cse AND (fsm_output(6)));
  mux_92_nl <= MUX_s_1_2_2(or_271_nl, nand_535_nl, fsm_output(5));
  nor_nl <= NOT((fsm_output(7)) OR mux_92_nl);
  and_2150_nl <= (fsm_output(7)) AND (fsm_output(5)) AND (fsm_output(2)) AND (fsm_output(1))
      AND (NOT (fsm_output(6)));
  mux_93_nl <= MUX_s_1_2_2(nor_nl, and_2150_nl, fsm_output(4));
  nor_2184_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10")));
  nor_2185_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(2)) OR nor_2186_cse OR
      (fsm_output(6)));
  mux_91_nl <= MUX_s_1_2_2(nor_2184_nl, nor_2185_nl, fsm_output(7));
  and_2151_nl <= (fsm_output(4)) AND mux_91_nl;
  mux_94_nl <= MUX_s_1_2_2(mux_93_nl, and_2151_nl, fsm_output(3));
  S1_OUTER_LOOP_k_asn_S2_COPY_LOOP_for_i_5_0_sva_2_4_S1_OUTER_LOOP_k_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      S1_OUTER_LOOP_k_mux1h_nl, mux_94_nl);
  not_9788_nl <= NOT mux_tmp_4069;
  S2_INNER_LOOP1_for_p_S2_INNER_LOOP1_for_p_and_nl <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"),
      (S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)), not_9788_nl);
  nor_1347_nl <= NOT(and_2141_cse OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01")));
  mux_3755_nl <= MUX_s_1_2_2(nor_1346_cse, nor_1347_nl, fsm_output(5));
  and_2138_nl <= (fsm_output(2)) AND (fsm_output(0)) AND (fsm_output(1)) AND (NOT
      (fsm_output(7))) AND (fsm_output(6));
  and_1301_nl <= (fsm_output(2)) AND (NOT(nor_1375_cse OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("10"))));
  mux_3754_nl <= MUX_s_1_2_2(and_2138_nl, and_1301_nl, fsm_output(5));
  mux_3756_nl <= MUX_s_1_2_2(mux_3755_nl, mux_3754_nl, fsm_output(4));
  nor_1352_nl <= NOT((fsm_output(2)) OR nor_2186_cse OR CONV_SL_1_1(fsm_output(7
      DOWNTO 6)/=STD_LOGIC_VECTOR'("10")));
  mux_3753_nl <= MUX_s_1_2_2(nor_1368_cse, nor_1352_nl, fsm_output(5));
  and_1302_nl <= (fsm_output(4)) AND mux_3753_nl;
  mux_3757_nl <= MUX_s_1_2_2(mux_3756_nl, and_1302_nl, fsm_output(3));
  mux_3772_nl <= MUX_s_1_2_2(not_tmp_1345, or_4854_cse, fsm_output(5));
  mux_3773_nl <= MUX_s_1_2_2(mux_3772_nl, mux_tmp_3769, or_3894_cse);
  mux_3774_nl <= MUX_s_1_2_2((NOT mux_3773_nl), or_tmp_3662, fsm_output(4));
  mux_3768_nl <= MUX_s_1_2_2((fsm_output(6)), (fsm_output(3)), fsm_output(5));
  mux_3770_nl <= MUX_s_1_2_2((NOT mux_tmp_3769), mux_3768_nl, fsm_output(1));
  mux_3766_nl <= MUX_s_1_2_2((NOT (fsm_output(6))), or_tmp_3661, fsm_output(5));
  mux_3767_nl <= MUX_s_1_2_2(or_tmp_3662, mux_3766_nl, and_1317_cse);
  mux_3771_nl <= MUX_s_1_2_2(mux_3770_nl, mux_3767_nl, fsm_output(4));
  mux_3775_nl <= MUX_s_1_2_2(mux_3774_nl, mux_3771_nl, fsm_output(2));
  mux_3764_nl <= MUX_s_1_2_2((fsm_output(6)), or_4854_cse, and_dcpl_113);
  or_3935_nl <= and_1317_cse OR (fsm_output(5));
  mux_3762_nl <= MUX_s_1_2_2(or_tmp_3661, (fsm_output(6)), or_3935_nl);
  mux_3759_nl <= MUX_s_1_2_2((fsm_output(6)), or_4854_cse, fsm_output(5));
  mux_3760_nl <= MUX_s_1_2_2(mux_3759_nl, or_tmp_3658, fsm_output(0));
  mux_3758_nl <= MUX_s_1_2_2(or_tmp_3658, or_dcpl_276, fsm_output(0));
  mux_3761_nl <= MUX_s_1_2_2(mux_3760_nl, mux_3758_nl, fsm_output(1));
  mux_3763_nl <= MUX_s_1_2_2(mux_3762_nl, mux_3761_nl, fsm_output(4));
  mux_3765_nl <= MUX_s_1_2_2(mux_3764_nl, mux_3763_nl, fsm_output(2));
  mux_3776_nl <= MUX_s_1_2_2(mux_3775_nl, (NOT mux_3765_nl), fsm_output(7));
  S2_COPY_LOOP_for_i_mux1h_2_rgt <= MUX1HOT_v_6_3_2(('0' & S1_OUTER_LOOP_k_asn_S2_COPY_LOOP_for_i_5_0_sva_2_4_S1_OUTER_LOOP_k_and_nl),
      z_out, (STD_LOGIC_VECTOR'( "000") & S2_INNER_LOOP1_for_p_S2_INNER_LOOP1_for_p_and_nl),
      STD_LOGIC_VECTOR'( mux_3757_nl & and_dcpl_88 & mux_3776_nl));
  nand_570_cse <= NOT((fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(0)) AND
      (fsm_output(1)) AND (fsm_output(2)));
  nand_569_cse <= NOT((fsm_output(5)) AND (fsm_output(1)) AND (fsm_output(2)));
  or_4769_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("10"));
  or_4781_cse <= (fsm_output(5)) OR (NOT (fsm_output(3)));
  nand_568_cse <= NOT((fsm_output(1)) AND (fsm_output(3)));
  or_4699_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"));
  operator_20_true_1_and_cse <= core_wen AND (NOT(or_tmp_301 OR or_dcpl_277));
  or_4378_cse <= (fsm_output(0)) OR (NOT (fsm_output(2)));
  S5_COPY_LOOP_for_acc_6_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(revArr_rsci_s_din_mxwt(9
      DOWNTO 5)) + UNSIGNED(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg & reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg),
      5));
  operator_20_true_1_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(reg_S2_COPY_LOOP_for_i_5_0_2_reg),
      3), 4) + UNSIGNED'( "0001"), 4));
  and_1193_nl <= (NOT mux_tmp_3812) AND and_dcpl_82 AND and_dcpl_79;
  mux_3825_nl <= MUX_s_1_2_2(nor_tmp_1200, (NOT mux_tmp_3819), fsm_output(6));
  mux_47_nl <= MUX_s_1_2_2(or_129_cse, or_2273_cse, fsm_output(0));
  mux_48_nl <= MUX_s_1_2_2(mux_47_nl, (fsm_output(4)), fsm_output(6));
  mux_3826_nl <= MUX_s_1_2_2(mux_3825_nl, mux_48_nl, fsm_output(5));
  mux_3820_nl <= MUX_s_1_2_2((NOT mux_tmp_3819), or_tmp_3706, fsm_output(6));
  mux_3822_nl <= MUX_s_1_2_2((NOT mux_45_cse), mux_3820_nl, fsm_output(5));
  mux_3827_nl <= MUX_s_1_2_2(mux_3826_nl, mux_3822_nl, fsm_output(3));
  mux_3816_nl <= MUX_s_1_2_2(or_2273_cse, or_tmp_3536, fsm_output(0));
  or_3984_nl <= (fsm_output(6)) OR (NOT mux_3816_nl);
  mux_3817_nl <= MUX_s_1_2_2(or_3984_nl, or_124_cse, fsm_output(5));
  mux_3815_nl <= MUX_s_1_2_2(or_124_cse, or_4376_cse, fsm_output(5));
  mux_3818_nl <= MUX_s_1_2_2(mux_3817_nl, mux_3815_nl, fsm_output(3));
  mux_3828_nl <= MUX_s_1_2_2(mux_3827_nl, (NOT mux_3818_nl), fsm_output(7));
  S34_OUTER_LOOP_for_a_mux1h_nl <= MUX1HOT_v_5_5_2(S34_OUTER_LOOP_for_a_acc_2_tmp,
      STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(S5_COPY_LOOP_for_acc_6_nl), 5)), (reg_S2_COPY_LOOP_for_i_5_0_1_reg
      & reg_S2_COPY_LOOP_for_i_5_0_2_reg), ('0' & STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(operator_20_true_1_acc_nl),
      4))), S6_OUTER_LOOP_for_acc_tmp, STD_LOGIC_VECTOR'( and_dcpl_1082 & and_dcpl_1088
      & and_1193_nl & mux_3828_nl & and_dcpl_1084));
  or_3982_nl <= (fsm_output(6)) OR (NOT and_2141_cse);
  or_3981_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(1));
  mux_3813_nl <= MUX_s_1_2_2(or_3982_nl, or_3981_nl, fsm_output(5));
  mux_3814_nl <= MUX_s_1_2_2(mux_3813_nl, mux_tmp_3812, fsm_output(3));
  S1_OUTER_LOOP_for_nand_nl <= NOT((NOT mux_3814_nl) AND and_dcpl_1086);
  S34_OUTER_LOOP_for_a_and_rgt <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), S34_OUTER_LOOP_for_a_mux1h_nl,
      S1_OUTER_LOOP_for_nand_nl);
  or_4805_cse <= (NOT (fsm_output(1))) OR (fsm_output(5));
  or_4797_cse <= (fsm_output(3)) OR (fsm_output(1));
  nor_2412_cse <= NOT((fsm_output(1)) OR (fsm_output(5)));
  nor_2411_cse <= NOT((NOT (fsm_output(1))) OR (fsm_output(5)));
  S1_OUTER_LOOP_for_and_1_cse <= core_wen AND (and_dcpl_1091 OR and_dcpl_93 OR and_dcpl_1084);
  S1_OUTER_LOOP_for_and_2_cse <= core_wen AND (and_dcpl_1091 OR and_dcpl_1092 OR
      and_dcpl_1084);
  S1_OUTER_LOOP_for_and_5_cse <= core_wen AND (and_dcpl_1082 OR and_dcpl_1084);
  S1_OUTER_LOOP_for_and_16_cse <= core_wen AND (and_dcpl_1091 OR and_dcpl_1088 OR
      and_dcpl_1092 OR and_dcpl_1084);
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_61_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11111"));
  or_4691_nl <= (fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(1))
      OR (fsm_output(4));
  or_4692_nl <= (NOT (fsm_output(6))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR (NOT (fsm_output(1))) OR (fsm_output(4));
  mux_3853_nl <= MUX_s_1_2_2(or_4691_nl, or_4692_nl, fsm_output(5));
  or_4020_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(4));
  mux_3852_nl <= MUX_s_1_2_2(or_4020_nl, or_tmp_3740, fsm_output(6));
  or_4693_nl <= (fsm_output(5)) OR mux_3852_nl;
  mux_3854_nl <= MUX_s_1_2_2(mux_3853_nl, or_4693_nl, fsm_output(3));
  S1_OUTER_LOOP_for_and_34_cse <= core_wen AND ((NOT(mux_3854_nl OR (fsm_output(7))))
      OR and_dcpl_1084);
  S1_OUTER_LOOP_for_and_39_cse <= core_wen AND (and_dcpl_1095 OR not_tmp_1436 OR
      and_dcpl_1092 OR and_dcpl_1084);
  S1_OUTER_LOOP_for_and_44_cse <= core_wen AND (and_dcpl_1095 OR and_dcpl_1092 OR
      and_dcpl_1084);
  S1_OUTER_LOOP_for_and_47_cse <= core_wen AND (and_dcpl_1095 OR and_dcpl_93 OR and_dcpl_1084);
  S6_OUTER_LOOP_for_nor_22_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  S1_OUTER_LOOP_for_and_55_cse <= core_wen AND (and_dcpl_1096 OR and_dcpl_1092 OR
      and_dcpl_77);
  S1_OUTER_LOOP_for_and_60_cse <= core_wen AND (and_dcpl_1096 OR and_dcpl_1097 OR
      and_dcpl_1092 OR and_dcpl_77);
  butterFly_4_f1_butterFly_4_f1_nor_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  nor_1311_cse <= NOT((fsm_output(3)) OR (NOT (fsm_output(5))) OR (fsm_output(1)));
  nor_1308_cse <= NOT((fsm_output(5)) OR (NOT (fsm_output(0))));
  nor_1303_cse <= NOT((fsm_output(4)) OR (fsm_output(7)));
  or_4162_cse <= (fsm_output(7)) OR (NOT (fsm_output(5)));
  or_4165_cse <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("10"));
  or_4376_cse <= (fsm_output(4)) OR (fsm_output(6));
  or_119_cse <= (fsm_output(2)) OR (NOT (fsm_output(4)));
  S2_INNER_LOOP1_tf_and_1_cse <= core_wen AND mux_tmp_4069;
  or_4342_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"));
  mux_4078_nl <= MUX_s_1_2_2(nor_tmp_1200, (NOT mux_tmp_4075), fsm_output(6));
  or_4296_nl <= (NOT((fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(1)))) OR (fsm_output(4));
  mux_4079_nl <= MUX_s_1_2_2(mux_4078_nl, or_4296_nl, fsm_output(5));
  mux_4076_nl <= MUX_s_1_2_2((NOT mux_tmp_4075), or_tmp_3706, fsm_output(6));
  mux_4077_nl <= MUX_s_1_2_2((NOT mux_45_cse), mux_4076_nl, fsm_output(5));
  mux_4080_nl <= MUX_s_1_2_2(mux_4079_nl, mux_4077_nl, fsm_output(3));
  mux_4071_nl <= MUX_s_1_2_2(or_tmp_3538, or_tmp_4014, fsm_output(5));
  mux_4070_nl <= MUX_s_1_2_2(or_tmp_4014, or_4376_cse, fsm_output(5));
  mux_4072_nl <= MUX_s_1_2_2(mux_4071_nl, mux_4070_nl, fsm_output(3));
  mux_4081_nl <= MUX_s_1_2_2(mux_4080_nl, (NOT mux_4072_nl), fsm_output(7));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_mux_6_rgt <= MUX_v_5_2_2((revArr_rsci_s_din_mxwt(4
      DOWNTO 0)), (STD_LOGIC_VECTOR'( "00") & operator_20_true_28_acc_tmp), mux_4081_nl);
  or_4818_cse <= (fsm_output(3)) OR (fsm_output(5));
  and_2881_cse <= (fsm_output(3)) AND (fsm_output(5));
  and_1274_cse <= (fsm_output(5)) AND (fsm_output(1));
  nor_2197_cse <= NOT((fsm_output(6)) OR (NOT (fsm_output(4))));
  butterFly_f1_and_cse <= core_wen AND (NOT(or_tmp_245 OR or_dcpl_277));
  butterFly_4_f1_and_cse <= core_wen AND (NOT(or_dcpl_286 OR or_tmp_3871 OR or_4679_cse));
  butterFly_8_f1_and_cse <= core_wen AND (NOT(or_dcpl_286 OR or_4165_cse OR or_2158_cse));
  operator_20_true_8_and_cse <= core_wen AND (NOT(or_tmp_3740 OR or_4165_cse OR or_4679_cse));
  butterFly_12_f1_and_cse <= core_wen AND (NOT(or_tmp_3540 OR (fsm_output(2)) OR
      (NOT (fsm_output(0))) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR
      or_2158_cse));
  butterFly_16_f1_and_cse <= core_wen AND (NOT(or_tmp_246 OR or_dcpl_276 OR (NOT
      (fsm_output(3))) OR (NOT (fsm_output(7)))));
  butterFly_20_f1_and_cse <= core_wen AND (NOT(or_tmp_246 OR or_dcpl_302));
  operator_20_true_15_and_cse <= core_wen AND (NOT((NOT nor_tmp_3) OR or_4378_cse
      OR or_dcpl_302));
  S6_OUTER_LOOP_for_nor_44_cse <= NOT((S6_OUTER_LOOP_for_acc_tmp(3)) OR (S6_OUTER_LOOP_for_acc_tmp(1)));
  or_261_cse <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1));
  nor_2169_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))));
  mux_108_cse <= MUX_s_1_2_2(nor_2411_cse, nor_2169_nl, fsm_output(6));
  or_309_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_324_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_338_cse <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_337_cse <= (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  or_336_cse <= (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(7));
  or_315_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00000"));
  nor_2142_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  or_394_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_401_cse <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  nor_2144_cse <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  or_387_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_395_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_448_cse <= (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_445_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_447_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00010"));
  nand_492_cse <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  or_501_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_549_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_555_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00100"));
  nor_2081_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 2)/=STD_LOGIC_VECTOR'("000"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01")));
  or_632_cse <= (fsm_output(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (fsm_output(1))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  or_618_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_634_cse <= (fsm_output(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (NOT
      (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  or_686_cse <= (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_682_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_684_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00110"));
  nand_479_cse <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(2 DOWNTO 0)=STD_LOGIC_VECTOR'("111")));
  or_735_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_789_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_795_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01000"));
  nor_2030_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  or_863_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  nor_2032_cse <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  or_856_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_864_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_911_cse <= (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_908_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_910_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01010"));
  or_955_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_1006_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_1012_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01100"));
  or_1073_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_1130_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_1133_cse <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01110"));
  nand_449_cse <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4));
  nor_1928_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  or_1309_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  nor_1930_cse <= NOT((NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  or_1310_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_1358_cse <= (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_1527_cse <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"));
  or_1547_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  nor_1822_cse <= NOT(CONV_SL_1_1(fsm_output(4 DOWNTO 1)/=STD_LOGIC_VECTOR'("0001"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110")));
  and_1812_cse <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg;
  or_1783_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  nand_520_cse <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4);
  or_1784_cse <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  nand_393_cse <= NOT((fsm_output(1)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  nand_517_cse <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 2)=STD_LOGIC_VECTOR'("11"))
      AND S1_OUTER_LOOP_for_acc_svs_4);
  nand_351_cse <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)=STD_LOGIC_VECTOR'("111"))
      AND S1_OUTER_LOOP_for_acc_svs_4);
  nand_336_cse <= NOT((fsm_output(1)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  and_1713_cse <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4;
  or_2161_cse <= (fsm_output(6)) OR (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7));
  or_2158_cse <= (fsm_output(3)) OR (fsm_output(7));
  or_2157_cse <= (fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(7));
  or_2147_cse <= (fsm_output(3)) OR (NOT (fsm_output(7)));
  nand_331_cse <= NOT((fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(1)) AND
      (fsm_output(3)) AND (NOT (fsm_output(7))));
  or_2199_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_2215_cse <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2)));
  or_2273_cse <= (NOT (fsm_output(2))) OR (fsm_output(4));
  or_2272_cse <= (fsm_output(2)) OR (fsm_output(4));
  or_2271_cse <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4));
  or_2396_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_2585_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  and_1532_cse <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01111"));
  or_2958_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_3159_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  and_1447_cse <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10111"));
  or_3377_cse <= (fsm_output(6)) OR (fsm_output(4)) OR (fsm_output(1)) OR (fsm_output(3))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  and_1403_cse <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11011"));
  and_1373_cse <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11101"));
  and_1344_cse <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11111"));
  tmp_37_lpi_3_dfm_mx0w0 <= MUX1HOT_v_32_32_2(S2_INNER_LOOP1_tf_sva, S2_INNER_LOOP1_tfh_sva,
      operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm, tmp_13_sva_4,
      tmp_16_sva_4, tmp_13_sva_5, tmp_13_sva_6, tmp_12_sva_2, tmp_16_sva_8, tmp_13_sva_7,
      tmp_22_sva_5, modulo_add_base_1_sva, tmp_12_sva_4, mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm,
      mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm, mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm,
      operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm, tmp_12_sva_5,
      tmp_12_sva_6, operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm,
      tmp_12_sva_7, tmp_1_sva_7, tmp_16_sva_22, tmp_16_sva_23, tmp_13_sva_2, tmp_10_sva_2,
      tmp_16_sva_26, tmp_10_sva_4, tmp_10_sva_5, tmp_10_sva_6, tmp_10_sva_7, tmp_16_sva_31,
      STD_LOGIC_VECTOR'( S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_26_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_60_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_61_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_8_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_9_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_1_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_18_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_19_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_2_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_20_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_21_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_22_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_23_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_24_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_25_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_27_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_28_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_29_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_30_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_4_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_45_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_53_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_57_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_59_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_6_itm));
  tmp_7_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_15_sva, tmp_15_sva_1, tmp_15_sva_2,
      tmp_15_sva_3, tmp_15_sva_4, tmp_15_sva_5, tmp_15_sva_6, tmp_15_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm
      & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm &
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm));
  S34_OUTER_LOOP_for_a_acc_2_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(reg_S2_COPY_LOOP_for_i_5_0_1_reg
      & reg_S2_COPY_LOOP_for_i_5_0_2_reg) + UNSIGNED(S1_OUTER_LOOP_for_p_sva_1(4
      DOWNTO 0)), 5));
  S6_OUTER_LOOP_for_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(S1_OUTER_LOOP_for_p_sva_1(4
      DOWNTO 0)) + UNSIGNED(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg & reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg),
      5));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_nor_itm_mx0w0 <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp/=STD_LOGIC_VECTOR'("00000")));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_9_itm_mx0w1 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))));
  S34_OUTER_LOOP_for_a_nor_itm_mx0w0 <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(4
      DOWNTO 1)/=STD_LOGIC_VECTOR'("0000")));
  S34_OUTER_LOOP_for_a_nor_1_itm_mx0w1 <= NOT((S34_OUTER_LOOP_for_a_acc_2_tmp(4))
      OR (S34_OUTER_LOOP_for_a_acc_2_tmp(3)) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(2))
      OR (S34_OUTER_LOOP_for_a_acc_2_tmp(0)));
  S34_OUTER_LOOP_for_a_nor_14_itm_mx0w1 <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(3
      DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("00011"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("00101"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("00110"));
  S1_OUTER_LOOP_for_nor_90_cse <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(4
      DOWNTO 3)/=STD_LOGIC_VECTOR'("00")));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND S1_OUTER_LOOP_for_nor_90_cse;
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01001"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01010"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01011"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01100"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01101"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("01110"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_5_itm_mx0w1 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_25_itm_mx0w2 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1010"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10001"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10010"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10011"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10100"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10101"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("10110"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_8_itm_mx0w1 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_27_itm_mx0w2 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1100"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11000"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11001"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11010"));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11100"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_nor_itm_mx0w1 <= NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000")));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_29_itm_mx0w0 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp=STD_LOGIC_VECTOR'("11110"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_4_itm_mx0w1 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))));
  S1_OUTER_LOOP_for_nor_76_cse <= NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_6_itm_mx0w0 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)=STD_LOGIC_VECTOR'("111")) AND S1_OUTER_LOOP_for_nor_76_cse;
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_10_itm_mx0w0 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)) AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))
      AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_12_itm_mx0w0 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))
      AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_13_itm_mx0w0 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)=STD_LOGIC_VECTOR'("111")) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_14_itm_mx0w0 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_18_itm_mx0w0 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0011"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_20_itm_mx0w0 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0101"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_21_itm_mx0w0 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0110"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_16_itm_mx0w1 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0001"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_24_itm_mx0w0 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1001"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_19_itm_mx0w1 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0100"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_2_itm_mx0w1 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("00"))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_23_itm_mx0w1 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1000"));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_11_itm_mx0w0 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 2)=STD_LOGIC_VECTOR'("11")) AND (NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
  S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_17_itm_mx0w0 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0010"));
  or_233_cse <= (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))) OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1));
  nand_508_cse <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg);
  modulo_add_base_3_sva_mx0w4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_6_lpi_4_dfm)
      + UNSIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_add_base_2_sva_mx0w5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_4_lpi_4_dfm)
      + UNSIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_base_1_sva_mx0w6 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_2_lpi_4_dfm)
      + UNSIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_add_base_sva_mx0w7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_lpi_4_dfm)
      + UNSIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_add_base_7_sva_mx0w9 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_34_lpi_4_dfm)
      + UNSIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_add_base_6_sva_mx0w10 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_32_lpi_4_dfm)
      + UNSIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_add_base_5_sva_mx0w11 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_30_lpi_4_dfm)
      + UNSIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_base_4_sva_mx0w12 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_28_lpi_4_dfm)
      + UNSIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_add_base_11_sva_mx0w14 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_14_lpi_3_dfm)
      + UNSIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_base_10_sva_mx0w15 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_12_lpi_3_dfm)
      + UNSIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_add_base_9_sva_mx0w16 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_10_lpi_3_dfm)
      + UNSIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_add_base_8_sva_mx0w17 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_8_lpi_3_dfm)
      + UNSIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_add_base_15_sva_mx0w21 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_44_lpi_4_dfm)
      + UNSIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_add_base_14_sva_mx0w22 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_42_lpi_4_dfm)
      + UNSIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_add_base_13_sva_mx0w23 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_40_lpi_4_dfm)
      + UNSIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_base_12_sva_mx0w24 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_38_lpi_4_dfm)
      + UNSIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_add_base_19_sva_mx0w26 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_23_lpi_4_dfm)
      + UNSIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_add_base_18_sva_mx0w27 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_21_lpi_4_dfm)
      + UNSIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_add_base_17_sva_mx0w28 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_19_lpi_4_dfm)
      + UNSIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_base_16_sva_mx0w29 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_17_lpi_4_dfm)
      + UNSIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_add_base_23_sva_mx0w30 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_52_lpi_3_dfm)
      + UNSIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_add_base_22_sva_mx0w31 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_50_lpi_3_dfm)
      + UNSIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_add_base_21_sva_mx0w32 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_48_lpi_3_dfm)
      + UNSIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_base_20_sva_mx0w33 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_46_lpi_3_dfm)
      + UNSIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  S2_INNER_LOOP1_tf_and_psp_sva_1 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg AND (operator_33_true_return_2_3_0_sva_3
      & operator_33_true_return_2_3_0_sva_2_0);
  operator_20_true_28_acc_tmp <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(reg_S2_COPY_LOOP_for_i_5_0_2_reg)
      + UNSIGNED'( "001"), 3));
  tmp_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_26_sva_26, tmp_26_sva_27, tmp_21_sva_2,
      tmp_26_sva_29, tmp_21_sva_4, tmp_21_sva_5, tmp_21_sva_6, tmp_21_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm));
  tmp_2_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_16_sva_22, tmp_16_sva_23, tmp_10_sva_2,
      tmp_16_sva_26, tmp_10_sva_4, tmp_10_sva_5, tmp_10_sva_6, tmp_10_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm));
  tmp_4_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_16_sva_31, tmp_16_sva_4, tmp_12_sva_2,
      tmp_16_sva_8, tmp_12_sva_4, tmp_12_sva_5, tmp_12_sva_6, tmp_12_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm));
  tmp_6_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_14_sva, tmp_14_sva_1, tmp_14_sva_2,
      tmp_14_sva_3, tmp_14_sva_4, tmp_14_sva_5, tmp_14_sva_6, tmp_14_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm
      & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm &
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm));
  tmp_1_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(modulo_add_base_1_sva, mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm,
      mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm, mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm,
      operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm, operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm,
      operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm, tmp_1_sva_7,
      STD_LOGIC_VECTOR'( S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm & butterFly_3_f1_asn_17
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm));
  tmp_3_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_26_sva, tmp_26_sva_1, tmp_13_sva_2,
      tmp_26_sva_10, tmp_13_sva_4, tmp_13_sva_5, tmp_13_sva_6, tmp_13_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm));
  tmp_5_lpi_4_dfm_mx0w0 <= MUX1HOT_v_32_8_2(tmp_26_sva_5, tmp_26_sva_6, tmp_22_sva_2,
      tmp_26_sva_8, tmp_22_sva_4, tmp_22_sva_5, tmp_22_sva_6, tmp_22_sva_7, STD_LOGIC_VECTOR'(
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm & butterFly_3_f1_asn_17 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
      & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm));
  butterFly_3_f1_asn_17 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND S6_OUTER_LOOP_for_nor_22_cse;
  modulo_sub_base_3_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_6_lpi_4_dfm)
      - SIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_2_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_4_lpi_4_dfm)
      - SIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_add_3_qr_lpi_4_dfm_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_1_sva)
      - UNSIGNED(m_sva), 32));
  modulo_sub_base_1_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_2_lpi_4_dfm)
      - SIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_lpi_4_dfm) - SIGNED(reg_mult_res_lpi_4_dfm_cse),
      32));
  S2_INNER_LOOP1_r_4_0_sva_2 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg),
      4), 5) + SIGNED'( "00001"), 5));
  modulo_sub_base_7_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_34_lpi_4_dfm)
      - SIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_6_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_32_lpi_4_dfm)
      - SIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_5_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_30_lpi_4_dfm)
      - SIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_4_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_28_lpi_4_dfm)
      - SIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_11_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_14_lpi_3_dfm)
      - SIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_10_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_12_lpi_3_dfm)
      - SIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_9_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_3_dfm)
      - SIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_8_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_8_lpi_3_dfm)
      - SIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  S1_OUTER_LOOP_k_5_0_sva_2 <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_UNSIGNED(UNSIGNED(reg_S2_COPY_LOOP_for_i_5_0_1_reg
      & reg_S2_COPY_LOOP_for_i_5_0_2_reg), 5), 6) + SIGNED'( "000001"), 6));
  modulo_sub_base_15_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_44_lpi_4_dfm)
      - SIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_14_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_42_lpi_4_dfm)
      - SIGNED(reg_mult_3_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_13_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_40_lpi_4_dfm)
      - SIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_12_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_38_lpi_4_dfm)
      - SIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_19_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_23_lpi_4_dfm)
      - SIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_17_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_19_lpi_4_dfm)
      - SIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_16_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_17_lpi_4_dfm)
      - SIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_23_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_52_lpi_3_dfm)
      - SIGNED(reg_mult_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_21_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_48_lpi_3_dfm)
      - SIGNED(reg_mult_2_res_lpi_4_dfm_cse), 32));
  modulo_sub_base_20_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_46_lpi_3_dfm)
      - SIGNED(reg_mult_1_res_lpi_4_dfm_cse), 32));
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))
      AND S1_OUTER_LOOP_for_nor_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      AND S1_OUTER_LOOP_for_nor_1_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))
      AND S1_OUTER_LOOP_for_nor_3_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      AND S1_OUTER_LOOP_for_nor_7_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND S1_OUTER_LOOP_for_nor_14_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58 <= (S1_OUTER_LOOP_for_acc_svs_3_0(2))
      AND S1_OUTER_LOOP_for_nor_28_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_66 <= (S1_OUTER_LOOP_for_acc_svs_3_0(3))
      AND S1_OUTER_LOOP_for_nor_32_itm;
  and_dcpl_42 <= S6_OUTER_LOOP_for_nor_22_cse AND (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  not_tmp_28 <= NOT((fsm_output(5)) AND (fsm_output(3)));
  nor_tmp_3 <= (fsm_output(4)) AND (fsm_output(1));
  nor_tmp_4 <= (fsm_output(2)) AND (fsm_output(4));
  or_tmp_35 <= (fsm_output(4)) OR (fsm_output(1));
  nor_tmp_8 <= (fsm_output(3)) AND (fsm_output(7));
  or_tmp_48 <= (fsm_output(5)) OR (fsm_output(7));
  or_tmp_59 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"))
      OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)));
  or_tmp_77 <= (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))) OR (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)));
  and_dcpl_53 <= (S2_INNER_LOOP1_r_4_0_sva_2(4)) AND S2_OUTER_LOOP_c_1_sva;
  and_dcpl_54 <= NOT((fsm_output(3)) OR (fsm_output(7)));
  or_4688_nl <= (fsm_output(6)) OR (NOT (fsm_output(1)));
  or_4689_nl <= (NOT (fsm_output(6))) OR (fsm_output(1));
  mux_100_cse <= MUX_s_1_2_2(or_4688_nl, or_4689_nl, fsm_output(5));
  and_dcpl_57 <= NOT(mux_100_cse OR (fsm_output(4)));
  and_dcpl_60 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_61 <= and_dcpl_60 AND nor_tmp_8;
  and_dcpl_64 <= nor_tmp_3 AND nor_1730_cse;
  and_dcpl_66 <= (NOT (fsm_output(2))) AND (fsm_output(0));
  and_dcpl_67 <= nor_tmp_3 AND and_dcpl_66;
  and_dcpl_69 <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00")));
  and_dcpl_70 <= and_dcpl_69 AND and_dcpl_54;
  and_dcpl_71 <= NOT((fsm_output(4)) OR (fsm_output(1)));
  and_dcpl_72 <= and_dcpl_71 AND nor_1730_cse;
  and_dcpl_74 <= (NOT (fsm_output(3))) AND (fsm_output(7));
  and_dcpl_75 <= and_dcpl_60 AND and_dcpl_74;
  and_dcpl_76 <= nor_tmp_3 AND and_2893_cse;
  and_dcpl_77 <= and_dcpl_76 AND and_dcpl_75;
  and_dcpl_79 <= (fsm_output(3)) AND (NOT (fsm_output(7)));
  and_dcpl_82 <= NOT((fsm_output(4)) OR (fsm_output(0)));
  nor_2165_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(5))) OR (fsm_output(2))
      OR (fsm_output(1)));
  nor_2166_nl <= NOT((fsm_output(3)) OR (fsm_output(5)) OR (NOT and_2141_cse));
  mux_112_nl <= MUX_s_1_2_2(nor_2165_nl, nor_2166_nl, fsm_output(7));
  and_dcpl_84 <= mux_112_nl AND and_dcpl_82 AND (NOT (fsm_output(6)));
  or_4696_nl <= (fsm_output(3)) OR (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(1))
      OR (fsm_output(4));
  or_4697_nl <= (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT and_1306_cse);
  mux_113_nl <= MUX_s_1_2_2(or_4696_nl, or_4697_nl, fsm_output(7));
  and_dcpl_86 <= NOT(mux_113_nl OR (fsm_output(0)) OR (fsm_output(5)));
  and_2095_nl <= (fsm_output(5)) AND (fsm_output(6)) AND (fsm_output(2)) AND (fsm_output(1));
  nor_2162_nl <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(2)) OR (fsm_output(1)));
  not_tmp_116 <= MUX_s_1_2_2(and_2095_nl, nor_2162_nl, fsm_output(3));
  and_dcpl_88 <= not_tmp_116 AND and_dcpl_82 AND (NOT (fsm_output(7)));
  and_dcpl_89 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_90 <= and_dcpl_89 AND and_dcpl_79;
  and_dcpl_91 <= (fsm_output(4)) AND (NOT (fsm_output(1)));
  and_dcpl_92 <= and_dcpl_91 AND and_dcpl_66;
  and_dcpl_93 <= and_dcpl_92 AND and_dcpl_90;
  or_tmp_131 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_134 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7)));
  or_320_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_318_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_121 <= MUX_s_1_2_2(or_320_nl, or_318_nl, fsm_output(1));
  or_331_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_329_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_127_nl <= MUX_s_1_2_2(or_tmp_131, or_329_nl, fsm_output(3));
  mux_tmp_128 <= MUX_s_1_2_2(or_331_nl, mux_127_nl, fsm_output(1));
  or_tmp_156 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_94 <= and_dcpl_69 AND and_dcpl_79;
  and_dcpl_95 <= (NOT (fsm_output(4))) AND (fsm_output(1));
  and_dcpl_96 <= and_dcpl_95 AND and_dcpl_66;
  and_dcpl_97 <= and_dcpl_96 AND and_dcpl_94;
  and_dcpl_98 <= NOT((fsm_output(2)) OR (fsm_output(5)));
  and_dcpl_99 <= and_dcpl_98 AND and_dcpl_54;
  or_tmp_166 <= (NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(4)));
  or_341_nl <= (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(4));
  mux_tmp_139 <= MUX_s_1_2_2(or_tmp_166, or_341_nl, fsm_output(6));
  and_dcpl_100 <= (NOT mux_tmp_139) AND and_dcpl_99;
  and_dcpl_101 <= and_dcpl_60 AND and_dcpl_79;
  and_dcpl_102 <= and_dcpl_64 AND and_dcpl_101;
  and_dcpl_103 <= (fsm_output(5)) AND (NOT (fsm_output(3)));
  and_dcpl_105 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND
      and_dcpl_103;
  or_tmp_169 <= (NOT (fsm_output(6))) OR (fsm_output(2)) OR (fsm_output(4));
  and_dcpl_107 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_108 <= and_dcpl_107 AND and_dcpl_54;
  and_dcpl_109 <= and_dcpl_96 AND and_dcpl_108;
  and_dcpl_110 <= (fsm_output(2)) AND (NOT (fsm_output(0)));
  and_dcpl_111 <= and_dcpl_95 AND and_dcpl_110;
  and_dcpl_112 <= and_dcpl_111 AND and_dcpl_108;
  and_dcpl_113 <= CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"));
  or_tmp_170 <= (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(2))
      OR (fsm_output(1));
  nand_502_nl <= NOT((fsm_output(3)) AND (fsm_output(6)) AND (fsm_output(0)) AND
      (fsm_output(2)) AND (fsm_output(1)));
  mux_141_nl <= MUX_s_1_2_2(nand_502_nl, or_tmp_170, fsm_output(7));
  and_dcpl_114 <= (NOT mux_141_nl) AND and_dcpl_113;
  and_dcpl_115 <= and_dcpl_69 AND nor_tmp_8;
  and_dcpl_116 <= and_dcpl_72 AND and_dcpl_115;
  and_dcpl_117 <= and_dcpl_103 AND (fsm_output(7));
  and_dcpl_119 <= and_dcpl_110 AND (NOT (fsm_output(6))) AND and_dcpl_117;
  and_dcpl_121 <= S6_OUTER_LOOP_for_nor_44_cse AND (NOT (S6_OUTER_LOOP_for_acc_tmp(0)));
  and_dcpl_123 <= nor_tmp_3 AND (NOT (S6_OUTER_LOOP_for_acc_tmp(4))) AND (NOT (S6_OUTER_LOOP_for_acc_tmp(2)));
  and_dcpl_125 <= and_dcpl_123 AND and_dcpl_121 AND and_dcpl_119;
  and_dcpl_126 <= and_dcpl_95 AND nor_1730_cse;
  and_dcpl_127 <= and_dcpl_126 AND and_dcpl_108;
  and_dcpl_128 <= and_dcpl_107 AND and_dcpl_79;
  and_dcpl_129 <= and_dcpl_76 AND and_dcpl_128;
  and_dcpl_130 <= and_dcpl_91 AND nor_1730_cse;
  and_dcpl_131 <= and_dcpl_130 AND and_dcpl_75;
  nor_tmp_31 <= (fsm_output(1)) AND (fsm_output(3)) AND (fsm_output(5));
  and_dcpl_135 <= (NOT (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2))) AND (fsm_output(5));
  and_dcpl_136 <= (fsm_output(4)) AND (NOT (reg_drf_revArr_ptr_1_smx_9_0_1_reg(1)));
  and_dcpl_137 <= and_dcpl_136 AND (NOT (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)));
  nor_2154_nl <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010")));
  mux_155_nl <= MUX_s_1_2_2(nor_2154_nl, and_2120_cse, fsm_output(6));
  nand_501_nl <= NOT((fsm_output(3)) AND mux_155_nl);
  mux_156_itm <= MUX_s_1_2_2(nand_501_nl, or_tmp_170, fsm_output(7));
  nor_tmp_35 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("11"));
  nor_tmp_36 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  and_dcpl_140 <= NOT((operator_20_true_28_acc_tmp(1)) OR (fsm_output(5)));
  and_dcpl_141 <= NOT((fsm_output(2)) OR (operator_20_true_28_acc_tmp(0)));
  and_dcpl_142 <= and_dcpl_141 AND (NOT (operator_20_true_28_acc_tmp(2)));
  nor_2150_nl <= NOT((fsm_output(3)) OR mux_tmp_139);
  nor_2151_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(0))
      OR (fsm_output(1)) OR (fsm_output(4)));
  not_tmp_149 <= MUX_s_1_2_2(nor_2150_nl, nor_2151_nl, fsm_output(7));
  or_dcpl_177 <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0));
  or_dcpl_178 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1));
  or_dcpl_179 <= or_dcpl_178 OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1));
  or_dcpl_180 <= or_dcpl_179 OR or_dcpl_177;
  or_tmp_207 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_405_nl <= (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_186 <= MUX_s_1_2_2(or_448_cse, or_405_nl, fsm_output(0));
  and_dcpl_148 <= and_dcpl_91 AND and_2893_cse;
  and_dcpl_149 <= and_dcpl_148 AND and_dcpl_101;
  and_dcpl_151 <= NOT((fsm_output(2)) OR (fsm_output(6)));
  and_dcpl_152 <= and_dcpl_151 AND and_dcpl_74;
  and_2083_cse <= (fsm_output(0)) AND (fsm_output(4));
  mux_tmp_193 <= MUX_s_1_2_2(and_dcpl_82, and_2083_cse, fsm_output(5));
  and_dcpl_154 <= mux_tmp_193 AND (fsm_output(1)) AND and_dcpl_152;
  and_dcpl_155 <= S6_OUTER_LOOP_for_nor_44_cse AND (S6_OUTER_LOOP_for_acc_tmp(0));
  and_dcpl_157 <= and_dcpl_123 AND and_dcpl_155 AND and_dcpl_119;
  and_dcpl_158 <= and_dcpl_69 AND and_dcpl_74;
  and_dcpl_162 <= NOT((reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) OR (fsm_output(6)));
  and_dcpl_164 <= S6_OUTER_LOOP_for_nor_22_cse AND and_dcpl_162;
  or_tmp_245 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (NOT nor_tmp_3);
  or_tmp_246 <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(4));
  and_2134_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 0)=STD_LOGIC_VECTOR'("111101"));
  mux_211_nl <= MUX_s_1_2_2(or_tmp_246, or_tmp_245, fsm_output(5));
  nor_2135_nl <= NOT((fsm_output(3)) OR mux_211_nl);
  not_tmp_169 <= MUX_s_1_2_2(and_2134_nl, nor_2135_nl, fsm_output(7));
  and_dcpl_168 <= not_tmp_149 AND and_dcpl_42 AND and_dcpl_98;
  or_dcpl_181 <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  or_dcpl_182 <= or_dcpl_179 OR or_dcpl_181;
  or_tmp_263 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_452_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_231 <= MUX_s_1_2_2(or_452_nl, or_435_cse, fsm_output(1));
  and_dcpl_170 <= and_dcpl_91 AND and_dcpl_110;
  and_dcpl_171 <= and_dcpl_170 AND and_dcpl_101;
  nor_2120_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(4)));
  nor_2121_nl <= NOT((fsm_output(0)) OR (NOT nor_tmp_3));
  mux_243_nl <= MUX_s_1_2_2(nor_2120_nl, nor_2121_nl, fsm_output(5));
  and_dcpl_173 <= mux_243_nl AND and_dcpl_152;
  and_dcpl_174 <= (S6_OUTER_LOOP_for_acc_tmp(1)) AND (NOT (S6_OUTER_LOOP_for_acc_tmp(3)));
  and_dcpl_175 <= and_dcpl_174 AND (NOT (S6_OUTER_LOOP_for_acc_tmp(0)));
  and_dcpl_177 <= and_dcpl_123 AND and_dcpl_175 AND and_dcpl_119;
  and_dcpl_178 <= and_dcpl_71 AND and_dcpl_66;
  and_dcpl_179 <= and_dcpl_178 AND and_dcpl_158;
  and_dcpl_180 <= and_dcpl_64 AND and_dcpl_75;
  or_tmp_301 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(4));
  nor_2117_nl <= NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("111100")));
  or_483_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT nor_tmp_3);
  mux_262_nl <= MUX_s_1_2_2(or_tmp_301, or_483_nl, fsm_output(5));
  nor_2118_nl <= NOT((fsm_output(3)) OR mux_262_nl);
  not_tmp_188 <= MUX_s_1_2_2(nor_2117_nl, nor_2118_nl, fsm_output(7));
  or_dcpl_183 <= or_dcpl_178 OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)));
  or_dcpl_184 <= or_dcpl_183 OR or_dcpl_177;
  or_tmp_317 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"));
  and_dcpl_184 <= and_dcpl_67 AND and_dcpl_101;
  and_dcpl_187 <= mux_tmp_193 AND (NOT (fsm_output(1))) AND and_dcpl_152;
  and_dcpl_188 <= and_dcpl_174 AND (S6_OUTER_LOOP_for_acc_tmp(0));
  and_dcpl_190 <= and_dcpl_123 AND and_dcpl_188 AND and_dcpl_119;
  and_dcpl_191 <= and_dcpl_72 AND and_dcpl_158;
  and_dcpl_192 <= and_dcpl_92 AND and_dcpl_75;
  mux_295_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_2881_cse);
  mux_296_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_2080_cse);
  mux_297_cse <= MUX_s_1_2_2(mux_296_cse, mux_295_cse, fsm_output(1));
  and_2057_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_2058_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_301_nl <= MUX_s_1_2_2(and_2057_nl, and_2058_nl, fsm_output(0));
  or_527_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_300_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_527_nl);
  mux_tmp_302 <= MUX_s_1_2_2(mux_301_nl, mux_300_nl, fsm_output(3));
  and_2054_nl <= (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(1))
      AND (fsm_output(4));
  or_534_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(4));
  mux_316_nl <= MUX_s_1_2_2(or_534_nl, or_tmp_166, fsm_output(5));
  nor_2101_nl <= NOT((fsm_output(3)) OR mux_316_nl);
  not_tmp_209 <= MUX_s_1_2_2(and_2054_nl, nor_2101_nl, fsm_output(7));
  or_dcpl_185 <= or_dcpl_183 OR or_dcpl_181;
  or_tmp_362 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_365 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7)));
  or_560_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_558_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_340 <= MUX_s_1_2_2(or_560_nl, or_558_nl, fsm_output(1));
  or_571_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_569_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_346_nl <= MUX_s_1_2_2(or_tmp_362, or_569_nl, fsm_output(3));
  mux_tmp_347 <= MUX_s_1_2_2(or_571_nl, mux_346_nl, fsm_output(1));
  or_tmp_386 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_199 <= nor_tmp_3 AND (NOT (S6_OUTER_LOOP_for_acc_tmp(4))) AND (S6_OUTER_LOOP_for_acc_tmp(2));
  and_dcpl_201 <= and_dcpl_199 AND and_dcpl_121 AND and_dcpl_119;
  and_dcpl_203 <= and_dcpl_136 AND (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0));
  nor_tmp_96 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  and_dcpl_206 <= (NOT (fsm_output(2))) AND (operator_20_true_28_acc_tmp(0));
  and_dcpl_207 <= and_dcpl_206 AND (NOT (operator_20_true_28_acc_tmp(2)));
  or_dcpl_186 <= (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))) OR (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1));
  or_dcpl_187 <= or_dcpl_186 OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1));
  or_dcpl_188 <= or_dcpl_187 OR or_dcpl_177;
  or_625_nl <= (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  or_623_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR (NOT (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  mux_tmp_391 <= MUX_s_1_2_2(or_625_nl, or_623_nl, reg_S2_COPY_LOOP_for_i_5_0_2_reg(2));
  or_648_nl <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  mux_tmp_403 <= MUX_s_1_2_2(or_686_cse, or_648_nl, fsm_output(0));
  and_dcpl_213 <= and_dcpl_199 AND and_dcpl_155 AND and_dcpl_119;
  and_dcpl_215 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (NOT (fsm_output(6)));
  and_dcpl_216 <= S6_OUTER_LOOP_for_nor_22_cse AND and_dcpl_215;
  and_dcpl_220 <= not_tmp_149 AND butterFly_3_f1_asn_17 AND and_dcpl_98;
  or_dcpl_189 <= or_dcpl_187 OR or_dcpl_181;
  or_tmp_493 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_693_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_445 <= MUX_s_1_2_2(or_693_nl, or_673_cse, fsm_output(1));
  and_dcpl_224 <= and_dcpl_199 AND and_dcpl_175 AND and_dcpl_119;
  or_dcpl_190 <= or_dcpl_186 OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)));
  or_dcpl_191 <= or_dcpl_190 OR or_dcpl_177;
  nand_480_cse <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  or_tmp_545 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR nand_480_cse;
  and_dcpl_230 <= and_dcpl_199 AND and_dcpl_188 AND and_dcpl_119;
  and_2014_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_2015_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0111"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_515_nl <= MUX_s_1_2_2(and_2014_nl, and_2015_nl, fsm_output(0));
  or_767_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_514_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_767_nl);
  mux_tmp_516 <= MUX_s_1_2_2(mux_515_nl, mux_514_nl, fsm_output(3));
  or_dcpl_192 <= or_dcpl_190 OR or_dcpl_181;
  or_tmp_595 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_598 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7)));
  or_800_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_798_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_549 <= MUX_s_1_2_2(or_800_nl, or_798_nl, fsm_output(1));
  or_811_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_809_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_555_nl <= MUX_s_1_2_2(or_tmp_595, or_809_nl, fsm_output(3));
  mux_tmp_556 <= MUX_s_1_2_2(or_811_nl, mux_555_nl, fsm_output(1));
  or_tmp_620 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_236 <= (NOT (S6_OUTER_LOOP_for_acc_tmp(1))) AND (S6_OUTER_LOOP_for_acc_tmp(3));
  and_dcpl_237 <= and_dcpl_236 AND (NOT (S6_OUTER_LOOP_for_acc_tmp(0)));
  and_dcpl_239 <= and_dcpl_123 AND and_dcpl_237 AND and_dcpl_119;
  and_dcpl_241 <= (fsm_output(4)) AND (reg_drf_revArr_ptr_1_smx_9_0_1_reg(1));
  and_dcpl_242 <= and_dcpl_241 AND (NOT (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)));
  nor_tmp_165 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  and_dcpl_245 <= (operator_20_true_28_acc_tmp(1)) AND (NOT (fsm_output(5)));
  or_dcpl_193 <= (NOT (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0));
  or_dcpl_194 <= or_dcpl_179 OR or_dcpl_193;
  or_874_nl <= (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_609 <= MUX_s_1_2_2(or_911_cse, or_874_nl, fsm_output(0));
  and_dcpl_250 <= and_dcpl_236 AND (S6_OUTER_LOOP_for_acc_tmp(0));
  and_dcpl_252 <= and_dcpl_123 AND and_dcpl_250 AND and_dcpl_119;
  and_dcpl_254 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_255 <= and_dcpl_254 AND and_dcpl_162;
  and_dcpl_257 <= and_dcpl_254 AND (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  and_dcpl_259 <= not_tmp_149 AND and_dcpl_257 AND and_dcpl_98;
  or_dcpl_195 <= NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  or_dcpl_196 <= or_dcpl_179 OR or_dcpl_195;
  or_915_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_651 <= MUX_s_1_2_2(or_915_nl, or_898_cse, fsm_output(1));
  and_dcpl_262 <= (S6_OUTER_LOOP_for_acc_tmp(1)) AND (S6_OUTER_LOOP_for_acc_tmp(3));
  and_dcpl_263 <= and_dcpl_262 AND (NOT (S6_OUTER_LOOP_for_acc_tmp(0)));
  and_dcpl_265 <= and_dcpl_123 AND and_dcpl_263 AND and_dcpl_119;
  or_dcpl_197 <= or_dcpl_183 OR or_dcpl_193;
  or_tmp_759 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"));
  and_dcpl_270 <= and_dcpl_262 AND (S6_OUTER_LOOP_for_acc_tmp(0));
  and_dcpl_272 <= and_dcpl_123 AND and_dcpl_270 AND and_dcpl_119;
  and_1972_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1973_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_718_nl <= MUX_s_1_2_2(and_1972_nl, and_1973_nl, fsm_output(0));
  or_988_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_717_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_988_nl);
  mux_tmp_719 <= MUX_s_1_2_2(mux_718_nl, mux_717_nl, fsm_output(3));
  or_dcpl_198 <= or_dcpl_183 OR or_dcpl_195;
  or_tmp_806 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_809 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7)));
  or_1017_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1015_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_755 <= MUX_s_1_2_2(or_1017_nl, or_1015_nl, fsm_output(1));
  or_1028_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1026_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(7));
  mux_761_nl <= MUX_s_1_2_2(or_tmp_806, or_1026_nl, fsm_output(3));
  mux_tmp_762 <= MUX_s_1_2_2(or_1028_nl, mux_761_nl, fsm_output(1));
  or_tmp_830 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_279 <= and_dcpl_199 AND and_dcpl_237 AND and_dcpl_119;
  and_dcpl_281 <= and_dcpl_241 AND (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0));
  nor_tmp_225 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  or_dcpl_199 <= or_dcpl_187 OR or_dcpl_193;
  or_tmp_875 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  not_tmp_389 <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  or_1097_nl <= (fsm_output(1)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  mux_tmp_815 <= MUX_s_1_2_2(or_1135_cse, or_1097_nl, fsm_output(0));
  and_dcpl_289 <= and_dcpl_199 AND and_dcpl_250 AND and_dcpl_119;
  and_dcpl_291 <= and_dcpl_254 AND and_dcpl_215;
  and_dcpl_293 <= and_dcpl_254 AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0));
  and_dcpl_295 <= not_tmp_149 AND and_dcpl_293 AND and_dcpl_98;
  or_dcpl_200 <= or_dcpl_187 OR or_dcpl_195;
  or_tmp_931 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_1142_nl <= (NOT (fsm_output(0))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR
      not_tmp_389;
  or_1140_nl <= (fsm_output(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  mux_tmp_857 <= MUX_s_1_2_2(or_1142_nl, or_1140_nl, fsm_output(1));
  and_dcpl_299 <= and_dcpl_199 AND and_dcpl_263 AND and_dcpl_119;
  or_dcpl_201 <= or_dcpl_190 OR or_dcpl_193;
  or_tmp_982 <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)) OR (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"))));
  and_dcpl_305 <= and_dcpl_199 AND and_dcpl_270 AND and_dcpl_119;
  and_1923_nl <= ((CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4) AND (fsm_output(5))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1925_nl <= ((CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) AND (fsm_output(5))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_927_nl <= MUX_s_1_2_2(and_1923_nl, and_1925_nl, fsm_output(0));
  nand_442_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4) AND (NOT (fsm_output(5))));
  mux_926_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_442_nl);
  mux_tmp_928 <= MUX_s_1_2_2(mux_927_nl, mux_926_nl, fsm_output(3));
  or_dcpl_202 <= or_dcpl_190 OR or_dcpl_195;
  or_tmp_1030 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_1033 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7)));
  or_1245_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1243_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_962 <= MUX_s_1_2_2(or_1245_nl, or_1243_nl, fsm_output(1));
  or_1255_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1253_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_968_nl <= MUX_s_1_2_2(or_tmp_1030, or_1253_nl, fsm_output(3));
  mux_tmp_969 <= MUX_s_1_2_2(or_1255_nl, mux_968_nl, fsm_output(1));
  or_tmp_1054 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  not_tmp_451 <= NOT((S6_OUTER_LOOP_for_acc_tmp(4)) OR (NOT (fsm_output(4))));
  and_dcpl_312 <= nor_tmp_3 AND (S6_OUTER_LOOP_for_acc_tmp(4)) AND (NOT (S6_OUTER_LOOP_for_acc_tmp(2)));
  and_dcpl_314 <= and_dcpl_312 AND and_dcpl_121 AND and_dcpl_119;
  or_tmp_1079 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  and_dcpl_316 <= (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2)) AND (fsm_output(5));
  nor_tmp_299 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  and_dcpl_319 <= and_dcpl_141 AND (operator_20_true_28_acc_tmp(2));
  or_dcpl_203 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)));
  or_dcpl_204 <= or_dcpl_203 OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1));
  or_dcpl_205 <= or_dcpl_204 OR or_dcpl_177;
  or_tmp_1110 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  or_1322_nl <= (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_1025 <= MUX_s_1_2_2(or_1358_cse, or_1322_nl, fsm_output(0));
  and_dcpl_325 <= and_dcpl_312 AND and_dcpl_155 AND and_dcpl_119;
  or_tmp_1133 <= (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  and_dcpl_327 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_328 <= and_dcpl_327 AND and_dcpl_162;
  and_dcpl_330 <= and_dcpl_327 AND (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  and_dcpl_332 <= not_tmp_149 AND and_dcpl_330 AND and_dcpl_98;
  or_dcpl_206 <= or_dcpl_204 OR or_dcpl_181;
  or_1362_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_1069 <= MUX_s_1_2_2(or_1362_nl, or_1344_cse, fsm_output(1));
  or_tmp_1162 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  and_dcpl_336 <= and_dcpl_312 AND and_dcpl_175 AND and_dcpl_119;
  or_tmp_1185 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  or_dcpl_207 <= or_dcpl_203 OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)));
  or_dcpl_208 <= or_dcpl_207 OR or_dcpl_177;
  or_tmp_1200 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  or_tmp_1212 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  and_dcpl_342 <= and_dcpl_312 AND and_dcpl_188 AND and_dcpl_119;
  and_1879_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1880_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1141_nl <= MUX_s_1_2_2(and_1879_nl, and_1880_nl, fsm_output(0));
  or_1439_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5));
  mux_1140_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1439_nl);
  mux_tmp_1142 <= MUX_s_1_2_2(mux_1141_nl, mux_1140_nl, fsm_output(3));
  or_tmp_1235 <= (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  or_dcpl_209 <= or_dcpl_207 OR or_dcpl_181;
  or_tmp_1248 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_1251 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7)));
  or_1470_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1468_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1179 <= MUX_s_1_2_2(or_1470_nl, or_1468_nl, fsm_output(1));
  or_1480_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1478_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1185_nl <= MUX_s_1_2_2(or_tmp_1248, or_1478_nl, fsm_output(3));
  mux_tmp_1186 <= MUX_s_1_2_2(or_1480_nl, mux_1185_nl, fsm_output(1));
  or_tmp_1271 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  not_tmp_542 <= (NOT((S6_OUTER_LOOP_for_acc_tmp(2)) AND (S6_OUTER_LOOP_for_acc_tmp(4))))
      AND (fsm_output(4));
  and_dcpl_349 <= nor_tmp_3 AND (S6_OUTER_LOOP_for_acc_tmp(4)) AND (S6_OUTER_LOOP_for_acc_tmp(2));
  and_dcpl_351 <= and_dcpl_349 AND and_dcpl_121 AND and_dcpl_119;
  not_tmp_551 <= NOT(S1_OUTER_LOOP_for_acc_svs_4 AND (S1_OUTER_LOOP_for_acc_svs_3_0(2)));
  or_tmp_1298 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR nand_508_cse;
  nor_tmp_366 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  and_dcpl_355 <= and_dcpl_206 AND (operator_20_true_28_acc_tmp(2));
  or_dcpl_210 <= NOT((reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) AND (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)));
  or_dcpl_211 <= or_dcpl_210 OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1));
  or_dcpl_212 <= or_dcpl_211 OR or_dcpl_177;
  or_tmp_1316 <= (NOT (fsm_output(1))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_tmp_1319 <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_tmp_1324 <= (or_1527_cse AND (fsm_output(1))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  or_tmp_1340 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  nand_546_nl <= NOT((fsm_output(1)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101")));
  or_1559_nl <= (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_tmp_1243 <= MUX_s_1_2_2(nand_546_nl, or_1559_nl, fsm_output(0));
  and_dcpl_361 <= and_dcpl_349 AND and_dcpl_155 AND and_dcpl_119;
  or_tmp_1363 <= (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR nand_508_cse;
  and_dcpl_363 <= and_dcpl_327 AND and_dcpl_215;
  and_dcpl_365 <= and_dcpl_327 AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0));
  and_dcpl_367 <= not_tmp_149 AND and_dcpl_365 AND and_dcpl_98;
  or_dcpl_213 <= or_dcpl_211 OR or_dcpl_181;
  or_tmp_1379 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  not_tmp_590 <= NOT((reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)));
  or_1604_nl <= (NOT (fsm_output(0))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR
      not_tmp_590;
  or_1602_nl <= (fsm_output(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR not_tmp_590;
  mux_tmp_1287 <= MUX_s_1_2_2(or_1604_nl, or_1602_nl, fsm_output(1));
  or_tmp_1397 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110")) OR (NOT
      S1_OUTER_LOOP_for_acc_svs_4);
  not_tmp_598 <= (NOT((S6_OUTER_LOOP_for_acc_tmp(1)) AND (S6_OUTER_LOOP_for_acc_tmp(2))
      AND (S6_OUTER_LOOP_for_acc_tmp(4)))) AND (fsm_output(4));
  and_dcpl_371 <= and_dcpl_349 AND and_dcpl_175 AND and_dcpl_119;
  or_tmp_1422 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR nand_508_cse;
  or_dcpl_214 <= or_dcpl_210 OR (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)));
  or_dcpl_215 <= or_dcpl_214 OR or_dcpl_177;
  or_tmp_1437 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR nand_480_cse;
  or_tmp_1452 <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"))
      AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111")) AND
      S1_OUTER_LOOP_for_acc_svs_4);
  and_dcpl_377 <= and_dcpl_349 AND and_dcpl_188 AND and_dcpl_119;
  and_1831_nl <= ((CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5))) OR (fsm_output(7))) AND
      (fsm_output(6));
  and_1833_nl <= ((CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("0111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (fsm_output(5))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1362_nl <= MUX_s_1_2_2(and_1831_nl, and_1833_nl, fsm_output(0));
  nand_408_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (NOT (fsm_output(5))));
  mux_1361_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_408_nl);
  mux_tmp_1363 <= MUX_s_1_2_2(mux_1362_nl, mux_1361_nl, fsm_output(3));
  or_tmp_1479 <= (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR nand_508_cse;
  or_dcpl_216 <= or_dcpl_214 OR or_dcpl_181;
  or_tmp_1492 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("01"));
  or_tmp_1495 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(7)));
  or_1721_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1719_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1397 <= MUX_s_1_2_2(or_1721_nl, or_1719_nl, fsm_output(1));
  or_1731_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1729_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1403_nl <= MUX_s_1_2_2(or_tmp_1492, or_1729_nl, fsm_output(3));
  mux_tmp_1404 <= MUX_s_1_2_2(or_1731_nl, mux_1403_nl, fsm_output(1));
  or_tmp_1516 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_384 <= and_dcpl_312 AND and_dcpl_237 AND and_dcpl_119;
  or_tmp_1540 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  nor_tmp_445 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  or_dcpl_217 <= or_dcpl_204 OR or_dcpl_193;
  or_tmp_1558 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_tmp_1572 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_520_cse;
  or_1796_nl <= (fsm_output(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_tmp_1460 <= MUX_s_1_2_2(nand_393_cse, or_1796_nl, fsm_output(0));
  and_dcpl_393 <= and_dcpl_312 AND and_dcpl_250 AND and_dcpl_119;
  or_tmp_1595 <= (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  and_dcpl_395 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_396 <= and_dcpl_395 AND and_dcpl_162;
  and_dcpl_398 <= and_dcpl_395 AND (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  and_dcpl_400 <= not_tmp_149 AND and_dcpl_398 AND and_dcpl_98;
  or_dcpl_218 <= or_dcpl_204 OR or_dcpl_195;
  or_tmp_1610 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  nand_396_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  mux_tmp_1504 <= MUX_s_1_2_2(nand_396_nl, or_1818_cse, fsm_output(1));
  or_tmp_1624 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("010"))
      OR nand_520_cse;
  and_dcpl_404 <= and_dcpl_312 AND and_dcpl_263 AND and_dcpl_119;
  or_tmp_1647 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  or_dcpl_219 <= or_dcpl_207 OR or_dcpl_193;
  or_tmp_1662 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  or_tmp_1677 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("011"))
      OR nand_520_cse;
  and_dcpl_410 <= and_dcpl_312 AND and_dcpl_270 AND and_dcpl_119;
  and_1777_nl <= ((CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1011"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5))) OR (fsm_output(7))) AND
      (fsm_output(6));
  and_1779_nl <= ((CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1011"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (fsm_output(5))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1576_nl <= MUX_s_1_2_2(and_1777_nl, and_1779_nl, fsm_output(0));
  nand_380_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1011"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (NOT (fsm_output(5))));
  mux_1575_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_380_nl);
  mux_tmp_1577 <= MUX_s_1_2_2(mux_1576_nl, mux_1575_nl, fsm_output(3));
  or_tmp_1703 <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))));
  or_dcpl_220 <= or_dcpl_207 OR or_dcpl_195;
  or_tmp_1716 <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01")));
  or_tmp_1719 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(7)));
  or_1949_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"));
  or_1947_nl <= (NOT (fsm_output(3))) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  mux_tmp_1614 <= MUX_s_1_2_2(or_1949_nl, or_1947_nl, fsm_output(1));
  nand_518_nl <= NOT((fsm_output(3)) AND CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10")));
  or_1957_nl <= (fsm_output(6)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7));
  mux_1620_nl <= MUX_s_1_2_2(or_tmp_1716, or_1957_nl, fsm_output(3));
  mux_tmp_1621 <= MUX_s_1_2_2(nand_518_nl, mux_1620_nl, fsm_output(1));
  or_tmp_1739 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("111"))
      OR CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  and_dcpl_417 <= and_dcpl_349 AND and_dcpl_237 AND and_dcpl_119;
  not_tmp_741 <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)));
  or_tmp_1765 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_741;
  nor_tmp_525 <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)))) OR (fsm_output(7))) AND (fsm_output(6));
  or_dcpl_221 <= or_dcpl_211 OR or_dcpl_193;
  or_tmp_1783 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) OR not_tmp_590;
  or_tmp_1796 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_517_cse;
  or_2025_nl <= (fsm_output(1)) OR nand_480_cse;
  mux_tmp_1677 <= MUX_s_1_2_2(nand_336_cse, or_2025_nl, fsm_output(0));
  and_dcpl_426 <= and_dcpl_349 AND and_dcpl_250 AND and_dcpl_119;
  or_tmp_1818 <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_741;
  and_dcpl_428 <= and_dcpl_395 AND and_dcpl_215;
  and_dcpl_430 <= and_dcpl_395 AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0));
  and_dcpl_432 <= not_tmp_149 AND and_dcpl_430 AND and_dcpl_98;
  or_dcpl_222 <= or_dcpl_211 OR or_dcpl_195;
  or_tmp_1833 <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  nand_353_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  or_2062_nl <= (fsm_output(0)) OR nand_480_cse;
  mux_tmp_1721 <= MUX_s_1_2_2(nand_353_nl, or_2062_nl, fsm_output(1));
  or_tmp_1845 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR nand_351_cse;
  and_dcpl_436 <= and_dcpl_349 AND and_dcpl_263 AND and_dcpl_119;
  or_tmp_1867 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))));
  or_dcpl_223 <= or_dcpl_214 OR or_dcpl_193;
  and_dcpl_442 <= and_dcpl_349 AND and_dcpl_270 AND and_dcpl_119;
  and_1699_nl <= ((CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5))) OR (fsm_output(7))) AND
      (fsm_output(6));
  and_1701_nl <= ((CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (fsm_output(5))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1792_nl <= MUX_s_1_2_2(and_1699_nl, and_1701_nl, fsm_output(0));
  nand_335_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (NOT (fsm_output(5))));
  mux_1791_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_335_nl);
  mux_tmp_1793 <= MUX_s_1_2_2(mux_1792_nl, mux_1791_nl, fsm_output(3));
  or_2140_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  or_2139_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_tmp_1820 <= MUX_s_1_2_2(or_2140_nl, or_2139_nl, fsm_output(0));
  or_2142_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  or_2141_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_1821 <= MUX_s_1_2_2(or_2142_nl, or_2141_nl, fsm_output(1));
  or_tmp_1918 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  or_tmp_1924 <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_1832 <= MUX_s_1_2_2(or_4679_cse, or_tmp_1924, fsm_output(1));
  or_tmp_1928 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  and_dcpl_447 <= and_dcpl_71 AND and_dcpl_110;
  and_dcpl_448 <= and_dcpl_447 AND and_dcpl_70;
  and_dcpl_449 <= and_dcpl_71 AND and_2893_cse;
  and_dcpl_450 <= and_dcpl_449 AND and_dcpl_70;
  and_dcpl_451 <= and_dcpl_72 AND and_dcpl_94;
  nor_1740_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(0)))
      OR (fsm_output(4)));
  nor_1741_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (fsm_output(0))
      OR (NOT (fsm_output(4))));
  not_tmp_833 <= MUX_s_1_2_2(nor_1740_nl, nor_1741_nl, fsm_output(7));
  and_dcpl_454 <= not_tmp_833 AND nor_2178_cse_1 AND (NOT (fsm_output(6)));
  mux_1845_nl <= MUX_s_1_2_2(nand_568_cse, or_4797_cse, fsm_output(7));
  and_dcpl_456 <= NOT(mux_1845_nl OR (fsm_output(4)));
  and_dcpl_457 <= and_dcpl_456 AND nor_1730_cse AND and_dcpl_60;
  and_dcpl_458 <= and_dcpl_89 AND and_dcpl_54;
  and_dcpl_459 <= and_dcpl_64 AND and_dcpl_458;
  and_dcpl_460 <= (NOT (fsm_output(5))) AND (fsm_output(3));
  and_dcpl_461 <= and_dcpl_460 AND (NOT (fsm_output(7)));
  and_dcpl_462 <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (fsm_output(0)));
  and_dcpl_464 <= and_dcpl_462 AND (fsm_output(6)) AND and_dcpl_461;
  and_dcpl_466 <= S1_OUTER_LOOP_for_nor_76_cse AND (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)));
  and_dcpl_467 <= NOT((fsm_output(2)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)));
  and_dcpl_468 <= and_dcpl_91 AND and_dcpl_467;
  and_dcpl_469 <= and_dcpl_468 AND and_dcpl_466;
  and_dcpl_470 <= and_dcpl_469 AND and_dcpl_464;
  and_dcpl_472 <= nor_1730_cse AND (fsm_output(6)) AND and_dcpl_461;
  and_dcpl_475 <= and_dcpl_178 AND and_dcpl_128;
  and_dcpl_476 <= and_dcpl_95 AND and_2893_cse;
  and_dcpl_477 <= and_dcpl_476 AND and_dcpl_128;
  and_dcpl_478 <= and_dcpl_60 AND and_dcpl_54;
  and_dcpl_479 <= and_dcpl_178 AND and_dcpl_478;
  and_dcpl_480 <= and_dcpl_130 AND and_dcpl_115;
  and_dcpl_483 <= NOT((reg_drf_revArr_ptr_1_smx_9_0_1_reg(2)) OR (fsm_output(2)));
  and_dcpl_484 <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  or_2184_nl <= (NOT (fsm_output(6))) OR (fsm_output(0)) OR (NOT nor_tmp_3);
  or_2182_nl <= (fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (fsm_output(4));
  mux_1863_nl <= MUX_s_1_2_2(or_2184_nl, or_2182_nl, fsm_output(5));
  nor_1732_nl <= NOT((fsm_output(3)) OR mux_1863_nl);
  nor_1733_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(0)) OR (fsm_output(1)) OR (NOT (fsm_output(4))));
  not_tmp_843 <= MUX_s_1_2_2(nor_1732_nl, nor_1733_nl, fsm_output(7));
  and_dcpl_488 <= and_dcpl_462 AND (NOT (fsm_output(6))) AND and_dcpl_461;
  and_dcpl_489 <= and_dcpl_71 AND and_dcpl_467;
  and_dcpl_490 <= and_dcpl_489 AND and_dcpl_466;
  and_dcpl_492 <= (NOT (operator_20_true_28_acc_tmp(1))) AND (fsm_output(5));
  and_dcpl_493 <= NOT((fsm_output(4)) OR (operator_20_true_28_acc_tmp(0)));
  and_dcpl_494 <= and_dcpl_493 AND (NOT (operator_20_true_28_acc_tmp(2)));
  and_dcpl_497 <= NOT((S34_OUTER_LOOP_for_a_acc_2_tmp(0)) OR (fsm_output(0)));
  and_dcpl_499 <= S1_OUTER_LOOP_for_nor_90_cse AND (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(1)));
  and_dcpl_501 <= and_dcpl_499 AND and_dcpl_497 AND and_dcpl_90;
  and_dcpl_503 <= and_dcpl_91 AND (NOT (fsm_output(2))) AND (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(2)));
  or_dcpl_225 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"));
  or_dcpl_226 <= (S34_OUTER_LOOP_for_a_acc_2_tmp(2)) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(4));
  or_dcpl_227 <= or_dcpl_226 OR (S34_OUTER_LOOP_for_a_acc_2_tmp(3));
  or_tmp_1976 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2204_cse <= (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_2208_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_2207_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1886_nl <= MUX_s_1_2_2(or_2208_nl, or_2207_nl, fsm_output(1));
  or_2209_nl <= (fsm_output(4)) OR mux_1886_nl;
  or_2206_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_1883_nl <= MUX_s_1_2_2(or_tmp_1976, or_2204_cse, fsm_output(0));
  nand_112_nl <= NOT((fsm_output(3)) AND (NOT mux_1883_nl));
  mux_1884_nl <= MUX_s_1_2_2(or_2206_nl, nand_112_nl, fsm_output(1));
  or_2203_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1885_nl <= MUX_s_1_2_2(mux_1884_nl, or_2203_nl, fsm_output(4));
  mux_tmp_1887 <= MUX_s_1_2_2(or_2209_nl, mux_1885_nl, fsm_output(6));
  or_tmp_1981 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_tmp_1983 <= (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_4685_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 0)/=STD_LOGIC_VECTOR'("100100"));
  or_4686_nl <= (NOT (fsm_output(3))) OR (fsm_output(5)) OR (NOT (fsm_output(0)))
      OR (fsm_output(2)) OR (NOT nor_tmp_3);
  mux_1903_nl <= MUX_s_1_2_2(or_4685_nl, or_4686_nl, fsm_output(7));
  and_dcpl_506 <= NOT(mux_1903_nl OR (fsm_output(6)));
  and_dcpl_507 <= and_dcpl_148 AND and_dcpl_458;
  and_dcpl_508 <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) AND (NOT (fsm_output(0)));
  and_dcpl_510 <= and_dcpl_508 AND (fsm_output(6)) AND and_dcpl_461;
  and_dcpl_511 <= and_dcpl_469 AND and_dcpl_510;
  nand_532_nl <= NOT((fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(2)) AND
      (NOT (fsm_output(1))) AND (fsm_output(4)));
  or_2238_nl <= (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(1))
      OR (fsm_output(4));
  mux_1915_nl <= MUX_s_1_2_2(nand_532_nl, or_2238_nl, fsm_output(5));
  nor_1717_nl <= NOT((fsm_output(3)) OR mux_1915_nl);
  nor_1718_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (fsm_output(6))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (NOT nor_tmp_3));
  not_tmp_865 <= MUX_s_1_2_2(nor_1717_nl, nor_1718_nl, fsm_output(7));
  and_dcpl_519 <= and_dcpl_508 AND (NOT (fsm_output(6))) AND and_dcpl_461;
  and_dcpl_521 <= (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))) AND (fsm_output(5));
  and_dcpl_522 <= NOT((fsm_output(4)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)));
  and_dcpl_523 <= and_dcpl_522 AND (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)));
  and_dcpl_525 <= (NOT mux_156_itm) AND and_dcpl_523 AND and_dcpl_521;
  and_dcpl_526 <= (S34_OUTER_LOOP_for_a_acc_2_tmp(0)) AND (NOT (fsm_output(0)));
  and_dcpl_528 <= and_dcpl_499 AND and_dcpl_526 AND and_dcpl_90;
  or_dcpl_229 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"));
  nor_1712_cse <= NOT((fsm_output(3)) OR (fsm_output(0)));
  or_2262_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_2261_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1937_nl <= MUX_s_1_2_2(or_2262_nl, or_2261_nl, fsm_output(1));
  or_2259_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_2258_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1935_nl <= MUX_s_1_2_2(or_2259_nl, or_2258_nl, fsm_output(3));
  nor_1713_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  nor_1714_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  mux_1934_nl <= MUX_s_1_2_2(nor_1713_nl, nor_1714_nl, fsm_output(0));
  nand_115_nl <= NOT((fsm_output(3)) AND mux_1934_nl);
  mux_1936_nl <= MUX_s_1_2_2(mux_1935_nl, nand_115_nl, fsm_output(1));
  mux_tmp_1938 <= MUX_s_1_2_2(mux_1937_nl, mux_1936_nl, fsm_output(6));
  or_tmp_2035 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  and_dcpl_533 <= not_tmp_833 AND (fsm_output(1)) AND (NOT (fsm_output(2))) AND (NOT
      (fsm_output(6)));
  and_dcpl_534 <= and_dcpl_170 AND and_dcpl_458;
  and_dcpl_535 <= S1_OUTER_LOOP_for_nor_76_cse AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1));
  and_dcpl_536 <= and_dcpl_468 AND and_dcpl_535;
  and_dcpl_537 <= and_dcpl_536 AND and_dcpl_464;
  and_dcpl_540 <= and_dcpl_96 AND and_dcpl_478;
  and_dcpl_541 <= and_dcpl_64 AND and_dcpl_115;
  and_1666_nl <= ((NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))) OR (NOT (fsm_output(3)))))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2277_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_1956_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2277_nl);
  or_2276_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_1955_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2276_nl);
  mux_1957_nl <= MUX_s_1_2_2(mux_1956_nl, mux_1955_nl, fsm_output(0));
  mux_tmp_1958 <= MUX_s_1_2_2(and_1666_nl, mux_1957_nl, fsm_output(2));
  or_2289_nl <= (NOT (fsm_output(6))) OR (fsm_output(0)) OR (NOT (fsm_output(2)))
      OR (fsm_output(1)) OR (NOT (fsm_output(4)));
  or_2287_nl <= (fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(2)) OR (NOT
      (fsm_output(1))) OR (fsm_output(4));
  mux_1973_nl <= MUX_s_1_2_2(or_2289_nl, or_2287_nl, fsm_output(5));
  nor_1706_nl <= NOT((fsm_output(3)) OR mux_1973_nl);
  nor_1707_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (fsm_output(6))
      OR (fsm_output(0)) OR (fsm_output(2)) OR (NOT nor_tmp_3));
  not_tmp_874 <= MUX_s_1_2_2(nor_1706_nl, nor_1707_nl, fsm_output(7));
  and_dcpl_544 <= and_dcpl_489 AND and_dcpl_535;
  and_dcpl_546 <= S1_OUTER_LOOP_for_nor_90_cse AND (S34_OUTER_LOOP_for_a_acc_2_tmp(1));
  and_dcpl_548 <= and_dcpl_546 AND and_dcpl_497 AND and_dcpl_90;
  or_dcpl_231 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("10"));
  or_tmp_2071 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  or_tmp_2075 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_tmp_2076 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_1993_nl <= MUX_s_1_2_2(or_tmp_2075, or_2204_cse, fsm_output(0));
  mux_1994_nl <= MUX_s_1_2_2(or_tmp_2076, mux_1993_nl, fsm_output(1));
  nand_117_nl <= NOT((fsm_output(3)) AND (NOT mux_1994_nl));
  mux_1995_nl <= MUX_s_1_2_2(or_395_cse, nand_117_nl, fsm_output(6));
  or_2306_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_1996 <= MUX_s_1_2_2(mux_1995_nl, or_2306_nl, fsm_output(4));
  or_2312_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_tmp_1999 <= MUX_s_1_2_2(or_2312_nl, or_tmp_2071, fsm_output(1));
  nor_1701_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(5))) OR (fsm_output(0))
      OR (NOT (fsm_output(1))) OR (fsm_output(4)));
  nor_1702_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (NOT (fsm_output(0)))
      OR (fsm_output(1)) OR (NOT (fsm_output(4))));
  mux_2011_nl <= MUX_s_1_2_2(nor_1701_nl, nor_1702_nl, fsm_output(7));
  and_dcpl_551 <= mux_2011_nl AND and_dcpl_151;
  and_dcpl_552 <= and_dcpl_67 AND and_dcpl_458;
  and_dcpl_553 <= and_dcpl_536 AND and_dcpl_510;
  and_dcpl_556 <= and_dcpl_126 AND and_dcpl_478;
  and_dcpl_557 <= and_dcpl_92 AND and_dcpl_115;
  and_1656_nl <= ((NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))) OR (NOT (fsm_output(3)))))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2323_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2017_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2323_nl);
  or_2322_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2016_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2322_nl);
  mux_2018_nl <= MUX_s_1_2_2(mux_2017_nl, mux_2016_nl, fsm_output(0));
  mux_tmp_2019 <= MUX_s_1_2_2(and_1656_nl, mux_2018_nl, fsm_output(2));
  and_dcpl_559 <= NOT((reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) OR (fsm_output(2)));
  nor_tmp_674 <= (fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(1)) AND (fsm_output(4));
  or_2333_nl <= (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(1))) OR (fsm_output(4));
  mux_2034_nl <= MUX_s_1_2_2((NOT nor_tmp_674), or_2333_nl, fsm_output(5));
  nor_1695_nl <= NOT((fsm_output(3)) OR mux_2034_nl);
  nor_1696_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(5)) OR (fsm_output(6))
      OR (NOT (fsm_output(0))) OR (fsm_output(1)) OR (NOT (fsm_output(4))));
  not_tmp_890 <= MUX_s_1_2_2(nor_1695_nl, nor_1696_nl, fsm_output(7));
  and_dcpl_564 <= and_dcpl_546 AND and_dcpl_526 AND and_dcpl_90;
  or_dcpl_233 <= NOT(CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11")));
  or_2349_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  or_2348_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_tmp_2052 <= MUX_s_1_2_2(or_2349_nl, or_2348_nl, fsm_output(0));
  or_2351_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  or_2350_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2053 <= MUX_s_1_2_2(or_2351_nl, or_2350_nl, fsm_output(1));
  or_tmp_2119 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  or_tmp_2122 <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2064 <= MUX_s_1_2_2(or_4679_cse, or_tmp_2122, fsm_output(1));
  or_tmp_2126 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  and_dcpl_567 <= (NOT (fsm_output(2))) AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2));
  and_dcpl_568 <= and_dcpl_91 AND and_dcpl_567;
  and_dcpl_569 <= and_dcpl_568 AND and_dcpl_466;
  and_dcpl_570 <= and_dcpl_569 AND and_dcpl_464;
  and_dcpl_574 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_577 <= and_dcpl_71 AND and_dcpl_567;
  and_dcpl_578 <= and_dcpl_577 AND and_dcpl_466;
  and_dcpl_580 <= (NOT (fsm_output(4))) AND (operator_20_true_28_acc_tmp(0));
  and_dcpl_581 <= and_dcpl_580 AND (NOT (operator_20_true_28_acc_tmp(2)));
  and_dcpl_585 <= and_dcpl_91 AND (NOT (fsm_output(2))) AND (S34_OUTER_LOOP_for_a_acc_2_tmp(2));
  or_dcpl_235 <= (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(2))) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(4));
  or_dcpl_236 <= or_dcpl_235 OR (S34_OUTER_LOOP_for_a_acc_2_tmp(3));
  or_tmp_2168 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2405_cse <= (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_2411_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_2409_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2114_nl <= MUX_s_1_2_2(or_2411_nl, or_2409_nl, fsm_output(1));
  or_2412_nl <= (fsm_output(4)) OR mux_2114_nl;
  or_2407_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_2111_nl <= MUX_s_1_2_2(or_tmp_2168, or_2405_cse, fsm_output(0));
  nand_121_nl <= NOT((fsm_output(3)) AND (NOT mux_2111_nl));
  mux_2112_nl <= MUX_s_1_2_2(or_2407_nl, nand_121_nl, fsm_output(1));
  or_2403_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2113_nl <= MUX_s_1_2_2(mux_2112_nl, or_2403_nl, fsm_output(4));
  mux_tmp_2115 <= MUX_s_1_2_2(or_2412_nl, mux_2113_nl, fsm_output(6));
  or_tmp_2176 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_tmp_2179 <= (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  and_dcpl_588 <= and_dcpl_569 AND and_dcpl_510;
  and_dcpl_594 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (fsm_output(5));
  and_dcpl_596 <= (NOT mux_156_itm) AND and_dcpl_523 AND and_dcpl_594;
  or_2462_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_2460_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_2162_nl <= MUX_s_1_2_2(or_2462_nl, or_2460_nl, fsm_output(1));
  or_2457_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_2455_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2160_nl <= MUX_s_1_2_2(or_2457_nl, or_2455_nl, fsm_output(3));
  nor_1673_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  nor_1674_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_2159_nl <= MUX_s_1_2_2(nor_1673_nl, nor_1674_nl, fsm_output(0));
  nand_124_nl <= NOT((fsm_output(3)) AND mux_2159_nl);
  mux_2161_nl <= MUX_s_1_2_2(mux_2160_nl, nand_124_nl, fsm_output(1));
  mux_tmp_2163 <= MUX_s_1_2_2(mux_2162_nl, mux_2161_nl, fsm_output(6));
  or_tmp_2228 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  and_dcpl_599 <= and_dcpl_568 AND and_dcpl_535;
  and_dcpl_600 <= and_dcpl_599 AND and_dcpl_464;
  and_1626_nl <= ((NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))) OR (NOT (fsm_output(3)))))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2480_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2185_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2480_nl);
  or_2479_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2184_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2479_nl);
  mux_2186_nl <= MUX_s_1_2_2(mux_2185_nl, mux_2184_nl, fsm_output(0));
  mux_tmp_2187 <= MUX_s_1_2_2(and_1626_nl, mux_2186_nl, fsm_output(2));
  and_dcpl_605 <= and_dcpl_577 AND and_dcpl_535;
  or_tmp_2259 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  or_tmp_2265 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_tmp_2266 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2216_nl <= MUX_s_1_2_2(or_tmp_2265, or_2405_cse, fsm_output(0));
  mux_2217_nl <= MUX_s_1_2_2(or_tmp_2266, mux_2216_nl, fsm_output(1));
  nand_126_nl <= NOT((fsm_output(3)) AND (NOT mux_2217_nl));
  mux_2218_nl <= MUX_s_1_2_2(or_634_cse, nand_126_nl, fsm_output(6));
  or_2502_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2219 <= MUX_s_1_2_2(mux_2218_nl, or_2502_nl, fsm_output(4));
  or_2511_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"));
  mux_tmp_2222 <= MUX_s_1_2_2(or_2511_nl, or_tmp_2259, fsm_output(1));
  and_dcpl_609 <= and_dcpl_599 AND and_dcpl_510;
  and_1615_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4) AND (fsm_output(5)) AND (fsm_output(3)))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2521_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2243_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2521_nl);
  or_2520_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0111"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2242_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2520_nl);
  mux_2244_nl <= MUX_s_1_2_2(mux_2243_nl, mux_2242_nl, fsm_output(0));
  mux_tmp_2245 <= MUX_s_1_2_2(and_1615_nl, mux_2244_nl, fsm_output(2));
  and_dcpl_613 <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (NOT (fsm_output(2)));
  or_2538_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  or_2537_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_tmp_2272 <= MUX_s_1_2_2(or_2538_nl, or_2537_nl, fsm_output(0));
  or_2540_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  or_2539_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_2273 <= MUX_s_1_2_2(or_2540_nl, or_2539_nl, fsm_output(1));
  or_tmp_2300 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  or_tmp_2306 <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_2284 <= MUX_s_1_2_2(or_4679_cse, or_tmp_2306, fsm_output(1));
  or_tmp_2310 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  and_dcpl_619 <= (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3));
  and_dcpl_620 <= and_dcpl_619 AND (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)));
  and_dcpl_621 <= and_dcpl_468 AND and_dcpl_620;
  and_dcpl_622 <= and_dcpl_621 AND and_dcpl_464;
  and_dcpl_626 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_629 <= and_dcpl_489 AND and_dcpl_620;
  and_dcpl_631 <= (operator_20_true_28_acc_tmp(1)) AND (fsm_output(5));
  and_dcpl_634 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(4 DOWNTO 3)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_635 <= and_dcpl_634 AND (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(1)));
  and_dcpl_637 <= and_dcpl_635 AND and_dcpl_497 AND and_dcpl_90;
  or_dcpl_241 <= or_dcpl_226 OR (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(3)));
  or_tmp_2348 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2590_cse <= (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_2594_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_2593_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2334_nl <= MUX_s_1_2_2(or_2594_nl, or_2593_nl, fsm_output(1));
  or_2595_nl <= (fsm_output(4)) OR mux_2334_nl;
  or_2592_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_2331_nl <= MUX_s_1_2_2(or_tmp_2348, or_2590_cse, fsm_output(0));
  nand_130_nl <= NOT((fsm_output(3)) AND (NOT mux_2331_nl));
  mux_2332_nl <= MUX_s_1_2_2(or_2592_nl, nand_130_nl, fsm_output(1));
  or_2589_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2333_nl <= MUX_s_1_2_2(mux_2332_nl, or_2589_nl, fsm_output(4));
  mux_tmp_2335 <= MUX_s_1_2_2(or_2595_nl, mux_2333_nl, fsm_output(6));
  or_tmp_2353 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_tmp_2355 <= (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  and_dcpl_640 <= and_dcpl_621 AND and_dcpl_510;
  and_dcpl_646 <= and_dcpl_522 AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1));
  and_dcpl_648 <= (NOT mux_156_itm) AND and_dcpl_646 AND and_dcpl_521;
  and_dcpl_650 <= and_dcpl_635 AND and_dcpl_526 AND and_dcpl_90;
  or_2638_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_2637_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_2382_nl <= MUX_s_1_2_2(or_2638_nl, or_2637_nl, fsm_output(1));
  or_2635_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_2634_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2380_nl <= MUX_s_1_2_2(or_2635_nl, or_2634_nl, fsm_output(3));
  nor_1640_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  nor_1641_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  mux_2379_nl <= MUX_s_1_2_2(nor_1640_nl, nor_1641_nl, fsm_output(0));
  nand_133_nl <= NOT((fsm_output(3)) AND mux_2379_nl);
  mux_2381_nl <= MUX_s_1_2_2(mux_2380_nl, nand_133_nl, fsm_output(1));
  mux_tmp_2383 <= MUX_s_1_2_2(mux_2382_nl, mux_2381_nl, fsm_output(6));
  or_tmp_2398 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  and_dcpl_653 <= and_dcpl_619 AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1));
  and_dcpl_654 <= and_dcpl_468 AND and_dcpl_653;
  and_dcpl_655 <= and_dcpl_654 AND and_dcpl_464;
  and_1585_nl <= ((NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))) OR (NOT (fsm_output(3)))))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2653_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2401_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2653_nl);
  or_2652_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2400_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2652_nl);
  mux_2402_nl <= MUX_s_1_2_2(mux_2401_nl, mux_2400_nl, fsm_output(0));
  mux_tmp_2403 <= MUX_s_1_2_2(and_1585_nl, mux_2402_nl, fsm_output(2));
  and_dcpl_660 <= and_dcpl_489 AND and_dcpl_653;
  and_dcpl_662 <= and_dcpl_634 AND (S34_OUTER_LOOP_for_a_acc_2_tmp(1));
  and_dcpl_664 <= and_dcpl_662 AND and_dcpl_497 AND and_dcpl_90;
  or_tmp_2428 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  or_tmp_2432 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_tmp_2433 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2436_nl <= MUX_s_1_2_2(or_tmp_2432, or_2590_cse, fsm_output(0));
  mux_2437_nl <= MUX_s_1_2_2(or_tmp_2433, mux_2436_nl, fsm_output(1));
  nand_135_nl <= NOT((fsm_output(3)) AND (NOT mux_2437_nl));
  mux_2438_nl <= MUX_s_1_2_2(or_864_cse, nand_135_nl, fsm_output(6));
  or_2675_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_2439 <= MUX_s_1_2_2(mux_2438_nl, or_2675_nl, fsm_output(4));
  or_2681_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_tmp_2442 <= MUX_s_1_2_2(or_2681_nl, or_tmp_2428, fsm_output(1));
  and_dcpl_667 <= and_dcpl_654 AND and_dcpl_510;
  and_1574_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1011"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4) AND (fsm_output(5)) AND (fsm_output(3)))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2689_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2459_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2689_nl);
  or_2688_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2458_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2688_nl);
  mux_2460_nl <= MUX_s_1_2_2(mux_2459_nl, mux_2458_nl, fsm_output(0));
  mux_tmp_2461 <= MUX_s_1_2_2(and_1574_nl, mux_2460_nl, fsm_output(2));
  and_dcpl_675 <= and_dcpl_662 AND and_dcpl_526 AND and_dcpl_90;
  or_2710_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  or_2709_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_tmp_2492 <= MUX_s_1_2_2(or_2710_nl, or_2709_nl, fsm_output(0));
  or_2712_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  or_2711_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  mux_tmp_2493 <= MUX_s_1_2_2(or_2712_nl, or_2711_nl, fsm_output(1));
  or_tmp_2469 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  or_tmp_2472 <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  mux_tmp_2504 <= MUX_s_1_2_2(or_4679_cse, or_tmp_2472, fsm_output(1));
  or_tmp_2476 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  and_dcpl_678 <= and_dcpl_568 AND and_dcpl_620;
  and_dcpl_679 <= and_dcpl_678 AND and_dcpl_464;
  and_dcpl_683 <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_686 <= and_dcpl_577 AND and_dcpl_620;
  or_dcpl_246 <= or_dcpl_235 OR (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(3)));
  or_tmp_2518 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_2765_cse <= (NOT (fsm_output(2))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR
      not_tmp_389;
  or_2771_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  or_2769_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  mux_2554_nl <= MUX_s_1_2_2(or_2771_nl, or_2769_nl, fsm_output(1));
  or_2772_nl <= (fsm_output(4)) OR mux_2554_nl;
  or_2767_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101")) OR
      S1_OUTER_LOOP_for_acc_svs_4;
  mux_2551_nl <= MUX_s_1_2_2(or_tmp_2518, or_2765_cse, fsm_output(0));
  nand_139_nl <= NOT((fsm_output(3)) AND (NOT mux_2551_nl));
  mux_2552_nl <= MUX_s_1_2_2(or_2767_nl, nand_139_nl, fsm_output(1));
  or_2763_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  mux_2553_nl <= MUX_s_1_2_2(mux_2552_nl, or_2763_nl, fsm_output(4));
  mux_tmp_2555 <= MUX_s_1_2_2(or_2772_nl, mux_2553_nl, fsm_output(6));
  or_tmp_2526 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  or_tmp_2529 <= (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  and_dcpl_692 <= and_dcpl_678 AND and_dcpl_510;
  and_dcpl_699 <= (NOT mux_156_itm) AND and_dcpl_646 AND and_dcpl_594;
  or_2822_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  or_2820_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  mux_2602_nl <= MUX_s_1_2_2(or_2822_nl, or_2820_nl, fsm_output(1));
  or_2817_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  or_2815_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_2600_nl <= MUX_s_1_2_2(or_2817_nl, or_2815_nl, fsm_output(3));
  nor_1608_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4);
  nor_1609_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389);
  mux_2599_nl <= MUX_s_1_2_2(nor_1608_nl, nor_1609_nl, fsm_output(0));
  nand_142_nl <= NOT((fsm_output(3)) AND mux_2599_nl);
  mux_2601_nl <= MUX_s_1_2_2(mux_2600_nl, nand_142_nl, fsm_output(1));
  mux_tmp_2603 <= MUX_s_1_2_2(mux_2602_nl, mux_2601_nl, fsm_output(6));
  or_tmp_2578 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  and_dcpl_702 <= and_dcpl_568 AND and_dcpl_653;
  and_dcpl_703 <= and_dcpl_702 AND and_dcpl_464;
  and_1542_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1110"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4) AND (fsm_output(5)) AND (fsm_output(3)))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2840_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2625_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2840_nl);
  or_2839_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2624_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2839_nl);
  mux_2626_nl <= MUX_s_1_2_2(mux_2625_nl, mux_2624_nl, fsm_output(0));
  mux_tmp_2627 <= MUX_s_1_2_2(and_1542_nl, mux_2626_nl, fsm_output(2));
  and_dcpl_708 <= and_dcpl_577 AND and_dcpl_653;
  or_tmp_2609 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  or_tmp_2615 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1111"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  or_tmp_2616 <= NOT((fsm_output(0)) AND (NOT (fsm_output(2))) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_2656_nl <= MUX_s_1_2_2(or_tmp_2615, or_2765_cse, fsm_output(0));
  mux_2657_nl <= MUX_s_1_2_2(or_tmp_2616, mux_2656_nl, fsm_output(1));
  nand_144_nl <= NOT((fsm_output(3)) AND (NOT mux_2657_nl));
  mux_2658_nl <= MUX_s_1_2_2(or_1085_cse, nand_144_nl, fsm_output(6));
  or_2862_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR not_tmp_389;
  mux_tmp_2659 <= MUX_s_1_2_2(mux_2658_nl, or_2862_nl, fsm_output(4));
  or_2871_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR not_tmp_389;
  mux_tmp_2662 <= MUX_s_1_2_2(or_2871_nl, or_tmp_2609, fsm_output(1));
  and_dcpl_712 <= and_dcpl_702 AND and_dcpl_510;
  and_1528_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND (NOT S1_OUTER_LOOP_for_acc_svs_4) AND (fsm_output(5)) AND (fsm_output(3)))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_2881_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1111"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5)) OR (fsm_output(3));
  mux_2683_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2881_nl);
  or_2880_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1111"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(5)) OR (fsm_output(3));
  mux_2682_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2880_nl);
  mux_2684_nl <= MUX_s_1_2_2(mux_2683_nl, mux_2682_nl, fsm_output(0));
  mux_tmp_2685 <= MUX_s_1_2_2(and_1528_nl, mux_2684_nl, fsm_output(2));
  or_2901_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_2899_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_tmp_2712 <= MUX_s_1_2_2(or_2901_nl, or_2899_nl, fsm_output(0));
  or_2905_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  or_2903_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_2713 <= MUX_s_1_2_2(or_2905_nl, or_2903_nl, fsm_output(1));
  or_tmp_2656 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  or_tmp_2663 <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_2723 <= MUX_s_1_2_2(or_4679_cse, or_tmp_2663, fsm_output(1));
  or_tmp_2666 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100"));
  and_dcpl_721 <= reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)));
  and_dcpl_722 <= and_dcpl_721 AND (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)));
  and_dcpl_723 <= and_dcpl_468 AND and_dcpl_722;
  and_dcpl_724 <= and_dcpl_723 AND and_dcpl_464;
  and_dcpl_728 <= (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2)) AND (NOT (fsm_output(2)));
  and_dcpl_731 <= and_dcpl_489 AND and_dcpl_722;
  and_dcpl_733 <= and_dcpl_493 AND (operator_20_true_28_acc_tmp(2));
  and_dcpl_736 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(4 DOWNTO 3)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_737 <= and_dcpl_736 AND (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(1)));
  and_dcpl_739 <= and_dcpl_737 AND and_dcpl_497 AND and_dcpl_90;
  or_dcpl_251 <= (S34_OUTER_LOOP_for_a_acc_2_tmp(2)) OR (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(4)));
  or_dcpl_252 <= or_dcpl_251 OR (S34_OUTER_LOOP_for_a_acc_2_tmp(3));
  or_tmp_2710 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_2962_cse <= (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_2968_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_2967_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2774_nl <= MUX_s_1_2_2(or_2968_nl, or_2967_nl, fsm_output(1));
  or_2969_nl <= (fsm_output(4)) OR mux_2774_nl;
  or_2966_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2771_nl <= MUX_s_1_2_2(or_tmp_2710, or_2962_cse, fsm_output(0));
  nand_148_nl <= NOT((fsm_output(3)) AND (NOT mux_2771_nl));
  mux_2772_nl <= MUX_s_1_2_2(or_2966_nl, nand_148_nl, fsm_output(1));
  or_2961_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2773_nl <= MUX_s_1_2_2(mux_2772_nl, or_2961_nl, fsm_output(4));
  mux_tmp_2775 <= MUX_s_1_2_2(or_2969_nl, mux_2773_nl, fsm_output(6));
  or_tmp_2716 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_tmp_2717 <= (NOT (fsm_output(0))) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  and_dcpl_742 <= and_dcpl_723 AND and_dcpl_510;
  and_dcpl_748 <= (NOT (fsm_output(4))) AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2));
  and_dcpl_749 <= and_dcpl_748 AND (NOT (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)));
  and_dcpl_751 <= (NOT mux_156_itm) AND and_dcpl_749 AND and_dcpl_521;
  and_dcpl_753 <= and_dcpl_737 AND and_dcpl_526 AND and_dcpl_90;
  or_3018_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_3017_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_2822_nl <= MUX_s_1_2_2(or_3018_nl, or_3017_nl, fsm_output(1));
  or_3015_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_3014_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2820_nl <= MUX_s_1_2_2(or_3015_nl, or_3014_nl, fsm_output(3));
  nor_1577_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  nor_1578_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100")));
  mux_2819_nl <= MUX_s_1_2_2(nor_1577_nl, nor_1578_nl, fsm_output(0));
  nand_151_nl <= NOT((fsm_output(3)) AND mux_2819_nl);
  mux_2821_nl <= MUX_s_1_2_2(mux_2820_nl, nand_151_nl, fsm_output(1));
  mux_tmp_2823 <= MUX_s_1_2_2(mux_2822_nl, mux_2821_nl, fsm_output(6));
  or_tmp_2765 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  and_dcpl_756 <= and_dcpl_721 AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1));
  and_dcpl_757 <= and_dcpl_468 AND and_dcpl_756;
  and_dcpl_758 <= and_dcpl_757 AND and_dcpl_464;
  and_1498_nl <= ((NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(3)))))
      OR (fsm_output(7))) AND (fsm_output(6));
  or_3036_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_2841_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3036_nl);
  or_3035_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_2840_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3035_nl);
  mux_2842_nl <= MUX_s_1_2_2(mux_2841_nl, mux_2840_nl, fsm_output(0));
  mux_tmp_2843 <= MUX_s_1_2_2(and_1498_nl, mux_2842_nl, fsm_output(2));
  and_dcpl_763 <= and_dcpl_489 AND and_dcpl_756;
  and_dcpl_765 <= and_dcpl_736 AND (S34_OUTER_LOOP_for_a_acc_2_tmp(1));
  and_dcpl_767 <= and_dcpl_765 AND and_dcpl_497 AND and_dcpl_90;
  or_tmp_2802 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  or_tmp_2806 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_tmp_2808 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2876_nl <= MUX_s_1_2_2(or_tmp_2806, or_2962_cse, fsm_output(0));
  mux_2877_nl <= MUX_s_1_2_2(or_tmp_2808, mux_2876_nl, fsm_output(1));
  nand_153_nl <= NOT((fsm_output(3)) AND (NOT mux_2877_nl));
  mux_2878_nl <= MUX_s_1_2_2(or_1310_cse, nand_153_nl, fsm_output(6));
  or_3059_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_2879 <= MUX_s_1_2_2(mux_2878_nl, or_3059_nl, fsm_output(4));
  or_3067_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_tmp_2880 <= MUX_s_1_2_2(or_3067_nl, or_tmp_2802, fsm_output(1));
  and_dcpl_770 <= and_dcpl_757 AND and_dcpl_510;
  and_1487_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0011"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  or_3077_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_2899_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3077_nl);
  or_3076_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_2898_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3076_nl);
  mux_2900_nl <= MUX_s_1_2_2(mux_2899_nl, mux_2898_nl, fsm_output(0));
  mux_tmp_2901 <= MUX_s_1_2_2(and_1487_nl, mux_2900_nl, fsm_output(2));
  and_dcpl_778 <= and_dcpl_765 AND and_dcpl_526 AND and_dcpl_90;
  or_3103_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_3101_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_tmp_2932 <= MUX_s_1_2_2(or_3103_nl, or_3101_nl, fsm_output(0));
  or_3107_nl <= (fsm_output(3)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  or_3105_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  mux_tmp_2933 <= MUX_s_1_2_2(or_3107_nl, or_3105_nl, fsm_output(1));
  or_tmp_2855 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  or_tmp_2858 <= (fsm_output(3)) OR (fsm_output(7)) OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  mux_tmp_2943 <= MUX_s_1_2_2(or_4679_cse, or_tmp_2858, fsm_output(1));
  or_tmp_2861 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101"));
  and_dcpl_781 <= and_dcpl_568 AND and_dcpl_722;
  and_dcpl_782 <= and_dcpl_781 AND and_dcpl_464;
  and_dcpl_788 <= and_dcpl_577 AND and_dcpl_722;
  and_dcpl_790 <= and_dcpl_580 AND (operator_20_true_28_acc_tmp(2));
  or_dcpl_257 <= NOT((S34_OUTER_LOOP_for_a_acc_2_tmp(2)) AND (S34_OUTER_LOOP_for_a_acc_2_tmp(4)));
  or_dcpl_258 <= or_dcpl_257 OR (S34_OUTER_LOOP_for_a_acc_2_tmp(3));
  or_tmp_2909 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  nand_542_cse <= NOT((fsm_output(2)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101")));
  or_3175_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  or_3173_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_2994_nl <= MUX_s_1_2_2(or_3175_nl, or_3173_nl, fsm_output(1));
  or_3176_nl <= (fsm_output(4)) OR mux_2994_nl;
  or_3171_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_2991_nl <= MUX_s_1_2_2(or_tmp_2909, nand_542_cse, fsm_output(0));
  nand_157_nl <= NOT((fsm_output(3)) AND (NOT mux_2991_nl));
  mux_2992_nl <= MUX_s_1_2_2(or_3171_nl, nand_157_nl, fsm_output(1));
  or_3165_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_2993_nl <= MUX_s_1_2_2(mux_2992_nl, or_3165_nl, fsm_output(4));
  mux_tmp_2995 <= MUX_s_1_2_2(or_3176_nl, mux_2993_nl, fsm_output(6));
  or_tmp_2918 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  or_tmp_2920 <= NOT((fsm_output(0)) AND (fsm_output(2)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101")));
  and_dcpl_795 <= and_dcpl_781 AND and_dcpl_510;
  and_dcpl_802 <= (NOT mux_156_itm) AND and_dcpl_749 AND and_dcpl_594;
  or_3232_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  or_3230_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_3042_nl <= MUX_s_1_2_2(or_3232_nl, or_3230_nl, fsm_output(1));
  or_3227_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  or_3225_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  mux_3040_nl <= MUX_s_1_2_2(or_3227_nl, or_3225_nl, fsm_output(3));
  nor_1543_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  nor_1544_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  mux_3039_nl <= MUX_s_1_2_2(nor_1543_nl, nor_1544_nl, fsm_output(0));
  nand_160_nl <= NOT((fsm_output(3)) AND mux_3039_nl);
  mux_3041_nl <= MUX_s_1_2_2(mux_3040_nl, nand_160_nl, fsm_output(1));
  mux_tmp_3043 <= MUX_s_1_2_2(mux_3042_nl, mux_3041_nl, fsm_output(6));
  or_tmp_2974 <= NOT((fsm_output(2)) AND (fsm_output(4)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101")));
  and_dcpl_805 <= and_dcpl_568 AND and_dcpl_756;
  and_dcpl_806 <= and_dcpl_805 AND and_dcpl_464;
  and_1457_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0110"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  or_3253_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3065_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3253_nl);
  or_3252_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3064_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3252_nl);
  mux_3066_nl <= MUX_s_1_2_2(mux_3065_nl, mux_3064_nl, fsm_output(0));
  mux_tmp_3067 <= MUX_s_1_2_2(and_1457_nl, mux_3066_nl, fsm_output(2));
  and_dcpl_811 <= and_dcpl_577 AND and_dcpl_756;
  or_tmp_3012 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  or_tmp_3018 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4);
  or_tmp_3020 <= NOT((fsm_output(0)) AND (NOT (fsm_output(2))) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND S1_OUTER_LOOP_for_acc_svs_4);
  mux_3096_nl <= MUX_s_1_2_2(or_tmp_3018, nand_542_cse, fsm_output(0));
  mux_3097_nl <= MUX_s_1_2_2(or_tmp_3020, mux_3096_nl, fsm_output(1));
  nand_162_nl <= NOT((fsm_output(3)) AND (NOT mux_3097_nl));
  mux_3098_nl <= MUX_s_1_2_2(or_1547_cse, nand_162_nl, fsm_output(6));
  or_3276_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_tmp_3099 <= MUX_s_1_2_2(mux_3098_nl, or_3276_nl, fsm_output(4));
  or_3287_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"));
  mux_tmp_3100 <= MUX_s_1_2_2(or_3287_nl, or_tmp_3012, fsm_output(1));
  and_dcpl_815 <= and_dcpl_805 AND and_dcpl_510;
  and_1444_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("0111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  or_3299_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3123_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3299_nl);
  or_3298_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3122_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3298_nl);
  mux_3124_nl <= MUX_s_1_2_2(mux_3123_nl, mux_3122_nl, fsm_output(0));
  mux_tmp_3125 <= MUX_s_1_2_2(and_1444_nl, mux_3124_nl, fsm_output(2));
  not_tmp_1143 <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11")));
  or_3321_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("000"))
      OR nand_520_cse;
  or_3319_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")) OR nand_520_cse;
  mux_tmp_3152 <= MUX_s_1_2_2(or_3321_nl, or_3319_nl, fsm_output(0));
  or_3325_nl <= (fsm_output(3)) OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)) OR not_tmp_1143;
  or_3323_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0))
      OR not_tmp_1143;
  mux_tmp_3153 <= MUX_s_1_2_2(or_3325_nl, or_3323_nl, fsm_output(1));
  or_tmp_3064 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0))
      OR not_tmp_1143;
  or_tmp_3071 <= (fsm_output(3)) OR (fsm_output(7)) OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0))
      OR not_tmp_1143;
  mux_tmp_3163 <= MUX_s_1_2_2(or_4679_cse, or_tmp_3071, fsm_output(1));
  or_tmp_3074 <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(7)))
      OR (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)) OR not_tmp_1143;
  and_dcpl_825 <= and_1812_cse AND (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)));
  and_dcpl_826 <= and_dcpl_468 AND and_dcpl_825;
  and_dcpl_827 <= and_dcpl_826 AND and_dcpl_464;
  and_dcpl_833 <= and_dcpl_489 AND and_dcpl_825;
  and_dcpl_837 <= CONV_SL_1_1(S34_OUTER_LOOP_for_a_acc_2_tmp(4 DOWNTO 3)=STD_LOGIC_VECTOR'("11"));
  and_dcpl_838 <= and_dcpl_837 AND (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(1)));
  and_dcpl_840 <= and_dcpl_838 AND and_dcpl_497 AND and_dcpl_90;
  or_dcpl_263 <= or_dcpl_251 OR (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(3)));
  or_tmp_3118 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("001")) OR nand_520_cse;
  nand_300_cse <= NOT((fsm_output(2)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  or_3387_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("01")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_3386_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_3214_nl <= MUX_s_1_2_2(or_3387_nl, or_3386_nl, fsm_output(1));
  or_3388_nl <= (fsm_output(4)) OR mux_3214_nl;
  or_3385_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("001"))
      OR nand_520_cse;
  mux_3211_nl <= MUX_s_1_2_2(or_tmp_3118, nand_300_cse, fsm_output(0));
  nand_166_nl <= NOT((fsm_output(3)) AND (NOT mux_3211_nl));
  mux_3212_nl <= MUX_s_1_2_2(or_3385_nl, nand_166_nl, fsm_output(1));
  or_3380_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_3213_nl <= MUX_s_1_2_2(mux_3212_nl, or_3380_nl, fsm_output(4));
  mux_tmp_3215 <= MUX_s_1_2_2(or_3388_nl, mux_3213_nl, fsm_output(6));
  or_tmp_3124 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_tmp_3125 <= NOT((fsm_output(0)) AND (fsm_output(2)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  and_dcpl_843 <= and_dcpl_826 AND and_dcpl_510;
  and_dcpl_849 <= and_dcpl_748 AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1));
  and_dcpl_851 <= (NOT mux_156_itm) AND and_dcpl_849 AND and_dcpl_521;
  and_dcpl_853 <= and_dcpl_838 AND and_dcpl_526 AND and_dcpl_90;
  or_3437_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_3436_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_3262_nl <= MUX_s_1_2_2(or_3437_nl, or_3436_nl, fsm_output(1));
  or_3434_nl <= (fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_3433_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR nand_520_cse;
  mux_3260_nl <= MUX_s_1_2_2(or_3434_nl, or_3433_nl, fsm_output(3));
  nor_1509_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("010")) OR nand_520_cse);
  nor_1510_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110")));
  mux_3259_nl <= MUX_s_1_2_2(nor_1509_nl, nor_1510_nl, fsm_output(0));
  nand_169_nl <= NOT((fsm_output(3)) AND mux_3259_nl);
  mux_3261_nl <= MUX_s_1_2_2(mux_3260_nl, nand_169_nl, fsm_output(1));
  mux_tmp_3263 <= MUX_s_1_2_2(mux_3262_nl, mux_3261_nl, fsm_output(6));
  or_tmp_3173 <= NOT((fsm_output(2)) AND (fsm_output(4)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  and_dcpl_856 <= and_1812_cse AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1));
  and_dcpl_857 <= and_dcpl_468 AND and_dcpl_856;
  and_dcpl_858 <= and_dcpl_857 AND and_dcpl_464;
  and_1413_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1010"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  or_3455_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3281_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3455_nl);
  or_3454_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3280_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3454_nl);
  mux_3282_nl <= MUX_s_1_2_2(mux_3281_nl, mux_3280_nl, fsm_output(0));
  mux_tmp_3283 <= MUX_s_1_2_2(and_1413_nl, mux_3282_nl, fsm_output(2));
  and_dcpl_863 <= and_dcpl_489 AND and_dcpl_856;
  and_dcpl_865 <= and_dcpl_837 AND (S34_OUTER_LOOP_for_a_acc_2_tmp(1));
  and_dcpl_867 <= and_dcpl_865 AND and_dcpl_497 AND and_dcpl_90;
  or_tmp_3210 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  or_tmp_3214 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2 DOWNTO
      0)/=STD_LOGIC_VECTOR'("011")) OR nand_520_cse;
  or_tmp_3216 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("011")) OR nand_520_cse;
  mux_3316_nl <= MUX_s_1_2_2(or_tmp_3214, nand_300_cse, fsm_output(0));
  mux_3317_nl <= MUX_s_1_2_2(or_tmp_3216, mux_3316_nl, fsm_output(1));
  nand_171_nl <= NOT((fsm_output(3)) AND (NOT mux_3317_nl));
  mux_3318_nl <= MUX_s_1_2_2(or_1784_cse, nand_171_nl, fsm_output(6));
  or_3478_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_tmp_3319 <= MUX_s_1_2_2(mux_3318_nl, or_3478_nl, fsm_output(4));
  or_3486_nl <= (fsm_output(0)) OR (NOT (fsm_output(2))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_tmp_3320 <= MUX_s_1_2_2(or_3486_nl, or_tmp_3210, fsm_output(1));
  and_dcpl_870 <= and_dcpl_857 AND and_dcpl_510;
  and_1400_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1011"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  or_3496_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3339_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3496_nl);
  or_3495_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3338_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3495_nl);
  mux_3340_nl <= MUX_s_1_2_2(mux_3339_nl, mux_3338_nl, fsm_output(0));
  mux_tmp_3341 <= MUX_s_1_2_2(and_1400_nl, mux_3340_nl, fsm_output(2));
  and_dcpl_878 <= and_dcpl_865 AND and_dcpl_526 AND and_dcpl_90;
  not_tmp_1199 <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg=STD_LOGIC_VECTOR'("111")));
  or_3522_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(3))) OR (fsm_output(7))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_517_cse;
  or_3520_nl <= (fsm_output(1)) OR (NOT (fsm_output(3))) OR (fsm_output(7)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")) OR nand_517_cse;
  mux_tmp_3372 <= MUX_s_1_2_2(or_3522_nl, or_3520_nl, fsm_output(0));
  or_3525_nl <= (fsm_output(3)) OR not_tmp_1199;
  or_3524_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR not_tmp_1199;
  mux_tmp_3373 <= MUX_s_1_2_2(or_3525_nl, or_3524_nl, fsm_output(1));
  or_tmp_3261 <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(7)) OR not_tmp_1199;
  or_tmp_3264 <= (fsm_output(3)) OR (fsm_output(7)) OR not_tmp_1199;
  mux_tmp_3383 <= MUX_s_1_2_2(or_4679_cse, or_tmp_3264, fsm_output(1));
  or_tmp_3266 <= (fsm_output(1)) OR (NOT((fsm_output(3)) AND (fsm_output(7)) AND
      CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg=STD_LOGIC_VECTOR'("111"))));
  and_dcpl_881 <= and_dcpl_568 AND and_dcpl_825;
  and_dcpl_882 <= and_dcpl_881 AND and_dcpl_464;
  and_dcpl_888 <= and_dcpl_577 AND and_dcpl_825;
  or_dcpl_268 <= or_dcpl_257 OR (NOT (S34_OUTER_LOOP_for_a_acc_2_tmp(3)));
  nor_tmp_1094 <= (fsm_output(2)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  or_tmp_3312 <= (fsm_output(2)) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO
      0)/=STD_LOGIC_VECTOR'("01")) OR nand_517_cse;
  or_3587_nl <= (fsm_output(3)) OR (NOT nor_tmp_1094);
  or_3586_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 2)/=STD_LOGIC_VECTOR'("10")) OR nand_480_cse;
  mux_3434_nl <= MUX_s_1_2_2(or_3587_nl, or_3586_nl, fsm_output(1));
  or_3588_nl <= (fsm_output(4)) OR mux_3434_nl;
  or_4398_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_517_cse;
  mux_3431_nl <= MUX_s_1_2_2((NOT or_tmp_3312), nor_tmp_1094, fsm_output(0));
  nand_277_nl <= NOT((fsm_output(3)) AND mux_3431_nl);
  mux_3432_nl <= MUX_s_1_2_2(or_4398_nl, nand_277_nl, fsm_output(1));
  or_3580_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000")) OR
      nand_480_cse;
  mux_3433_nl <= MUX_s_1_2_2(mux_3432_nl, or_3580_nl, fsm_output(4));
  mux_tmp_3435 <= MUX_s_1_2_2(or_3588_nl, mux_3433_nl, fsm_output(6));
  or_tmp_3320 <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT nor_tmp_1094);
  not_tmp_1218 <= NOT((fsm_output(0)) AND (fsm_output(2)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  and_dcpl_894 <= and_dcpl_881 AND and_dcpl_510;
  and_dcpl_901 <= (NOT mux_156_itm) AND and_dcpl_849 AND and_dcpl_594;
  not_tmp_1235 <= NOT((fsm_output(4)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  or_3642_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(4))
      OR nand_480_cse;
  or_3640_nl <= nor_1712_cse OR (fsm_output(2)) OR (fsm_output(4)) OR nand_480_cse;
  mux_3482_nl <= MUX_s_1_2_2(or_3642_nl, or_3640_nl, fsm_output(1));
  or_3637_nl <= (fsm_output(0)) OR (fsm_output(2)) OR not_tmp_1235;
  or_3635_nl <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(0))
      OR nand_351_cse;
  mux_3480_nl <= MUX_s_1_2_2(or_3637_nl, or_3635_nl, fsm_output(3));
  nor_1476_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(0))
      OR nand_351_cse);
  nor_1477_nl <= NOT((NOT (fsm_output(2))) OR (fsm_output(4)) OR nand_480_cse);
  mux_3479_nl <= MUX_s_1_2_2(nor_1476_nl, nor_1477_nl, fsm_output(0));
  nand_177_nl <= NOT((fsm_output(3)) AND mux_3479_nl);
  mux_3481_nl <= MUX_s_1_2_2(mux_3480_nl, nand_177_nl, fsm_output(1));
  mux_tmp_3483 <= MUX_s_1_2_2(mux_3482_nl, mux_3481_nl, fsm_output(6));
  not_tmp_1239 <= NOT((fsm_output(2)) AND (fsm_output(4)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111")));
  and_dcpl_904 <= and_dcpl_568 AND and_dcpl_856;
  and_dcpl_905 <= and_dcpl_904 AND and_dcpl_464;
  and_1359_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1110"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  or_3661_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3505_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3661_nl);
  or_3660_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3504_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3660_nl);
  mux_3506_nl <= MUX_s_1_2_2(mux_3505_nl, mux_3504_nl, fsm_output(0));
  mux_tmp_3507 <= MUX_s_1_2_2(and_1359_nl, mux_3506_nl, fsm_output(2));
  and_dcpl_910 <= and_dcpl_577 AND and_dcpl_856;
  or_tmp_3410 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR nand_480_cse;
  not_tmp_1250 <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4);
  or_tmp_3413 <= (fsm_output(2)) OR not_tmp_1250;
  or_tmp_3415 <= (NOT (fsm_output(0))) OR (fsm_output(2)) OR not_tmp_1250;
  or_4389_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")) OR nand_480_cse;
  mux_3536_nl <= MUX_s_1_2_2((NOT or_tmp_3413), nor_tmp_1094, fsm_output(0));
  mux_3537_nl <= MUX_s_1_2_2((NOT or_tmp_3415), mux_3536_nl, fsm_output(1));
  nand_259_nl <= NOT((fsm_output(3)) AND mux_3537_nl);
  mux_3538_nl <= MUX_s_1_2_2(or_4389_nl, nand_259_nl, fsm_output(6));
  or_3684_nl <= (NOT (fsm_output(6))) OR (fsm_output(3)) OR (fsm_output(1)) OR (fsm_output(0))
      OR (fsm_output(2)) OR nand_480_cse;
  mux_tmp_3539 <= MUX_s_1_2_2(mux_3538_nl, or_3684_nl, fsm_output(4));
  or_3691_nl <= (fsm_output(0)) OR (NOT nor_tmp_1094);
  mux_tmp_3540 <= MUX_s_1_2_2(or_3691_nl, or_tmp_3410, fsm_output(1));
  nor_tmp_1140 <= (fsm_output(2)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4;
  and_dcpl_914 <= and_dcpl_904 AND and_dcpl_510;
  or_dcpl_273 <= not_tmp_741 OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("11"));
  and_1341_nl <= (((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5)) AND (fsm_output(3))) OR
      (fsm_output(7))) AND (fsm_output(6));
  nand_256_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1111"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (NOT (fsm_output(5))) AND (NOT (fsm_output(3))));
  mux_3563_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_256_nl);
  nand_257_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (NOT (fsm_output(5))) AND (NOT (fsm_output(3))));
  mux_3562_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_257_nl);
  mux_3564_nl <= MUX_s_1_2_2(mux_3563_nl, mux_3562_nl, fsm_output(0));
  mux_tmp_3565 <= MUX_s_1_2_2(and_1341_nl, mux_3564_nl, fsm_output(2));
  and_dcpl_924 <= nor_1711_cse AND (NOT (fsm_output(7)));
  and_dcpl_925 <= NOT((fsm_output(4)) OR (fsm_output(2)));
  and_dcpl_927 <= and_dcpl_925 AND (NOT (fsm_output(6))) AND and_dcpl_924;
  and_dcpl_932 <= and_dcpl_91 AND and_dcpl_151 AND and_2881_cse AND (fsm_output(7));
  and_dcpl_934 <= and_dcpl_126 AND and_dcpl_70;
  and_dcpl_935 <= and_dcpl_92 AND and_dcpl_61;
  not_tmp_1278 <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(2)) AND (fsm_output(1)));
  not_tmp_1311 <= NOT(S1_OUTER_LOOP_for_acc_svs_4 AND (S1_OUTER_LOOP_for_acc_svs_3_0(2))
      AND (fsm_output(1)));
  not_tmp_1328 <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4
      AND (S1_OUTER_LOOP_for_acc_svs_3_0(2)) AND (fsm_output(1)));
  and_dcpl_1000 <= (fsm_output(0)) AND (NOT (fsm_output(6)));
  and_dcpl_1007 <= and_dcpl_67 AND and_dcpl_90;
  and_dcpl_1008 <= and_dcpl_76 AND and_dcpl_458;
  and_dcpl_1010 <= and_dcpl_449 AND and_dcpl_108;
  or_tmp_3536 <= nor_2178_cse_1 OR (fsm_output(4));
  or_tmp_3537 <= (fsm_output(6)) OR or_tmp_3536;
  or_tmp_3538 <= (fsm_output(6)) OR (NOT (fsm_output(4)));
  or_tmp_3540 <= (fsm_output(1)) OR (NOT (fsm_output(4)));
  mux_tmp_3659 <= MUX_s_1_2_2(or_tmp_3540, (fsm_output(4)), fsm_output(2));
  or_tmp_3550 <= (fsm_output(7)) OR (fsm_output(2)) OR (NOT((fsm_output(0)) AND (fsm_output(4))));
  and_dcpl_1011 <= NOT((fsm_output(5)) OR (fsm_output(7)));
  and_dcpl_1012 <= NOT((fsm_output(0)) OR (fsm_output(6)));
  and_dcpl_1013 <= and_dcpl_1012 AND and_dcpl_1011;
  xor_dcpl_1 <= (fsm_output(2)) XOR (fsm_output(3));
  and_dcpl_1014 <= and_dcpl_91 AND xor_dcpl_1;
  not_tmp_1345 <= NOT((fsm_output(3)) AND (fsm_output(6)));
  nor_1388_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(6)))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))));
  nor_1389_nl <= NOT((NOT (fsm_output(7))) OR (NOT (fsm_output(3))) OR (fsm_output(6))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))));
  mux_3682_nl <= MUX_s_1_2_2(nor_1388_nl, nor_1389_nl, fsm_output(5));
  or_3846_nl <= (NOT (fsm_output(3))) OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT
      (fsm_output(2)));
  or_3844_nl <= (fsm_output(3)) OR (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(2)));
  mux_3681_nl <= MUX_s_1_2_2(or_3846_nl, or_3844_nl, fsm_output(7));
  nor_1390_nl <= NOT((fsm_output(5)) OR mux_3681_nl);
  mux_3683_nl <= MUX_s_1_2_2(mux_3682_nl, nor_1390_nl, fsm_output(4));
  or_3841_nl <= (fsm_output(6)) OR (fsm_output(0)) OR (NOT (fsm_output(2)));
  or_3839_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR (fsm_output(2));
  mux_3680_nl <= MUX_s_1_2_2(or_3841_nl, or_3839_nl, fsm_output(3));
  nor_1391_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR mux_3680_nl);
  not_tmp_1349 <= MUX_s_1_2_2(mux_3683_nl, nor_1391_nl, fsm_output(1));
  and_dcpl_1022 <= (fsm_output(5)) AND (NOT (fsm_output(7)));
  and_dcpl_1023 <= and_dcpl_1000 AND and_dcpl_1022;
  mux_3695_itm <= MUX_s_1_2_2(or_119_cse, or_2273_cse, fsm_output(3));
  and_dcpl_1024 <= NOT(mux_3695_itm OR (fsm_output(1)));
  and_dcpl_1027 <= (NOT mux_3695_itm) AND (fsm_output(1));
  and_dcpl_1031 <= (fsm_output(0)) AND (fsm_output(6));
  and_dcpl_1032 <= and_dcpl_1031 AND and_dcpl_1011;
  and_dcpl_1033 <= and_dcpl_71 AND xor_dcpl_1;
  and_dcpl_1035 <= (NOT (fsm_output(0))) AND (fsm_output(6));
  and_dcpl_1037 <= and_dcpl_95 AND xor_dcpl_1;
  and_dcpl_1041 <= and_dcpl_64 AND and_dcpl_90;
  and_dcpl_1044 <= and_dcpl_103 AND (NOT (fsm_output(7)));
  and_dcpl_1052 <= and_dcpl_95 AND and_dcpl_1000;
  and_dcpl_1054 <= (NOT (fsm_output(5))) AND (fsm_output(7));
  mux_tmp_3698 <= MUX_s_1_2_2((NOT nor_tmp_3), or_tmp_3540, fsm_output(2));
  mux_tmp_3714 <= MUX_s_1_2_2((NOT (fsm_output(2))), (fsm_output(2)), fsm_output(1));
  and_dcpl_1070 <= NOT((fsm_output(7)) OR (S1_OUTER_LOOP_k_5_0_sva_2(5)));
  mux_tmp_3730 <= MUX_s_1_2_2((fsm_output(6)), (fsm_output(7)), fsm_output(5));
  or_tmp_3658 <= (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(3));
  or_tmp_3661 <= (fsm_output(6)) OR (NOT (fsm_output(3)));
  or_tmp_3662 <= (fsm_output(5)) OR not_tmp_1345;
  mux_tmp_3769 <= MUX_s_1_2_2((NOT (fsm_output(6))), (fsm_output(6)), fsm_output(5));
  nor_1343_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(4)));
  nor_1344_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(0)) OR (NOT (fsm_output(4))));
  mux_3798_nl <= MUX_s_1_2_2(nor_1343_nl, nor_1344_nl, fsm_output(3));
  and_dcpl_1082 <= mux_3798_nl AND nor_2178_cse_1 AND and_dcpl_1011;
  nand_242_cse <= NOT((fsm_output(7)) AND (fsm_output(5)));
  and_dcpl_1083 <= nor_tmp_3 AND and_dcpl_110;
  and_dcpl_1084 <= and_dcpl_1083 AND and_dcpl_75;
  or_dcpl_276 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("00"));
  or_dcpl_277 <= or_dcpl_276 OR or_2158_cse;
  and_dcpl_1085 <= (NOT (fsm_output(4))) AND (fsm_output(0));
  and_dcpl_1086 <= and_dcpl_1085 AND (NOT (fsm_output(7)));
  or_3980_nl <= (fsm_output(6)) OR (NOT (fsm_output(2))) OR (fsm_output(1));
  or_3979_nl <= (NOT (fsm_output(6))) OR (fsm_output(2)) OR (NOT (fsm_output(1)));
  mux_tmp_3812 <= MUX_s_1_2_2(or_3980_nl, or_3979_nl, fsm_output(5));
  and_dcpl_1088 <= not_tmp_116 AND and_dcpl_1086;
  or_tmp_3706 <= and_2120_cse OR (fsm_output(4));
  mux_tmp_3819 <= MUX_s_1_2_2(and_dcpl_71, nor_tmp_3, fsm_output(2));
  nor_tmp_1200 <= or_4342_cse AND (fsm_output(4));
  and_dcpl_1091 <= and_dcpl_178 AND and_dcpl_70;
  and_dcpl_1092 <= and_dcpl_130 AND and_dcpl_90;
  or_tmp_3740 <= (fsm_output(0)) OR (fsm_output(2)) OR (fsm_output(1)) OR (NOT (fsm_output(4)));
  nor_1326_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(0))) OR (fsm_output(2))
      OR (fsm_output(1)));
  nor_1327_nl <= NOT((NOT (fsm_output(6))) OR (fsm_output(0)) OR (NOT and_2141_cse));
  mux_3855_nl <= MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output(5));
  nor_1328_nl <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(2))
      OR (fsm_output(1)));
  mux_3856_nl <= MUX_s_1_2_2(mux_3855_nl, nor_1328_nl, fsm_output(3));
  and_dcpl_1095 <= mux_3856_nl AND nor_1303_cse;
  mux_3859_nl <= MUX_s_1_2_2((fsm_output(5)), (NOT (fsm_output(5))), fsm_output(3));
  nand_197_nl <= NOT((NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("10"))))
      AND mux_3859_nl);
  or_99_nl <= (fsm_output(7)) OR not_tmp_28;
  or_100_nl <= (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(3));
  mux_3858_nl <= MUX_s_1_2_2(or_99_nl, or_100_nl, fsm_output(6));
  mux_3860_nl <= MUX_s_1_2_2(nand_197_nl, mux_3858_nl, fsm_output(1));
  nor_1323_nl <= NOT((fsm_output(2)) OR (fsm_output(4)) OR mux_3860_nl);
  nor_1324_nl <= NOT((NOT (fsm_output(4))) OR (fsm_output(1)) OR (fsm_output(6))
      OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(5)));
  nor_1325_nl <= NOT((fsm_output(4)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(6)))
      OR (fsm_output(7)) OR not_tmp_28);
  mux_3857_nl <= MUX_s_1_2_2(nor_1324_nl, nor_1325_nl, fsm_output(2));
  not_tmp_1436 <= MUX_s_1_2_2(nor_1323_nl, mux_3857_nl, fsm_output(0));
  nor_1321_nl <= NOT((fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(2)) OR (NOT
      (fsm_output(1))));
  and_1289_nl <= (fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(1));
  mux_3874_nl <= MUX_s_1_2_2(nor_1321_nl, and_1289_nl, fsm_output(5));
  nor_1322_nl <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (NOT (fsm_output(0)))
      OR (fsm_output(2)) OR (fsm_output(1)));
  mux_3875_nl <= MUX_s_1_2_2(mux_3874_nl, nor_1322_nl, fsm_output(3));
  and_dcpl_1096 <= mux_3875_nl AND nor_1303_cse;
  or_tmp_3812 <= (NOT (fsm_output(1))) OR (fsm_output(7)) OR (NOT (fsm_output(0)))
      OR (fsm_output(4));
  or_tmp_3814 <= (fsm_output(1)) OR (NOT (fsm_output(7))) OR (NOT (fsm_output(0)))
      OR (fsm_output(4));
  or_4095_nl <= (NOT (fsm_output(1))) OR (fsm_output(7)) OR (fsm_output(0)) OR (NOT
      (fsm_output(4)));
  mux_3896_nl <= MUX_s_1_2_2(or_4095_nl, or_tmp_3814, fsm_output(5));
  mux_3895_nl <= MUX_s_1_2_2(or_tmp_3814, or_tmp_3812, fsm_output(5));
  mux_3897_nl <= MUX_s_1_2_2(mux_3896_nl, mux_3895_nl, fsm_output(3));
  or_4090_nl <= (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(0)) OR (NOT (fsm_output(4)));
  mux_3894_nl <= MUX_s_1_2_2(or_tmp_3812, or_4090_nl, fsm_output(5));
  or_4092_nl <= (fsm_output(3)) OR mux_3894_nl;
  mux_3898_nl <= MUX_s_1_2_2(mux_3897_nl, or_4092_nl, fsm_output(6));
  and_dcpl_1097 <= NOT(mux_3898_nl OR (fsm_output(2)));
  and_dcpl_1101 <= nor_2178_cse_1 AND mux_45_cse AND (fsm_output(0)) AND (NOT (fsm_output(5)))
      AND and_dcpl_79;
  nor_1312_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(4))));
  nor_1313_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(4)));
  mux_3907_nl <= MUX_s_1_2_2(nor_1312_nl, nor_1313_nl, fsm_output(6));
  and_dcpl_1103 <= mux_3907_nl AND (fsm_output(1)) AND and_dcpl_99;
  and_dcpl_1105 <= and_dcpl_456 AND and_dcpl_66 AND and_dcpl_60;
  or_4112_nl <= (NOT (fsm_output(6))) OR (fsm_output(4));
  mux_3908_nl <= MUX_s_1_2_2(or_4112_nl, or_tmp_3538, fsm_output(7));
  and_dcpl_1108 <= (NOT mux_3908_nl) AND (fsm_output(1)) AND and_2893_cse AND and_dcpl_103;
  and_dcpl_1109 <= and_dcpl_130 AND and_dcpl_108;
  and_dcpl_1110 <= and_dcpl_178 AND and_dcpl_115;
  and_dcpl_1112 <= and_dcpl_95 AND and_dcpl_151 AND and_dcpl_924;
  and_dcpl_1113 <= and_dcpl_178 AND and_dcpl_94;
  and_dcpl_1114 <= and_dcpl_64 AND and_dcpl_70;
  and_dcpl_1115 <= and_dcpl_96 AND and_dcpl_458;
  and_dcpl_1116 <= and_dcpl_476 AND and_dcpl_108;
  or_tmp_3871 <= CONV_SL_1_1(fsm_output(6 DOWNTO 5)/=STD_LOGIC_VECTOR'("01"));
  or_4288_nl <= CONV_SL_1_1(fsm_output(6 DOWNTO 3)/=STD_LOGIC_VECTOR'("0010"));
  or_4287_nl <= (fsm_output(4)) OR not_tmp_28;
  or_4286_nl <= CONV_SL_1_1(fsm_output(5 DOWNTO 3)/=STD_LOGIC_VECTOR'("000"));
  mux_4055_nl <= MUX_s_1_2_2(or_4287_nl, or_4286_nl, fsm_output(6));
  mux_4056_nl <= MUX_s_1_2_2(or_4288_nl, mux_4055_nl, fsm_output(0));
  nor_1269_nl <= NOT((fsm_output(2)) OR (fsm_output(7)) OR mux_4056_nl);
  nor_1270_nl <= NOT((fsm_output(0)) OR (NOT (fsm_output(6))) OR (fsm_output(4))
      OR not_tmp_28);
  mux_4053_nl <= MUX_s_1_2_2(or_4818_cse, or_4781_cse, fsm_output(4));
  nor_1271_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(6)) OR mux_4053_nl);
  mux_4054_nl <= MUX_s_1_2_2(nor_1270_nl, nor_1271_nl, fsm_output(7));
  and_1275_nl <= (fsm_output(2)) AND mux_4054_nl;
  not_tmp_1520 <= MUX_s_1_2_2(nor_1269_nl, and_1275_nl, fsm_output(1));
  mux_73_nl <= MUX_s_1_2_2(and_1306_cse, nor_tmp_4, fsm_output(0));
  or_tmp_4011 <= (fsm_output(6)) OR mux_73_nl;
  nor_1268_nl <= NOT((fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(4)));
  mux_tmp_4062 <= MUX_s_1_2_2(nor_1268_nl, mux_tmp_3819, fsm_output(0));
  mux_4066_nl <= MUX_s_1_2_2(nor_tmp_1200, (NOT mux_tmp_4062), fsm_output(6));
  mux_4065_nl <= MUX_s_1_2_2(or_129_cse, (fsm_output(4)), fsm_output(6));
  mux_4067_nl <= MUX_s_1_2_2(mux_4066_nl, mux_4065_nl, fsm_output(5));
  mux_4063_nl <= MUX_s_1_2_2((NOT mux_tmp_4062), or_tmp_3706, fsm_output(6));
  mux_4064_nl <= MUX_s_1_2_2((NOT mux_45_cse), mux_4063_nl, fsm_output(5));
  mux_4068_nl <= MUX_s_1_2_2(mux_4067_nl, mux_4064_nl, fsm_output(3));
  or_4291_nl <= (fsm_output(6)) OR (NOT or_2273_cse);
  mux_4060_nl <= MUX_s_1_2_2(or_4291_nl, or_tmp_4011, fsm_output(5));
  mux_4059_nl <= MUX_s_1_2_2(or_tmp_4011, or_4376_cse, fsm_output(5));
  mux_4061_nl <= MUX_s_1_2_2(mux_4060_nl, mux_4059_nl, fsm_output(3));
  mux_tmp_4069 <= MUX_s_1_2_2((NOT mux_4068_nl), mux_4061_nl, fsm_output(7));
  and_dcpl_1136 <= and_dcpl_96 AND and_dcpl_70;
  or_tmp_4014 <= (fsm_output(6)) OR nor_tmp_1200;
  mux_4074_nl <= MUX_s_1_2_2(and_dcpl_71, (fsm_output(4)), fsm_output(2));
  mux_4073_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), or_4699_cse);
  mux_tmp_4075 <= MUX_s_1_2_2(mux_4074_nl, mux_4073_nl, fsm_output(0));
  mux_tmp_4094 <= MUX_s_1_2_2(or_tmp_48, (fsm_output(7)), fsm_output(4));
  or_dcpl_286 <= or_tmp_35 OR or_4378_cse;
  or_dcpl_302 <= or_tmp_3871 OR (fsm_output(3)) OR (NOT (fsm_output(7)));
  nor_2307_cse <= NOT((NOT (fsm_output(6))) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(4)));
  mux_3731_cse <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), fsm_output(5));
  nor_1346_cse <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00")));
  or_3962_nl <= (fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(6)) OR (fsm_output(7))
      OR (fsm_output(5));
  or_3971_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("011"));
  or_3969_nl <= CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("000"));
  mux_3809_nl <= MUX_s_1_2_2(or_3971_nl, or_3969_nl, fsm_output(1));
  mux_3802_nl <= MUX_s_1_2_2(or_3962_nl, mux_3809_nl, fsm_output(2));
  nor_1339_nl <= NOT((fsm_output(3)) OR mux_3802_nl);
  nor_1340_nl <= NOT((fsm_output(6)) OR nand_242_cse);
  nor_1251_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 5)/=STD_LOGIC_VECTOR'("010")));
  mux_3799_nl <= MUX_s_1_2_2(nor_1340_nl, nor_1251_nl, fsm_output(1));
  and_1294_nl <= (fsm_output(2)) AND (fsm_output(0)) AND mux_3799_nl;
  nor_1342_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(6))
      OR nand_242_cse);
  mux_3800_nl <= MUX_s_1_2_2(and_1294_nl, nor_1342_nl, fsm_output(3));
  S1_OUTER_LOOP_for_p_sva_1_mx0c1 <= MUX_s_1_2_2(nor_1339_nl, mux_3800_nl, fsm_output(4));
  nor_1304_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(4)))
      OR (NOT (fsm_output(5))) OR (fsm_output(7)) OR (fsm_output(3)) OR (fsm_output(6)));
  or_4127_nl <= (NOT (fsm_output(4))) OR (NOT (fsm_output(5))) OR (fsm_output(7))
      OR not_tmp_1345;
  or_4125_nl <= (fsm_output(7)) OR not_tmp_1345;
  or_4087_nl <= (NOT (fsm_output(3))) OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  mux_3916_nl <= MUX_s_1_2_2(or_4125_nl, or_4087_nl, fsm_output(5));
  mux_3915_nl <= MUX_s_1_2_2(or_tmp_3661, or_4854_cse, fsm_output(7));
  or_4123_nl <= (fsm_output(5)) OR mux_3915_nl;
  mux_3917_nl <= MUX_s_1_2_2(mux_3916_nl, or_4123_nl, fsm_output(4));
  mux_3918_nl <= MUX_s_1_2_2(or_4127_nl, mux_3917_nl, fsm_output(0));
  nor_1305_nl <= NOT((fsm_output(2)) OR mux_3918_nl);
  modulo_add_base_1_sva_mx0c3 <= MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output(1));
  modulo_add_base_1_sva_mx0c4 <= and_dcpl_72 AND and_dcpl_478;
  modulo_add_base_1_sva_mx0c9 <= and_dcpl_92 AND and_dcpl_101;
  modulo_add_base_1_sva_mx0c14 <= and_dcpl_92 AND and_dcpl_458;
  modulo_add_base_1_sva_mx0c18 <= and_dcpl_148 AND and_dcpl_90;
  modulo_add_base_1_sva_mx0c21 <= and_dcpl_1083 AND and_dcpl_128;
  modulo_add_base_1_sva_mx0c26 <= and_dcpl_76 AND and_dcpl_158;
  modulo_add_base_1_sva_mx0c30 <= and_dcpl_476 AND and_dcpl_61;
  nor_1299_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(0))) OR (fsm_output(6))
      OR (NOT (fsm_output(4))) OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  nor_1300_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 3)/=STD_LOGIC_VECTOR'("01110")));
  mux_3946_nl <= MUX_s_1_2_2((fsm_output(3)), (NOT (fsm_output(3))), fsm_output(5));
  and_1283_nl <= (fsm_output(7)) AND mux_3946_nl;
  nor_2195_nl <= NOT((fsm_output(5)) OR (fsm_output(3)) OR (fsm_output(7)));
  mux_3947_nl <= MUX_s_1_2_2(and_1283_nl, nor_2195_nl, fsm_output(4));
  nor_1302_nl <= NOT((fsm_output(4)) OR (fsm_output(7)) OR (fsm_output(5)) OR (fsm_output(3)));
  mux_3948_nl <= MUX_s_1_2_2(mux_3947_nl, nor_1302_nl, fsm_output(6));
  mux_3949_nl <= MUX_s_1_2_2(nor_1300_nl, mux_3948_nl, fsm_output(0));
  and_1282_nl <= (fsm_output(2)) AND mux_3949_nl;
  mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 <= MUX_s_1_2_2(nor_1299_nl, and_1282_nl,
      fsm_output(1));
  mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c7 <= and_dcpl_1083 AND and_dcpl_90;
  nor_1298_nl <= NOT((fsm_output(1)) OR (NOT (fsm_output(5))) OR (fsm_output(2))
      OR (NOT (fsm_output(4))) OR (fsm_output(7)) OR not_tmp_1345);
  mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 <= MUX_s_1_2_2(mux_3678_cse, nor_1298_nl,
      fsm_output(0));
  nor_1289_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111100")));
  nor_1290_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(7))) OR (fsm_output(3))
      OR (NOT (fsm_output(4))) OR (fsm_output(1)));
  or_4198_nl <= (fsm_output(3)) OR (NOT((fsm_output(4)) AND (fsm_output(1))));
  mux_3989_nl <= MUX_s_1_2_2(or_4198_nl, or_3852_cse, fsm_output(7));
  nor_1291_nl <= NOT((fsm_output(6)) OR mux_3989_nl);
  mux_3990_nl <= MUX_s_1_2_2(nor_1290_nl, nor_1291_nl, fsm_output(5));
  or_4195_nl <= (fsm_output(7)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(4)))
      OR (fsm_output(1));
  or_4194_nl <= (fsm_output(7)) OR (NOT (fsm_output(3))) OR (fsm_output(4)) OR (fsm_output(1));
  mux_3988_nl <= MUX_s_1_2_2(or_4195_nl, or_4194_nl, fsm_output(6));
  nor_1292_nl <= NOT((fsm_output(5)) OR mux_3988_nl);
  mux_3991_nl <= MUX_s_1_2_2(mux_3990_nl, nor_1292_nl, fsm_output(2));
  mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 <= MUX_s_1_2_2(nor_1289_nl, mux_3991_nl,
      fsm_output(0));
  nor_1283_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(6))) OR (fsm_output(0))
      OR (fsm_output(2)));
  nor_1284_nl <= NOT((fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(0)) OR (fsm_output(2)));
  mux_4007_nl <= MUX_s_1_2_2(nor_1283_nl, nor_1284_nl, fsm_output(4));
  and_1279_nl <= (fsm_output(3)) AND mux_4007_nl;
  mux_4006_nl <= MUX_s_1_2_2(nor_1730_cse, and_2893_cse, fsm_output(6));
  nor_1285_nl <= NOT((fsm_output(3)) OR (NOT(CONV_SL_1_1(fsm_output(5 DOWNTO 4)=STD_LOGIC_VECTOR'("11"))
      AND mux_4006_nl)));
  mux_4008_nl <= MUX_s_1_2_2(and_1279_nl, nor_1285_nl, fsm_output(1));
  or_4220_nl <= (NOT (fsm_output(4))) OR (fsm_output(5)) OR (fsm_output(6)) OR (fsm_output(0))
      OR (fsm_output(2));
  or_4219_nl <= (fsm_output(4)) OR (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(0))
      OR (fsm_output(2));
  mux_4005_nl <= MUX_s_1_2_2(or_4220_nl, or_4219_nl, fsm_output(3));
  nor_1287_nl <= NOT((fsm_output(1)) OR mux_4005_nl);
  operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm_mx0c3 <=
      MUX_s_1_2_2(mux_4008_nl, nor_1287_nl, fsm_output(7));
  nor_1278_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 2)/=STD_LOGIC_VECTOR'("001100")));
  nor_1279_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(2))) OR (fsm_output(7))
      OR (NOT (fsm_output(4))));
  nor_1280_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(7)))
      OR (fsm_output(4)));
  mux_4023_nl <= MUX_s_1_2_2(nor_1279_nl, nor_1280_nl, fsm_output(5));
  or_4243_nl <= (NOT (fsm_output(2))) OR (NOT (fsm_output(7))) OR (fsm_output(4));
  or_4131_nl <= (fsm_output(2)) OR (fsm_output(4)) OR (fsm_output(7));
  mux_4022_nl <= MUX_s_1_2_2(or_4243_nl, or_4131_nl, fsm_output(6));
  nor_1281_nl <= NOT((fsm_output(5)) OR mux_4022_nl);
  mux_4024_nl <= MUX_s_1_2_2(mux_4023_nl, nor_1281_nl, fsm_output(3));
  mux_4025_nl <= MUX_s_1_2_2(nor_1278_nl, mux_4024_nl, fsm_output(1));
  nor_1282_nl <= NOT(CONV_SL_1_1(fsm_output(7 DOWNTO 1)/=STD_LOGIC_VECTOR'("0111010")));
  operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm_mx0c3 <=
      MUX_s_1_2_2(mux_4025_nl, nor_1282_nl, fsm_output(0));
  mux_4041_nl <= MUX_s_1_2_2((fsm_output(6)), (NOT (fsm_output(6))), fsm_output(4));
  and_1277_nl <= nor_673_cse AND mux_4041_nl;
  nor_1274_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(5))) OR (fsm_output(0))
      OR (NOT((fsm_output(4)) AND (fsm_output(6)))));
  mux_4042_nl <= MUX_s_1_2_2(and_1277_nl, nor_1274_nl, fsm_output(2));
  nor_1275_nl <= NOT((NOT (fsm_output(2))) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(5)))
      OR (NOT (fsm_output(0))) OR (fsm_output(4)) OR (fsm_output(6)));
  mux_4043_nl <= MUX_s_1_2_2(mux_4042_nl, nor_1275_nl, fsm_output(1));
  nor_1276_nl <= NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR (fsm_output(4))
      OR (fsm_output(6)));
  nor_1277_nl <= NOT((fsm_output(5)) OR (NOT (fsm_output(0))) OR (fsm_output(4))
      OR (fsm_output(6)));
  mux_4040_nl <= MUX_s_1_2_2(nor_1276_nl, nor_1277_nl, fsm_output(3));
  and_1278_nl <= nor_2247_cse AND mux_4040_nl;
  operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm_mx0c3 <=
      MUX_s_1_2_2(mux_4043_nl, and_1278_nl, fsm_output(7));
  S2_OUTER_LOOP_c_1_sva_mx0c1 <= and_dcpl_76 AND and_dcpl_101;
  S2_OUTER_LOOP_c_1_sva_mx0c2 <= and_dcpl_148 AND and_dcpl_115;
  or_345_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_315_cse AND (fsm_output(4))));
  mux_140_nl <= MUX_s_1_2_2(or_tmp_169, or_345_nl, fsm_output(7));
  and_116_ssc <= (NOT mux_140_nl) AND and_dcpl_105;
  or_412_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00001")))
      AND (fsm_output(4))));
  mux_192_nl <= MUX_s_1_2_2(or_tmp_169, or_412_nl, fsm_output(7));
  and_164_ssc <= (NOT mux_192_nl) AND and_dcpl_105;
  or_470_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_447_cse AND (fsm_output(4))));
  mux_242_nl <= MUX_s_1_2_2(or_tmp_169, or_470_nl, fsm_output(7));
  and_191_ssc <= (NOT mux_242_nl) AND and_dcpl_105;
  or_525_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00011")))
      AND (fsm_output(4))));
  mux_294_nl <= MUX_s_1_2_2(or_tmp_169, or_525_nl, fsm_output(7));
  and_207_ssc <= (NOT mux_294_nl) AND and_dcpl_105;
  or_581_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_555_cse AND (fsm_output(4))));
  mux_358_nl <= MUX_s_1_2_2(or_tmp_169, or_581_nl, fsm_output(7));
  and_221_ssc <= (NOT mux_358_nl) AND and_dcpl_105;
  or_657_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00101")))
      AND (fsm_output(4))));
  mux_409_nl <= MUX_s_1_2_2(or_tmp_169, or_657_nl, fsm_output(7));
  and_237_ssc <= (NOT mux_409_nl) AND and_dcpl_105;
  or_713_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_684_cse AND (fsm_output(4))));
  mux_456_nl <= MUX_s_1_2_2(or_tmp_169, or_713_nl, fsm_output(7));
  and_253_ssc <= (NOT mux_456_nl) AND and_dcpl_105;
  or_766_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00111")))
      AND (fsm_output(4))));
  mux_505_nl <= MUX_s_1_2_2(or_tmp_169, or_766_nl, fsm_output(7));
  and_262_ssc <= (NOT mux_505_nl) AND and_dcpl_105;
  or_822_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_795_cse AND (fsm_output(4))));
  mux_567_nl <= MUX_s_1_2_2(or_tmp_169, or_822_nl, fsm_output(7));
  and_271_ssc <= (NOT mux_567_nl) AND and_dcpl_105;
  or_881_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01001")))
      AND (fsm_output(4))));
  mux_615_nl <= MUX_s_1_2_2(or_tmp_169, or_881_nl, fsm_output(7));
  and_288_ssc <= (NOT mux_615_nl) AND and_dcpl_105;
  or_933_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_910_cse AND (fsm_output(4))));
  mux_662_nl <= MUX_s_1_2_2(or_tmp_169, or_933_nl, fsm_output(7));
  and_305_ssc <= (NOT mux_662_nl) AND and_dcpl_105;
  or_986_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01011")))
      AND (fsm_output(4))));
  mux_711_nl <= MUX_s_1_2_2(or_tmp_169, or_986_nl, fsm_output(7));
  and_316_ssc <= (NOT mux_711_nl) AND and_dcpl_105;
  or_1038_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_1012_cse AND (fsm_output(4))));
  mux_773_nl <= MUX_s_1_2_2(or_tmp_169, or_1038_nl, fsm_output(7));
  and_326_ssc <= (NOT mux_773_nl) AND and_dcpl_105;
  or_1105_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01101")))
      AND (fsm_output(4))));
  mux_821_nl <= MUX_s_1_2_2(or_tmp_169, or_1105_nl, fsm_output(7));
  and_339_ssc <= (NOT mux_821_nl) AND and_dcpl_105;
  or_1162_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND or_1133_cse AND (fsm_output(4))));
  mux_868_nl <= MUX_s_1_2_2(or_tmp_169, or_1162_nl, fsm_output(7));
  and_354_ssc <= (NOT mux_868_nl) AND and_dcpl_105;
  or_1212_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01111"))))
      AND (fsm_output(4))));
  mux_917_nl <= MUX_s_1_2_2(or_tmp_169, or_1212_nl, fsm_output(7));
  and_363_ssc <= (NOT mux_917_nl) AND and_dcpl_105;
  or_1265_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_980_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1265_nl);
  or_1267_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_980_nl));
  mux_981_nl <= MUX_s_1_2_2(or_tmp_169, or_1267_nl, fsm_output(7));
  and_372_ssc <= (NOT mux_981_nl) AND and_dcpl_105;
  or_1330_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0001"));
  mux_1031_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1330_nl);
  or_1331_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1031_nl));
  mux_1032_nl <= MUX_s_1_2_2(or_tmp_169, or_1331_nl, fsm_output(7));
  and_387_ssc <= (NOT mux_1032_nl) AND and_dcpl_105;
  or_1383_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0010"));
  mux_1081_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1383_nl);
  or_1384_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1081_nl));
  mux_1082_nl <= MUX_s_1_2_2(or_tmp_169, or_1384_nl, fsm_output(7));
  and_402_ssc <= (NOT mux_1082_nl) AND and_dcpl_105;
  or_1436_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0011"));
  mux_1133_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1436_nl);
  or_1437_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1133_nl));
  mux_1134_nl <= MUX_s_1_2_2(or_tmp_169, or_1437_nl, fsm_output(7));
  and_410_ssc <= (NOT mux_1134_nl) AND and_dcpl_105;
  or_1489_nl <= (S6_OUTER_LOOP_for_acc_tmp(0)) OR (S6_OUTER_LOOP_for_acc_tmp(3))
      OR (S6_OUTER_LOOP_for_acc_tmp(1));
  mux_1197_nl <= MUX_s_1_2_2(not_tmp_542, (fsm_output(4)), or_1489_nl);
  or_1491_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1197_nl));
  mux_1198_nl <= MUX_s_1_2_2(or_tmp_169, or_1491_nl, fsm_output(7));
  and_419_ssc <= (NOT mux_1198_nl) AND and_dcpl_105;
  or_1568_nl <= (NOT (S6_OUTER_LOOP_for_acc_tmp(0))) OR (S6_OUTER_LOOP_for_acc_tmp(3))
      OR (S6_OUTER_LOOP_for_acc_tmp(1));
  mux_1249_nl <= MUX_s_1_2_2(not_tmp_542, (fsm_output(4)), or_1568_nl);
  or_1569_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1249_nl));
  mux_1250_nl <= MUX_s_1_2_2(or_tmp_169, or_1569_nl, fsm_output(7));
  and_433_ssc <= (NOT mux_1250_nl) AND and_dcpl_105;
  or_1627_nl <= (S6_OUTER_LOOP_for_acc_tmp(0)) OR (S6_OUTER_LOOP_for_acc_tmp(3));
  mux_1299_nl <= MUX_s_1_2_2(not_tmp_598, (fsm_output(4)), or_1627_nl);
  or_1629_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1299_nl));
  mux_1300_nl <= MUX_s_1_2_2(or_tmp_169, or_1629_nl, fsm_output(7));
  and_447_ssc <= (NOT mux_1300_nl) AND and_dcpl_105;
  or_1686_nl <= (NOT (S6_OUTER_LOOP_for_acc_tmp(0))) OR (S6_OUTER_LOOP_for_acc_tmp(3));
  mux_1351_nl <= MUX_s_1_2_2(not_tmp_598, (fsm_output(4)), or_1686_nl);
  or_1687_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1351_nl));
  mux_1352_nl <= MUX_s_1_2_2(or_tmp_169, or_1687_nl, fsm_output(7));
  and_455_ssc <= (NOT mux_1352_nl) AND and_dcpl_105;
  or_1741_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1000"));
  mux_1415_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1741_nl);
  or_1742_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1415_nl));
  mux_1416_nl <= MUX_s_1_2_2(or_tmp_169, or_1742_nl, fsm_output(7));
  and_464_ssc <= (NOT mux_1416_nl) AND and_dcpl_105;
  or_1804_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1001"));
  mux_1466_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1804_nl);
  or_1805_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1466_nl));
  mux_1467_nl <= MUX_s_1_2_2(or_tmp_169, or_1805_nl, fsm_output(7));
  and_475_ssc <= (NOT mux_1467_nl) AND and_dcpl_105;
  or_1857_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("1010"));
  mux_1516_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), or_1857_nl);
  or_1858_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1516_nl));
  mux_1517_nl <= MUX_s_1_2_2(or_tmp_169, or_1858_nl, fsm_output(7));
  and_490_ssc <= (NOT mux_1517_nl) AND and_dcpl_105;
  nand_382_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO 0)=STD_LOGIC_VECTOR'("1011")));
  mux_1568_nl <= MUX_s_1_2_2(not_tmp_451, (fsm_output(4)), nand_382_nl);
  or_1916_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1568_nl));
  mux_1569_nl <= MUX_s_1_2_2(or_tmp_169, or_1916_nl, fsm_output(7));
  and_498_ssc <= (NOT mux_1569_nl) AND and_dcpl_105;
  or_1968_nl <= (S6_OUTER_LOOP_for_acc_tmp(0)) OR (NOT (S6_OUTER_LOOP_for_acc_tmp(3)))
      OR (S6_OUTER_LOOP_for_acc_tmp(1));
  mux_1632_nl <= MUX_s_1_2_2(not_tmp_542, (fsm_output(4)), or_1968_nl);
  or_1969_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1632_nl));
  mux_1633_nl <= MUX_s_1_2_2(or_tmp_169, or_1969_nl, fsm_output(7));
  and_507_ssc <= (NOT mux_1633_nl) AND and_dcpl_105;
  or_2032_nl <= (NOT (S6_OUTER_LOOP_for_acc_tmp(0))) OR (NOT (S6_OUTER_LOOP_for_acc_tmp(3)))
      OR (S6_OUTER_LOOP_for_acc_tmp(1));
  mux_1683_nl <= MUX_s_1_2_2(not_tmp_542, (fsm_output(4)), or_2032_nl);
  or_2033_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1683_nl));
  mux_1684_nl <= MUX_s_1_2_2(or_tmp_169, or_2033_nl, fsm_output(7));
  and_518_ssc <= (NOT mux_1684_nl) AND and_dcpl_105;
  and_2137_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO 1)=STD_LOGIC_VECTOR'("1111"))))
      AND (fsm_output(4));
  mux_1733_nl <= MUX_s_1_2_2(and_2137_nl, (fsm_output(4)), S6_OUTER_LOOP_for_acc_tmp(0));
  or_2084_nl <= (fsm_output(6)) OR (NOT((fsm_output(2)) AND mux_1733_nl));
  mux_1734_nl <= MUX_s_1_2_2(or_tmp_169, or_2084_nl, fsm_output(7));
  and_532_ssc <= (NOT mux_1734_nl) AND and_dcpl_105;
  nand_109_nl <= NOT((NOT((fsm_output(6)) OR (NOT (fsm_output(2))))) AND (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11111"))))
      AND (fsm_output(4)));
  mux_1782_nl <= MUX_s_1_2_2(or_tmp_169, nand_109_nl, fsm_output(7));
  and_540_ssc <= (NOT mux_1782_nl) AND and_dcpl_105;
  and_173_ssc <= and_dcpl_126 AND and_dcpl_158;
  and_174_ssc <= and_dcpl_67 AND and_dcpl_75;
  and_615_ssc <= and_dcpl_447 AND and_dcpl_478;
  and_616_ssc <= and_dcpl_67 AND and_dcpl_115;
  butterFly_7_or_ssc_31 <= and_dcpl_102 OR and_dcpl_114;
  butterFly_7_or_201_cse <= butterFly_7_or_ssc_31 OR and_116_ssc OR and_dcpl_125;
  butterFly_7_or_ssc_30 <= and_dcpl_149 OR and_dcpl_154;
  butterFly_7_or_204_cse <= butterFly_7_or_ssc_30 OR and_164_ssc OR and_dcpl_157;
  butterFly_7_or_ssc_29 <= and_dcpl_171 OR and_dcpl_173;
  butterFly_7_or_207_cse <= butterFly_7_or_ssc_29 OR and_191_ssc OR and_dcpl_177;
  butterFly_7_or_ssc_28 <= and_dcpl_184 OR and_dcpl_187;
  butterFly_7_or_210_cse <= butterFly_7_or_ssc_28 OR and_207_ssc OR and_dcpl_190;
  butterFly_7_or_213_cse <= butterFly_7_or_ssc_31 OR and_221_ssc OR and_dcpl_201;
  butterFly_7_or_216_cse <= butterFly_7_or_ssc_30 OR and_237_ssc OR and_dcpl_213;
  butterFly_7_or_219_cse <= butterFly_7_or_ssc_29 OR and_253_ssc OR and_dcpl_224;
  butterFly_7_or_222_cse <= butterFly_7_or_ssc_28 OR and_262_ssc OR and_dcpl_230;
  butterFly_7_or_225_cse <= butterFly_7_or_ssc_31 OR and_271_ssc OR and_dcpl_239;
  butterFly_7_or_228_cse <= butterFly_7_or_ssc_30 OR and_288_ssc OR and_dcpl_252;
  butterFly_7_or_231_cse <= butterFly_7_or_ssc_29 OR and_305_ssc OR and_dcpl_265;
  butterFly_7_or_234_cse <= butterFly_7_or_ssc_28 OR and_316_ssc OR and_dcpl_272;
  butterFly_7_or_237_cse <= butterFly_7_or_ssc_31 OR and_326_ssc OR and_dcpl_279;
  butterFly_7_or_240_cse <= butterFly_7_or_ssc_30 OR and_339_ssc OR and_dcpl_289;
  butterFly_7_or_243_cse <= butterFly_7_or_ssc_29 OR and_354_ssc OR and_dcpl_299;
  butterFly_7_or_246_cse <= butterFly_7_or_ssc_28 OR and_363_ssc OR and_dcpl_305;
  butterFly_7_or_249_cse <= butterFly_7_or_ssc_31 OR and_372_ssc OR and_dcpl_314;
  butterFly_7_or_252_cse <= butterFly_7_or_ssc_30 OR and_387_ssc OR and_dcpl_325;
  butterFly_7_or_255_cse <= butterFly_7_or_ssc_29 OR and_402_ssc OR and_dcpl_336;
  butterFly_7_or_258_cse <= butterFly_7_or_ssc_28 OR and_410_ssc OR and_dcpl_342;
  butterFly_7_or_261_cse <= butterFly_7_or_ssc_31 OR and_419_ssc OR and_dcpl_351;
  butterFly_7_or_264_cse <= butterFly_7_or_ssc_30 OR and_433_ssc OR and_dcpl_361;
  butterFly_7_or_267_cse <= butterFly_7_or_ssc_29 OR and_447_ssc OR and_dcpl_371;
  butterFly_7_or_270_cse <= butterFly_7_or_ssc_28 OR and_455_ssc OR and_dcpl_377;
  butterFly_7_or_273_cse <= butterFly_7_or_ssc_31 OR and_464_ssc OR and_dcpl_384;
  butterFly_7_or_276_cse <= butterFly_7_or_ssc_30 OR and_475_ssc OR and_dcpl_393;
  butterFly_7_or_279_cse <= butterFly_7_or_ssc_29 OR and_490_ssc OR and_dcpl_404;
  butterFly_7_or_282_cse <= butterFly_7_or_ssc_28 OR and_498_ssc OR and_dcpl_410;
  butterFly_7_or_285_cse <= butterFly_7_or_ssc_31 OR and_507_ssc OR and_dcpl_417;
  butterFly_7_or_288_cse <= butterFly_7_or_ssc_30 OR and_518_ssc OR and_dcpl_426;
  butterFly_7_or_291_cse <= butterFly_7_or_ssc_29 OR and_532_ssc OR and_dcpl_436;
  butterFly_7_or_294_cse <= butterFly_7_or_ssc_28 OR and_540_ssc OR and_dcpl_442;
  butterFly_3_or_264_cse <= and_dcpl_457 OR and_dcpl_477;
  butterFly_3_butterFly_3_mux_rmff <= MUX_v_3_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), butterFly_3_or_264_cse);
  butterFly_3_butterFly_3_or_rmff <= ((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) AND
      (NOT and_dcpl_457)) OR and_dcpl_477;
  butterFly_3_or_201_cse <= and_dcpl_450 OR and_dcpl_470;
  butterFly_3_or_203_cse <= and_dcpl_450 OR and_dcpl_511;
  butterFly_3_or_205_cse <= and_dcpl_450 OR and_dcpl_537;
  butterFly_3_or_207_cse <= and_dcpl_450 OR and_dcpl_553;
  butterFly_3_or_209_cse <= and_dcpl_450 OR and_dcpl_570;
  butterFly_3_or_211_cse <= and_dcpl_450 OR and_dcpl_588;
  butterFly_3_or_213_cse <= and_dcpl_450 OR and_dcpl_600;
  butterFly_3_or_215_cse <= and_dcpl_450 OR and_dcpl_609;
  butterFly_3_or_217_cse <= and_dcpl_450 OR and_dcpl_622;
  butterFly_3_or_219_cse <= and_dcpl_450 OR and_dcpl_640;
  butterFly_3_or_221_cse <= and_dcpl_450 OR and_dcpl_655;
  butterFly_3_or_223_cse <= and_dcpl_450 OR and_dcpl_667;
  butterFly_3_or_225_cse <= and_dcpl_450 OR and_dcpl_679;
  butterFly_3_or_227_cse <= and_dcpl_450 OR and_dcpl_692;
  butterFly_3_or_229_cse <= and_dcpl_450 OR and_dcpl_703;
  butterFly_3_or_231_cse <= and_dcpl_450 OR and_dcpl_712;
  butterFly_3_or_233_cse <= and_dcpl_450 OR and_dcpl_724;
  butterFly_3_or_235_cse <= and_dcpl_450 OR and_dcpl_742;
  butterFly_3_or_237_cse <= and_dcpl_450 OR and_dcpl_758;
  butterFly_3_or_239_cse <= and_dcpl_450 OR and_dcpl_770;
  butterFly_3_or_241_cse <= and_dcpl_450 OR and_dcpl_782;
  butterFly_3_or_243_cse <= and_dcpl_450 OR and_dcpl_795;
  butterFly_3_or_245_cse <= and_dcpl_450 OR and_dcpl_806;
  butterFly_3_or_247_cse <= and_dcpl_450 OR and_dcpl_815;
  butterFly_3_or_249_cse <= and_dcpl_450 OR and_dcpl_827;
  butterFly_3_or_251_cse <= and_dcpl_450 OR and_dcpl_843;
  butterFly_3_or_253_cse <= and_dcpl_450 OR and_dcpl_858;
  butterFly_3_or_255_cse <= and_dcpl_450 OR and_dcpl_870;
  butterFly_3_or_257_cse <= and_dcpl_450 OR and_dcpl_882;
  butterFly_3_or_259_cse <= and_dcpl_450 OR and_dcpl_894;
  butterFly_3_or_261_cse <= and_dcpl_450 OR and_dcpl_905;
  butterFly_3_or_263_cse <= and_dcpl_450 OR and_dcpl_914;
  butterFly_3_or_296_cse <= and_dcpl_448 OR and_dcpl_454 OR and_dcpl_459;
  butterFly_3_or_301_cse <= and_dcpl_448 OR and_dcpl_506 OR and_dcpl_507;
  butterFly_3_or_306_cse <= and_dcpl_448 OR and_dcpl_533 OR and_dcpl_534;
  butterFly_3_or_311_cse <= and_dcpl_448 OR and_dcpl_551 OR and_dcpl_552;
  nor_2160_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (NOT nor_tmp_31));
  and_2091_nl <= (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(3))
      AND (fsm_output(5));
  mux_145_nl <= MUX_s_1_2_2(nor_2160_nl, and_2091_nl, fsm_output(6));
  mux_143_nl <= MUX_s_1_2_2(nor_1311_cse, nor_tmp_31, fsm_output(2));
  mux_144_nl <= MUX_s_1_2_2(mux_143_nl, and_1665_cse, fsm_output(0));
  or_352_nl <= (fsm_output(6)) OR mux_144_nl;
  mux_146_cse <= MUX_s_1_2_2(mux_145_nl, or_352_nl, fsm_output(7));
  and_2092_nl <= (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(3)) AND (fsm_output(5));
  mux_142_nl <= MUX_s_1_2_2(and_2092_nl, and_1665_cse, fsm_output(0));
  and_142_cse <= (fsm_output(7)) AND ((fsm_output(6)) OR mux_142_nl);
  nor_2158_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_148_nl <= MUX_s_1_2_2(nor_2157_cse, nor_2158_nl, fsm_output(0));
  mux_149_nl <= MUX_s_1_2_2(nor_2156_cse, mux_148_nl, fsm_output(6));
  nor_2159_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_150_nl <= MUX_s_1_2_2(mux_149_nl, nor_2159_nl, or_309_cse);
  mux_151_nl <= MUX_s_1_2_2(mux_150_nl, (fsm_output(6)), fsm_output(7));
  mux_147_nl <= MUX_s_1_2_2(mux_146_cse, and_142_cse, or_348_cse);
  butterFly_7_butterFly_7_or_rmff <= MUX_s_1_2_2(mux_151_nl, mux_147_nl, fsm_output(4));
  mux_204_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_435_cse);
  or_420_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_203_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_420_nl);
  mux_205_nl <= MUX_s_1_2_2(mux_204_nl, mux_203_nl, fsm_output(3));
  and_2078_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4)) OR (fsm_output(7))) AND (fsm_output(6));
  and_2079_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)) OR (fsm_output(7))) AND (fsm_output(6));
  mux_200_nl <= MUX_s_1_2_2(and_2078_nl, and_2079_nl, fsm_output(0));
  mux_201_nl <= MUX_s_1_2_2(mux_200_nl, nor_tmp_35, fsm_output(3));
  mux_206_nl <= MUX_s_1_2_2(mux_205_nl, mux_201_nl, fsm_output(5));
  mux_207_nl <= MUX_s_1_2_2(nor_tmp_35, mux_206_nl, nor_44_cse);
  or_415_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(3))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_198_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_415_nl);
  mux_195_nl <= MUX_s_1_2_2(or_324_cse, (fsm_output(7)), or_2242_cse);
  mux_196_nl <= MUX_s_1_2_2(nor_tmp_35, mux_195_nl, and_2080_cse);
  mux_197_nl <= MUX_s_1_2_2(mux_196_nl, mux_295_cse, fsm_output(1));
  mux_199_nl <= MUX_s_1_2_2(mux_198_nl, mux_197_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_2_rmff <= MUX_s_1_2_2(mux_207_nl, mux_199_nl, fsm_output(4));
  or_478_nl <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_256_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_478_nl);
  and_2069_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_2070_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_254_nl <= MUX_s_1_2_2(and_2069_nl, and_2070_nl, fsm_output(0));
  or_475_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_253_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_475_nl);
  mux_255_nl <= MUX_s_1_2_2(mux_254_nl, mux_253_nl, fsm_output(3));
  mux_257_nl <= MUX_s_1_2_2(mux_256_nl, mux_255_nl, fsm_output(1));
  mux_258_nl <= MUX_s_1_2_2(mux_257_nl, nor_tmp_35, fsm_output(2));
  or_474_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_251_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_474_nl);
  or_473_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_247_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_473_nl);
  mux_248_nl <= MUX_s_1_2_2(mux_247_nl, mux_3731_cse, fsm_output(0));
  mux_249_nl <= MUX_s_1_2_2(nor_tmp_35, mux_248_nl, fsm_output(3));
  mux_250_nl <= MUX_s_1_2_2(mux_249_nl, mux_295_cse, fsm_output(1));
  mux_252_nl <= MUX_s_1_2_2(mux_251_nl, mux_250_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_4_rmff <= MUX_s_1_2_2(mux_258_nl, mux_252_nl, fsm_output(4));
  or_530_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (fsm_output(5));
  mux_309_cse <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_530_nl);
  mux_298_cse <= MUX_s_1_2_2(nor_tmp_35, mux_297_cse, fsm_output(2));
  nor_78_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5))));
  mux_306_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_78_nl);
  mux_305_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, and_2080_cse);
  mux_307_nl <= MUX_s_1_2_2(mux_306_nl, mux_305_nl, fsm_output(1));
  mux_308_cse <= MUX_s_1_2_2(mux_307_nl, mux_297_cse, fsm_output(2));
  mux_310_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_302, fsm_output(1));
  mux_311_nl <= MUX_s_1_2_2(mux_310_nl, nor_tmp_35, fsm_output(2));
  mux_312_nl <= MUX_s_1_2_2(mux_311_nl, mux_308_cse, fsm_output(4));
  mux_303_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_302, nor_44_cse);
  mux_304_nl <= MUX_s_1_2_2(mux_303_nl, mux_298_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_6_rmff <= MUX_s_1_2_2(mux_312_nl, mux_304_nl, or_2242_cse);
  nor_2094_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_365_nl <= MUX_s_1_2_2(nor_2157_cse, nor_2094_nl, fsm_output(0));
  mux_366_nl <= MUX_s_1_2_2(nor_2156_cse, mux_365_nl, fsm_output(6));
  nor_2095_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_367_nl <= MUX_s_1_2_2(mux_366_nl, nor_2095_nl, or_549_cse);
  mux_368_nl <= MUX_s_1_2_2(mux_367_nl, (fsm_output(6)), fsm_output(7));
  mux_364_nl <= MUX_s_1_2_2(mux_146_cse, and_142_cse, or_582_cse);
  butterFly_7_butterFly_7_or_8_rmff <= MUX_s_1_2_2(mux_368_nl, mux_364_nl, fsm_output(4));
  mux_420_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_132_cse);
  or_663_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_419_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_663_nl);
  mux_421_nl <= MUX_s_1_2_2(mux_420_nl, mux_419_nl, fsm_output(3));
  and_2036_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4)) OR (fsm_output(7))) AND (fsm_output(6));
  and_2037_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)) OR (fsm_output(7))) AND (fsm_output(6));
  mux_416_nl <= MUX_s_1_2_2(and_2036_nl, and_2037_nl, fsm_output(0));
  mux_417_nl <= MUX_s_1_2_2(mux_416_nl, nor_tmp_35, fsm_output(3));
  mux_422_nl <= MUX_s_1_2_2(mux_421_nl, mux_417_nl, fsm_output(5));
  mux_423_nl <= MUX_s_1_2_2(nor_tmp_35, mux_422_nl, nor_44_cse);
  nor_105_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(3))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_414_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_105_nl);
  mux_411_nl <= MUX_s_1_2_2((fsm_output(7)), or_324_cse, nor_701_cse);
  mux_412_nl <= MUX_s_1_2_2(nor_tmp_35, mux_411_nl, and_2080_cse);
  mux_413_nl <= MUX_s_1_2_2(mux_412_nl, mux_295_cse, fsm_output(1));
  mux_415_nl <= MUX_s_1_2_2(mux_414_nl, mux_413_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_10_rmff <= MUX_s_1_2_2(mux_423_nl, mux_415_nl, fsm_output(4));
  nor_126_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_469_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_126_nl);
  and_2027_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_2028_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_467_nl <= MUX_s_1_2_2(and_2027_nl, and_2028_nl, fsm_output(0));
  or_714_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_466_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_714_nl);
  mux_468_nl <= MUX_s_1_2_2(mux_467_nl, mux_466_nl, fsm_output(3));
  mux_470_nl <= MUX_s_1_2_2(mux_469_nl, mux_468_nl, fsm_output(1));
  mux_471_nl <= MUX_s_1_2_2(mux_470_nl, nor_tmp_35, fsm_output(2));
  nor_121_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_464_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_121_nl);
  nor_120_nl <= NOT((NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001")));
  mux_460_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, nor_120_nl);
  mux_461_nl <= MUX_s_1_2_2(mux_460_nl, mux_3731_cse, fsm_output(0));
  mux_462_nl <= MUX_s_1_2_2(nor_tmp_35, mux_461_nl, fsm_output(3));
  mux_463_nl <= MUX_s_1_2_2(mux_462_nl, mux_295_cse, fsm_output(1));
  mux_465_nl <= MUX_s_1_2_2(mux_464_nl, mux_463_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_12_rmff <= MUX_s_1_2_2(mux_471_nl, mux_465_nl, fsm_output(4));
  mux_522_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_516, nor_44_cse);
  mux_523_nl <= MUX_s_1_2_2(mux_522_nl, mux_298_cse, fsm_output(4));
  mux_518_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_516, fsm_output(1));
  mux_519_nl <= MUX_s_1_2_2(mux_518_nl, nor_tmp_35, fsm_output(2));
  mux_520_nl <= MUX_s_1_2_2(mux_519_nl, mux_308_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_14_rmff <= MUX_s_1_2_2(mux_523_nl, mux_520_nl, nor_701_cse);
  nor_2043_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_574_nl <= MUX_s_1_2_2(nor_2157_cse, nor_2043_nl, fsm_output(0));
  mux_575_nl <= MUX_s_1_2_2(nor_2156_cse, mux_574_nl, fsm_output(6));
  nor_2044_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_576_nl <= MUX_s_1_2_2(mux_575_nl, nor_2044_nl, or_789_cse);
  mux_577_nl <= MUX_s_1_2_2(mux_576_nl, (fsm_output(6)), fsm_output(7));
  mux_573_nl <= MUX_s_1_2_2(mux_146_cse, and_142_cse, or_823_cse);
  butterFly_7_butterFly_7_or_16_rmff <= MUX_s_1_2_2(mux_577_nl, mux_573_nl, fsm_output(4));
  mux_626_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_898_cse);
  or_889_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_625_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_889_nl);
  mux_627_nl <= MUX_s_1_2_2(mux_626_nl, mux_625_nl, fsm_output(3));
  and_1994_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4)) OR (fsm_output(7))) AND (fsm_output(6));
  and_1995_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)) OR (fsm_output(7))) AND (fsm_output(6));
  mux_622_nl <= MUX_s_1_2_2(and_1994_nl, and_1995_nl, fsm_output(0));
  mux_623_nl <= MUX_s_1_2_2(mux_622_nl, nor_tmp_35, fsm_output(3));
  mux_628_nl <= MUX_s_1_2_2(mux_627_nl, mux_623_nl, fsm_output(5));
  mux_629_nl <= MUX_s_1_2_2(nor_tmp_35, mux_628_nl, nor_44_cse);
  or_884_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(3))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_620_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_884_nl);
  mux_617_nl <= MUX_s_1_2_2(or_324_cse, (fsm_output(7)), or_2619_cse);
  mux_618_nl <= MUX_s_1_2_2(nor_tmp_35, mux_617_nl, and_2080_cse);
  mux_619_nl <= MUX_s_1_2_2(mux_618_nl, mux_295_cse, fsm_output(1));
  mux_621_nl <= MUX_s_1_2_2(mux_620_nl, mux_619_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_18_rmff <= MUX_s_1_2_2(mux_629_nl, mux_621_nl, fsm_output(4));
  or_939_nl <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_675_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_939_nl);
  and_1985_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1986_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_673_nl <= MUX_s_1_2_2(and_1985_nl, and_1986_nl, fsm_output(0));
  or_936_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_672_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_936_nl);
  mux_674_nl <= MUX_s_1_2_2(mux_673_nl, mux_672_nl, fsm_output(3));
  mux_676_nl <= MUX_s_1_2_2(mux_675_nl, mux_674_nl, fsm_output(1));
  mux_677_nl <= MUX_s_1_2_2(mux_676_nl, nor_tmp_35, fsm_output(2));
  or_935_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_670_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_935_nl);
  or_934_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"));
  mux_666_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_934_nl);
  mux_667_nl <= MUX_s_1_2_2(mux_666_nl, mux_3731_cse, fsm_output(0));
  mux_668_nl <= MUX_s_1_2_2(nor_tmp_35, mux_667_nl, fsm_output(3));
  mux_669_nl <= MUX_s_1_2_2(mux_668_nl, mux_295_cse, fsm_output(1));
  mux_671_nl <= MUX_s_1_2_2(mux_670_nl, mux_669_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_20_rmff <= MUX_s_1_2_2(mux_677_nl, mux_671_nl, fsm_output(4));
  mux_727_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_719, fsm_output(1));
  mux_728_nl <= MUX_s_1_2_2(mux_727_nl, nor_tmp_35, fsm_output(2));
  mux_729_nl <= MUX_s_1_2_2(mux_728_nl, mux_308_cse, fsm_output(4));
  mux_720_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_719, nor_44_cse);
  mux_721_nl <= MUX_s_1_2_2(mux_720_nl, mux_298_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_22_rmff <= MUX_s_1_2_2(mux_729_nl, mux_721_nl, or_2619_cse);
  nor_1991_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_780_nl <= MUX_s_1_2_2(nor_2157_cse, nor_1991_nl, fsm_output(0));
  mux_781_nl <= MUX_s_1_2_2(nor_2156_cse, mux_780_nl, fsm_output(6));
  nor_1992_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_782_nl <= MUX_s_1_2_2(mux_781_nl, nor_1992_nl, or_1006_cse);
  mux_783_nl <= MUX_s_1_2_2(mux_782_nl, (fsm_output(6)), fsm_output(7));
  mux_779_nl <= MUX_s_1_2_2(mux_146_cse, and_142_cse, or_1039_cse);
  butterFly_7_butterFly_7_or_24_rmff <= MUX_s_1_2_2(mux_783_nl, mux_779_nl, fsm_output(4));
  mux_832_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_245_cse);
  or_1111_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4;
  mux_831_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1111_nl);
  mux_833_nl <= MUX_s_1_2_2(mux_832_nl, mux_831_nl, fsm_output(3));
  and_1950_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4)) OR (fsm_output(7))) AND (fsm_output(6));
  and_1951_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)) OR (fsm_output(7))) AND (fsm_output(6));
  mux_828_nl <= MUX_s_1_2_2(and_1950_nl, and_1951_nl, fsm_output(0));
  mux_829_nl <= MUX_s_1_2_2(mux_828_nl, nor_tmp_35, fsm_output(3));
  mux_834_nl <= MUX_s_1_2_2(mux_833_nl, mux_829_nl, fsm_output(5));
  mux_835_nl <= MUX_s_1_2_2(nor_tmp_35, mux_834_nl, nor_44_cse);
  and_1952_nl <= (fsm_output(1)) AND (fsm_output(5)) AND (NOT (fsm_output(3))) AND
      (fsm_output(0)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("011"));
  mux_826_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1952_nl);
  mux_823_nl <= MUX_s_1_2_2((fsm_output(7)), or_324_cse, nor_817_cse);
  mux_824_nl <= MUX_s_1_2_2(nor_tmp_35, mux_823_nl, and_2080_cse);
  mux_825_nl <= MUX_s_1_2_2(mux_824_nl, mux_295_cse, fsm_output(1));
  mux_827_nl <= MUX_s_1_2_2(mux_826_nl, mux_825_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_26_rmff <= MUX_s_1_2_2(mux_835_nl, mux_827_nl, fsm_output(4));
  nor_257_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011")));
  mux_881_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_257_nl);
  and_1939_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1940_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_879_nl <= MUX_s_1_2_2(and_1939_nl, and_1940_nl, fsm_output(0));
  or_1163_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1110"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(5));
  mux_878_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1163_nl);
  mux_880_nl <= MUX_s_1_2_2(mux_879_nl, mux_878_nl, fsm_output(3));
  mux_882_nl <= MUX_s_1_2_2(mux_881_nl, mux_880_nl, fsm_output(1));
  mux_883_nl <= MUX_s_1_2_2(mux_882_nl, nor_tmp_35, fsm_output(2));
  nor_252_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011")));
  mux_876_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_252_nl);
  and_1941_nl <= (fsm_output(5)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("011"));
  mux_872_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, and_1941_nl);
  mux_873_nl <= MUX_s_1_2_2(mux_872_nl, mux_3731_cse, fsm_output(0));
  mux_874_nl <= MUX_s_1_2_2(nor_tmp_35, mux_873_nl, fsm_output(3));
  mux_875_nl <= MUX_s_1_2_2(mux_874_nl, mux_295_cse, fsm_output(1));
  mux_877_nl <= MUX_s_1_2_2(mux_876_nl, mux_875_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_28_rmff <= MUX_s_1_2_2(mux_883_nl, mux_877_nl, fsm_output(4));
  mux_934_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_928, nor_44_cse);
  mux_935_nl <= MUX_s_1_2_2(mux_934_nl, mux_298_cse, fsm_output(4));
  mux_930_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_928, fsm_output(1));
  mux_931_nl <= MUX_s_1_2_2(mux_930_nl, nor_tmp_35, fsm_output(2));
  mux_932_nl <= MUX_s_1_2_2(mux_931_nl, mux_308_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_30_rmff <= MUX_s_1_2_2(mux_935_nl, mux_932_nl, nor_817_cse);
  nor_1940_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  nor_1943_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_988_nl <= MUX_s_1_2_2(nor_2157_cse, nor_1943_nl, fsm_output(0));
  mux_989_nl <= MUX_s_1_2_2(nor_2156_cse, mux_988_nl, fsm_output(6));
  nor_296_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_990_nl <= MUX_s_1_2_2(nor_1940_nl, mux_989_nl, nor_296_nl);
  mux_991_nl <= MUX_s_1_2_2(mux_990_nl, (fsm_output(6)), fsm_output(7));
  mux_987_nl <= MUX_s_1_2_2(and_142_cse, mux_146_cse, nor_291_cse);
  butterFly_7_butterFly_7_or_32_rmff <= MUX_s_1_2_2(mux_991_nl, mux_987_nl, fsm_output(4));
  mux_1043_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1344_cse);
  nor_310_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1042_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, nor_310_nl);
  mux_1044_nl <= MUX_s_1_2_2(mux_1043_nl, mux_1042_nl, fsm_output(3));
  and_1900_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1901_nl <= (nor_885_cse OR (fsm_output(7))) AND (fsm_output(6));
  mux_1039_nl <= MUX_s_1_2_2(and_1900_nl, and_1901_nl, fsm_output(0));
  mux_1040_nl <= MUX_s_1_2_2(mux_1039_nl, nor_tmp_35, fsm_output(3));
  mux_1045_nl <= MUX_s_1_2_2(mux_1044_nl, mux_1040_nl, fsm_output(5));
  mux_1046_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1045_nl, nor_44_cse);
  or_1334_nl <= (NOT (fsm_output(1))) OR (NOT (fsm_output(5))) OR (fsm_output(3))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1037_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1334_nl);
  mux_1034_nl <= MUX_s_1_2_2(or_324_cse, (fsm_output(7)), or_2999_cse);
  mux_1035_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1034_nl, and_2080_cse);
  mux_1036_nl <= MUX_s_1_2_2(mux_1035_nl, mux_295_cse, fsm_output(1));
  mux_1038_nl <= MUX_s_1_2_2(mux_1037_nl, mux_1036_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_34_rmff <= MUX_s_1_2_2(mux_1046_nl, mux_1038_nl, fsm_output(4));
  or_1390_nl <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1095_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1390_nl);
  and_1891_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1892_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1093_nl <= MUX_s_1_2_2(and_1891_nl, and_1892_nl, fsm_output(0));
  or_1387_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5));
  mux_1092_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1387_nl);
  mux_1094_nl <= MUX_s_1_2_2(mux_1093_nl, mux_1092_nl, fsm_output(3));
  mux_1096_nl <= MUX_s_1_2_2(mux_1095_nl, mux_1094_nl, fsm_output(1));
  mux_1097_nl <= MUX_s_1_2_2(mux_1096_nl, nor_tmp_35, fsm_output(2));
  or_1386_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1090_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1386_nl);
  or_1385_nl <= (NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1086_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1385_nl);
  mux_1087_nl <= MUX_s_1_2_2(mux_1086_nl, mux_3731_cse, fsm_output(0));
  mux_1088_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1087_nl, fsm_output(3));
  mux_1089_nl <= MUX_s_1_2_2(mux_1088_nl, mux_295_cse, fsm_output(1));
  mux_1091_nl <= MUX_s_1_2_2(mux_1090_nl, mux_1089_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_36_rmff <= MUX_s_1_2_2(mux_1097_nl, mux_1091_nl, fsm_output(4));
  mux_1150_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_1142, fsm_output(1));
  mux_1151_nl <= MUX_s_1_2_2(mux_1150_nl, nor_tmp_35, fsm_output(2));
  mux_1152_nl <= MUX_s_1_2_2(mux_1151_nl, mux_308_cse, fsm_output(4));
  mux_1143_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_1142, nor_44_cse);
  mux_1144_nl <= MUX_s_1_2_2(mux_1143_nl, mux_298_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_38_rmff <= MUX_s_1_2_2(mux_1152_nl, mux_1144_nl, or_2999_cse);
  nor_1887_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  nor_1890_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_1205_nl <= MUX_s_1_2_2(nor_2157_cse, nor_1890_nl, fsm_output(0));
  mux_1206_nl <= MUX_s_1_2_2(nor_2156_cse, mux_1205_nl, fsm_output(6));
  nor_361_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1207_nl <= MUX_s_1_2_2(nor_1887_nl, mux_1206_nl, nor_361_nl);
  mux_1208_nl <= MUX_s_1_2_2(mux_1207_nl, (fsm_output(6)), fsm_output(7));
  mux_1204_nl <= MUX_s_1_2_2(and_142_cse, mux_146_cse, nor_356_cse);
  butterFly_7_butterFly_7_or_40_rmff <= MUX_s_1_2_2(mux_1208_nl, mux_1204_nl, fsm_output(4));
  mux_1261_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_389_cse);
  nor_381_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1260_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, nor_381_nl);
  mux_1262_nl <= MUX_s_1_2_2(mux_1261_nl, mux_1260_nl, fsm_output(3));
  and_1856_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1857_nl <= (nor_951_cse OR (fsm_output(7))) AND (fsm_output(6));
  mux_1257_nl <= MUX_s_1_2_2(and_1856_nl, and_1857_nl, fsm_output(0));
  mux_1258_nl <= MUX_s_1_2_2(mux_1257_nl, nor_tmp_35, fsm_output(3));
  mux_1263_nl <= MUX_s_1_2_2(mux_1262_nl, mux_1258_nl, fsm_output(5));
  mux_1264_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1263_nl, nor_44_cse);
  and_1858_nl <= (fsm_output(1)) AND (fsm_output(5)) AND (NOT (fsm_output(3))) AND
      (fsm_output(0)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101"));
  mux_1255_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1858_nl);
  mux_1252_nl <= MUX_s_1_2_2((fsm_output(7)), or_324_cse, nor_947_cse);
  mux_1253_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1252_nl, and_2080_cse);
  mux_1254_nl <= MUX_s_1_2_2(mux_1253_nl, mux_295_cse, fsm_output(1));
  mux_1256_nl <= MUX_s_1_2_2(mux_1255_nl, mux_1254_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_42_rmff <= MUX_s_1_2_2(mux_1264_nl, mux_1256_nl, fsm_output(4));
  nor_401_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  mux_1313_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_401_nl);
  and_1845_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1846_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1311_nl <= MUX_s_1_2_2(and_1845_nl, and_1846_nl, fsm_output(0));
  or_1630_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5));
  mux_1310_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1630_nl);
  mux_1312_nl <= MUX_s_1_2_2(mux_1311_nl, mux_1310_nl, fsm_output(3));
  mux_1314_nl <= MUX_s_1_2_2(mux_1313_nl, mux_1312_nl, fsm_output(1));
  mux_1315_nl <= MUX_s_1_2_2(mux_1314_nl, nor_tmp_35, fsm_output(2));
  nor_396_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR
      (NOT (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101")));
  mux_1308_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_396_nl);
  and_1847_nl <= (fsm_output(5)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("101"));
  mux_1304_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, and_1847_nl);
  mux_1305_nl <= MUX_s_1_2_2(mux_1304_nl, mux_3731_cse, fsm_output(0));
  mux_1306_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1305_nl, fsm_output(3));
  mux_1307_nl <= MUX_s_1_2_2(mux_1306_nl, mux_295_cse, fsm_output(1));
  mux_1309_nl <= MUX_s_1_2_2(mux_1308_nl, mux_1307_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_44_rmff <= MUX_s_1_2_2(mux_1315_nl, mux_1309_nl, fsm_output(4));
  mux_1369_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_1363, nor_44_cse);
  mux_1370_nl <= MUX_s_1_2_2(mux_1369_nl, mux_298_cse, fsm_output(4));
  mux_1365_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_1363, fsm_output(1));
  mux_1366_nl <= MUX_s_1_2_2(mux_1365_nl, nor_tmp_35, fsm_output(2));
  mux_1367_nl <= MUX_s_1_2_2(mux_1366_nl, mux_308_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_46_rmff <= MUX_s_1_2_2(mux_1370_nl, mux_1367_nl, nor_947_cse);
  nor_1834_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  nor_1837_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_1423_nl <= MUX_s_1_2_2(nor_2157_cse, nor_1837_nl, fsm_output(0));
  mux_1424_nl <= MUX_s_1_2_2(nor_2156_cse, mux_1423_nl, fsm_output(6));
  nor_442_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1425_nl <= MUX_s_1_2_2(nor_1834_nl, mux_1424_nl, nor_442_nl);
  mux_1426_nl <= MUX_s_1_2_2(mux_1425_nl, (fsm_output(6)), fsm_output(7));
  mux_1422_nl <= MUX_s_1_2_2(and_142_cse, mux_146_cse, nor_437_cse);
  butterFly_7_butterFly_7_or_48_rmff <= MUX_s_1_2_2(mux_1426_nl, mux_1422_nl, fsm_output(4));
  mux_1478_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1818_cse);
  nor_460_nl <= NOT((NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1477_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, nor_460_nl);
  mux_1479_nl <= MUX_s_1_2_2(mux_1478_nl, mux_1477_nl, fsm_output(3));
  and_1805_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1806_nl <= (nor_1025_cse OR (fsm_output(7))) AND (fsm_output(6));
  mux_1474_nl <= MUX_s_1_2_2(and_1805_nl, and_1806_nl, fsm_output(0));
  mux_1475_nl <= MUX_s_1_2_2(mux_1474_nl, nor_tmp_35, fsm_output(3));
  mux_1480_nl <= MUX_s_1_2_2(mux_1479_nl, mux_1475_nl, fsm_output(5));
  mux_1481_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1480_nl, nor_44_cse);
  nand_399_nl <= NOT((fsm_output(1)) AND (fsm_output(5)) AND (NOT (fsm_output(3)))
      AND (fsm_output(0)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  mux_1472_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, nand_399_nl);
  mux_1469_nl <= MUX_s_1_2_2(or_324_cse, (fsm_output(7)), or_3418_cse);
  mux_1470_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1469_nl, and_2080_cse);
  mux_1471_nl <= MUX_s_1_2_2(mux_1470_nl, mux_295_cse, fsm_output(1));
  mux_1473_nl <= MUX_s_1_2_2(mux_1472_nl, mux_1471_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_50_rmff <= MUX_s_1_2_2(mux_1481_nl, mux_1473_nl, fsm_output(4));
  or_1864_nl <= (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_1530_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1864_nl);
  and_1793_nl <= ((NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1794_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(5))))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1528_nl <= MUX_s_1_2_2(and_1793_nl, and_1794_nl, fsm_output(0));
  or_1861_nl <= (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(5));
  mux_1527_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_1861_nl);
  mux_1529_nl <= MUX_s_1_2_2(mux_1528_nl, mux_1527_nl, fsm_output(3));
  mux_1531_nl <= MUX_s_1_2_2(mux_1530_nl, mux_1529_nl, fsm_output(1));
  mux_1532_nl <= MUX_s_1_2_2(mux_1531_nl, nor_tmp_35, fsm_output(2));
  or_1860_nl <= (NOT (fsm_output(1))) OR (fsm_output(3)) OR (fsm_output(0)) OR (NOT
      (fsm_output(5))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"));
  mux_1525_nl <= MUX_s_1_2_2((fsm_output(7)), nor_tmp_35, or_1860_nl);
  nand_390_nl <= NOT((fsm_output(5)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("110")));
  mux_1521_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_390_nl);
  mux_1522_nl <= MUX_s_1_2_2(mux_1521_nl, mux_3731_cse, fsm_output(0));
  mux_1523_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1522_nl, fsm_output(3));
  mux_1524_nl <= MUX_s_1_2_2(mux_1523_nl, mux_295_cse, fsm_output(1));
  mux_1526_nl <= MUX_s_1_2_2(mux_1525_nl, mux_1524_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_52_rmff <= MUX_s_1_2_2(mux_1532_nl, mux_1526_nl, fsm_output(4));
  mux_1585_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_1577, fsm_output(1));
  mux_1586_nl <= MUX_s_1_2_2(mux_1585_nl, nor_tmp_35, fsm_output(2));
  mux_1587_nl <= MUX_s_1_2_2(mux_1586_nl, mux_308_cse, fsm_output(4));
  mux_1578_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_1577, nor_44_cse);
  mux_1579_nl <= MUX_s_1_2_2(mux_1578_nl, mux_298_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_54_rmff <= MUX_s_1_2_2(mux_1587_nl, mux_1579_nl, or_3418_cse);
  nor_1783_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  nor_1786_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3)) OR (NOT (fsm_output(5))));
  mux_1640_nl <= MUX_s_1_2_2(nor_2157_cse, nor_1786_nl, fsm_output(0));
  mux_1641_nl <= MUX_s_1_2_2(nor_2156_cse, mux_1640_nl, fsm_output(6));
  nor_520_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4));
  mux_1642_nl <= MUX_s_1_2_2(nor_1783_nl, mux_1641_nl, nor_520_nl);
  mux_1643_nl <= MUX_s_1_2_2(mux_1642_nl, (fsm_output(6)), fsm_output(7));
  mux_1639_nl <= MUX_s_1_2_2(and_142_cse, mux_146_cse, and_1765_cse);
  butterFly_7_butterFly_7_or_56_rmff <= MUX_s_1_2_2(mux_1643_nl, mux_1639_nl, fsm_output(4));
  mux_1695_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1737_cse);
  and_1744_nl <= (fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1101"))
      AND S1_OUTER_LOOP_for_acc_svs_4;
  mux_1694_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, and_1744_nl);
  mux_1696_nl <= MUX_s_1_2_2(mux_1695_nl, mux_1694_nl, fsm_output(3));
  and_1745_nl <= ((CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1101"))
      AND S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(7))) AND (fsm_output(6));
  and_1747_nl <= (and_1366_cse OR (fsm_output(7))) AND (fsm_output(6));
  mux_1691_nl <= MUX_s_1_2_2(and_1745_nl, and_1747_nl, fsm_output(0));
  mux_1692_nl <= MUX_s_1_2_2(mux_1691_nl, nor_tmp_35, fsm_output(3));
  mux_1697_nl <= MUX_s_1_2_2(mux_1696_nl, mux_1692_nl, fsm_output(5));
  mux_1698_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1697_nl, nor_44_cse);
  and_1749_nl <= (fsm_output(1)) AND (fsm_output(5)) AND (NOT (fsm_output(3))) AND
      (fsm_output(0)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  mux_1689_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1749_nl);
  mux_1686_nl <= MUX_s_1_2_2((fsm_output(7)), or_324_cse, and_1369_cse);
  mux_1687_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1686_nl, and_2080_cse);
  mux_1688_nl <= MUX_s_1_2_2(mux_1687_nl, mux_295_cse, fsm_output(1));
  mux_1690_nl <= MUX_s_1_2_2(mux_1689_nl, mux_1688_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_58_rmff <= MUX_s_1_2_2(mux_1698_nl, mux_1690_nl, fsm_output(4));
  nor_574_nl <= NOT((fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(5)) OR
      CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("111")));
  mux_1747_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_574_nl);
  and_1724_nl <= ((CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1110"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(5))) OR (fsm_output(7))) AND
      (fsm_output(6));
  and_1726_nl <= ((CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1110"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (fsm_output(5))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_1745_nl <= MUX_s_1_2_2(and_1724_nl, and_1726_nl, fsm_output(0));
  nand_346_nl <= NOT((fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1110"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (NOT (fsm_output(5))));
  mux_1744_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, nand_346_nl);
  mux_1746_nl <= MUX_s_1_2_2(mux_1745_nl, mux_1744_nl, fsm_output(3));
  mux_1748_nl <= MUX_s_1_2_2(mux_1747_nl, mux_1746_nl, fsm_output(1));
  mux_1749_nl <= MUX_s_1_2_2(mux_1748_nl, nor_tmp_35, fsm_output(2));
  and_1728_nl <= (fsm_output(1)) AND (NOT (fsm_output(3))) AND (NOT (fsm_output(0)))
      AND (fsm_output(5)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  mux_1742_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1728_nl);
  and_1729_nl <= (fsm_output(5)) AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"));
  mux_1738_nl <= MUX_s_1_2_2(nor_tmp_35, mux_167_cse, and_1729_nl);
  mux_1739_nl <= MUX_s_1_2_2(mux_1738_nl, mux_3731_cse, fsm_output(0));
  mux_1740_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1739_nl, fsm_output(3));
  mux_1741_nl <= MUX_s_1_2_2(mux_1740_nl, mux_295_cse, fsm_output(1));
  mux_1743_nl <= MUX_s_1_2_2(mux_1742_nl, mux_1741_nl, fsm_output(2));
  butterFly_7_butterFly_7_or_60_rmff <= MUX_s_1_2_2(mux_1749_nl, mux_1743_nl, fsm_output(4));
  mux_1799_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_1793, nor_44_cse);
  mux_1800_nl <= MUX_s_1_2_2(mux_1799_nl, mux_298_cse, fsm_output(4));
  mux_1795_nl <= MUX_s_1_2_2(mux_309_cse, mux_tmp_1793, fsm_output(1));
  mux_1796_nl <= MUX_s_1_2_2(mux_1795_nl, nor_tmp_35, fsm_output(2));
  mux_1797_nl <= MUX_s_1_2_2(mux_1796_nl, mux_308_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_62_rmff <= MUX_s_1_2_2(mux_1800_nl, mux_1797_nl, and_1369_cse);
  and_1680_nl <= ((NOT((NOT (fsm_output(1))) OR (fsm_output(0)) OR (NOT (fsm_output(4)))))
      OR (fsm_output(7))) AND (fsm_output(6));
  nor_630_nl <= NOT((fsm_output(1)) OR (fsm_output(0)) OR (NOT (fsm_output(4))));
  mux_1856_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_630_nl);
  mux_1857_cse <= MUX_s_1_2_2(and_1680_nl, mux_1856_nl, fsm_output(3));
  or_2175_nl <= (fsm_output(1)) OR (NOT (fsm_output(0))) OR (fsm_output(4));
  mux_1854_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2175_nl);
  and_1683_nl <= or_3894_cse AND (fsm_output(4));
  mux_1846_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1683_nl);
  mux_1847_cse <= MUX_s_1_2_2(nor_tmp_35, mux_1846_nl, fsm_output(3));
  and_1681_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND (fsm_output(6));
  mux_1855_nl <= MUX_s_1_2_2(mux_1854_cse, and_1681_nl, fsm_output(3));
  mux_1858_nl <= MUX_s_1_2_2(mux_1857_cse, mux_1855_nl, fsm_output(5));
  and_1682_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND
      (fsm_output(6));
  mux_1859_nl <= MUX_s_1_2_2(mux_1858_nl, and_1682_nl, or_348_cse);
  or_2169_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4));
  mux_1850_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2169_nl);
  or_2168_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(4));
  mux_1849_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2168_nl);
  mux_1851_nl <= MUX_s_1_2_2(mux_1850_nl, mux_1849_nl, fsm_output(0));
  mux_1852_nl <= MUX_s_1_2_2(mux_1851_nl, nor_tmp_35, or_4797_cse);
  mux_1853_nl <= MUX_s_1_2_2(mux_1852_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_64_rmff <= MUX_s_1_2_2(mux_1859_nl, mux_1853_nl, fsm_output(2));
  or_2224_cse <= and_1674_cse OR (fsm_output(6));
  or_2231_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_2230_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_1908_nl <= MUX_s_1_2_2(or_2231_nl, or_2230_nl, fsm_output(0));
  or_2229_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_1909_nl <= MUX_s_1_2_2(mux_1908_nl, or_2229_nl, fsm_output(5));
  or_2228_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_1910_nl <= MUX_s_1_2_2(mux_1909_nl, or_2228_nl, fsm_output(3));
  nor_1722_nl <= NOT((fsm_output(1)) OR mux_1910_nl);
  nor_1723_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR nand_330_cse);
  mux_1911_nl <= MUX_s_1_2_2(nor_1722_nl, nor_1723_nl, fsm_output(4));
  or_2223_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_1904_nl <= MUX_s_1_2_2(or_2223_nl, or_3918_cse, fsm_output(5));
  mux_1905_nl <= MUX_s_1_2_2((fsm_output(6)), mux_1904_nl, fsm_output(3));
  mux_1906_nl <= MUX_s_1_2_2(or_2224_cse, mux_1905_nl, fsm_output(1));
  mux_1907_nl <= MUX_s_1_2_2((fsm_output(6)), mux_1906_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_65_rmff <= MUX_s_1_2_2(mux_1911_nl, mux_1907_nl, fsm_output(7));
  mux_1952_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1674_cse);
  mux_1951_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1665_cse);
  mux_1953_cse <= MUX_s_1_2_2(mux_1952_nl, mux_1951_nl, fsm_output(1));
  or_2281_nl <= (fsm_output(2)) OR (NOT (fsm_output(0))) OR (NOT (fsm_output(5)))
      OR (fsm_output(3));
  mux_1967_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2281_nl);
  and_1663_nl <= (nor_1711_cse OR (fsm_output(7))) AND (fsm_output(6));
  mux_1964_nl <= MUX_s_1_2_2(and_1663_nl, mux_295_cse, fsm_output(0));
  mux_1965_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1964_nl, fsm_output(2));
  nor_655_nl <= NOT((fsm_output(0)) OR (fsm_output(5)) OR (NOT (fsm_output(3))));
  mux_1962_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_655_nl);
  mux_1963_nl <= MUX_s_1_2_2(mux_1962_nl, mux_295_cse, fsm_output(2));
  mux_1966_cse <= MUX_s_1_2_2(mux_1965_nl, mux_1963_nl, fsm_output(1));
  mux_1968_nl <= MUX_s_1_2_2(mux_tmp_1958, mux_1967_cse, fsm_output(1));
  mux_1969_nl <= MUX_s_1_2_2(mux_1968_nl, mux_1966_cse, fsm_output(4));
  mux_1959_nl <= MUX_s_1_2_2(mux_tmp_1958, nor_tmp_35, fsm_output(1));
  mux_1960_nl <= MUX_s_1_2_2(mux_1959_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_66_rmff <= MUX_s_1_2_2(mux_1969_nl, mux_1960_nl, or_2242_cse);
  or_2327_nl <= (fsm_output(2)) OR (fsm_output(0)) OR (NOT (fsm_output(5))) OR (fsm_output(3));
  mux_2028_cse <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2327_nl);
  mux_2025_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_673_cse);
  mux_2026_nl <= MUX_s_1_2_2(mux_2025_nl, mux_296_cse, fsm_output(2));
  and_1652_nl <= ((NOT((NOT (fsm_output(0))) OR (fsm_output(5)) OR (fsm_output(3))))
      OR (fsm_output(7))) AND (fsm_output(6));
  mux_2023_nl <= MUX_s_1_2_2(and_1652_nl, mux_295_cse, fsm_output(2));
  mux_2027_cse <= MUX_s_1_2_2(mux_2026_nl, mux_2023_nl, fsm_output(1));
  mux_2029_nl <= MUX_s_1_2_2(mux_tmp_2019, mux_2028_cse, fsm_output(1));
  mux_2030_nl <= MUX_s_1_2_2(mux_2029_nl, mux_2027_cse, fsm_output(4));
  mux_2020_nl <= MUX_s_1_2_2(mux_tmp_2019, nor_tmp_35, fsm_output(1));
  mux_2021_nl <= MUX_s_1_2_2(mux_2020_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_67_rmff <= MUX_s_1_2_2(mux_2030_nl, mux_2021_nl, or_2242_cse);
  and_1641_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND (fsm_output(6));
  mux_2085_nl <= MUX_s_1_2_2(mux_1854_cse, and_1641_nl, fsm_output(3));
  mux_2088_nl <= MUX_s_1_2_2(mux_1857_cse, mux_2085_nl, fsm_output(5));
  and_1642_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND
      (fsm_output(6));
  mux_2089_nl <= MUX_s_1_2_2(mux_2088_nl, and_1642_nl, or_582_cse);
  or_2373_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4));
  mux_2080_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2373_nl);
  or_2372_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(4));
  mux_2079_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2372_nl);
  mux_2081_nl <= MUX_s_1_2_2(mux_2080_nl, mux_2079_nl, fsm_output(0));
  mux_2082_nl <= MUX_s_1_2_2(mux_2081_nl, nor_tmp_35, or_4797_cse);
  mux_2083_nl <= MUX_s_1_2_2(mux_2082_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_68_rmff <= MUX_s_1_2_2(mux_2089_nl, mux_2083_nl, fsm_output(2));
  or_2433_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_2432_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2135_nl <= MUX_s_1_2_2(or_2433_nl, or_2432_nl, fsm_output(0));
  or_2431_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2136_nl <= MUX_s_1_2_2(mux_2135_nl, or_2431_nl, fsm_output(5));
  or_2430_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_2137_nl <= MUX_s_1_2_2(mux_2136_nl, or_2430_nl, fsm_output(3));
  nor_1680_nl <= NOT((fsm_output(1)) OR mux_2137_nl);
  nor_1681_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("00")) OR nand_327_cse);
  mux_2138_nl <= MUX_s_1_2_2(nor_1680_nl, nor_1681_nl, fsm_output(4));
  or_2425_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_2131_nl <= MUX_s_1_2_2(or_2425_nl, or_3918_cse, fsm_output(5));
  mux_2132_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2131_nl, fsm_output(3));
  mux_2133_nl <= MUX_s_1_2_2(or_2224_cse, mux_2132_nl, fsm_output(1));
  mux_2134_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2133_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_69_rmff <= MUX_s_1_2_2(mux_2138_nl, mux_2134_nl, fsm_output(7));
  mux_2193_nl <= MUX_s_1_2_2(mux_tmp_2187, nor_tmp_35, fsm_output(1));
  mux_2194_nl <= MUX_s_1_2_2(mux_2193_nl, mux_1953_cse, fsm_output(4));
  mux_2188_nl <= MUX_s_1_2_2(mux_tmp_2187, mux_1967_cse, fsm_output(1));
  mux_2189_nl <= MUX_s_1_2_2(mux_2188_nl, mux_1966_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_70_rmff <= MUX_s_1_2_2(mux_2194_nl, mux_2189_nl, nor_701_cse);
  mux_2251_nl <= MUX_s_1_2_2(mux_tmp_2245, nor_tmp_35, fsm_output(1));
  mux_2252_nl <= MUX_s_1_2_2(mux_2251_nl, mux_1953_cse, fsm_output(4));
  mux_2246_nl <= MUX_s_1_2_2(mux_tmp_2245, mux_2028_cse, fsm_output(1));
  mux_2247_nl <= MUX_s_1_2_2(mux_2246_nl, mux_2027_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_71_rmff <= MUX_s_1_2_2(mux_2252_nl, mux_2247_nl, nor_701_cse);
  and_1600_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND (fsm_output(6));
  mux_2305_nl <= MUX_s_1_2_2(mux_1854_cse, and_1600_nl, fsm_output(3));
  mux_2308_nl <= MUX_s_1_2_2(mux_1857_cse, mux_2305_nl, fsm_output(5));
  and_1601_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND
      (fsm_output(6));
  mux_2309_nl <= MUX_s_1_2_2(mux_2308_nl, and_1601_nl, or_823_cse);
  or_2563_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4));
  mux_2300_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2563_nl);
  or_2562_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(4));
  mux_2299_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2562_nl);
  mux_2301_nl <= MUX_s_1_2_2(mux_2300_nl, mux_2299_nl, fsm_output(0));
  mux_2302_nl <= MUX_s_1_2_2(mux_2301_nl, nor_tmp_35, or_4797_cse);
  mux_2303_nl <= MUX_s_1_2_2(mux_2302_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_72_rmff <= MUX_s_1_2_2(mux_2309_nl, mux_2303_nl, fsm_output(2));
  or_2614_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_2613_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2355_nl <= MUX_s_1_2_2(or_2614_nl, or_2613_nl, fsm_output(0));
  or_2612_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2356_nl <= MUX_s_1_2_2(mux_2355_nl, or_2612_nl, fsm_output(5));
  or_2611_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_2357_nl <= MUX_s_1_2_2(mux_2356_nl, or_2611_nl, fsm_output(3));
  nor_1647_nl <= NOT((fsm_output(1)) OR mux_2357_nl);
  nor_1648_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))
      OR nand_330_cse);
  mux_2358_nl <= MUX_s_1_2_2(nor_1647_nl, nor_1648_nl, fsm_output(4));
  or_2606_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_2351_nl <= MUX_s_1_2_2(or_2606_nl, or_3918_cse, fsm_output(5));
  mux_2352_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2351_nl, fsm_output(3));
  mux_2353_nl <= MUX_s_1_2_2(or_2224_cse, mux_2352_nl, fsm_output(1));
  mux_2354_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2353_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_73_rmff <= MUX_s_1_2_2(mux_2358_nl, mux_2354_nl, fsm_output(7));
  mux_2413_nl <= MUX_s_1_2_2(mux_tmp_2403, mux_1967_cse, fsm_output(1));
  mux_2414_nl <= MUX_s_1_2_2(mux_2413_nl, mux_1966_cse, fsm_output(4));
  mux_2404_nl <= MUX_s_1_2_2(mux_tmp_2403, nor_tmp_35, fsm_output(1));
  mux_2405_nl <= MUX_s_1_2_2(mux_2404_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_74_rmff <= MUX_s_1_2_2(mux_2414_nl, mux_2405_nl, or_2619_cse);
  mux_2471_nl <= MUX_s_1_2_2(mux_tmp_2461, mux_2028_cse, fsm_output(1));
  mux_2472_nl <= MUX_s_1_2_2(mux_2471_nl, mux_2027_cse, fsm_output(4));
  mux_2462_nl <= MUX_s_1_2_2(mux_tmp_2461, nor_tmp_35, fsm_output(1));
  mux_2463_nl <= MUX_s_1_2_2(mux_2462_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_75_rmff <= MUX_s_1_2_2(mux_2472_nl, mux_2463_nl, or_2619_cse);
  and_1559_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100")) OR
      S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND (fsm_output(6));
  mux_2525_nl <= MUX_s_1_2_2(mux_1854_cse, and_1559_nl, fsm_output(3));
  mux_2528_nl <= MUX_s_1_2_2(mux_1857_cse, mux_2525_nl, fsm_output(5));
  and_1560_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4)))) OR (fsm_output(7))) AND
      (fsm_output(6));
  mux_2529_nl <= MUX_s_1_2_2(mux_2528_nl, and_1560_nl, or_1039_cse);
  or_2734_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(4));
  mux_2520_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2734_nl);
  or_2733_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(4));
  mux_2519_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2733_nl);
  mux_2521_nl <= MUX_s_1_2_2(mux_2520_nl, mux_2519_nl, fsm_output(0));
  mux_2522_nl <= MUX_s_1_2_2(mux_2521_nl, nor_tmp_35, or_4797_cse);
  mux_2523_nl <= MUX_s_1_2_2(mux_2522_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_76_rmff <= MUX_s_1_2_2(mux_2529_nl, mux_2523_nl, fsm_output(2));
  or_2793_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_2792_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2575_nl <= MUX_s_1_2_2(or_2793_nl, or_2792_nl, fsm_output(0));
  or_2791_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2576_nl <= MUX_s_1_2_2(mux_2575_nl, or_2791_nl, fsm_output(5));
  or_2790_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1101"))
      OR S1_OUTER_LOOP_for_acc_svs_4 OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_2577_nl <= MUX_s_1_2_2(mux_2576_nl, or_2790_nl, fsm_output(3));
  nor_1614_nl <= NOT((fsm_output(1)) OR mux_2577_nl);
  nor_1615_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      OR (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(6)))));
  mux_2578_nl <= MUX_s_1_2_2(nor_1614_nl, nor_1615_nl, fsm_output(4));
  or_2785_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_2571_nl <= MUX_s_1_2_2(or_2785_nl, or_3918_cse, fsm_output(5));
  mux_2572_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2571_nl, fsm_output(3));
  mux_2573_nl <= MUX_s_1_2_2(or_2224_cse, mux_2572_nl, fsm_output(1));
  mux_2574_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2573_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_77_rmff <= MUX_s_1_2_2(mux_2578_nl, mux_2574_nl, fsm_output(7));
  mux_2633_nl <= MUX_s_1_2_2(mux_tmp_2627, nor_tmp_35, fsm_output(1));
  mux_2634_nl <= MUX_s_1_2_2(mux_2633_nl, mux_1953_cse, fsm_output(4));
  mux_2628_nl <= MUX_s_1_2_2(mux_tmp_2627, mux_1967_cse, fsm_output(1));
  mux_2629_nl <= MUX_s_1_2_2(mux_2628_nl, mux_1966_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_78_rmff <= MUX_s_1_2_2(mux_2634_nl, mux_2629_nl, nor_817_cse);
  mux_2691_nl <= MUX_s_1_2_2(mux_tmp_2685, nor_tmp_35, fsm_output(1));
  mux_2692_nl <= MUX_s_1_2_2(mux_2691_nl, mux_1953_cse, fsm_output(4));
  mux_2686_nl <= MUX_s_1_2_2(mux_tmp_2685, mux_2028_cse, fsm_output(1));
  mux_2687_nl <= MUX_s_1_2_2(mux_2686_nl, mux_2027_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_79_rmff <= MUX_s_1_2_2(mux_2692_nl, mux_2687_nl, nor_817_cse);
  and_1512_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1514_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2745_nl <= MUX_s_1_2_2(mux_1854_cse, and_1514_nl, fsm_output(3));
  mux_2748_nl <= MUX_s_1_2_2(mux_1857_cse, mux_2745_nl, fsm_output(5));
  mux_2749_nl <= MUX_s_1_2_2(and_1512_nl, mux_2748_nl, nor_291_cse);
  or_2934_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4));
  mux_2740_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2934_nl);
  or_2933_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(4));
  mux_2739_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_2933_nl);
  mux_2741_nl <= MUX_s_1_2_2(mux_2740_nl, mux_2739_nl, fsm_output(0));
  mux_2742_nl <= MUX_s_1_2_2(mux_2741_nl, nor_tmp_35, or_4797_cse);
  mux_2743_nl <= MUX_s_1_2_2(mux_2742_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_80_rmff <= MUX_s_1_2_2(mux_2749_nl, mux_2743_nl, fsm_output(2));
  or_2991_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_2990_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2795_nl <= MUX_s_1_2_2(or_2991_nl, or_2990_nl, fsm_output(0));
  or_2989_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_2796_nl <= MUX_s_1_2_2(mux_2795_nl, or_2989_nl, fsm_output(5));
  or_2988_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_2797_nl <= MUX_s_1_2_2(mux_2796_nl, or_2988_nl, fsm_output(3));
  nor_1584_nl <= NOT((fsm_output(1)) OR mux_2797_nl);
  nor_1585_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR nand_330_cse);
  mux_2798_nl <= MUX_s_1_2_2(nor_1584_nl, nor_1585_nl, fsm_output(4));
  or_2983_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_2791_nl <= MUX_s_1_2_2(or_2983_nl, or_3918_cse, fsm_output(5));
  mux_2792_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2791_nl, fsm_output(3));
  mux_2793_nl <= MUX_s_1_2_2(or_2224_cse, mux_2792_nl, fsm_output(1));
  mux_2794_nl <= MUX_s_1_2_2((fsm_output(6)), mux_2793_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_81_rmff <= MUX_s_1_2_2(mux_2798_nl, mux_2794_nl, fsm_output(7));
  mux_2853_nl <= MUX_s_1_2_2(mux_tmp_2843, mux_1967_cse, fsm_output(1));
  mux_2854_nl <= MUX_s_1_2_2(mux_2853_nl, mux_1966_cse, fsm_output(4));
  mux_2844_nl <= MUX_s_1_2_2(mux_tmp_2843, nor_tmp_35, fsm_output(1));
  mux_2845_nl <= MUX_s_1_2_2(mux_2844_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_82_rmff <= MUX_s_1_2_2(mux_2854_nl, mux_2845_nl, or_2999_cse);
  mux_2911_nl <= MUX_s_1_2_2(mux_tmp_2901, mux_2028_cse, fsm_output(1));
  mux_2912_nl <= MUX_s_1_2_2(mux_2911_nl, mux_2027_cse, fsm_output(4));
  mux_2902_nl <= MUX_s_1_2_2(mux_tmp_2901, nor_tmp_35, fsm_output(1));
  mux_2903_nl <= MUX_s_1_2_2(mux_2902_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_83_rmff <= MUX_s_1_2_2(mux_2912_nl, mux_2903_nl, or_2999_cse);
  and_1472_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1474_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_2965_nl <= MUX_s_1_2_2(mux_1854_cse, and_1474_nl, fsm_output(3));
  mux_2968_nl <= MUX_s_1_2_2(mux_1857_cse, mux_2965_nl, fsm_output(5));
  mux_2969_nl <= MUX_s_1_2_2(and_1472_nl, mux_2968_nl, nor_356_cse);
  or_3135_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4));
  mux_2960_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3135_nl);
  or_3134_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(4));
  mux_2959_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3134_nl);
  mux_2961_nl <= MUX_s_1_2_2(mux_2960_nl, mux_2959_nl, fsm_output(0));
  mux_2962_nl <= MUX_s_1_2_2(mux_2961_nl, nor_tmp_35, or_4797_cse);
  mux_2963_nl <= MUX_s_1_2_2(mux_2962_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_84_rmff <= MUX_s_1_2_2(mux_2969_nl, mux_2963_nl, fsm_output(2));
  or_3200_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_3199_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_3015_nl <= MUX_s_1_2_2(or_3200_nl, or_3199_nl, fsm_output(0));
  or_3198_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_3016_nl <= MUX_s_1_2_2(mux_3015_nl, or_3198_nl, fsm_output(5));
  or_3197_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_3017_nl <= MUX_s_1_2_2(mux_3016_nl, or_3197_nl, fsm_output(3));
  nor_1550_nl <= NOT((fsm_output(1)) OR mux_3017_nl);
  nor_1551_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("10")) OR nand_327_cse);
  mux_3018_nl <= MUX_s_1_2_2(nor_1550_nl, nor_1551_nl, fsm_output(4));
  or_3192_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_3011_nl <= MUX_s_1_2_2(or_3192_nl, or_3918_cse, fsm_output(5));
  mux_3012_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3011_nl, fsm_output(3));
  mux_3013_nl <= MUX_s_1_2_2(or_2224_cse, mux_3012_nl, fsm_output(1));
  mux_3014_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3013_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_85_rmff <= MUX_s_1_2_2(mux_3018_nl, mux_3014_nl, fsm_output(7));
  mux_3073_nl <= MUX_s_1_2_2(mux_tmp_3067, nor_tmp_35, fsm_output(1));
  mux_3074_nl <= MUX_s_1_2_2(mux_3073_nl, mux_1953_cse, fsm_output(4));
  mux_3068_nl <= MUX_s_1_2_2(mux_tmp_3067, mux_1967_cse, fsm_output(1));
  mux_3069_nl <= MUX_s_1_2_2(mux_3068_nl, mux_1966_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_86_rmff <= MUX_s_1_2_2(mux_3074_nl, mux_3069_nl, nor_947_cse);
  mux_3131_nl <= MUX_s_1_2_2(mux_tmp_3125, nor_tmp_35, fsm_output(1));
  mux_3132_nl <= MUX_s_1_2_2(mux_3131_nl, mux_1953_cse, fsm_output(4));
  mux_3126_nl <= MUX_s_1_2_2(mux_tmp_3125, mux_2028_cse, fsm_output(1));
  mux_3127_nl <= MUX_s_1_2_2(mux_3126_nl, mux_2027_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_87_rmff <= MUX_s_1_2_2(mux_3132_nl, mux_3127_nl, nor_947_cse);
  and_1428_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1430_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3185_nl <= MUX_s_1_2_2(mux_1854_cse, and_1430_nl, fsm_output(3));
  mux_3188_nl <= MUX_s_1_2_2(mux_1857_cse, mux_3185_nl, fsm_output(5));
  mux_3189_nl <= MUX_s_1_2_2(and_1428_nl, mux_3188_nl, nor_437_cse);
  or_3354_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4));
  mux_3180_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3354_nl);
  or_3353_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1000"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(4));
  mux_3179_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3353_nl);
  mux_3181_nl <= MUX_s_1_2_2(mux_3180_nl, mux_3179_nl, fsm_output(0));
  mux_3182_nl <= MUX_s_1_2_2(mux_3181_nl, nor_tmp_35, or_4797_cse);
  mux_3183_nl <= MUX_s_1_2_2(mux_3182_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_88_rmff <= MUX_s_1_2_2(mux_3189_nl, mux_3183_nl, fsm_output(2));
  or_3410_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  or_3409_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_3235_nl <= MUX_s_1_2_2(or_3410_nl, or_3409_nl, fsm_output(0));
  or_3408_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_3236_nl <= MUX_s_1_2_2(mux_3235_nl, or_3408_nl, fsm_output(5));
  or_3407_nl <= (NOT (fsm_output(5))) OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(2)) OR (NOT (fsm_output(6)));
  mux_3237_nl <= MUX_s_1_2_2(mux_3236_nl, or_3407_nl, fsm_output(3));
  nor_1516_nl <= NOT((fsm_output(1)) OR mux_3237_nl);
  nor_1517_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))
      OR nand_330_cse);
  mux_3238_nl <= MUX_s_1_2_2(nor_1516_nl, nor_1517_nl, fsm_output(4));
  or_3402_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))
      OR (NOT (fsm_output(0))) OR (fsm_output(2)))) OR (fsm_output(6));
  mux_3231_nl <= MUX_s_1_2_2(or_3402_nl, or_3918_cse, fsm_output(5));
  mux_3232_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3231_nl, fsm_output(3));
  mux_3233_nl <= MUX_s_1_2_2(or_2224_cse, mux_3232_nl, fsm_output(1));
  mux_3234_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3233_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_89_rmff <= MUX_s_1_2_2(mux_3238_nl, mux_3234_nl, fsm_output(7));
  mux_3293_nl <= MUX_s_1_2_2(mux_tmp_3283, mux_1967_cse, fsm_output(1));
  mux_3294_nl <= MUX_s_1_2_2(mux_3293_nl, mux_1966_cse, fsm_output(4));
  mux_3284_nl <= MUX_s_1_2_2(mux_tmp_3283, nor_tmp_35, fsm_output(1));
  mux_3285_nl <= MUX_s_1_2_2(mux_3284_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_90_rmff <= MUX_s_1_2_2(mux_3294_nl, mux_3285_nl, or_3418_cse);
  mux_3351_nl <= MUX_s_1_2_2(mux_tmp_3341, mux_2028_cse, fsm_output(1));
  mux_3352_nl <= MUX_s_1_2_2(mux_3351_nl, mux_2027_cse, fsm_output(4));
  mux_3342_nl <= MUX_s_1_2_2(mux_tmp_3341, nor_tmp_35, fsm_output(1));
  mux_3343_nl <= MUX_s_1_2_2(mux_3342_nl, mux_1953_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_91_rmff <= MUX_s_1_2_2(mux_3352_nl, mux_3343_nl, or_3418_cse);
  and_1382_nl <= ((NOT((NOT (fsm_output(5))) OR (NOT (fsm_output(3))) OR (fsm_output(1))
      OR (NOT (fsm_output(0))) OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  and_1384_nl <= ((NOT(CONV_SL_1_1(fsm_output(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100")) OR
      (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4)))) OR (fsm_output(7)))
      AND (fsm_output(6));
  mux_3405_nl <= MUX_s_1_2_2(mux_1854_cse, and_1384_nl, fsm_output(3));
  mux_3408_nl <= MUX_s_1_2_2(mux_1857_cse, mux_3405_nl, fsm_output(5));
  mux_3409_nl <= MUX_s_1_2_2(and_1382_nl, mux_3408_nl, and_1765_cse);
  or_3551_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT S1_OUTER_LOOP_for_acc_svs_4) OR (fsm_output(4));
  mux_3400_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3551_nl);
  or_3550_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1100"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(4));
  mux_3399_nl <= MUX_s_1_2_2(mux_167_cse, nor_tmp_35, or_3550_nl);
  mux_3401_nl <= MUX_s_1_2_2(mux_3400_nl, mux_3399_nl, fsm_output(0));
  mux_3402_nl <= MUX_s_1_2_2(mux_3401_nl, nor_tmp_35, or_4797_cse);
  mux_3403_nl <= MUX_s_1_2_2(mux_3402_nl, mux_1847_cse, fsm_output(5));
  butterFly_7_butterFly_7_or_92_rmff <= MUX_s_1_2_2(mux_3409_nl, mux_3403_nl, fsm_output(2));
  nand_271_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1101"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (fsm_output(2)) AND (NOT (fsm_output(6))));
  nand_272_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1101"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (fsm_output(2)) AND (NOT (fsm_output(6))));
  mux_3455_nl <= MUX_s_1_2_2(nand_271_nl, nand_272_nl, fsm_output(0));
  or_3608_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("111"))
      OR (fsm_output(0)) OR (NOT (fsm_output(2))) OR (fsm_output(6));
  mux_3456_nl <= MUX_s_1_2_2(mux_3455_nl, or_3608_nl, fsm_output(5));
  nand_273_nl <= NOT((fsm_output(5)) AND (fsm_output(0)) AND CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0=STD_LOGIC_VECTOR'("1101"))
      AND S1_OUTER_LOOP_for_acc_svs_4 AND (NOT (fsm_output(2))) AND (fsm_output(6)));
  mux_3457_nl <= MUX_s_1_2_2(mux_3456_nl, nand_273_nl, fsm_output(3));
  nor_1483_nl <= NOT((fsm_output(1)) OR mux_3457_nl);
  nor_1484_nl <= NOT((fsm_output(1)) OR (fsm_output(3)) OR (fsm_output(5)) OR (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(6)))));
  mux_3458_nl <= MUX_s_1_2_2(nor_1483_nl, nor_1484_nl, fsm_output(4));
  or_3602_nl <= (CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"))
      AND (fsm_output(0)) AND (NOT (fsm_output(2)))) OR (fsm_output(6));
  mux_3451_nl <= MUX_s_1_2_2(or_3602_nl, or_3918_cse, fsm_output(5));
  mux_3452_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3451_nl, fsm_output(3));
  mux_3453_nl <= MUX_s_1_2_2(or_2224_cse, mux_3452_nl, fsm_output(1));
  mux_3454_nl <= MUX_s_1_2_2((fsm_output(6)), mux_3453_nl, fsm_output(4));
  butterFly_7_butterFly_7_or_93_rmff <= MUX_s_1_2_2(mux_3458_nl, mux_3454_nl, fsm_output(7));
  mux_3513_nl <= MUX_s_1_2_2(mux_tmp_3507, nor_tmp_35, fsm_output(1));
  mux_3514_nl <= MUX_s_1_2_2(mux_3513_nl, mux_1953_cse, fsm_output(4));
  mux_3508_nl <= MUX_s_1_2_2(mux_tmp_3507, mux_1967_cse, fsm_output(1));
  mux_3509_nl <= MUX_s_1_2_2(mux_3508_nl, mux_1966_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_94_rmff <= MUX_s_1_2_2(mux_3514_nl, mux_3509_nl, and_1369_cse);
  mux_3571_nl <= MUX_s_1_2_2(mux_tmp_3565, nor_tmp_35, fsm_output(1));
  mux_3572_nl <= MUX_s_1_2_2(mux_3571_nl, mux_1953_cse, fsm_output(4));
  mux_3566_nl <= MUX_s_1_2_2(mux_tmp_3565, mux_2028_cse, fsm_output(1));
  mux_3567_nl <= MUX_s_1_2_2(mux_3566_nl, mux_2027_cse, fsm_output(4));
  butterFly_7_butterFly_7_or_95_rmff <= MUX_s_1_2_2(mux_3572_nl, mux_3567_nl, and_1369_cse);
  and_151_seb <= (NOT mux_156_itm) AND and_dcpl_137 AND and_dcpl_135;
  nor_2156_cse <= NOT((NOT (fsm_output(0))) OR (fsm_output(2)) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(3))) OR (fsm_output(5)));
  nor_2157_cse <= NOT((fsm_output(2)) OR (NOT (fsm_output(1))) OR (fsm_output(3))
      OR (NOT (fsm_output(5))));
  or_348_cse <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("000"));
  and_179_seb <= not_tmp_169 AND and_dcpl_164;
  and_2080_cse <= (fsm_output(5)) AND (fsm_output(3)) AND (fsm_output(0));
  nor_44_cse <= NOT(CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01")));
  and_201_seb <= not_tmp_188 AND and_dcpl_164;
  and_217_seb <= not_tmp_209 AND and_dcpl_42 AND and_dcpl_151;
  and_230_seb <= (NOT mux_156_itm) AND and_dcpl_203 AND and_dcpl_135;
  or_582_cse <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("001"));
  and_243_seb <= not_tmp_169 AND and_dcpl_216;
  and_257_seb <= not_tmp_188 AND and_dcpl_216;
  and_267_seb <= not_tmp_209 AND butterFly_3_f1_asn_17 AND and_dcpl_151;
  and_281_seb <= (NOT mux_156_itm) AND and_dcpl_242 AND and_dcpl_135;
  or_823_cse <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("010"));
  and_295_seb <= not_tmp_169 AND and_dcpl_255;
  and_311_seb <= not_tmp_188 AND and_dcpl_255;
  and_322_seb <= not_tmp_209 AND and_dcpl_257 AND and_dcpl_151;
  and_333_seb <= (NOT mux_156_itm) AND and_dcpl_281 AND and_dcpl_135;
  or_1039_cse <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("011"));
  and_344_seb <= not_tmp_169 AND and_dcpl_291;
  and_358_seb <= not_tmp_188 AND and_dcpl_291;
  and_368_seb <= not_tmp_209 AND and_dcpl_293 AND and_dcpl_151;
  and_381_seb <= (NOT mux_156_itm) AND and_dcpl_137 AND and_dcpl_316;
  nor_291_cse <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("100")));
  and_393_seb <= not_tmp_169 AND and_dcpl_328;
  and_406_seb <= not_tmp_188 AND and_dcpl_328;
  and_415_seb <= not_tmp_209 AND and_dcpl_330 AND and_dcpl_151;
  and_427_seb <= (NOT mux_156_itm) AND and_dcpl_203 AND and_dcpl_316;
  nor_356_cse <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("101")));
  and_438_seb <= not_tmp_169 AND and_dcpl_363;
  and_451_seb <= not_tmp_188 AND and_dcpl_363;
  and_460_seb <= not_tmp_209 AND and_dcpl_365 AND and_dcpl_151;
  and_470_seb <= (NOT mux_156_itm) AND and_dcpl_242 AND and_dcpl_316;
  nor_437_cse <= NOT(CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg/=STD_LOGIC_VECTOR'("110")));
  and_481_seb <= not_tmp_169 AND and_dcpl_396;
  and_494_seb <= not_tmp_188 AND and_dcpl_396;
  and_503_seb <= not_tmp_209 AND and_dcpl_398 AND and_dcpl_151;
  and_513_seb <= (NOT mux_156_itm) AND and_dcpl_281 AND and_dcpl_316;
  and_1765_cse <= CONV_SL_1_1(reg_drf_revArr_ptr_1_smx_9_0_1_reg=STD_LOGIC_VECTOR'("111"));
  and_523_seb <= not_tmp_169 AND and_dcpl_428;
  and_536_seb <= not_tmp_188 AND and_dcpl_428;
  and_546_seb <= not_tmp_209 AND and_dcpl_430 AND and_dcpl_151;
  and_587_seb <= not_tmp_843 AND and_dcpl_484 AND and_dcpl_483;
  and_618_seb <= not_tmp_865 AND and_dcpl_42;
  and_1674_cse <= (fsm_output(3)) AND (fsm_output(5)) AND (fsm_output(0)) AND (fsm_output(2));
  nand_330_cse <= NOT((fsm_output(0)) AND (fsm_output(2)) AND (fsm_output(6)));
  and_644_seb <= not_tmp_874 AND and_dcpl_42;
  and_1665_cse <= (fsm_output(2)) AND (fsm_output(5)) AND (fsm_output(3));
  nor_1711_cse <= NOT((fsm_output(5)) OR (fsm_output(3)));
  and_662_seb <= not_tmp_890 AND S6_OUTER_LOOP_for_nor_22_cse AND and_dcpl_559;
  nor_673_cse <= NOT((NOT (fsm_output(0))) OR (fsm_output(5)) OR (NOT (fsm_output(3))));
  and_677_seb <= not_tmp_843 AND and_dcpl_574 AND and_dcpl_483;
  and_693_seb <= not_tmp_865 AND butterFly_3_f1_asn_17;
  nand_327_cse <= NOT((reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (fsm_output(0)) AND
      (fsm_output(2)) AND (fsm_output(6)));
  and_705_seb <= not_tmp_874 AND butterFly_3_f1_asn_17;
  and_716_seb <= not_tmp_890 AND S6_OUTER_LOOP_for_nor_22_cse AND and_dcpl_613;
  and_729_seb <= not_tmp_843 AND and_dcpl_626 AND and_dcpl_483;
  and_745_seb <= not_tmp_865 AND and_dcpl_257;
  and_760_seb <= not_tmp_874 AND and_dcpl_257;
  and_773_seb <= not_tmp_890 AND and_dcpl_254 AND and_dcpl_559;
  and_786_seb <= not_tmp_843 AND and_dcpl_683 AND and_dcpl_483;
  and_797_seb <= not_tmp_865 AND and_dcpl_293;
  and_808_seb <= not_tmp_874 AND and_dcpl_293;
  and_818_seb <= not_tmp_890 AND and_dcpl_254 AND and_dcpl_613;
  and_831_seb <= not_tmp_843 AND and_dcpl_484 AND and_dcpl_728;
  and_847_seb <= not_tmp_865 AND and_dcpl_330;
  and_863_seb <= not_tmp_874 AND and_dcpl_330;
  and_876_seb <= not_tmp_890 AND and_dcpl_327 AND and_dcpl_559;
  and_888_seb <= not_tmp_843 AND and_dcpl_574 AND and_dcpl_728;
  and_900_seb <= not_tmp_865 AND and_dcpl_365;
  and_911_seb <= not_tmp_874 AND and_dcpl_365;
  and_921_seb <= not_tmp_890 AND and_dcpl_327 AND and_dcpl_613;
  and_933_seb <= not_tmp_843 AND and_dcpl_626 AND and_dcpl_728;
  and_948_seb <= not_tmp_865 AND and_dcpl_398;
  and_963_seb <= not_tmp_874 AND and_dcpl_398;
  and_976_seb <= not_tmp_890 AND and_dcpl_395 AND and_dcpl_559;
  and_988_seb <= not_tmp_843 AND and_dcpl_683 AND and_dcpl_728;
  and_1000_seb <= not_tmp_865 AND and_dcpl_430;
  and_1011_seb <= not_tmp_874 AND and_dcpl_430;
  and_1022_seb <= not_tmp_890 AND and_dcpl_395 AND and_dcpl_613;
  twiddle_rsci_adrb_d <= twiddle_rsci_adrb_d_reg;
  twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d_reg;
  twiddle_h_rsci_adrb_d <= twiddle_h_rsci_adrb_d_reg;
  twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d <= twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d_reg;
  butterFly_7_or_360_cse <= and_dcpl_100 OR and_dcpl_116;
  butterFly_7_butterFly_7_mux_31_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_125);
  butterFly_7_or_168_nl <= (butterFly_7_butterFly_7_mux_31_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2274_nl <= NOT(and_dcpl_125 OR butterFly_7_or_360_cse);
  mux1h_62_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2274_nl & and_dcpl_125 & butterFly_7_or_360_cse));
  butterFly_7_mux_93_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_125);
  butterFly_7_butterFly_7_or_191_nl <= (butterFly_7_mux_93_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_169_nl <= and_116_ssc OR and_dcpl_125;
  butterFly_7_mux1h_230_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_169_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_72_nl <= (butterFly_7_mux1h_230_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_63_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_201_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_264_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_201_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_202_nl <= (butterFly_7_mux1h_264_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_0_0_i_adra_d <= butterFly_7_or_168_nl & mux1h_62_nl & butterFly_7_butterFly_7_or_191_nl
      & butterFly_7_or_72_nl & mux1h_63_nl & butterFly_7_or_202_nl;
  butterFly_7_or_38_nl <= ((NOT reg_modulo_add_7_slc_32_svs_st_cse) AND and_dcpl_129)
      OR ((NOT reg_modulo_add_7_slc_32_svs_st_cse) AND and_dcpl_131);
  butterFly_7_or_39_nl <= (reg_modulo_add_7_slc_32_svs_st_cse AND and_dcpl_129) OR
      (reg_modulo_add_7_slc_32_svs_st_cse AND and_dcpl_131);
  butterFly_7_mux1h_1_nl <= MUX1HOT_v_32_3_2(modulo_sub_7_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, STD_LOGIC_VECTOR'( and_dcpl_102 & butterFly_7_or_38_nl
      & butterFly_7_or_39_nl));
  butterFly_7_and_149_nl <= (NOT reg_modulo_add_7_slc_32_svs_st_cse) AND and_dcpl_102;
  butterFly_7_and_150_nl <= reg_modulo_add_7_slc_32_svs_st_cse AND and_dcpl_102;
  butterFly_7_mux1h_167_nl <= MUX1HOT_v_32_7_2(reg_tmp_54_lpi_3_dfm_cse, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, reg_mult_2_res_lpi_4_dfm_cse, reg_mult_1_res_lpi_4_dfm_cse,
      modulo_sub_15_qr_lpi_4_dfm, modulo_sub_23_qr_lpi_3_dfm, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_and_149_nl & butterFly_7_and_150_nl & and_dcpl_127
      & and_dcpl_109 & and_dcpl_129 & and_dcpl_131));
  xx_rsc_0_0_i_da_d_pff <= butterFly_7_mux1h_1_nl & butterFly_7_mux1h_167_nl;
  xx_rsc_0_0_i_wea_d <= STD_LOGIC_VECTOR'( and_151_seb & butterFly_7_butterFly_7_or_rmff);
  butterFly_7_butterFly_7_or_1_nl <= and_dcpl_125 OR (not_tmp_149 AND and_dcpl_142
      AND and_dcpl_140);
  or_373_nl <= (fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("000"));
  mux_172_nl <= MUX_s_1_2_2(mux_171_cse, nor_tmp_35, or_373_nl);
  mux_164_nl <= MUX_s_1_2_2(nor_tmp_36, mux_163_cse, fsm_output(4));
  or_370_nl <= nor_2152_cse OR (fsm_output(3));
  mux_158_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_370_nl);
  mux_159_nl <= MUX_s_1_2_2(nor_tmp_35, mux_158_nl, fsm_output(1));
  mux_160_nl <= MUX_s_1_2_2(mux_159_nl, mux_213_cse, fsm_output(0));
  mux_161_nl <= MUX_s_1_2_2(nor_tmp_36, mux_160_nl, fsm_output(4));
  or_368_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_165_nl <= MUX_s_1_2_2(mux_164_nl, mux_161_nl, or_368_nl);
  mux_166_nl <= MUX_s_1_2_2(nor_tmp_35, mux_165_nl, fsm_output(5));
  mux_173_nl <= MUX_s_1_2_2(mux_172_nl, mux_166_nl, fsm_output(2));
  butterFly_7_and_311_nl <= (NOT(or_dcpl_180 AND and_dcpl_125)) AND mux_173_nl;
  xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_1_nl
      & butterFly_7_and_311_nl);
  xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_151_seb
      & butterFly_7_butterFly_7_or_rmff);
  butterFly_7_butterFly_7_mux_30_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_157);
  butterFly_7_or_165_nl <= (butterFly_7_butterFly_7_mux_30_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2275_nl <= NOT(and_dcpl_157 OR butterFly_7_or_360_cse);
  mux1h_60_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2275_nl & and_dcpl_157 & butterFly_7_or_360_cse));
  butterFly_7_mux_92_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_157);
  butterFly_7_butterFly_7_or_190_nl <= (butterFly_7_mux_92_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_170_nl <= and_164_ssc OR and_dcpl_157;
  butterFly_7_mux1h_228_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_170_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_71_nl <= (butterFly_7_mux1h_228_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_61_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_204_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_265_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_204_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_205_nl <= (butterFly_7_mux1h_265_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_1_0_i_adra_d <= butterFly_7_or_165_nl & mux1h_60_nl & butterFly_7_butterFly_7_or_190_nl
      & butterFly_7_or_71_nl & mux1h_61_nl & butterFly_7_or_205_nl;
  butterFly_7_or_36_nl <= ((NOT reg_modulo_add_2_slc_32_svs_st_cse) AND and_173_ssc)
      OR ((NOT reg_modulo_add_3_slc_32_svs_st_cse) AND and_174_ssc);
  butterFly_7_or_37_nl <= (reg_modulo_add_2_slc_32_svs_st_cse AND and_173_ssc) OR
      (reg_modulo_add_3_slc_32_svs_st_cse AND and_174_ssc);
  butterFly_7_mux1h_5_nl <= MUX1HOT_v_32_3_2(modulo_sub_4_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, STD_LOGIC_VECTOR'( and_dcpl_149 & butterFly_7_or_36_nl
      & butterFly_7_or_37_nl));
  butterFly_7_and_143_nl <= (NOT reg_modulo_add_5_slc_32_svs_st_cse) AND and_dcpl_149;
  butterFly_7_and_144_nl <= reg_modulo_add_5_slc_32_svs_st_cse AND and_dcpl_149;
  butterFly_7_mux1h_166_nl <= MUX1HOT_v_32_7_2(reg_tmp_54_lpi_3_dfm_cse, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, reg_mult_2_res_lpi_4_dfm_cse, reg_mult_1_res_lpi_4_dfm_cse,
      modulo_sub_12_qr_lpi_4_dfm, modulo_sub_20_qr_lpi_3_dfm, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_and_143_nl & butterFly_7_and_144_nl & and_dcpl_127
      & and_dcpl_109 & and_173_ssc & and_174_ssc));
  xx_rsc_1_0_i_da_d_pff <= butterFly_7_mux1h_5_nl & butterFly_7_mux1h_166_nl;
  xx_rsc_1_0_i_wea_d <= STD_LOGIC_VECTOR'( and_179_seb & butterFly_7_butterFly_7_or_2_rmff);
  butterFly_7_butterFly_7_or_3_nl <= and_dcpl_157 OR and_dcpl_168;
  and_2075_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_49_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00001"))
      OR (NOT (fsm_output(1))));
  mux_215_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_49_nl);
  or_432_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))))
      OR (fsm_output(3));
  mux_216_nl <= MUX_s_1_2_2(mux_215_nl, mux_162_cse, or_432_nl);
  mux_217_nl <= MUX_s_1_2_2(mux_216_nl, mux_213_cse, fsm_output(0));
  mux_218_nl <= MUX_s_1_2_2(and_2075_nl, mux_217_nl, fsm_output(4));
  mux_219_nl <= MUX_s_1_2_2(nor_tmp_35, mux_218_nl, fsm_output(5));
  mux_227_nl <= MUX_s_1_2_2(mux_226_cse, mux_219_nl, fsm_output(2));
  butterFly_7_and_312_nl <= (NOT(or_dcpl_182 AND and_dcpl_157)) AND mux_227_nl;
  xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_3_nl
      & butterFly_7_and_312_nl);
  xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_179_seb
      & butterFly_7_butterFly_7_or_2_rmff);
  butterFly_7_butterFly_7_mux_29_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_177);
  butterFly_7_or_162_nl <= (butterFly_7_butterFly_7_mux_29_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2276_nl <= NOT(and_dcpl_177 OR butterFly_7_or_360_cse);
  mux1h_58_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2276_nl & and_dcpl_177 & butterFly_7_or_360_cse));
  butterFly_7_mux_91_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_177);
  butterFly_7_butterFly_7_or_189_nl <= (butterFly_7_mux_91_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_171_nl <= and_191_ssc OR and_dcpl_177;
  butterFly_7_mux1h_226_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_171_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_70_nl <= (butterFly_7_mux1h_226_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_59_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_207_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_266_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_207_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_208_nl <= (butterFly_7_mux1h_266_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_2_0_i_adra_d <= butterFly_7_or_162_nl & mux1h_58_nl & butterFly_7_butterFly_7_or_189_nl
      & butterFly_7_or_70_nl & mux1h_59_nl & butterFly_7_or_208_nl;
  butterFly_7_or_34_nl <= ((NOT modulo_add_13_slc_32_svs_st) AND and_dcpl_179) OR
      ((NOT reg_modulo_add_11_slc_32_svs_st_cse) AND and_dcpl_180);
  butterFly_7_or_35_nl <= (modulo_add_13_slc_32_svs_st AND and_dcpl_179) OR (reg_modulo_add_11_slc_32_svs_st_cse
      AND and_dcpl_180);
  butterFly_7_mux1h_9_nl <= MUX1HOT_v_32_3_2(modulo_sub_5_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, STD_LOGIC_VECTOR'( and_dcpl_171 & butterFly_7_or_34_nl
      & butterFly_7_or_35_nl));
  butterFly_7_and_137_nl <= (NOT reg_modulo_add_5_slc_32_svs_st_cse) AND and_dcpl_171;
  butterFly_7_and_138_nl <= reg_modulo_add_5_slc_32_svs_st_cse AND and_dcpl_171;
  butterFly_7_mux1h_165_nl <= MUX1HOT_v_32_7_2(reg_tmp_54_lpi_3_dfm_cse, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, reg_mult_2_res_lpi_4_dfm_cse, reg_mult_1_res_lpi_4_dfm_cse,
      modulo_sub_13_qr_lpi_4_dfm, modulo_sub_21_qr_lpi_3_dfm, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_and_137_nl & butterFly_7_and_138_nl & and_dcpl_127
      & and_dcpl_109 & and_dcpl_179 & and_dcpl_180));
  xx_rsc_2_0_i_da_d_pff <= butterFly_7_mux1h_9_nl & butterFly_7_mux1h_165_nl;
  xx_rsc_2_0_i_wea_d <= STD_LOGIC_VECTOR'( and_201_seb & butterFly_7_butterFly_7_or_4_rmff);
  butterFly_7_butterFly_7_or_5_nl <= and_dcpl_177 OR and_dcpl_168;
  and_2066_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_62_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00010"))
      OR (NOT (fsm_output(1))));
  mux_266_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_62_nl);
  or_489_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))))
      OR (fsm_output(3));
  mux_267_nl <= MUX_s_1_2_2(mux_266_nl, mux_162_cse, or_489_nl);
  mux_268_nl <= MUX_s_1_2_2(mux_267_nl, mux_213_cse, fsm_output(0));
  mux_269_nl <= MUX_s_1_2_2(and_2066_nl, mux_268_nl, fsm_output(4));
  mux_270_nl <= MUX_s_1_2_2(nor_tmp_35, mux_269_nl, fsm_output(5));
  mux_278_nl <= MUX_s_1_2_2(mux_226_cse, mux_270_nl, fsm_output(2));
  butterFly_7_and_313_nl <= (NOT(or_dcpl_184 AND and_dcpl_177)) AND mux_278_nl;
  xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_5_nl
      & butterFly_7_and_313_nl);
  xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_201_seb
      & butterFly_7_butterFly_7_or_4_rmff);
  butterFly_7_butterFly_7_mux_28_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_190);
  butterFly_7_or_159_nl <= (butterFly_7_butterFly_7_mux_28_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2277_nl <= NOT(and_dcpl_190 OR butterFly_7_or_360_cse);
  mux1h_56_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2277_nl & and_dcpl_190 & butterFly_7_or_360_cse));
  butterFly_7_mux_90_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_190);
  butterFly_7_butterFly_7_or_188_nl <= (butterFly_7_mux_90_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_172_nl <= and_207_ssc OR and_dcpl_190;
  butterFly_7_mux1h_224_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_172_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_69_nl <= (butterFly_7_mux1h_224_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_57_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_210_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_267_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_210_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_211_nl <= (butterFly_7_mux1h_267_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_3_0_i_adra_d <= butterFly_7_or_159_nl & mux1h_56_nl & butterFly_7_butterFly_7_or_188_nl
      & butterFly_7_or_69_nl & mux1h_57_nl & butterFly_7_or_211_nl;
  butterFly_7_or_32_nl <= ((NOT reg_modulo_add_6_slc_32_svs_st_cse) AND and_dcpl_191)
      OR ((NOT reg_modulo_add_1_slc_32_svs_st_cse) AND and_dcpl_192);
  butterFly_7_or_33_nl <= (reg_modulo_add_6_slc_32_svs_st_cse AND and_dcpl_191) OR
      (reg_modulo_add_1_slc_32_svs_st_cse AND and_dcpl_192);
  butterFly_7_mux1h_13_nl <= MUX1HOT_v_32_3_2(modulo_sub_6_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, STD_LOGIC_VECTOR'( and_dcpl_184 & butterFly_7_or_32_nl
      & butterFly_7_or_33_nl));
  butterFly_7_and_131_nl <= (NOT reg_modulo_add_6_slc_32_svs_st_cse) AND and_dcpl_184;
  butterFly_7_and_132_nl <= reg_modulo_add_6_slc_32_svs_st_cse AND and_dcpl_184;
  butterFly_7_mux1h_164_nl <= MUX1HOT_v_32_7_2(reg_tmp_54_lpi_3_dfm_cse, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, reg_mult_2_res_lpi_4_dfm_cse, reg_mult_1_res_lpi_4_dfm_cse,
      modulo_sub_14_qr_lpi_4_dfm, reg_modulo_sub_18_qr_lpi_4_dfm_cse, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_and_131_nl & butterFly_7_and_132_nl & and_dcpl_127
      & and_dcpl_109 & and_dcpl_191 & and_dcpl_192));
  xx_rsc_3_0_i_da_d_pff <= butterFly_7_mux1h_13_nl & butterFly_7_mux1h_164_nl;
  xx_rsc_3_0_i_wea_d <= STD_LOGIC_VECTOR'( and_217_seb & butterFly_7_butterFly_7_or_6_rmff);
  butterFly_7_butterFly_7_or_7_nl <= and_dcpl_190 OR and_dcpl_168;
  and_2052_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_82_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00011"))
      OR (NOT (fsm_output(1))));
  mux_320_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_82_nl);
  or_537_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))))
      OR (fsm_output(3));
  mux_321_nl <= MUX_s_1_2_2(mux_320_nl, mux_162_cse, or_537_nl);
  mux_322_nl <= MUX_s_1_2_2(mux_321_nl, mux_213_cse, fsm_output(0));
  mux_323_nl <= MUX_s_1_2_2(and_2052_nl, mux_322_nl, fsm_output(4));
  mux_324_nl <= MUX_s_1_2_2(nor_tmp_35, mux_323_nl, fsm_output(5));
  mux_332_nl <= MUX_s_1_2_2(mux_226_cse, mux_324_nl, fsm_output(2));
  butterFly_7_and_314_nl <= (NOT(or_dcpl_185 AND and_dcpl_190)) AND mux_332_nl;
  xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_7_nl
      & butterFly_7_and_314_nl);
  xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_217_seb
      & butterFly_7_butterFly_7_or_6_rmff);
  butterFly_7_butterFly_7_mux_27_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_201);
  butterFly_7_or_156_nl <= (butterFly_7_butterFly_7_mux_27_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2278_nl <= NOT(and_dcpl_201 OR butterFly_7_or_360_cse);
  mux1h_54_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2278_nl & and_dcpl_201 & butterFly_7_or_360_cse));
  butterFly_7_mux_89_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_201);
  butterFly_7_butterFly_7_or_187_nl <= (butterFly_7_mux_89_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_173_nl <= and_221_ssc OR and_dcpl_201;
  butterFly_7_mux1h_222_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_173_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_68_nl <= (butterFly_7_mux1h_222_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_55_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_213_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_268_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_213_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_214_nl <= (butterFly_7_mux1h_268_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_4_0_i_adra_d <= butterFly_7_or_156_nl & mux1h_54_nl & butterFly_7_butterFly_7_or_187_nl
      & butterFly_7_or_68_nl & mux1h_55_nl & butterFly_7_or_214_nl;
  xx_rsc_4_0_i_wea_d <= STD_LOGIC_VECTOR'( and_230_seb & butterFly_7_butterFly_7_or_8_rmff);
  butterFly_7_butterFly_7_or_9_nl <= and_dcpl_201 OR (not_tmp_149 AND and_dcpl_207
      AND and_dcpl_140);
  nor_97_nl <= NOT((fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("001")));
  mux_387_nl <= MUX_s_1_2_2(nor_tmp_35, mux_171_cse, nor_97_nl);
  mux_379_nl <= MUX_s_1_2_2(nor_tmp_96, mux_163_cse, fsm_output(4));
  or_605_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00100"))))
      OR (fsm_output(3));
  mux_373_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_605_nl);
  mux_374_nl <= MUX_s_1_2_2(nor_tmp_35, mux_373_nl, fsm_output(1));
  mux_375_nl <= MUX_s_1_2_2(mux_374_nl, mux_213_cse, fsm_output(0));
  mux_376_nl <= MUX_s_1_2_2(nor_tmp_96, mux_375_nl, fsm_output(4));
  or_603_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_380_nl <= MUX_s_1_2_2(mux_379_nl, mux_376_nl, or_603_nl);
  mux_381_nl <= MUX_s_1_2_2(nor_tmp_35, mux_380_nl, fsm_output(5));
  mux_388_nl <= MUX_s_1_2_2(mux_387_nl, mux_381_nl, fsm_output(2));
  butterFly_7_and_315_nl <= (NOT(or_dcpl_188 AND and_dcpl_201)) AND mux_388_nl;
  xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_9_nl
      & butterFly_7_and_315_nl);
  xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_230_seb
      & butterFly_7_butterFly_7_or_8_rmff);
  butterFly_7_butterFly_7_mux_26_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_213);
  butterFly_7_or_153_nl <= (butterFly_7_butterFly_7_mux_26_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2279_nl <= NOT(and_dcpl_213 OR butterFly_7_or_360_cse);
  mux1h_52_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2279_nl & and_dcpl_213 & butterFly_7_or_360_cse));
  butterFly_7_mux_88_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_213);
  butterFly_7_butterFly_7_or_186_nl <= (butterFly_7_mux_88_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_174_nl <= and_237_ssc OR and_dcpl_213;
  butterFly_7_mux1h_220_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_174_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_67_nl <= (butterFly_7_mux1h_220_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_53_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_216_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_269_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_216_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_217_nl <= (butterFly_7_mux1h_269_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_5_0_i_adra_d <= butterFly_7_or_153_nl & mux1h_52_nl & butterFly_7_butterFly_7_or_186_nl
      & butterFly_7_or_67_nl & mux1h_53_nl & butterFly_7_or_217_nl;
  xx_rsc_5_0_i_wea_d <= STD_LOGIC_VECTOR'( and_243_seb & butterFly_7_butterFly_7_or_10_rmff);
  butterFly_7_butterFly_7_or_11_nl <= and_dcpl_213 OR and_dcpl_220;
  and_2033_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_113_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00101"))
      OR (NOT (fsm_output(1))));
  mux_429_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_113_nl);
  or_670_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))))
      OR (fsm_output(3));
  mux_430_nl <= MUX_s_1_2_2(mux_429_nl, mux_162_cse, or_670_nl);
  mux_431_nl <= MUX_s_1_2_2(mux_430_nl, mux_213_cse, fsm_output(0));
  mux_432_nl <= MUX_s_1_2_2(and_2033_nl, mux_431_nl, fsm_output(4));
  mux_433_nl <= MUX_s_1_2_2(nor_tmp_35, mux_432_nl, fsm_output(5));
  mux_441_nl <= MUX_s_1_2_2(mux_440_cse, mux_433_nl, fsm_output(2));
  butterFly_7_and_316_nl <= (NOT(or_dcpl_189 AND and_dcpl_213)) AND mux_441_nl;
  xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_11_nl
      & butterFly_7_and_316_nl);
  xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_243_seb
      & butterFly_7_butterFly_7_or_10_rmff);
  butterFly_7_butterFly_7_mux_25_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_224);
  butterFly_7_or_150_nl <= (butterFly_7_butterFly_7_mux_25_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2280_nl <= NOT(and_dcpl_224 OR butterFly_7_or_360_cse);
  mux1h_50_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2280_nl & and_dcpl_224 & butterFly_7_or_360_cse));
  butterFly_7_mux_87_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_224);
  butterFly_7_butterFly_7_or_185_nl <= (butterFly_7_mux_87_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_175_nl <= and_253_ssc OR and_dcpl_224;
  butterFly_7_mux1h_218_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_175_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_66_nl <= (butterFly_7_mux1h_218_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_51_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_219_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_270_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_219_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_220_nl <= (butterFly_7_mux1h_270_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_6_0_i_adra_d <= butterFly_7_or_150_nl & mux1h_50_nl & butterFly_7_butterFly_7_or_185_nl
      & butterFly_7_or_66_nl & mux1h_51_nl & butterFly_7_or_220_nl;
  xx_rsc_6_0_i_wea_d <= STD_LOGIC_VECTOR'( and_257_seb & butterFly_7_butterFly_7_or_12_rmff);
  butterFly_7_butterFly_7_or_13_nl <= and_dcpl_224 OR and_dcpl_220;
  mux_486_nl <= MUX_s_1_2_2(nor_tmp_35, mux_223_cse, nor_132_cse);
  mux_487_nl <= MUX_s_1_2_2(mux_486_nl, mux_435_cse, fsm_output(4));
  mux_488_nl <= MUX_s_1_2_2(mux_487_nl, nor_tmp_35, fsm_output(5));
  and_2024_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_129_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00110"))
      OR (NOT (fsm_output(1))));
  mux_477_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_129_nl);
  or_724_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))))
      OR (fsm_output(3));
  mux_478_nl <= MUX_s_1_2_2(mux_477_nl, mux_162_cse, or_724_nl);
  mux_479_nl <= MUX_s_1_2_2(mux_478_nl, mux_213_cse, fsm_output(0));
  mux_480_nl <= MUX_s_1_2_2(and_2024_nl, mux_479_nl, fsm_output(4));
  mux_481_nl <= MUX_s_1_2_2(nor_tmp_35, mux_480_nl, fsm_output(5));
  mux_489_nl <= MUX_s_1_2_2(mux_488_nl, mux_481_nl, fsm_output(2));
  butterFly_7_and_317_nl <= (NOT(or_dcpl_191 AND and_dcpl_224)) AND mux_489_nl;
  xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_13_nl
      & butterFly_7_and_317_nl);
  xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_257_seb
      & butterFly_7_butterFly_7_or_12_rmff);
  butterFly_7_butterFly_7_mux_24_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_230);
  butterFly_7_or_147_nl <= (butterFly_7_butterFly_7_mux_24_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2281_nl <= NOT(and_dcpl_230 OR butterFly_7_or_360_cse);
  mux1h_48_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2281_nl & and_dcpl_230 & butterFly_7_or_360_cse));
  butterFly_7_mux_86_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_230);
  butterFly_7_butterFly_7_or_184_nl <= (butterFly_7_mux_86_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_176_nl <= and_262_ssc OR and_dcpl_230;
  butterFly_7_mux1h_216_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_176_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_65_nl <= (butterFly_7_mux1h_216_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_49_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_222_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_271_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_222_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_223_nl <= (butterFly_7_mux1h_271_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_7_0_i_adra_d <= butterFly_7_or_147_nl & mux1h_48_nl & butterFly_7_butterFly_7_or_184_nl
      & butterFly_7_or_65_nl & mux1h_49_nl & butterFly_7_or_223_nl;
  xx_rsc_7_0_i_wea_d <= STD_LOGIC_VECTOR'( and_267_seb & butterFly_7_butterFly_7_or_14_rmff);
  butterFly_7_butterFly_7_or_15_nl <= and_dcpl_230 OR and_dcpl_220;
  and_2010_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0111"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_152_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("00111"))
      OR (NOT (fsm_output(1))));
  mux_529_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_152_nl);
  or_777_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("111"))))
      OR (fsm_output(3));
  mux_530_nl <= MUX_s_1_2_2(mux_529_nl, mux_162_cse, or_777_nl);
  mux_531_nl <= MUX_s_1_2_2(mux_530_nl, mux_213_cse, fsm_output(0));
  mux_532_nl <= MUX_s_1_2_2(and_2010_nl, mux_531_nl, fsm_output(4));
  mux_533_nl <= MUX_s_1_2_2(nor_tmp_35, mux_532_nl, fsm_output(5));
  mux_541_nl <= MUX_s_1_2_2(mux_440_cse, mux_533_nl, fsm_output(2));
  butterFly_7_and_318_nl <= (NOT(or_dcpl_192 AND and_dcpl_230)) AND mux_541_nl;
  xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_15_nl
      & butterFly_7_and_318_nl);
  xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_267_seb
      & butterFly_7_butterFly_7_or_14_rmff);
  butterFly_7_butterFly_7_mux_23_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_239);
  butterFly_7_or_144_nl <= (butterFly_7_butterFly_7_mux_23_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2282_nl <= NOT(and_dcpl_239 OR butterFly_7_or_360_cse);
  mux1h_46_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2282_nl & and_dcpl_239 & butterFly_7_or_360_cse));
  butterFly_7_mux_85_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_239);
  butterFly_7_butterFly_7_or_183_nl <= (butterFly_7_mux_85_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_177_nl <= and_271_ssc OR and_dcpl_239;
  butterFly_7_mux1h_214_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_177_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_64_nl <= (butterFly_7_mux1h_214_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_47_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_225_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_272_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_225_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_226_nl <= (butterFly_7_mux1h_272_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_8_0_i_adra_d <= butterFly_7_or_144_nl & mux1h_46_nl & butterFly_7_butterFly_7_or_183_nl
      & butterFly_7_or_64_nl & mux1h_47_nl & butterFly_7_or_226_nl;
  xx_rsc_8_0_i_wea_d <= STD_LOGIC_VECTOR'( and_281_seb & butterFly_7_butterFly_7_or_16_rmff);
  butterFly_7_butterFly_7_or_17_nl <= and_dcpl_239 OR (not_tmp_149 AND and_dcpl_142
      AND and_dcpl_245);
  or_846_nl <= (fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("010"));
  mux_596_nl <= MUX_s_1_2_2(mux_171_cse, nor_tmp_35, or_846_nl);
  mux_588_nl <= MUX_s_1_2_2(nor_tmp_165, mux_163_cse, fsm_output(4));
  or_843_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01000"))))
      OR (fsm_output(3));
  mux_582_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_843_nl);
  mux_583_nl <= MUX_s_1_2_2(nor_tmp_35, mux_582_nl, fsm_output(1));
  mux_584_nl <= MUX_s_1_2_2(mux_583_nl, mux_213_cse, fsm_output(0));
  mux_585_nl <= MUX_s_1_2_2(nor_tmp_165, mux_584_nl, fsm_output(4));
  or_841_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_589_nl <= MUX_s_1_2_2(mux_588_nl, mux_585_nl, or_841_nl);
  mux_590_nl <= MUX_s_1_2_2(nor_tmp_35, mux_589_nl, fsm_output(5));
  mux_597_nl <= MUX_s_1_2_2(mux_596_nl, mux_590_nl, fsm_output(2));
  butterFly_7_and_319_nl <= (NOT(or_dcpl_194 AND and_dcpl_239)) AND mux_597_nl;
  xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_17_nl
      & butterFly_7_and_319_nl);
  xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_281_seb
      & butterFly_7_butterFly_7_or_16_rmff);
  butterFly_7_butterFly_7_mux_22_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_252);
  butterFly_7_or_141_nl <= (butterFly_7_butterFly_7_mux_22_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2283_nl <= NOT(and_dcpl_252 OR butterFly_7_or_360_cse);
  mux1h_44_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2283_nl & and_dcpl_252 & butterFly_7_or_360_cse));
  butterFly_7_mux_84_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_252);
  butterFly_7_butterFly_7_or_182_nl <= (butterFly_7_mux_84_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_178_nl <= and_288_ssc OR and_dcpl_252;
  butterFly_7_mux1h_212_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_178_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_63_nl <= (butterFly_7_mux1h_212_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_45_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_228_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_273_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_228_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_229_nl <= (butterFly_7_mux1h_273_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_9_0_i_adra_d <= butterFly_7_or_141_nl & mux1h_44_nl & butterFly_7_butterFly_7_or_182_nl
      & butterFly_7_or_63_nl & mux1h_45_nl & butterFly_7_or_229_nl;
  xx_rsc_9_0_i_wea_d <= STD_LOGIC_VECTOR'( and_295_seb & butterFly_7_butterFly_7_or_18_rmff);
  butterFly_7_butterFly_7_or_19_nl <= and_dcpl_252 OR and_dcpl_259;
  and_1991_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_177_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01001"))
      OR (NOT (fsm_output(1))));
  mux_635_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_177_nl);
  or_895_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))))
      OR (fsm_output(3));
  mux_636_nl <= MUX_s_1_2_2(mux_635_nl, mux_162_cse, or_895_nl);
  mux_637_nl <= MUX_s_1_2_2(mux_636_nl, mux_213_cse, fsm_output(0));
  mux_638_nl <= MUX_s_1_2_2(and_1991_nl, mux_637_nl, fsm_output(4));
  mux_639_nl <= MUX_s_1_2_2(nor_tmp_35, mux_638_nl, fsm_output(5));
  mux_647_nl <= MUX_s_1_2_2(mux_646_cse, mux_639_nl, fsm_output(2));
  butterFly_7_and_320_nl <= (NOT(or_dcpl_196 AND and_dcpl_252)) AND mux_647_nl;
  xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_19_nl
      & butterFly_7_and_320_nl);
  xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_295_seb
      & butterFly_7_butterFly_7_or_18_rmff);
  butterFly_7_butterFly_7_mux_21_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_265);
  butterFly_7_or_138_nl <= (butterFly_7_butterFly_7_mux_21_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2284_nl <= NOT(and_dcpl_265 OR butterFly_7_or_360_cse);
  mux1h_42_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2284_nl & and_dcpl_265 & butterFly_7_or_360_cse));
  butterFly_7_mux_83_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_265);
  butterFly_7_butterFly_7_or_181_nl <= (butterFly_7_mux_83_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_179_nl <= and_305_ssc OR and_dcpl_265;
  butterFly_7_mux1h_210_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_179_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_62_nl <= (butterFly_7_mux1h_210_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_43_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_231_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_274_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_231_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_232_nl <= (butterFly_7_mux1h_274_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_10_0_i_adra_d <= butterFly_7_or_138_nl & mux1h_42_nl & butterFly_7_butterFly_7_or_181_nl
      & butterFly_7_or_62_nl & mux1h_43_nl & butterFly_7_or_232_nl;
  xx_rsc_10_0_i_wea_d <= STD_LOGIC_VECTOR'( and_311_seb & butterFly_7_butterFly_7_or_20_rmff);
  butterFly_7_butterFly_7_or_21_nl <= and_dcpl_265 OR and_dcpl_259;
  and_1982_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_190_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01010"))
      OR (NOT (fsm_output(1))));
  mux_683_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_190_nl);
  or_944_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))))
      OR (fsm_output(3));
  mux_684_nl <= MUX_s_1_2_2(mux_683_nl, mux_162_cse, or_944_nl);
  mux_685_nl <= MUX_s_1_2_2(mux_684_nl, mux_213_cse, fsm_output(0));
  mux_686_nl <= MUX_s_1_2_2(and_1982_nl, mux_685_nl, fsm_output(4));
  mux_687_nl <= MUX_s_1_2_2(nor_tmp_35, mux_686_nl, fsm_output(5));
  mux_695_nl <= MUX_s_1_2_2(mux_646_cse, mux_687_nl, fsm_output(2));
  butterFly_7_and_321_nl <= (NOT(or_dcpl_197 AND and_dcpl_265)) AND mux_695_nl;
  xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_21_nl
      & butterFly_7_and_321_nl);
  xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_311_seb
      & butterFly_7_butterFly_7_or_20_rmff);
  butterFly_7_butterFly_7_mux_20_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_272);
  butterFly_7_or_135_nl <= (butterFly_7_butterFly_7_mux_20_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2285_nl <= NOT(and_dcpl_272 OR butterFly_7_or_360_cse);
  mux1h_40_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2285_nl & and_dcpl_272 & butterFly_7_or_360_cse));
  butterFly_7_mux_82_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_272);
  butterFly_7_butterFly_7_or_180_nl <= (butterFly_7_mux_82_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_180_nl <= and_316_ssc OR and_dcpl_272;
  butterFly_7_mux1h_208_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_180_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_61_nl <= (butterFly_7_mux1h_208_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_41_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_234_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_275_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_234_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_235_nl <= (butterFly_7_mux1h_275_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_11_0_i_adra_d <= butterFly_7_or_135_nl & mux1h_40_nl & butterFly_7_butterFly_7_or_180_nl
      & butterFly_7_or_61_nl & mux1h_41_nl & butterFly_7_or_235_nl;
  xx_rsc_11_0_i_wea_d <= STD_LOGIC_VECTOR'( and_322_seb & butterFly_7_butterFly_7_or_22_rmff);
  butterFly_7_butterFly_7_or_23_nl <= and_dcpl_272 OR and_dcpl_259;
  nor_213_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010")));
  mux_744_nl <= MUX_s_1_2_2(nor_tmp_35, mux_223_cse, nor_213_nl);
  mux_745_nl <= MUX_s_1_2_2(mux_744_nl, mux_641_cse, fsm_output(4));
  mux_746_nl <= MUX_s_1_2_2(mux_745_nl, nor_tmp_35, fsm_output(5));
  and_1968_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1011"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_210_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01011"))
      OR (NOT (fsm_output(1))));
  mux_735_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_210_nl);
  or_995_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))))
      OR (fsm_output(3));
  mux_736_nl <= MUX_s_1_2_2(mux_735_nl, mux_162_cse, or_995_nl);
  mux_737_nl <= MUX_s_1_2_2(mux_736_nl, mux_213_cse, fsm_output(0));
  mux_738_nl <= MUX_s_1_2_2(and_1968_nl, mux_737_nl, fsm_output(4));
  mux_739_nl <= MUX_s_1_2_2(nor_tmp_35, mux_738_nl, fsm_output(5));
  mux_747_nl <= MUX_s_1_2_2(mux_746_nl, mux_739_nl, fsm_output(2));
  butterFly_7_and_322_nl <= (NOT(or_dcpl_198 AND and_dcpl_272)) AND mux_747_nl;
  xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_23_nl
      & butterFly_7_and_322_nl);
  xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_322_seb
      & butterFly_7_butterFly_7_or_22_rmff);
  butterFly_7_butterFly_7_mux_19_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_279);
  butterFly_7_or_132_nl <= (butterFly_7_butterFly_7_mux_19_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2286_nl <= NOT(and_dcpl_279 OR butterFly_7_or_360_cse);
  mux1h_38_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2286_nl & and_dcpl_279 & butterFly_7_or_360_cse));
  butterFly_7_mux_81_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_279);
  butterFly_7_butterFly_7_or_179_nl <= (butterFly_7_mux_81_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_181_nl <= and_326_ssc OR and_dcpl_279;
  butterFly_7_mux1h_206_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_181_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_60_nl <= (butterFly_7_mux1h_206_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_39_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_237_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_276_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_237_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_238_nl <= (butterFly_7_mux1h_276_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_12_0_i_adra_d <= butterFly_7_or_132_nl & mux1h_38_nl & butterFly_7_butterFly_7_or_179_nl
      & butterFly_7_or_60_nl & mux1h_39_nl & butterFly_7_or_238_nl;
  xx_rsc_12_0_i_wea_d <= STD_LOGIC_VECTOR'( and_333_seb & butterFly_7_butterFly_7_or_24_rmff);
  butterFly_7_butterFly_7_or_25_nl <= and_dcpl_279 OR (not_tmp_149 AND and_dcpl_207
      AND and_dcpl_245);
  nor_226_nl <= NOT((fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("011")));
  mux_802_nl <= MUX_s_1_2_2(nor_tmp_35, mux_171_cse, nor_226_nl);
  mux_794_nl <= MUX_s_1_2_2(nor_tmp_225, mux_163_cse, fsm_output(4));
  or_1062_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01100"))))
      OR (fsm_output(3));
  mux_788_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_1062_nl);
  mux_789_nl <= MUX_s_1_2_2(nor_tmp_35, mux_788_nl, fsm_output(1));
  mux_790_nl <= MUX_s_1_2_2(mux_789_nl, mux_213_cse, fsm_output(0));
  mux_791_nl <= MUX_s_1_2_2(nor_tmp_225, mux_790_nl, fsm_output(4));
  or_1060_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_795_nl <= MUX_s_1_2_2(mux_794_nl, mux_791_nl, or_1060_nl);
  mux_796_nl <= MUX_s_1_2_2(nor_tmp_35, mux_795_nl, fsm_output(5));
  mux_803_nl <= MUX_s_1_2_2(mux_802_nl, mux_796_nl, fsm_output(2));
  butterFly_7_and_323_nl <= (NOT(or_dcpl_199 AND and_dcpl_279)) AND mux_803_nl;
  xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_25_nl
      & butterFly_7_and_323_nl);
  xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_333_seb
      & butterFly_7_butterFly_7_or_24_rmff);
  butterFly_7_butterFly_7_mux_18_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_289);
  butterFly_7_or_129_nl <= (butterFly_7_butterFly_7_mux_18_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2287_nl <= NOT(and_dcpl_289 OR butterFly_7_or_360_cse);
  mux1h_36_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2287_nl & and_dcpl_289 & butterFly_7_or_360_cse));
  butterFly_7_mux_80_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_289);
  butterFly_7_butterFly_7_or_178_nl <= (butterFly_7_mux_80_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_182_nl <= and_339_ssc OR and_dcpl_289;
  butterFly_7_mux1h_204_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_182_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_59_nl <= (butterFly_7_mux1h_204_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_37_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_240_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_277_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_240_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_241_nl <= (butterFly_7_mux1h_277_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_13_0_i_adra_d <= butterFly_7_or_129_nl & mux1h_36_nl & butterFly_7_butterFly_7_or_178_nl
      & butterFly_7_or_59_nl & mux1h_37_nl & butterFly_7_or_241_nl;
  xx_rsc_13_0_i_wea_d <= STD_LOGIC_VECTOR'( and_344_seb & butterFly_7_butterFly_7_or_26_rmff);
  butterFly_7_butterFly_7_or_27_nl <= and_dcpl_289 OR and_dcpl_295;
  and_1947_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1101"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_242_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01101"))
      OR (NOT (fsm_output(1))));
  mux_841_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_242_nl);
  or_1119_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))))
      OR (fsm_output(3));
  mux_842_nl <= MUX_s_1_2_2(mux_841_nl, mux_162_cse, or_1119_nl);
  mux_843_nl <= MUX_s_1_2_2(mux_842_nl, mux_213_cse, fsm_output(0));
  mux_844_nl <= MUX_s_1_2_2(and_1947_nl, mux_843_nl, fsm_output(4));
  mux_845_nl <= MUX_s_1_2_2(nor_tmp_35, mux_844_nl, fsm_output(5));
  mux_853_nl <= MUX_s_1_2_2(mux_852_cse, mux_845_nl, fsm_output(2));
  butterFly_7_and_324_nl <= (NOT(or_dcpl_200 AND and_dcpl_289)) AND mux_853_nl;
  xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_27_nl
      & butterFly_7_and_324_nl);
  xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_344_seb
      & butterFly_7_butterFly_7_or_26_rmff);
  butterFly_7_butterFly_7_mux_17_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_299);
  butterFly_7_or_126_nl <= (butterFly_7_butterFly_7_mux_17_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2288_nl <= NOT(and_dcpl_299 OR butterFly_7_or_360_cse);
  mux1h_34_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2288_nl & and_dcpl_299 & butterFly_7_or_360_cse));
  butterFly_7_mux_79_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_299);
  butterFly_7_butterFly_7_or_177_nl <= (butterFly_7_mux_79_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_183_nl <= and_354_ssc OR and_dcpl_299;
  butterFly_7_mux1h_202_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_183_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_58_nl <= (butterFly_7_mux1h_202_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_35_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_243_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_278_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_243_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_244_nl <= (butterFly_7_mux1h_278_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_14_0_i_adra_d <= butterFly_7_or_126_nl & mux1h_34_nl & butterFly_7_butterFly_7_or_177_nl
      & butterFly_7_or_58_nl & mux1h_35_nl & butterFly_7_or_244_nl;
  xx_rsc_14_0_i_wea_d <= STD_LOGIC_VECTOR'( and_358_seb & butterFly_7_butterFly_7_or_28_rmff);
  butterFly_7_butterFly_7_or_29_nl <= and_dcpl_299 OR and_dcpl_295;
  and_1936_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1110"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_260_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("01110"))
      OR (NOT (fsm_output(1))));
  mux_889_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_260_nl);
  or_1173_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("01"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))))
      OR (fsm_output(3));
  mux_890_nl <= MUX_s_1_2_2(mux_889_nl, mux_162_cse, or_1173_nl);
  mux_891_nl <= MUX_s_1_2_2(mux_890_nl, mux_213_cse, fsm_output(0));
  mux_892_nl <= MUX_s_1_2_2(and_1936_nl, mux_891_nl, fsm_output(4));
  mux_893_nl <= MUX_s_1_2_2(nor_tmp_35, mux_892_nl, fsm_output(5));
  mux_901_nl <= MUX_s_1_2_2(mux_852_cse, mux_893_nl, fsm_output(2));
  butterFly_7_and_325_nl <= (NOT(or_dcpl_201 AND and_dcpl_299)) AND mux_901_nl;
  xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_29_nl
      & butterFly_7_and_325_nl);
  xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_358_seb
      & butterFly_7_butterFly_7_or_28_rmff);
  butterFly_7_butterFly_7_mux_16_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_305);
  butterFly_7_or_123_nl <= (butterFly_7_butterFly_7_mux_16_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2289_nl <= NOT(and_dcpl_305 OR butterFly_7_or_360_cse);
  mux1h_32_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2289_nl & and_dcpl_305 & butterFly_7_or_360_cse));
  butterFly_7_mux_78_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_305);
  butterFly_7_butterFly_7_or_176_nl <= (butterFly_7_mux_78_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_184_nl <= and_363_ssc OR and_dcpl_305;
  butterFly_7_mux1h_200_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_184_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_57_nl <= (butterFly_7_mux1h_200_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_33_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_246_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_279_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_246_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_247_nl <= (butterFly_7_mux1h_279_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_15_0_i_adra_d <= butterFly_7_or_123_nl & mux1h_32_nl & butterFly_7_butterFly_7_or_176_nl
      & butterFly_7_or_57_nl & mux1h_33_nl & butterFly_7_or_247_nl;
  xx_rsc_15_0_i_wea_d <= STD_LOGIC_VECTOR'( and_368_seb & butterFly_7_butterFly_7_or_30_rmff);
  butterFly_7_butterFly_7_or_31_nl <= and_dcpl_305 OR and_dcpl_295;
  or_1226_nl <= (fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"));
  mux_950_nl <= MUX_s_1_2_2(mux_223_cse, nor_tmp_35, or_1226_nl);
  mux_951_nl <= MUX_s_1_2_2(mux_950_nl, mux_847_cse, fsm_output(4));
  mux_952_nl <= MUX_s_1_2_2(mux_951_nl, nor_tmp_35, fsm_output(5));
  and_1917_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1111"))
      OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1918_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01111"))
      AND (fsm_output(1));
  mux_941_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1918_nl);
  or_1223_nl <= and_1919_cse OR (fsm_output(3));
  mux_942_nl <= MUX_s_1_2_2(mux_941_nl, mux_162_cse, or_1223_nl);
  mux_943_nl <= MUX_s_1_2_2(mux_942_nl, mux_213_cse, fsm_output(0));
  mux_944_nl <= MUX_s_1_2_2(and_1917_nl, mux_943_nl, fsm_output(4));
  mux_945_nl <= MUX_s_1_2_2(nor_tmp_35, mux_944_nl, fsm_output(5));
  mux_953_nl <= MUX_s_1_2_2(mux_952_nl, mux_945_nl, fsm_output(2));
  butterFly_7_and_326_nl <= (NOT(or_dcpl_202 AND and_dcpl_305)) AND mux_953_nl;
  xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_31_nl
      & butterFly_7_and_326_nl);
  xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_368_seb
      & butterFly_7_butterFly_7_or_30_rmff);
  butterFly_7_butterFly_7_mux_15_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_314);
  butterFly_7_or_120_nl <= (butterFly_7_butterFly_7_mux_15_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2290_nl <= NOT(and_dcpl_314 OR butterFly_7_or_360_cse);
  mux1h_30_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2290_nl & and_dcpl_314 & butterFly_7_or_360_cse));
  butterFly_7_mux_77_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_314);
  butterFly_7_butterFly_7_or_175_nl <= (butterFly_7_mux_77_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_185_nl <= and_372_ssc OR and_dcpl_314;
  butterFly_7_mux1h_198_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_185_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_56_nl <= (butterFly_7_mux1h_198_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_31_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_249_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_280_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_249_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_250_nl <= (butterFly_7_mux1h_280_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_16_0_i_adra_d <= butterFly_7_or_120_nl & mux1h_30_nl & butterFly_7_butterFly_7_or_175_nl
      & butterFly_7_or_56_nl & mux1h_31_nl & butterFly_7_or_250_nl;
  xx_rsc_16_0_i_wea_d <= STD_LOGIC_VECTOR'( and_381_seb & butterFly_7_butterFly_7_or_32_rmff);
  butterFly_7_butterFly_7_or_33_nl <= and_dcpl_314 OR (not_tmp_149 AND and_dcpl_319
      AND and_dcpl_140);
  or_1289_nl <= (fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("100"));
  mux_1010_nl <= MUX_s_1_2_2(mux_171_cse, nor_tmp_35, or_1289_nl);
  mux_1002_nl <= MUX_s_1_2_2(nor_tmp_299, mux_163_cse, fsm_output(4));
  or_1286_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10000"))))
      OR (fsm_output(3));
  mux_996_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_1286_nl);
  mux_997_nl <= MUX_s_1_2_2(nor_tmp_35, mux_996_nl, fsm_output(1));
  mux_998_nl <= MUX_s_1_2_2(mux_997_nl, mux_213_cse, fsm_output(0));
  mux_999_nl <= MUX_s_1_2_2(nor_tmp_299, mux_998_nl, fsm_output(4));
  or_1284_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1003_nl <= MUX_s_1_2_2(mux_1002_nl, mux_999_nl, or_1284_nl);
  mux_1004_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1003_nl, fsm_output(5));
  mux_1011_nl <= MUX_s_1_2_2(mux_1010_nl, mux_1004_nl, fsm_output(2));
  butterFly_7_and_327_nl <= (NOT(or_dcpl_205 AND and_dcpl_314)) AND mux_1011_nl;
  xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_33_nl
      & butterFly_7_and_327_nl);
  xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_381_seb
      & butterFly_7_butterFly_7_or_32_rmff);
  butterFly_7_butterFly_7_mux_14_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_325);
  butterFly_7_or_117_nl <= (butterFly_7_butterFly_7_mux_14_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2291_nl <= NOT(and_dcpl_325 OR butterFly_7_or_360_cse);
  mux1h_28_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2291_nl & and_dcpl_325 & butterFly_7_or_360_cse));
  butterFly_7_mux_76_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_325);
  butterFly_7_butterFly_7_or_174_nl <= (butterFly_7_mux_76_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_186_nl <= and_387_ssc OR and_dcpl_325;
  butterFly_7_mux1h_196_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_186_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_55_nl <= (butterFly_7_mux1h_196_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_29_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_252_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_281_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_252_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_253_nl <= (butterFly_7_mux1h_281_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_17_0_i_adra_d <= butterFly_7_or_117_nl & mux1h_28_nl & butterFly_7_butterFly_7_or_174_nl
      & butterFly_7_or_55_nl & mux1h_29_nl & butterFly_7_or_253_nl;
  xx_rsc_17_0_i_wea_d <= STD_LOGIC_VECTOR'( and_393_seb & butterFly_7_butterFly_7_or_34_rmff);
  butterFly_7_butterFly_7_or_35_nl <= and_dcpl_325 OR and_dcpl_332;
  and_1897_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0001"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_314_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10001"))
      OR (NOT (fsm_output(1))));
  mux_1052_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_314_nl);
  or_1341_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))))
      OR (fsm_output(3));
  mux_1053_nl <= MUX_s_1_2_2(mux_1052_nl, mux_162_cse, or_1341_nl);
  mux_1054_nl <= MUX_s_1_2_2(mux_1053_nl, mux_213_cse, fsm_output(0));
  mux_1055_nl <= MUX_s_1_2_2(and_1897_nl, mux_1054_nl, fsm_output(4));
  mux_1056_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1055_nl, fsm_output(5));
  mux_1064_nl <= MUX_s_1_2_2(mux_1063_cse, mux_1056_nl, fsm_output(2));
  butterFly_7_and_328_nl <= (NOT(or_dcpl_206 AND and_dcpl_325)) AND mux_1064_nl;
  xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_35_nl
      & butterFly_7_and_328_nl);
  xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_393_seb
      & butterFly_7_butterFly_7_or_34_rmff);
  butterFly_7_butterFly_7_mux_13_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_336);
  butterFly_7_or_114_nl <= (butterFly_7_butterFly_7_mux_13_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2292_nl <= NOT(and_dcpl_336 OR butterFly_7_or_360_cse);
  mux1h_26_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2292_nl & and_dcpl_336 & butterFly_7_or_360_cse));
  butterFly_7_mux_75_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_336);
  butterFly_7_butterFly_7_or_173_nl <= (butterFly_7_mux_75_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_187_nl <= and_402_ssc OR and_dcpl_336;
  butterFly_7_mux1h_194_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_187_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_54_nl <= (butterFly_7_mux1h_194_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_27_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_255_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_282_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_255_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_256_nl <= (butterFly_7_mux1h_282_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_18_0_i_adra_d <= butterFly_7_or_114_nl & mux1h_26_nl & butterFly_7_butterFly_7_or_173_nl
      & butterFly_7_or_54_nl & mux1h_27_nl & butterFly_7_or_256_nl;
  xx_rsc_18_0_i_wea_d <= STD_LOGIC_VECTOR'( and_406_seb & butterFly_7_butterFly_7_or_36_rmff);
  butterFly_7_butterFly_7_or_37_nl <= and_dcpl_336 OR and_dcpl_332;
  and_1888_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_327_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10010"))
      OR (NOT (fsm_output(1))));
  mux_1103_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_327_nl);
  or_1394_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))))
      OR (fsm_output(3));
  mux_1104_nl <= MUX_s_1_2_2(mux_1103_nl, mux_162_cse, or_1394_nl);
  mux_1105_nl <= MUX_s_1_2_2(mux_1104_nl, mux_213_cse, fsm_output(0));
  mux_1106_nl <= MUX_s_1_2_2(and_1888_nl, mux_1105_nl, fsm_output(4));
  mux_1107_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1106_nl, fsm_output(5));
  mux_1115_nl <= MUX_s_1_2_2(mux_1063_cse, mux_1107_nl, fsm_output(2));
  butterFly_7_and_329_nl <= (NOT(or_dcpl_208 AND and_dcpl_336)) AND mux_1115_nl;
  xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_37_nl
      & butterFly_7_and_329_nl);
  xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_406_seb
      & butterFly_7_butterFly_7_or_36_rmff);
  butterFly_7_butterFly_7_mux_12_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_342);
  butterFly_7_or_111_nl <= (butterFly_7_butterFly_7_mux_12_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2293_nl <= NOT(and_dcpl_342 OR butterFly_7_or_360_cse);
  mux1h_24_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2293_nl & and_dcpl_342 & butterFly_7_or_360_cse));
  butterFly_7_mux_74_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_342);
  butterFly_7_butterFly_7_or_172_nl <= (butterFly_7_mux_74_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_188_nl <= and_410_ssc OR and_dcpl_342;
  butterFly_7_mux1h_192_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_188_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_53_nl <= (butterFly_7_mux1h_192_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_25_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_258_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_283_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_258_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_259_nl <= (butterFly_7_mux1h_283_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_19_0_i_adra_d <= butterFly_7_or_111_nl & mux1h_24_nl & butterFly_7_butterFly_7_or_172_nl
      & butterFly_7_or_53_nl & mux1h_25_nl & butterFly_7_or_259_nl;
  xx_rsc_19_0_i_wea_d <= STD_LOGIC_VECTOR'( and_415_seb & butterFly_7_butterFly_7_or_38_rmff);
  butterFly_7_butterFly_7_or_39_nl <= and_dcpl_342 OR and_dcpl_332;
  and_1875_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0011"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_347_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10011"))
      OR (NOT (fsm_output(1))));
  mux_1158_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_347_nl);
  or_1446_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("011"))))
      OR (fsm_output(3));
  mux_1159_nl <= MUX_s_1_2_2(mux_1158_nl, mux_162_cse, or_1446_nl);
  mux_1160_nl <= MUX_s_1_2_2(mux_1159_nl, mux_213_cse, fsm_output(0));
  mux_1161_nl <= MUX_s_1_2_2(and_1875_nl, mux_1160_nl, fsm_output(4));
  mux_1162_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1161_nl, fsm_output(5));
  mux_1170_nl <= MUX_s_1_2_2(mux_1063_cse, mux_1162_nl, fsm_output(2));
  butterFly_7_and_330_nl <= (NOT(or_dcpl_209 AND and_dcpl_342)) AND mux_1170_nl;
  xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_39_nl
      & butterFly_7_and_330_nl);
  xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_415_seb
      & butterFly_7_butterFly_7_or_38_rmff);
  butterFly_7_butterFly_7_mux_11_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_351);
  butterFly_7_or_108_nl <= (butterFly_7_butterFly_7_mux_11_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2294_nl <= NOT(and_dcpl_351 OR butterFly_7_or_360_cse);
  mux1h_22_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2294_nl & and_dcpl_351 & butterFly_7_or_360_cse));
  butterFly_7_mux_73_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_351);
  butterFly_7_butterFly_7_or_171_nl <= (butterFly_7_mux_73_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_189_nl <= and_419_ssc OR and_dcpl_351;
  butterFly_7_mux1h_190_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_189_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_52_nl <= (butterFly_7_mux1h_190_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_23_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_261_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_284_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_261_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_262_nl <= (butterFly_7_mux1h_284_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_20_0_i_adra_d <= butterFly_7_or_108_nl & mux1h_22_nl & butterFly_7_butterFly_7_or_171_nl
      & butterFly_7_or_52_nl & mux1h_23_nl & butterFly_7_or_262_nl;
  xx_rsc_20_0_i_wea_d <= STD_LOGIC_VECTOR'( and_427_seb & butterFly_7_butterFly_7_or_40_rmff);
  butterFly_7_butterFly_7_or_41_nl <= and_dcpl_351 OR (not_tmp_149 AND and_dcpl_355
      AND and_dcpl_140);
  nor_367_nl <= NOT((fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("101")));
  mux_1227_nl <= MUX_s_1_2_2(nor_tmp_35, mux_171_cse, nor_367_nl);
  mux_1219_nl <= MUX_s_1_2_2(nor_tmp_366, mux_163_cse, fsm_output(4));
  or_1513_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10100"))))
      OR (fsm_output(3));
  mux_1213_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_1513_nl);
  mux_1214_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1213_nl, fsm_output(1));
  mux_1215_nl <= MUX_s_1_2_2(mux_1214_nl, mux_213_cse, fsm_output(0));
  mux_1216_nl <= MUX_s_1_2_2(nor_tmp_366, mux_1215_nl, fsm_output(4));
  or_1511_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1220_nl <= MUX_s_1_2_2(mux_1219_nl, mux_1216_nl, or_1511_nl);
  mux_1221_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1220_nl, fsm_output(5));
  mux_1228_nl <= MUX_s_1_2_2(mux_1227_nl, mux_1221_nl, fsm_output(2));
  butterFly_7_and_331_nl <= (NOT(or_dcpl_212 AND and_dcpl_351)) AND mux_1228_nl;
  xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_41_nl
      & butterFly_7_and_331_nl);
  xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_427_seb
      & butterFly_7_butterFly_7_or_40_rmff);
  butterFly_7_butterFly_7_mux_10_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_361);
  butterFly_7_or_105_nl <= (butterFly_7_butterFly_7_mux_10_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2295_nl <= NOT(and_dcpl_361 OR butterFly_7_or_360_cse);
  mux1h_20_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2295_nl & and_dcpl_361 & butterFly_7_or_360_cse));
  butterFly_7_mux_72_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_361);
  butterFly_7_butterFly_7_or_170_nl <= (butterFly_7_mux_72_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_190_nl <= and_433_ssc OR and_dcpl_361;
  butterFly_7_mux1h_188_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_190_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_51_nl <= (butterFly_7_mux1h_188_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_21_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_264_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_285_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_264_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_265_nl <= (butterFly_7_mux1h_285_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_21_0_i_adra_d <= butterFly_7_or_105_nl & mux1h_20_nl & butterFly_7_butterFly_7_or_170_nl
      & butterFly_7_or_51_nl & mux1h_21_nl & butterFly_7_or_265_nl;
  xx_rsc_21_0_i_wea_d <= STD_LOGIC_VECTOR'( and_438_seb & butterFly_7_butterFly_7_or_42_rmff);
  butterFly_7_butterFly_7_or_43_nl <= and_dcpl_361 OR and_dcpl_367;
  and_1853_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0101"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_386_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10101"))
      OR (NOT (fsm_output(1))));
  mux_1270_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_386_nl);
  or_1579_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("101"))))
      OR (fsm_output(3));
  mux_1271_nl <= MUX_s_1_2_2(mux_1270_nl, mux_162_cse, or_1579_nl);
  mux_1272_nl <= MUX_s_1_2_2(mux_1271_nl, mux_213_cse, fsm_output(0));
  mux_1273_nl <= MUX_s_1_2_2(and_1853_nl, mux_1272_nl, fsm_output(4));
  mux_1274_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1273_nl, fsm_output(5));
  mux_1282_nl <= MUX_s_1_2_2(mux_1281_cse, mux_1274_nl, fsm_output(2));
  butterFly_7_and_332_nl <= (NOT(or_dcpl_213 AND and_dcpl_361)) AND mux_1282_nl;
  xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_43_nl
      & butterFly_7_and_332_nl);
  xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_438_seb
      & butterFly_7_butterFly_7_or_42_rmff);
  butterFly_7_butterFly_7_mux_9_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_371);
  butterFly_7_or_102_nl <= (butterFly_7_butterFly_7_mux_9_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2296_nl <= NOT(and_dcpl_371 OR butterFly_7_or_360_cse);
  mux1h_18_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2296_nl & and_dcpl_371 & butterFly_7_or_360_cse));
  butterFly_7_mux_71_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_371);
  butterFly_7_butterFly_7_or_169_nl <= (butterFly_7_mux_71_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_191_nl <= and_447_ssc OR and_dcpl_371;
  butterFly_7_mux1h_186_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_191_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_50_nl <= (butterFly_7_mux1h_186_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_19_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_267_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_286_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_267_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_268_nl <= (butterFly_7_mux1h_286_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_22_0_i_adra_d <= butterFly_7_or_102_nl & mux1h_18_nl & butterFly_7_butterFly_7_or_169_nl
      & butterFly_7_or_50_nl & mux1h_19_nl & butterFly_7_or_268_nl;
  xx_rsc_22_0_i_wea_d <= STD_LOGIC_VECTOR'( and_451_seb & butterFly_7_butterFly_7_or_44_rmff);
  butterFly_7_butterFly_7_or_45_nl <= and_dcpl_371 OR and_dcpl_367;
  and_1842_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0110"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_405_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("10110"))
      OR (NOT (fsm_output(1))));
  mux_1321_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_405_nl);
  or_1639_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("10"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110"))))
      OR (fsm_output(3));
  mux_1322_nl <= MUX_s_1_2_2(mux_1321_nl, mux_162_cse, or_1639_nl);
  mux_1323_nl <= MUX_s_1_2_2(mux_1322_nl, mux_213_cse, fsm_output(0));
  mux_1324_nl <= MUX_s_1_2_2(and_1842_nl, mux_1323_nl, fsm_output(4));
  mux_1325_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1324_nl, fsm_output(5));
  mux_1333_nl <= MUX_s_1_2_2(mux_1281_cse, mux_1325_nl, fsm_output(2));
  butterFly_7_and_333_nl <= (NOT(or_dcpl_215 AND and_dcpl_371)) AND mux_1333_nl;
  xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_45_nl
      & butterFly_7_and_333_nl);
  xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_451_seb
      & butterFly_7_butterFly_7_or_44_rmff);
  butterFly_7_butterFly_7_mux_8_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_377);
  butterFly_7_or_99_nl <= (butterFly_7_butterFly_7_mux_8_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2297_nl <= NOT(and_dcpl_377 OR butterFly_7_or_360_cse);
  mux1h_16_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2297_nl & and_dcpl_377 & butterFly_7_or_360_cse));
  butterFly_7_mux_70_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_377);
  butterFly_7_butterFly_7_or_168_nl <= (butterFly_7_mux_70_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_192_nl <= and_455_ssc OR and_dcpl_377;
  butterFly_7_mux1h_184_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_192_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_49_nl <= (butterFly_7_mux1h_184_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_17_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_270_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_287_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_270_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_271_nl <= (butterFly_7_mux1h_287_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_23_0_i_adra_d <= butterFly_7_or_99_nl & mux1h_16_nl & butterFly_7_butterFly_7_or_168_nl
      & butterFly_7_or_49_nl & mux1h_17_nl & butterFly_7_or_271_nl;
  xx_rsc_23_0_i_wea_d <= STD_LOGIC_VECTOR'( and_460_seb & butterFly_7_butterFly_7_or_46_rmff);
  butterFly_7_butterFly_7_or_47_nl <= and_dcpl_377 OR and_dcpl_367;
  and_1825_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0111"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1826_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10111"))
      AND (fsm_output(1));
  mux_1376_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1826_nl);
  or_1698_nl <= and_1827_cse OR (fsm_output(3));
  mux_1377_nl <= MUX_s_1_2_2(mux_1376_nl, mux_162_cse, or_1698_nl);
  mux_1378_nl <= MUX_s_1_2_2(mux_1377_nl, mux_213_cse, fsm_output(0));
  mux_1379_nl <= MUX_s_1_2_2(and_1825_nl, mux_1378_nl, fsm_output(4));
  mux_1380_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1379_nl, fsm_output(5));
  mux_1388_nl <= MUX_s_1_2_2(mux_1281_cse, mux_1380_nl, fsm_output(2));
  butterFly_7_and_334_nl <= (NOT(or_dcpl_216 AND and_dcpl_377)) AND mux_1388_nl;
  xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_47_nl
      & butterFly_7_and_334_nl);
  xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_460_seb
      & butterFly_7_butterFly_7_or_46_rmff);
  butterFly_7_butterFly_7_mux_7_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_384);
  butterFly_7_or_96_nl <= (butterFly_7_butterFly_7_mux_7_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2298_nl <= NOT(and_dcpl_384 OR butterFly_7_or_360_cse);
  mux1h_14_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2298_nl & and_dcpl_384 & butterFly_7_or_360_cse));
  butterFly_7_mux_69_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_384);
  butterFly_7_butterFly_7_or_167_nl <= (butterFly_7_mux_69_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_193_nl <= and_464_ssc OR and_dcpl_384;
  butterFly_7_mux1h_182_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_193_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_48_nl <= (butterFly_7_mux1h_182_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_15_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_273_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_288_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_273_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_274_nl <= (butterFly_7_mux1h_288_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_24_0_i_adra_d <= butterFly_7_or_96_nl & mux1h_14_nl & butterFly_7_butterFly_7_or_167_nl
      & butterFly_7_or_48_nl & mux1h_15_nl & butterFly_7_or_274_nl;
  xx_rsc_24_0_i_wea_d <= STD_LOGIC_VECTOR'( and_470_seb & butterFly_7_butterFly_7_or_48_rmff);
  butterFly_7_butterFly_7_or_49_nl <= and_dcpl_384 OR (not_tmp_149 AND and_dcpl_319
      AND and_dcpl_245);
  or_1764_nl <= (fsm_output(5)) OR CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("110"));
  mux_1445_nl <= MUX_s_1_2_2(mux_171_cse, nor_tmp_35, or_1764_nl);
  mux_1437_nl <= MUX_s_1_2_2(nor_tmp_445, mux_163_cse, fsm_output(4));
  or_1761_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11000"))))
      OR (fsm_output(3));
  mux_1431_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_1761_nl);
  mux_1432_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1431_nl, fsm_output(1));
  mux_1433_nl <= MUX_s_1_2_2(mux_1432_nl, mux_213_cse, fsm_output(0));
  mux_1434_nl <= MUX_s_1_2_2(nor_tmp_445, mux_1433_nl, fsm_output(4));
  or_1759_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000"));
  mux_1438_nl <= MUX_s_1_2_2(mux_1437_nl, mux_1434_nl, or_1759_nl);
  mux_1439_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1438_nl, fsm_output(5));
  mux_1446_nl <= MUX_s_1_2_2(mux_1445_nl, mux_1439_nl, fsm_output(2));
  butterFly_7_and_335_nl <= (NOT(or_dcpl_217 AND and_dcpl_384)) AND mux_1446_nl;
  xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_49_nl
      & butterFly_7_and_335_nl);
  xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_470_seb
      & butterFly_7_butterFly_7_or_48_rmff);
  butterFly_7_butterFly_7_mux_6_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_393);
  butterFly_7_or_93_nl <= (butterFly_7_butterFly_7_mux_6_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2299_nl <= NOT(and_dcpl_393 OR butterFly_7_or_360_cse);
  mux1h_12_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2299_nl & and_dcpl_393 & butterFly_7_or_360_cse));
  butterFly_7_mux_68_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_393);
  butterFly_7_butterFly_7_or_166_nl <= (butterFly_7_mux_68_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_194_nl <= and_475_ssc OR and_dcpl_393;
  butterFly_7_mux1h_180_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_194_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_47_nl <= (butterFly_7_mux1h_180_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_13_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_276_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_289_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_276_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_277_nl <= (butterFly_7_mux1h_289_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_25_0_i_adra_d <= butterFly_7_or_93_nl & mux1h_12_nl & butterFly_7_butterFly_7_or_166_nl
      & butterFly_7_or_47_nl & mux1h_13_nl & butterFly_7_or_277_nl;
  xx_rsc_25_0_i_wea_d <= STD_LOGIC_VECTOR'( and_481_seb & butterFly_7_butterFly_7_or_50_rmff);
  butterFly_7_butterFly_7_or_51_nl <= and_dcpl_393 OR and_dcpl_400;
  and_1802_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1001"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_464_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11001"))
      OR (NOT (fsm_output(1))));
  mux_1487_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_464_nl);
  or_1815_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("001"))))
      OR (fsm_output(3));
  mux_1488_nl <= MUX_s_1_2_2(mux_1487_nl, mux_162_cse, or_1815_nl);
  mux_1489_nl <= MUX_s_1_2_2(mux_1488_nl, mux_213_cse, fsm_output(0));
  mux_1490_nl <= MUX_s_1_2_2(and_1802_nl, mux_1489_nl, fsm_output(4));
  mux_1491_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1490_nl, fsm_output(5));
  mux_1499_nl <= MUX_s_1_2_2(mux_1498_cse, mux_1491_nl, fsm_output(2));
  butterFly_7_and_336_nl <= (NOT(or_dcpl_218 AND and_dcpl_393)) AND mux_1499_nl;
  xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_51_nl
      & butterFly_7_and_336_nl);
  xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_481_seb
      & butterFly_7_butterFly_7_or_50_rmff);
  butterFly_7_butterFly_7_mux_5_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_404);
  butterFly_7_or_90_nl <= (butterFly_7_butterFly_7_mux_5_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2300_nl <= NOT(and_dcpl_404 OR butterFly_7_or_360_cse);
  mux1h_10_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2300_nl & and_dcpl_404 & butterFly_7_or_360_cse));
  butterFly_7_mux_67_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_404);
  butterFly_7_butterFly_7_or_165_nl <= (butterFly_7_mux_67_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_195_nl <= and_490_ssc OR and_dcpl_404;
  butterFly_7_mux1h_178_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_195_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_46_nl <= (butterFly_7_mux1h_178_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_11_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_279_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_290_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_279_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_280_nl <= (butterFly_7_mux1h_290_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_26_0_i_adra_d <= butterFly_7_or_90_nl & mux1h_10_nl & butterFly_7_butterFly_7_or_165_nl
      & butterFly_7_or_46_nl & mux1h_11_nl & butterFly_7_or_280_nl;
  xx_rsc_26_0_i_wea_d <= STD_LOGIC_VECTOR'( and_494_seb & butterFly_7_butterFly_7_or_52_rmff);
  butterFly_7_butterFly_7_or_53_nl <= and_dcpl_404 OR and_dcpl_400;
  nor_483_nl <= NOT((fsm_output(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("110")));
  mux_1547_nl <= MUX_s_1_2_2(nor_tmp_35, mux_223_cse, nor_483_nl);
  mux_1548_nl <= MUX_s_1_2_2(mux_1547_nl, mux_1493_cse, fsm_output(4));
  mux_1549_nl <= MUX_s_1_2_2(mux_1548_nl, nor_tmp_35, fsm_output(5));
  and_1790_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1010"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  nor_480_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11010"))
      OR (NOT (fsm_output(1))));
  mux_1538_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), nor_480_nl);
  or_1869_nl <= (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("010"))))
      OR (fsm_output(3));
  mux_1539_nl <= MUX_s_1_2_2(mux_1538_nl, mux_162_cse, or_1869_nl);
  mux_1540_nl <= MUX_s_1_2_2(mux_1539_nl, mux_213_cse, fsm_output(0));
  mux_1541_nl <= MUX_s_1_2_2(and_1790_nl, mux_1540_nl, fsm_output(4));
  mux_1542_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1541_nl, fsm_output(5));
  mux_1550_nl <= MUX_s_1_2_2(mux_1549_nl, mux_1542_nl, fsm_output(2));
  butterFly_7_and_337_nl <= (NOT(or_dcpl_219 AND and_dcpl_404)) AND mux_1550_nl;
  xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_53_nl
      & butterFly_7_and_337_nl);
  xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_494_seb
      & butterFly_7_butterFly_7_or_52_rmff);
  butterFly_7_butterFly_7_mux_4_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_410);
  butterFly_7_or_87_nl <= (butterFly_7_butterFly_7_mux_4_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2301_nl <= NOT(and_dcpl_410 OR butterFly_7_or_360_cse);
  mux1h_8_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2301_nl & and_dcpl_410 & butterFly_7_or_360_cse));
  butterFly_7_mux_66_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_410);
  butterFly_7_butterFly_7_or_164_nl <= (butterFly_7_mux_66_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_196_nl <= and_498_ssc OR and_dcpl_410;
  butterFly_7_mux1h_176_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_196_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_45_nl <= (butterFly_7_mux1h_176_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_9_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_282_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_291_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_282_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_283_nl <= (butterFly_7_mux1h_291_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_27_0_i_adra_d <= butterFly_7_or_87_nl & mux1h_8_nl & butterFly_7_butterFly_7_or_164_nl
      & butterFly_7_or_45_nl & mux1h_9_nl & butterFly_7_or_283_nl;
  xx_rsc_27_0_i_wea_d <= STD_LOGIC_VECTOR'( and_503_seb & butterFly_7_butterFly_7_or_54_rmff);
  butterFly_7_butterFly_7_or_55_nl <= and_dcpl_410 OR and_dcpl_400;
  and_1771_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1011"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1772_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11011"))
      AND (fsm_output(1));
  mux_1593_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1772_nl);
  or_1925_nl <= and_1773_cse OR (fsm_output(3));
  mux_1594_nl <= MUX_s_1_2_2(mux_1593_nl, mux_162_cse, or_1925_nl);
  mux_1595_nl <= MUX_s_1_2_2(mux_1594_nl, mux_213_cse, fsm_output(0));
  mux_1596_nl <= MUX_s_1_2_2(and_1771_nl, mux_1595_nl, fsm_output(4));
  mux_1597_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1596_nl, fsm_output(5));
  mux_1605_nl <= MUX_s_1_2_2(mux_1498_cse, mux_1597_nl, fsm_output(2));
  butterFly_7_and_338_nl <= (NOT(or_dcpl_220 AND and_dcpl_410)) AND mux_1605_nl;
  xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_55_nl
      & butterFly_7_and_338_nl);
  xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_503_seb
      & butterFly_7_butterFly_7_or_54_rmff);
  butterFly_7_butterFly_7_mux_3_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_417);
  butterFly_7_or_84_nl <= (butterFly_7_butterFly_7_mux_3_nl AND (NOT and_dcpl_114))
      OR and_dcpl_102;
  nor_2302_nl <= NOT(and_dcpl_417 OR butterFly_7_or_360_cse);
  mux1h_6_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2302_nl & and_dcpl_417 & butterFly_7_or_360_cse));
  butterFly_7_mux_65_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_417);
  butterFly_7_butterFly_7_or_163_nl <= (butterFly_7_mux_65_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_197_nl <= and_507_ssc OR and_dcpl_417;
  butterFly_7_mux1h_174_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_197_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_44_nl <= (butterFly_7_mux1h_174_nl AND (NOT and_dcpl_102)) OR and_dcpl_114;
  mux1h_7_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_285_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_292_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_285_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_286_nl <= (butterFly_7_mux1h_292_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_28_0_i_adra_d <= butterFly_7_or_84_nl & mux1h_6_nl & butterFly_7_butterFly_7_or_163_nl
      & butterFly_7_or_44_nl & mux1h_7_nl & butterFly_7_or_286_nl;
  xx_rsc_28_0_i_wea_d <= STD_LOGIC_VECTOR'( and_513_seb & butterFly_7_butterFly_7_or_56_rmff);
  butterFly_7_butterFly_7_or_57_nl <= and_dcpl_417 OR (not_tmp_149 AND and_dcpl_355
      AND and_dcpl_245);
  and_1759_nl <= (NOT (fsm_output(5))) AND CONV_SL_1_1(operator_20_true_28_acc_tmp=STD_LOGIC_VECTOR'("111"));
  mux_1662_nl <= MUX_s_1_2_2(nor_tmp_35, mux_171_cse, and_1759_nl);
  mux_1654_nl <= MUX_s_1_2_2(nor_tmp_525, mux_163_cse, fsm_output(4));
  or_1991_nl <= (NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp/=STD_LOGIC_VECTOR'("11100"))))
      OR (fsm_output(3));
  mux_1648_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), or_1991_nl);
  mux_1649_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1648_nl, fsm_output(1));
  mux_1650_nl <= MUX_s_1_2_2(mux_1649_nl, mux_213_cse, fsm_output(0));
  mux_1651_nl <= MUX_s_1_2_2(nor_tmp_525, mux_1650_nl, fsm_output(4));
  or_1989_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("11"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("100"));
  mux_1655_nl <= MUX_s_1_2_2(mux_1654_nl, mux_1651_nl, or_1989_nl);
  mux_1656_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1655_nl, fsm_output(5));
  mux_1663_nl <= MUX_s_1_2_2(mux_1662_nl, mux_1656_nl, fsm_output(2));
  butterFly_7_and_339_nl <= (NOT(or_dcpl_221 AND and_dcpl_417)) AND mux_1663_nl;
  xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_57_nl
      & butterFly_7_and_339_nl);
  xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_513_seb
      & butterFly_7_butterFly_7_or_56_rmff);
  butterFly_7_butterFly_7_mux_2_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_426);
  butterFly_7_or_81_nl <= (butterFly_7_butterFly_7_mux_2_nl AND (NOT and_dcpl_154))
      OR and_dcpl_149;
  nor_2303_nl <= NOT(and_dcpl_426 OR butterFly_7_or_360_cse);
  mux1h_4_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2303_nl & and_dcpl_426 & butterFly_7_or_360_cse));
  butterFly_7_mux_64_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_426);
  butterFly_7_butterFly_7_or_162_nl <= (butterFly_7_mux_64_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_198_nl <= and_518_ssc OR and_dcpl_426;
  butterFly_7_mux1h_172_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_198_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_43_nl <= (butterFly_7_mux1h_172_nl AND (NOT and_dcpl_149)) OR and_dcpl_154;
  mux1h_5_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_288_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_293_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_288_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_289_nl <= (butterFly_7_mux1h_293_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_29_0_i_adra_d <= butterFly_7_or_81_nl & mux1h_4_nl & butterFly_7_butterFly_7_or_162_nl
      & butterFly_7_or_43_nl & mux1h_5_nl & butterFly_7_or_289_nl;
  xx_rsc_29_0_i_wea_d <= STD_LOGIC_VECTOR'( and_523_seb & butterFly_7_butterFly_7_or_58_rmff);
  butterFly_7_butterFly_7_or_59_nl <= and_dcpl_426 OR and_dcpl_432;
  and_1738_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1101"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1739_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11101"))
      AND (fsm_output(1));
  mux_1704_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1739_nl);
  or_2043_nl <= and_1740_cse OR (fsm_output(3));
  mux_1705_nl <= MUX_s_1_2_2(mux_1704_nl, mux_162_cse, or_2043_nl);
  mux_1706_nl <= MUX_s_1_2_2(mux_1705_nl, mux_213_cse, fsm_output(0));
  mux_1707_nl <= MUX_s_1_2_2(and_1738_nl, mux_1706_nl, fsm_output(4));
  mux_1708_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1707_nl, fsm_output(5));
  mux_1716_nl <= MUX_s_1_2_2(mux_1715_cse, mux_1708_nl, fsm_output(2));
  butterFly_7_and_340_nl <= (NOT(or_dcpl_222 AND and_dcpl_426)) AND mux_1716_nl;
  xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_59_nl
      & butterFly_7_and_340_nl);
  xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_523_seb
      & butterFly_7_butterFly_7_or_58_rmff);
  butterFly_7_butterFly_7_mux_1_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_436);
  butterFly_7_or_78_nl <= (butterFly_7_butterFly_7_mux_1_nl AND (NOT and_dcpl_173))
      OR and_dcpl_171;
  nor_2304_nl <= NOT(and_dcpl_436 OR butterFly_7_or_360_cse);
  mux1h_2_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2304_nl & and_dcpl_436 & butterFly_7_or_360_cse));
  butterFly_7_mux_63_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), and_dcpl_436);
  butterFly_7_butterFly_7_or_161_nl <= (butterFly_7_mux_63_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_199_nl <= and_532_ssc OR and_dcpl_436;
  butterFly_7_mux1h_170_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_199_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_42_nl <= (butterFly_7_mux1h_170_nl AND (NOT and_dcpl_171)) OR and_dcpl_173;
  mux1h_3_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_291_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_294_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_291_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_292_nl <= (butterFly_7_mux1h_294_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_30_0_i_adra_d <= butterFly_7_or_78_nl & mux1h_2_nl & butterFly_7_butterFly_7_or_161_nl
      & butterFly_7_or_42_nl & mux1h_3_nl & butterFly_7_or_292_nl;
  xx_rsc_30_0_i_wea_d <= STD_LOGIC_VECTOR'( and_536_seb & butterFly_7_butterFly_7_or_60_rmff);
  butterFly_7_butterFly_7_or_61_nl <= and_dcpl_436 OR and_dcpl_432;
  and_1719_nl <= ((NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("1110"))
      OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg) OR (fsm_output(0)) OR (fsm_output(3))
      OR (NOT (fsm_output(1))))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1720_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11110"))
      AND (fsm_output(1));
  mux_1755_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1720_nl);
  or_2092_nl <= and_1721_cse OR (fsm_output(3));
  mux_1756_nl <= MUX_s_1_2_2(mux_1755_nl, mux_162_cse, or_2092_nl);
  mux_1757_nl <= MUX_s_1_2_2(mux_1756_nl, mux_213_cse, fsm_output(0));
  mux_1758_nl <= MUX_s_1_2_2(and_1719_nl, mux_1757_nl, fsm_output(4));
  mux_1759_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1758_nl, fsm_output(5));
  mux_1767_nl <= MUX_s_1_2_2(mux_1715_cse, mux_1759_nl, fsm_output(2));
  butterFly_7_and_341_nl <= (NOT(or_dcpl_223 AND and_dcpl_436)) AND mux_1767_nl;
  xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_61_nl
      & butterFly_7_and_341_nl);
  xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_536_seb
      & butterFly_7_butterFly_7_or_60_rmff);
  butterFly_7_butterFly_7_mux_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), and_dcpl_442);
  butterFly_7_or_75_nl <= (butterFly_7_butterFly_7_mux_nl AND (NOT and_dcpl_187))
      OR and_dcpl_184;
  nor_2305_nl <= NOT(and_dcpl_442 OR butterFly_7_or_360_cse);
  mux1h_nl <= MUX1HOT_v_3_3_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)),
      ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      nor_2305_nl & and_dcpl_442 & butterFly_7_or_360_cse));
  butterFly_7_mux_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      and_dcpl_442);
  butterFly_7_butterFly_7_or_160_nl <= (butterFly_7_mux_nl AND (NOT and_dcpl_100))
      OR and_dcpl_116;
  butterFly_7_or_200_nl <= and_540_ssc OR and_dcpl_442;
  butterFly_7_mux1h_168_nl <= MUX1HOT_s_1_5_2((reg_drf_revArr_ptr_1_smx_9_0_reg(1)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)), reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_360_cse & butterFly_7_or_200_nl & and_dcpl_109
      & and_dcpl_112));
  butterFly_7_or_41_nl <= (butterFly_7_mux1h_168_nl AND (NOT and_dcpl_184)) OR and_dcpl_187;
  mux1h_1_nl <= MUX1HOT_v_3_5_2(((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3 DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3
      DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2 DOWNTO 0)), STD_LOGIC_VECTOR'(
      and_dcpl_97 & butterFly_7_or_294_cse & and_dcpl_109 & and_dcpl_112 & butterFly_7_or_360_cse));
  butterFly_7_mux1h_295_nl <= MUX1HOT_s_1_4_2((reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)),
      (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)), (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)),
      (S1_OUTER_LOOP_for_acc_svs_3_0(0)), STD_LOGIC_VECTOR'( and_dcpl_97 & butterFly_7_or_294_cse
      & and_dcpl_109 & and_dcpl_112));
  butterFly_7_or_295_nl <= (butterFly_7_mux1h_295_nl AND (NOT and_dcpl_116)) OR and_dcpl_100;
  xx_rsc_31_0_i_adra_d <= butterFly_7_or_75_nl & mux1h_nl & butterFly_7_butterFly_7_or_160_nl
      & butterFly_7_or_41_nl & mux1h_1_nl & butterFly_7_or_295_nl;
  xx_rsc_31_0_i_wea_d <= STD_LOGIC_VECTOR'( and_546_seb & butterFly_7_butterFly_7_or_62_rmff);
  butterFly_7_butterFly_7_or_63_nl <= and_dcpl_442 OR and_dcpl_432;
  and_1689_nl <= ((CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg=STD_LOGIC_VECTOR'("1111"))
      AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg AND (NOT (fsm_output(0))) AND (NOT (fsm_output(3)))
      AND (fsm_output(1))) OR (fsm_output(7))) AND (fsm_output(6));
  and_1691_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11111"))
      AND (fsm_output(1));
  mux_1806_nl <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(7)), and_1691_nl);
  or_2130_nl <= and_1692_cse OR (fsm_output(3));
  mux_1807_nl <= MUX_s_1_2_2(mux_1806_nl, mux_162_cse, or_2130_nl);
  mux_1808_nl <= MUX_s_1_2_2(mux_1807_nl, mux_213_cse, fsm_output(0));
  mux_1809_nl <= MUX_s_1_2_2(and_1689_nl, mux_1808_nl, fsm_output(4));
  mux_1810_nl <= MUX_s_1_2_2(nor_tmp_35, mux_1809_nl, fsm_output(5));
  mux_1818_nl <= MUX_s_1_2_2(mux_1715_cse, mux_1810_nl, fsm_output(2));
  butterFly_7_and_342_nl <= (NOT((or_dcpl_214 OR or_dcpl_195) AND and_dcpl_442))
      AND mux_1818_nl;
  xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_butterFly_7_or_63_nl
      & butterFly_7_and_342_nl);
  xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_546_seb
      & butterFly_7_butterFly_7_or_62_rmff);
  butterFly_3_or_137_nl <= and_dcpl_470 OR (or_2189_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_1_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_137_nl);
  butterFly_3_or_70_nl <= (butterFly_3_butterFly_3_mux_1_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_103_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_201_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_134_nl <= (butterFly_3_mux1h_103_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_135_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_201_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_136_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_201_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_298_nl <= (butterFly_3_mux1h_136_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_0_0_i_adra_d <= butterFly_3_or_70_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_134_nl & butterFly_3_mux1h_135_nl
      & butterFly_3_or_298_nl;
  butterFly_3_or_456_cse <= and_dcpl_448 OR and_dcpl_475;
  butterFly_3_and_18_nl <= (NOT reg_modulo_add_11_slc_32_svs_st_cse) AND and_dcpl_459;
  butterFly_3_and_19_nl <= reg_modulo_add_11_slc_32_svs_st_cse AND and_dcpl_459;
  butterFly_3_mux1h_1_nl <= MUX1HOT_v_32_4_2(modulo_sub_3_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_19_qr_lpi_4_dfm, STD_LOGIC_VECTOR'(
      and_dcpl_479 & butterFly_3_and_18_nl & butterFly_3_and_19_nl & and_dcpl_480));
  butterFly_3_or_6_nl <= ((NOT reg_modulo_add_3_slc_32_svs_st_cse) AND and_dcpl_479)
      OR ((NOT reg_modulo_add_6_slc_32_svs_st_cse) AND and_dcpl_480);
  butterFly_3_or_7_nl <= (reg_modulo_add_3_slc_32_svs_st_cse AND and_dcpl_479) OR
      (reg_modulo_add_6_slc_32_svs_st_cse AND and_dcpl_480);
  butterFly_3_mux1h_39_nl <= MUX1HOT_v_32_5_2(reg_tmp_54_lpi_3_dfm_cse, tmp_55_lpi_3_dfm,
      modulo_add_base_1_sva, modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_11_qr_lpi_3_dfm,
      STD_LOGIC_VECTOR'( butterFly_3_or_456_cse & and_dcpl_450 & butterFly_3_or_6_nl
      & butterFly_3_or_7_nl & and_dcpl_459));
  yy_rsc_0_0_i_da_d_pff <= butterFly_3_mux1h_1_nl & butterFly_3_mux1h_39_nl;
  yy_rsc_0_0_i_wea_d <= STD_LOGIC_VECTOR'( and_587_seb & butterFly_7_butterFly_7_or_64_rmff);
  butterFly_7_or_nl <= ((NOT(or_dcpl_227 OR or_dcpl_225 OR (and_dcpl_490 AND and_dcpl_488)))
      AND mux_1880_seb) OR ((NOT mux_156_itm) AND and_dcpl_494 AND and_dcpl_492);
  butterFly_7_and_343_nl <= (NOT(or_2189_cse AND and_dcpl_503 AND and_dcpl_501))
      AND mux_1880_seb;
  yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_nl
      & butterFly_7_and_343_nl);
  yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_587_seb
      & butterFly_7_butterFly_7_or_64_rmff);
  butterFly_3_or_139_nl <= and_dcpl_511 OR (or_2245_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_3_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_139_nl);
  butterFly_3_or_68_nl <= (butterFly_3_butterFly_3_mux_3_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_101_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_203_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_132_nl <= (butterFly_3_mux1h_101_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_134_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_203_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_137_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_203_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_303_nl <= (butterFly_3_mux1h_137_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_1_0_i_adra_d <= butterFly_3_or_68_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_132_nl & butterFly_3_mux1h_134_nl
      & butterFly_3_or_303_nl;
  butterFly_3_and_12_nl <= (NOT reg_modulo_add_5_slc_32_svs_st_cse) AND and_dcpl_507;
  butterFly_3_and_13_nl <= reg_modulo_add_5_slc_32_svs_st_cse AND and_dcpl_507;
  butterFly_3_mux1h_3_nl <= MUX1HOT_v_32_4_2(modulo_sub_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_16_qr_lpi_4_dfm, STD_LOGIC_VECTOR'(
      and_615_ssc & butterFly_3_and_12_nl & butterFly_3_and_13_nl & and_616_ssc));
  butterFly_3_or_4_nl <= ((NOT reg_modulo_add_3_slc_32_svs_st_cse) AND and_615_ssc)
      OR ((NOT reg_modulo_add_2_slc_32_svs_st_cse) AND and_616_ssc);
  butterFly_3_or_5_nl <= (reg_modulo_add_3_slc_32_svs_st_cse AND and_615_ssc) OR
      (reg_modulo_add_2_slc_32_svs_st_cse AND and_616_ssc);
  butterFly_3_mux1h_38_nl <= MUX1HOT_v_32_5_2(reg_tmp_54_lpi_3_dfm_cse, tmp_55_lpi_3_dfm,
      modulo_add_base_1_sva, modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_8_qr_lpi_3_dfm,
      STD_LOGIC_VECTOR'( butterFly_3_or_456_cse & and_dcpl_450 & butterFly_3_or_4_nl
      & butterFly_3_or_5_nl & and_dcpl_507));
  yy_rsc_1_0_i_da_d_pff <= butterFly_3_mux1h_3_nl & butterFly_3_mux1h_38_nl;
  yy_rsc_1_0_i_wea_d <= STD_LOGIC_VECTOR'( and_618_seb & butterFly_7_butterFly_7_or_65_rmff);
  butterFly_7_or_1_nl <= ((NOT(or_dcpl_227 OR or_dcpl_229 OR (and_dcpl_490 AND and_dcpl_519)))
      AND mux_1932_seb) OR and_dcpl_525;
  butterFly_7_and_344_nl <= (NOT(or_2245_cse AND and_dcpl_503 AND and_dcpl_528))
      AND mux_1932_seb;
  yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_1_nl
      & butterFly_7_and_344_nl);
  yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_618_seb
      & butterFly_7_butterFly_7_or_65_rmff);
  butterFly_3_or_141_nl <= and_dcpl_537 OR (or_2294_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_5_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_141_nl);
  butterFly_3_or_66_nl <= (butterFly_3_butterFly_3_mux_5_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_99_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_205_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_130_nl <= (butterFly_3_mux1h_99_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_133_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_205_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_138_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_205_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_308_nl <= (butterFly_3_mux1h_138_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_2_0_i_adra_d <= butterFly_3_or_66_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_130_nl & butterFly_3_mux1h_133_nl
      & butterFly_3_or_308_nl;
  butterFly_3_and_6_nl <= (NOT reg_modulo_add_6_slc_32_svs_st_cse) AND and_dcpl_534;
  butterFly_3_and_7_nl <= reg_modulo_add_6_slc_32_svs_st_cse AND and_dcpl_534;
  butterFly_3_mux1h_5_nl <= MUX1HOT_v_32_4_2(modulo_sub_1_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_17_qr_lpi_4_dfm, STD_LOGIC_VECTOR'(
      and_dcpl_540 & butterFly_3_and_6_nl & butterFly_3_and_7_nl & and_dcpl_541));
  butterFly_3_or_2_nl <= ((NOT reg_modulo_add_1_slc_32_svs_st_cse) AND and_dcpl_540)
      OR ((NOT reg_modulo_add_11_slc_32_svs_st_cse) AND and_dcpl_541);
  butterFly_3_or_3_nl <= (reg_modulo_add_1_slc_32_svs_st_cse AND and_dcpl_540) OR
      (reg_modulo_add_11_slc_32_svs_st_cse AND and_dcpl_541);
  butterFly_3_mux1h_37_nl <= MUX1HOT_v_32_5_2(reg_tmp_54_lpi_3_dfm_cse, tmp_55_lpi_3_dfm,
      modulo_add_base_1_sva, modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_9_qr_lpi_3_dfm,
      STD_LOGIC_VECTOR'( butterFly_3_or_456_cse & and_dcpl_450 & butterFly_3_or_2_nl
      & butterFly_3_or_3_nl & and_dcpl_534));
  yy_rsc_2_0_i_da_d_pff <= butterFly_3_mux1h_5_nl & butterFly_3_mux1h_37_nl;
  yy_rsc_2_0_i_wea_d <= STD_LOGIC_VECTOR'( and_644_seb & butterFly_7_butterFly_7_or_66_rmff);
  butterFly_7_or_2_nl <= ((NOT(or_dcpl_227 OR or_dcpl_231 OR (and_dcpl_544 AND and_dcpl_488)))
      AND mux_1990_seb) OR and_dcpl_525;
  butterFly_7_and_345_nl <= (NOT(or_2294_cse AND and_dcpl_503 AND and_dcpl_548))
      AND mux_1990_seb;
  yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_2_nl
      & butterFly_7_and_345_nl);
  yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_644_seb
      & butterFly_7_butterFly_7_or_66_rmff);
  butterFly_3_or_143_nl <= and_dcpl_553 OR (or_2338_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_7_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_143_nl);
  butterFly_3_or_64_nl <= (butterFly_3_butterFly_3_mux_7_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_97_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_207_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_128_nl <= (butterFly_3_mux1h_97_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_132_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_207_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_139_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_207_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_313_nl <= (butterFly_3_mux1h_139_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_3_0_i_adra_d <= butterFly_3_or_64_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_128_nl & butterFly_3_mux1h_132_nl
      & butterFly_3_or_313_nl;
  butterFly_3_and_nl <= (NOT reg_modulo_add_1_slc_32_svs_st_cse) AND and_dcpl_552;
  butterFly_3_and_1_nl <= reg_modulo_add_1_slc_32_svs_st_cse AND and_dcpl_552;
  butterFly_3_mux1h_7_nl <= MUX1HOT_v_32_4_2(modulo_sub_2_qr_lpi_4_dfm, modulo_add_base_1_sva,
      modulo_add_3_qr_lpi_4_dfm_mx0w0, reg_modulo_sub_18_qr_lpi_4_dfm_cse, STD_LOGIC_VECTOR'(
      and_dcpl_556 & butterFly_3_and_nl & butterFly_3_and_1_nl & and_dcpl_557));
  butterFly_3_or_nl <= ((NOT reg_modulo_add_2_slc_32_svs_st_cse) AND and_dcpl_556)
      OR ((NOT reg_modulo_add_1_slc_32_svs_st_cse) AND and_dcpl_557);
  butterFly_3_or_1_nl <= (reg_modulo_add_2_slc_32_svs_st_cse AND and_dcpl_556) OR
      (reg_modulo_add_1_slc_32_svs_st_cse AND and_dcpl_557);
  butterFly_3_mux1h_36_nl <= MUX1HOT_v_32_5_2(reg_tmp_54_lpi_3_dfm_cse, tmp_55_lpi_3_dfm,
      modulo_add_base_1_sva, modulo_add_3_qr_lpi_4_dfm_mx0w0, modulo_sub_10_qr_lpi_3_dfm,
      STD_LOGIC_VECTOR'( butterFly_3_or_456_cse & and_dcpl_450 & butterFly_3_or_nl
      & butterFly_3_or_1_nl & and_dcpl_552));
  yy_rsc_3_0_i_da_d_pff <= butterFly_3_mux1h_7_nl & butterFly_3_mux1h_36_nl;
  yy_rsc_3_0_i_wea_d <= STD_LOGIC_VECTOR'( and_662_seb & butterFly_7_butterFly_7_or_67_rmff);
  butterFly_7_or_3_nl <= ((NOT(or_dcpl_227 OR or_dcpl_233 OR (and_dcpl_544 AND and_dcpl_519)))
      AND mux_2051_seb) OR and_dcpl_525;
  butterFly_7_and_346_nl <= (NOT(or_2338_cse AND and_dcpl_503 AND and_dcpl_564))
      AND mux_2051_seb;
  yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_3_nl
      & butterFly_7_and_346_nl);
  yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_662_seb
      & butterFly_7_butterFly_7_or_67_rmff);
  butterFly_3_or_145_nl <= and_dcpl_570 OR (or_2386_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_9_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_145_nl);
  butterFly_3_or_62_nl <= (butterFly_3_butterFly_3_mux_9_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_95_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_209_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_126_nl <= (butterFly_3_mux1h_95_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_131_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_209_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_140_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_209_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_318_nl <= (butterFly_3_mux1h_140_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_4_0_i_adra_d <= butterFly_3_or_62_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_126_nl & butterFly_3_mux1h_131_nl
      & butterFly_3_or_318_nl;
  yy_rsc_4_0_i_wea_d <= STD_LOGIC_VECTOR'( and_677_seb & butterFly_7_butterFly_7_or_68_rmff);
  butterFly_7_or_4_nl <= ((NOT(or_dcpl_236 OR or_dcpl_225 OR (and_dcpl_578 AND and_dcpl_488)))
      AND mux_2108_seb) OR ((NOT mux_156_itm) AND and_dcpl_581 AND and_dcpl_492);
  butterFly_7_and_347_nl <= (NOT(or_2386_cse AND and_dcpl_585 AND and_dcpl_501))
      AND mux_2108_seb;
  yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_4_nl
      & butterFly_7_and_347_nl);
  yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_677_seb
      & butterFly_7_butterFly_7_or_68_rmff);
  butterFly_3_or_147_nl <= and_dcpl_588 OR (or_2440_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_11_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_147_nl);
  butterFly_3_or_60_nl <= (butterFly_3_butterFly_3_mux_11_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_93_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_211_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_124_nl <= (butterFly_3_mux1h_93_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_130_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_211_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_141_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_211_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_323_nl <= (butterFly_3_mux1h_141_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_5_0_i_adra_d <= butterFly_3_or_60_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_124_nl & butterFly_3_mux1h_130_nl
      & butterFly_3_or_323_nl;
  yy_rsc_5_0_i_wea_d <= STD_LOGIC_VECTOR'( and_693_seb & butterFly_7_butterFly_7_or_69_rmff);
  butterFly_7_or_5_nl <= ((NOT(or_dcpl_236 OR or_dcpl_229 OR (and_dcpl_578 AND and_dcpl_519)))
      AND mux_2157_seb) OR and_dcpl_596;
  butterFly_7_and_348_nl <= (NOT(or_2440_cse AND and_dcpl_585 AND and_dcpl_528))
      AND mux_2157_seb;
  yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_5_nl
      & butterFly_7_and_348_nl);
  yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_693_seb
      & butterFly_7_butterFly_7_or_69_rmff);
  butterFly_3_or_149_nl <= and_dcpl_600 OR (or_2487_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_13_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_149_nl);
  butterFly_3_or_58_nl <= (butterFly_3_butterFly_3_mux_13_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_91_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_213_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_122_nl <= (butterFly_3_mux1h_91_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_129_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_213_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_142_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_213_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_328_nl <= (butterFly_3_mux1h_142_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_6_0_i_adra_d <= butterFly_3_or_58_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_122_nl & butterFly_3_mux1h_129_nl
      & butterFly_3_or_328_nl;
  yy_rsc_6_0_i_wea_d <= STD_LOGIC_VECTOR'( and_705_seb & butterFly_7_butterFly_7_or_70_rmff);
  butterFly_7_or_6_nl <= ((NOT(or_dcpl_236 OR or_dcpl_231 OR (and_dcpl_605 AND and_dcpl_488)))
      AND mux_2213_seb) OR and_dcpl_596;
  butterFly_7_and_349_nl <= (NOT(or_2487_cse AND and_dcpl_585 AND and_dcpl_548))
      AND mux_2213_seb;
  yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_6_nl
      & butterFly_7_and_349_nl);
  yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_705_seb
      & butterFly_7_butterFly_7_or_70_rmff);
  butterFly_3_or_151_nl <= and_dcpl_609 OR (or_2528_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_15_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_151_nl);
  butterFly_3_or_56_nl <= (butterFly_3_butterFly_3_mux_15_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_89_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_215_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_120_nl <= (butterFly_3_mux1h_89_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_128_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_215_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_143_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_215_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_333_nl <= (butterFly_3_mux1h_143_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_7_0_i_adra_d <= butterFly_3_or_56_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_120_nl & butterFly_3_mux1h_128_nl
      & butterFly_3_or_333_nl;
  yy_rsc_7_0_i_wea_d <= STD_LOGIC_VECTOR'( and_716_seb & butterFly_7_butterFly_7_or_71_rmff);
  butterFly_7_or_7_nl <= ((NOT(or_dcpl_236 OR or_dcpl_233 OR (and_dcpl_605 AND and_dcpl_519)))
      AND mux_2271_seb) OR and_dcpl_596;
  butterFly_7_and_350_nl <= (NOT(or_2528_cse AND and_dcpl_585 AND and_dcpl_564))
      AND mux_2271_seb;
  yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_7_nl
      & butterFly_7_and_350_nl);
  yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_716_seb
      & butterFly_7_butterFly_7_or_71_rmff);
  butterFly_3_or_153_nl <= and_dcpl_622 OR (or_2577_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_17_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_153_nl);
  butterFly_3_or_54_nl <= (butterFly_3_butterFly_3_mux_17_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_87_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_217_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_118_nl <= (butterFly_3_mux1h_87_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_127_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_217_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_144_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_217_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_338_nl <= (butterFly_3_mux1h_144_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_8_0_i_adra_d <= butterFly_3_or_54_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_118_nl & butterFly_3_mux1h_127_nl
      & butterFly_3_or_338_nl;
  yy_rsc_8_0_i_wea_d <= STD_LOGIC_VECTOR'( and_729_seb & butterFly_7_butterFly_7_or_72_rmff);
  butterFly_7_or_8_nl <= ((NOT(or_dcpl_241 OR or_dcpl_225 OR (and_dcpl_629 AND and_dcpl_488)))
      AND mux_2328_seb) OR ((NOT mux_156_itm) AND and_dcpl_494 AND and_dcpl_631);
  butterFly_7_and_351_nl <= (NOT(or_2577_cse AND and_dcpl_503 AND and_dcpl_637))
      AND mux_2328_seb;
  yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_8_nl
      & butterFly_7_and_351_nl);
  yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_729_seb
      & butterFly_7_butterFly_7_or_72_rmff);
  butterFly_3_or_155_nl <= and_dcpl_640 OR (or_2622_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_19_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_155_nl);
  butterFly_3_or_52_nl <= (butterFly_3_butterFly_3_mux_19_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_85_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_219_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_116_nl <= (butterFly_3_mux1h_85_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_126_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_219_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_145_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_219_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_343_nl <= (butterFly_3_mux1h_145_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_9_0_i_adra_d <= butterFly_3_or_52_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_116_nl & butterFly_3_mux1h_126_nl
      & butterFly_3_or_343_nl;
  yy_rsc_9_0_i_wea_d <= STD_LOGIC_VECTOR'( and_745_seb & butterFly_7_butterFly_7_or_73_rmff);
  butterFly_7_or_9_nl <= ((NOT(or_dcpl_241 OR or_dcpl_229 OR (and_dcpl_629 AND and_dcpl_519)))
      AND mux_2377_seb) OR and_dcpl_648;
  butterFly_7_and_352_nl <= (NOT(or_2622_cse AND and_dcpl_503 AND and_dcpl_650))
      AND mux_2377_seb;
  yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_9_nl
      & butterFly_7_and_352_nl);
  yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_745_seb
      & butterFly_7_butterFly_7_or_73_rmff);
  butterFly_3_or_157_nl <= and_dcpl_655 OR (or_2664_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_21_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_157_nl);
  butterFly_3_or_50_nl <= (butterFly_3_butterFly_3_mux_21_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_83_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_221_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_114_nl <= (butterFly_3_mux1h_83_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_125_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_221_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_146_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_221_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_348_nl <= (butterFly_3_mux1h_146_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_10_0_i_adra_d <= butterFly_3_or_50_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_114_nl & butterFly_3_mux1h_125_nl
      & butterFly_3_or_348_nl;
  yy_rsc_10_0_i_wea_d <= STD_LOGIC_VECTOR'( and_760_seb & butterFly_7_butterFly_7_or_74_rmff);
  butterFly_7_or_10_nl <= ((NOT(or_dcpl_241 OR or_dcpl_231 OR (and_dcpl_660 AND and_dcpl_488)))
      AND mux_2433_seb) OR and_dcpl_648;
  butterFly_7_and_353_nl <= (NOT(or_2664_cse AND and_dcpl_503 AND and_dcpl_664))
      AND mux_2433_seb;
  yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_10_nl
      & butterFly_7_and_353_nl);
  yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_760_seb
      & butterFly_7_butterFly_7_or_74_rmff);
  butterFly_3_or_159_nl <= and_dcpl_667 OR (or_2700_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_23_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_159_nl);
  butterFly_3_or_48_nl <= (butterFly_3_butterFly_3_mux_23_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_81_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_223_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_112_nl <= (butterFly_3_mux1h_81_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_124_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_223_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_147_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_223_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_353_nl <= (butterFly_3_mux1h_147_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_11_0_i_adra_d <= butterFly_3_or_48_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_112_nl & butterFly_3_mux1h_124_nl
      & butterFly_3_or_353_nl;
  yy_rsc_11_0_i_wea_d <= STD_LOGIC_VECTOR'( and_773_seb & butterFly_7_butterFly_7_or_75_rmff);
  butterFly_7_or_11_nl <= ((NOT(or_dcpl_241 OR or_dcpl_233 OR (and_dcpl_660 AND and_dcpl_519)))
      AND mux_2491_seb) OR and_dcpl_648;
  butterFly_7_and_354_nl <= (NOT(or_2700_cse AND and_dcpl_503 AND and_dcpl_675))
      AND mux_2491_seb;
  yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_11_nl
      & butterFly_7_and_354_nl);
  yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_773_seb
      & butterFly_7_butterFly_7_or_75_rmff);
  butterFly_3_or_161_nl <= and_dcpl_679 OR (or_2747_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_25_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_161_nl);
  butterFly_3_or_46_nl <= (butterFly_3_butterFly_3_mux_25_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_79_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_225_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_110_nl <= (butterFly_3_mux1h_79_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_123_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_225_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_148_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_225_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_358_nl <= (butterFly_3_mux1h_148_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_12_0_i_adra_d <= butterFly_3_or_46_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_110_nl & butterFly_3_mux1h_123_nl
      & butterFly_3_or_358_nl;
  yy_rsc_12_0_i_wea_d <= STD_LOGIC_VECTOR'( and_786_seb & butterFly_7_butterFly_7_or_76_rmff);
  butterFly_7_or_12_nl <= ((NOT(or_dcpl_246 OR or_dcpl_225 OR (and_dcpl_686 AND and_dcpl_488)))
      AND mux_2548_seb) OR ((NOT mux_156_itm) AND and_dcpl_581 AND and_dcpl_631);
  butterFly_7_and_355_nl <= (NOT(or_2747_cse AND and_dcpl_585 AND and_dcpl_637))
      AND mux_2548_seb;
  yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_12_nl
      & butterFly_7_and_355_nl);
  yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_786_seb
      & butterFly_7_butterFly_7_or_76_rmff);
  butterFly_3_or_163_nl <= and_dcpl_692 OR (or_2800_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_27_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_163_nl);
  butterFly_3_or_44_nl <= (butterFly_3_butterFly_3_mux_27_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_77_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_227_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_108_nl <= (butterFly_3_mux1h_77_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_122_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_227_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_149_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_227_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_363_nl <= (butterFly_3_mux1h_149_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_13_0_i_adra_d <= butterFly_3_or_44_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_108_nl & butterFly_3_mux1h_122_nl
      & butterFly_3_or_363_nl;
  yy_rsc_13_0_i_wea_d <= STD_LOGIC_VECTOR'( and_797_seb & butterFly_7_butterFly_7_or_77_rmff);
  butterFly_7_or_13_nl <= ((NOT(or_dcpl_246 OR or_dcpl_229 OR (and_dcpl_686 AND and_dcpl_519)))
      AND mux_2597_seb) OR and_dcpl_699;
  butterFly_7_and_356_nl <= (NOT(or_2800_cse AND and_dcpl_585 AND and_dcpl_650))
      AND mux_2597_seb;
  yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_13_nl
      & butterFly_7_and_356_nl);
  yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_797_seb
      & butterFly_7_butterFly_7_or_77_rmff);
  butterFly_3_or_165_nl <= and_dcpl_703 OR (or_2847_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_29_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_165_nl);
  butterFly_3_or_42_nl <= (butterFly_3_butterFly_3_mux_29_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_75_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_229_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_106_nl <= (butterFly_3_mux1h_75_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_121_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_229_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_150_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_229_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_368_nl <= (butterFly_3_mux1h_150_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_14_0_i_adra_d <= butterFly_3_or_42_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_106_nl & butterFly_3_mux1h_121_nl
      & butterFly_3_or_368_nl;
  yy_rsc_14_0_i_wea_d <= STD_LOGIC_VECTOR'( and_808_seb & butterFly_7_butterFly_7_or_78_rmff);
  butterFly_7_or_14_nl <= ((NOT(or_dcpl_246 OR or_dcpl_231 OR (and_dcpl_708 AND and_dcpl_488)))
      AND mux_2653_seb) OR and_dcpl_699;
  butterFly_7_and_357_nl <= (NOT(or_2847_cse AND and_dcpl_585 AND and_dcpl_664))
      AND mux_2653_seb;
  yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_14_nl
      & butterFly_7_and_357_nl);
  yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_808_seb
      & butterFly_7_butterFly_7_or_78_rmff);
  butterFly_3_or_167_nl <= and_dcpl_712 OR (nand_317_cse AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_31_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_167_nl);
  butterFly_3_or_40_nl <= (butterFly_3_butterFly_3_mux_31_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_73_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_231_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_104_nl <= (butterFly_3_mux1h_73_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_120_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_231_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_151_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_231_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_373_nl <= (butterFly_3_mux1h_151_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_15_0_i_adra_d <= butterFly_3_or_40_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_104_nl & butterFly_3_mux1h_120_nl
      & butterFly_3_or_373_nl;
  yy_rsc_15_0_i_wea_d <= STD_LOGIC_VECTOR'( and_818_seb & butterFly_7_butterFly_7_or_79_rmff);
  butterFly_7_or_15_nl <= ((NOT(or_dcpl_246 OR or_dcpl_233 OR (and_dcpl_708 AND and_dcpl_519)))
      AND mux_2711_seb) OR and_dcpl_699;
  butterFly_7_and_358_nl <= (NOT(nand_317_cse AND and_dcpl_585 AND and_dcpl_675))
      AND mux_2711_seb;
  yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_15_nl
      & butterFly_7_and_358_nl);
  yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_818_seb
      & butterFly_7_butterFly_7_or_79_rmff);
  butterFly_3_or_169_nl <= and_dcpl_724 OR (or_tmp_1079 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_33_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_169_nl);
  butterFly_3_or_38_nl <= (butterFly_3_butterFly_3_mux_33_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_71_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_233_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_102_nl <= (butterFly_3_mux1h_71_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_119_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_233_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_152_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_233_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_378_nl <= (butterFly_3_mux1h_152_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_16_0_i_adra_d <= butterFly_3_or_38_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_102_nl & butterFly_3_mux1h_119_nl
      & butterFly_3_or_378_nl;
  yy_rsc_16_0_i_wea_d <= STD_LOGIC_VECTOR'( and_831_seb & butterFly_7_butterFly_7_or_80_rmff);
  butterFly_7_or_16_nl <= ((NOT(or_dcpl_252 OR or_dcpl_225 OR (and_dcpl_731 AND and_dcpl_488)))
      AND mux_2768_seb) OR ((NOT mux_156_itm) AND and_dcpl_733 AND and_dcpl_492);
  butterFly_7_and_359_nl <= (NOT(or_tmp_1079 AND and_dcpl_503 AND and_dcpl_739))
      AND mux_2768_seb;
  yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_16_nl
      & butterFly_7_and_359_nl);
  yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_831_seb
      & butterFly_7_butterFly_7_or_80_rmff);
  butterFly_3_or_171_nl <= and_dcpl_742 OR (or_tmp_1133 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_35_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_171_nl);
  butterFly_3_or_36_nl <= (butterFly_3_butterFly_3_mux_35_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_69_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_235_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_100_nl <= (butterFly_3_mux1h_69_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_118_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_235_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_153_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_235_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_383_nl <= (butterFly_3_mux1h_153_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_17_0_i_adra_d <= butterFly_3_or_36_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_100_nl & butterFly_3_mux1h_118_nl
      & butterFly_3_or_383_nl;
  yy_rsc_17_0_i_wea_d <= STD_LOGIC_VECTOR'( and_847_seb & butterFly_7_butterFly_7_or_81_rmff);
  butterFly_7_or_17_nl <= ((NOT(or_dcpl_252 OR or_dcpl_229 OR (and_dcpl_731 AND and_dcpl_519)))
      AND mux_2817_seb) OR and_dcpl_751;
  butterFly_7_and_360_nl <= (NOT(or_tmp_1133 AND and_dcpl_503 AND and_dcpl_753))
      AND mux_2817_seb;
  yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_17_nl
      & butterFly_7_and_360_nl);
  yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_847_seb
      & butterFly_7_butterFly_7_or_81_rmff);
  butterFly_3_or_173_nl <= and_dcpl_758 OR (or_tmp_1185 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_37_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_173_nl);
  butterFly_3_or_34_nl <= (butterFly_3_butterFly_3_mux_37_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_67_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_237_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_98_nl <= (butterFly_3_mux1h_67_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_117_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_237_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_154_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_237_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_388_nl <= (butterFly_3_mux1h_154_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_18_0_i_adra_d <= butterFly_3_or_34_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_98_nl & butterFly_3_mux1h_117_nl
      & butterFly_3_or_388_nl;
  yy_rsc_18_0_i_wea_d <= STD_LOGIC_VECTOR'( and_863_seb & butterFly_7_butterFly_7_or_82_rmff);
  butterFly_7_or_18_nl <= ((NOT(or_dcpl_252 OR or_dcpl_231 OR (and_dcpl_763 AND and_dcpl_488)))
      AND mux_2873_seb) OR and_dcpl_751;
  butterFly_7_and_361_nl <= (NOT(or_tmp_1185 AND and_dcpl_503 AND and_dcpl_767))
      AND mux_2873_seb;
  yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_18_nl
      & butterFly_7_and_361_nl);
  yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_863_seb
      & butterFly_7_butterFly_7_or_82_rmff);
  butterFly_3_or_175_nl <= and_dcpl_770 OR (or_tmp_1235 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_39_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_175_nl);
  butterFly_3_or_32_nl <= (butterFly_3_butterFly_3_mux_39_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_65_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_239_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_96_nl <= (butterFly_3_mux1h_65_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_116_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_239_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_155_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_239_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_393_nl <= (butterFly_3_mux1h_155_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_19_0_i_adra_d <= butterFly_3_or_32_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_96_nl & butterFly_3_mux1h_116_nl
      & butterFly_3_or_393_nl;
  yy_rsc_19_0_i_wea_d <= STD_LOGIC_VECTOR'( and_876_seb & butterFly_7_butterFly_7_or_83_rmff);
  butterFly_7_or_19_nl <= ((NOT(or_dcpl_252 OR or_dcpl_233 OR (and_dcpl_763 AND and_dcpl_519)))
      AND mux_2931_seb) OR and_dcpl_751;
  butterFly_7_and_362_nl <= (NOT(or_tmp_1235 AND and_dcpl_503 AND and_dcpl_778))
      AND mux_2931_seb;
  yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_19_nl
      & butterFly_7_and_362_nl);
  yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_876_seb
      & butterFly_7_butterFly_7_or_83_rmff);
  butterFly_3_or_177_nl <= and_dcpl_782 OR (or_tmp_1298 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_41_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_177_nl);
  butterFly_3_or_30_nl <= (butterFly_3_butterFly_3_mux_41_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_63_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_241_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_94_nl <= (butterFly_3_mux1h_63_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_115_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_241_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_156_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_241_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_398_nl <= (butterFly_3_mux1h_156_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_20_0_i_adra_d <= butterFly_3_or_30_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_94_nl & butterFly_3_mux1h_115_nl
      & butterFly_3_or_398_nl;
  yy_rsc_20_0_i_wea_d <= STD_LOGIC_VECTOR'( and_888_seb & butterFly_7_butterFly_7_or_84_rmff);
  butterFly_7_or_20_nl <= ((NOT(or_dcpl_258 OR or_dcpl_225 OR (and_dcpl_788 AND and_dcpl_488)))
      AND mux_2988_seb) OR ((NOT mux_156_itm) AND and_dcpl_790 AND and_dcpl_492);
  butterFly_7_and_363_nl <= (NOT(or_tmp_1298 AND and_dcpl_585 AND and_dcpl_739))
      AND mux_2988_seb;
  yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_20_nl
      & butterFly_7_and_363_nl);
  yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_888_seb
      & butterFly_7_butterFly_7_or_84_rmff);
  butterFly_3_or_179_nl <= and_dcpl_795 OR (or_tmp_1363 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_43_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_179_nl);
  butterFly_3_or_28_nl <= (butterFly_3_butterFly_3_mux_43_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_61_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_243_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_92_nl <= (butterFly_3_mux1h_61_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_114_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_243_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_157_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_243_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_403_nl <= (butterFly_3_mux1h_157_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_21_0_i_adra_d <= butterFly_3_or_28_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_92_nl & butterFly_3_mux1h_114_nl
      & butterFly_3_or_403_nl;
  yy_rsc_21_0_i_wea_d <= STD_LOGIC_VECTOR'( and_900_seb & butterFly_7_butterFly_7_or_85_rmff);
  butterFly_7_or_21_nl <= ((NOT(or_dcpl_258 OR or_dcpl_229 OR (and_dcpl_788 AND and_dcpl_519)))
      AND mux_3037_seb) OR and_dcpl_802;
  butterFly_7_and_364_nl <= (NOT(or_tmp_1363 AND and_dcpl_585 AND and_dcpl_753))
      AND mux_3037_seb;
  yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_21_nl
      & butterFly_7_and_364_nl);
  yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_900_seb
      & butterFly_7_butterFly_7_or_85_rmff);
  butterFly_3_or_181_nl <= and_dcpl_806 OR (or_tmp_1422 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_45_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_181_nl);
  butterFly_3_or_26_nl <= (butterFly_3_butterFly_3_mux_45_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_59_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_245_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_90_nl <= (butterFly_3_mux1h_59_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_113_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_245_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_158_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_245_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_408_nl <= (butterFly_3_mux1h_158_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_22_0_i_adra_d <= butterFly_3_or_26_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_90_nl & butterFly_3_mux1h_113_nl
      & butterFly_3_or_408_nl;
  yy_rsc_22_0_i_wea_d <= STD_LOGIC_VECTOR'( and_911_seb & butterFly_7_butterFly_7_or_86_rmff);
  butterFly_7_or_22_nl <= ((NOT(or_dcpl_258 OR or_dcpl_231 OR (and_dcpl_811 AND and_dcpl_488)))
      AND mux_3093_seb) OR and_dcpl_802;
  butterFly_7_and_365_nl <= (NOT(or_tmp_1422 AND and_dcpl_585 AND and_dcpl_767))
      AND mux_3093_seb;
  yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_22_nl
      & butterFly_7_and_365_nl);
  yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_911_seb
      & butterFly_7_butterFly_7_or_86_rmff);
  butterFly_3_or_183_nl <= and_dcpl_815 OR (or_tmp_1479 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_47_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_183_nl);
  butterFly_3_or_24_nl <= (butterFly_3_butterFly_3_mux_47_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_57_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_247_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_88_nl <= (butterFly_3_mux1h_57_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_112_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_247_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_159_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_247_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_413_nl <= (butterFly_3_mux1h_159_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_23_0_i_adra_d <= butterFly_3_or_24_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_88_nl & butterFly_3_mux1h_112_nl
      & butterFly_3_or_413_nl;
  yy_rsc_23_0_i_wea_d <= STD_LOGIC_VECTOR'( and_921_seb & butterFly_7_butterFly_7_or_87_rmff);
  butterFly_7_or_23_nl <= ((NOT(or_dcpl_258 OR or_dcpl_233 OR (and_dcpl_811 AND and_dcpl_519)))
      AND mux_3151_seb) OR and_dcpl_802;
  butterFly_7_and_366_nl <= (NOT(or_tmp_1479 AND and_dcpl_585 AND and_dcpl_778))
      AND mux_3151_seb;
  yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_23_nl
      & butterFly_7_and_366_nl);
  yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_921_seb
      & butterFly_7_butterFly_7_or_87_rmff);
  butterFly_3_or_185_nl <= and_dcpl_827 OR (or_tmp_1540 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_49_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_185_nl);
  butterFly_3_or_22_nl <= (butterFly_3_butterFly_3_mux_49_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_55_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_249_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_86_nl <= (butterFly_3_mux1h_55_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_111_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_249_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_160_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_249_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_418_nl <= (butterFly_3_mux1h_160_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_24_0_i_adra_d <= butterFly_3_or_22_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_86_nl & butterFly_3_mux1h_111_nl
      & butterFly_3_or_418_nl;
  yy_rsc_24_0_i_wea_d <= STD_LOGIC_VECTOR'( and_933_seb & butterFly_7_butterFly_7_or_88_rmff);
  butterFly_7_or_24_nl <= ((NOT(or_dcpl_263 OR or_dcpl_225 OR (and_dcpl_833 AND and_dcpl_488)))
      AND mux_3208_seb) OR ((NOT mux_156_itm) AND and_dcpl_733 AND and_dcpl_631);
  butterFly_7_and_367_nl <= (NOT(or_tmp_1540 AND and_dcpl_503 AND and_dcpl_840))
      AND mux_3208_seb;
  yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_24_nl
      & butterFly_7_and_367_nl);
  yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_933_seb
      & butterFly_7_butterFly_7_or_88_rmff);
  butterFly_3_or_187_nl <= and_dcpl_843 OR (or_tmp_1595 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_51_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_187_nl);
  butterFly_3_or_20_nl <= (butterFly_3_butterFly_3_mux_51_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_53_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_251_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_84_nl <= (butterFly_3_mux1h_53_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_110_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_251_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_161_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_251_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_423_nl <= (butterFly_3_mux1h_161_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_25_0_i_adra_d <= butterFly_3_or_20_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_84_nl & butterFly_3_mux1h_110_nl
      & butterFly_3_or_423_nl;
  yy_rsc_25_0_i_wea_d <= STD_LOGIC_VECTOR'( and_948_seb & butterFly_7_butterFly_7_or_89_rmff);
  butterFly_7_or_25_nl <= ((NOT(or_dcpl_263 OR or_dcpl_229 OR (and_dcpl_833 AND and_dcpl_519)))
      AND mux_3257_seb) OR and_dcpl_851;
  butterFly_7_and_368_nl <= (NOT(or_tmp_1595 AND and_dcpl_503 AND and_dcpl_853))
      AND mux_3257_seb;
  yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_25_nl
      & butterFly_7_and_368_nl);
  yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_948_seb
      & butterFly_7_butterFly_7_or_89_rmff);
  butterFly_3_or_189_nl <= and_dcpl_858 OR (or_tmp_1647 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_53_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_189_nl);
  butterFly_3_or_18_nl <= (butterFly_3_butterFly_3_mux_53_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_51_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_253_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_82_nl <= (butterFly_3_mux1h_51_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_109_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_253_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_162_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_253_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_428_nl <= (butterFly_3_mux1h_162_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_26_0_i_adra_d <= butterFly_3_or_18_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_82_nl & butterFly_3_mux1h_109_nl
      & butterFly_3_or_428_nl;
  yy_rsc_26_0_i_wea_d <= STD_LOGIC_VECTOR'( and_963_seb & butterFly_7_butterFly_7_or_90_rmff);
  butterFly_7_or_26_nl <= ((NOT(or_dcpl_263 OR or_dcpl_231 OR (and_dcpl_863 AND and_dcpl_488)))
      AND mux_3313_seb) OR and_dcpl_851;
  butterFly_7_and_369_nl <= (NOT(or_tmp_1647 AND and_dcpl_503 AND and_dcpl_867))
      AND mux_3313_seb;
  yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_26_nl
      & butterFly_7_and_369_nl);
  yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_963_seb
      & butterFly_7_butterFly_7_or_90_rmff);
  butterFly_3_or_191_nl <= and_dcpl_870 OR (or_tmp_1703 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_55_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_191_nl);
  butterFly_3_or_16_nl <= (butterFly_3_butterFly_3_mux_55_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_49_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_255_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_80_nl <= (butterFly_3_mux1h_49_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_108_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_255_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_163_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_255_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_433_nl <= (butterFly_3_mux1h_163_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_27_0_i_adra_d <= butterFly_3_or_16_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_80_nl & butterFly_3_mux1h_108_nl
      & butterFly_3_or_433_nl;
  yy_rsc_27_0_i_wea_d <= STD_LOGIC_VECTOR'( and_976_seb & butterFly_7_butterFly_7_or_91_rmff);
  butterFly_7_or_27_nl <= ((NOT(or_dcpl_263 OR or_dcpl_233 OR (and_dcpl_863 AND and_dcpl_519)))
      AND mux_3371_seb) OR and_dcpl_851;
  butterFly_7_and_370_nl <= (NOT(or_tmp_1703 AND and_dcpl_503 AND and_dcpl_878))
      AND mux_3371_seb;
  yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_27_nl
      & butterFly_7_and_370_nl);
  yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_976_seb
      & butterFly_7_butterFly_7_or_91_rmff);
  butterFly_3_or_193_nl <= and_dcpl_882 OR (or_tmp_1765 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_57_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_193_nl);
  butterFly_3_or_14_nl <= (butterFly_3_butterFly_3_mux_57_nl AND (NOT and_dcpl_459))
      OR and_dcpl_454;
  butterFly_3_mux1h_47_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_257_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_78_nl <= (butterFly_3_mux1h_47_nl AND (NOT and_dcpl_454)) OR and_dcpl_459;
  butterFly_3_mux1h_107_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse & butterFly_3_or_257_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_164_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_296_cse
      & butterFly_3_or_257_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_438_nl <= (butterFly_3_mux1h_164_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_28_0_i_adra_d <= butterFly_3_or_14_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_78_nl & butterFly_3_mux1h_107_nl
      & butterFly_3_or_438_nl;
  yy_rsc_28_0_i_wea_d <= STD_LOGIC_VECTOR'( and_988_seb & butterFly_7_butterFly_7_or_92_rmff);
  butterFly_7_or_28_nl <= ((NOT(or_dcpl_268 OR or_dcpl_225 OR (and_dcpl_888 AND and_dcpl_488)))
      AND mux_3428_seb) OR ((NOT mux_156_itm) AND and_dcpl_790 AND and_dcpl_631);
  butterFly_7_and_371_nl <= (NOT(or_tmp_1765 AND and_dcpl_585 AND and_dcpl_840))
      AND mux_3428_seb;
  yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_28_nl
      & butterFly_7_and_371_nl);
  yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_988_seb
      & butterFly_7_butterFly_7_or_92_rmff);
  butterFly_3_or_195_nl <= and_dcpl_894 OR (or_tmp_1818 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_59_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_195_nl);
  butterFly_3_or_12_nl <= (butterFly_3_butterFly_3_mux_59_nl AND (NOT and_dcpl_507))
      OR and_dcpl_506;
  butterFly_3_mux1h_45_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_259_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_76_nl <= (butterFly_3_mux1h_45_nl AND (NOT and_dcpl_506)) OR and_dcpl_507;
  butterFly_3_mux1h_106_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse & butterFly_3_or_259_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_165_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_301_cse
      & butterFly_3_or_259_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_443_nl <= (butterFly_3_mux1h_165_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_29_0_i_adra_d <= butterFly_3_or_12_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_76_nl & butterFly_3_mux1h_106_nl
      & butterFly_3_or_443_nl;
  yy_rsc_29_0_i_wea_d <= STD_LOGIC_VECTOR'( and_1000_seb & butterFly_7_butterFly_7_or_93_rmff);
  butterFly_7_or_29_nl <= ((NOT(or_dcpl_268 OR or_dcpl_229 OR (and_dcpl_888 AND and_dcpl_519)))
      AND mux_3477_seb) OR and_dcpl_901;
  butterFly_7_and_372_nl <= (NOT(or_tmp_1818 AND and_dcpl_585 AND and_dcpl_853))
      AND mux_3477_seb;
  yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_29_nl
      & butterFly_7_and_372_nl);
  yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_1000_seb
      & butterFly_7_butterFly_7_or_93_rmff);
  butterFly_3_or_197_nl <= and_dcpl_905 OR (or_tmp_1867 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_61_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_197_nl);
  butterFly_3_or_10_nl <= (butterFly_3_butterFly_3_mux_61_nl AND (NOT and_dcpl_534))
      OR and_dcpl_533;
  butterFly_3_mux1h_43_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_261_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_74_nl <= (butterFly_3_mux1h_43_nl AND (NOT and_dcpl_533)) OR and_dcpl_534;
  butterFly_3_mux1h_105_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse & butterFly_3_or_261_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_166_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_306_cse
      & butterFly_3_or_261_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_448_nl <= (butterFly_3_mux1h_166_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_30_0_i_adra_d <= butterFly_3_or_10_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_74_nl & butterFly_3_mux1h_105_nl
      & butterFly_3_or_448_nl;
  yy_rsc_30_0_i_wea_d <= STD_LOGIC_VECTOR'( and_1011_seb & butterFly_7_butterFly_7_or_94_rmff);
  butterFly_7_or_30_nl <= ((NOT(or_dcpl_268 OR or_dcpl_231 OR (and_dcpl_910 AND and_dcpl_488)))
      AND mux_3533_seb) OR and_dcpl_901;
  butterFly_7_and_373_nl <= (NOT(or_tmp_1867 AND and_dcpl_585 AND and_dcpl_867))
      AND mux_3533_seb;
  yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_30_nl
      & butterFly_7_and_373_nl);
  yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_1011_seb
      & butterFly_7_butterFly_7_or_94_rmff);
  butterFly_3_or_199_nl <= and_dcpl_914 OR (or_dcpl_273 AND and_dcpl_91 AND and_dcpl_472);
  butterFly_3_butterFly_3_mux_63_nl <= MUX_s_1_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg, butterFly_3_or_199_nl);
  butterFly_3_or_8_nl <= (butterFly_3_butterFly_3_mux_63_nl AND (NOT and_dcpl_552))
      OR and_dcpl_551;
  butterFly_3_mux1h_41_nl <= MUX1HOT_s_1_5_2(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)), S1_OUTER_LOOP_for_acc_svs_4, (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)),
      (reg_drf_revArr_ptr_1_smx_9_0_reg(1)), STD_LOGIC_VECTOR'( and_dcpl_448 & butterFly_3_or_263_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_or_72_nl <= (butterFly_3_mux1h_41_nl AND (NOT and_dcpl_551)) OR and_dcpl_552;
  butterFly_3_mux1h_104_nl <= MUX1HOT_v_3_5_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)), ((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) & (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1))), (S1_OUTER_LOOP_for_acc_svs_3_0(3 DOWNTO 1)), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)), ((reg_drf_revArr_ptr_1_smx_9_0_reg(0)) & (reg_drf_revArr_ptr_1_smx_9_0_1_reg(2
      DOWNTO 1))), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse & butterFly_3_or_263_cse
      & and_dcpl_451 & butterFly_3_or_264_cse & and_dcpl_475));
  butterFly_3_mux1h_167_nl <= MUX1HOT_s_1_4_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)),
      (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)), (S1_OUTER_LOOP_for_acc_svs_3_0(0)),
      (reg_drf_revArr_ptr_1_smx_9_0_1_reg(0)), STD_LOGIC_VECTOR'( butterFly_3_or_311_cse
      & butterFly_3_or_263_cse & and_dcpl_451 & and_dcpl_475));
  butterFly_3_or_453_nl <= (butterFly_3_mux1h_167_nl AND (NOT and_dcpl_477)) OR and_dcpl_457;
  yy_rsc_31_0_i_adra_d <= butterFly_3_or_8_nl & butterFly_3_butterFly_3_mux_rmff
      & butterFly_3_butterFly_3_or_rmff & butterFly_3_or_72_nl & butterFly_3_mux1h_104_nl
      & butterFly_3_or_453_nl;
  yy_rsc_31_0_i_wea_d <= STD_LOGIC_VECTOR'( and_1022_seb & butterFly_7_butterFly_7_or_95_rmff);
  butterFly_7_or_31_nl <= ((NOT(or_dcpl_268 OR or_dcpl_233 OR (and_dcpl_910 AND and_dcpl_519)))
      AND mux_3591_seb) OR and_dcpl_901;
  butterFly_7_and_374_nl <= (NOT(or_dcpl_273 AND and_dcpl_585 AND and_dcpl_878))
      AND mux_3591_seb;
  yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= STD_LOGIC_VECTOR'( butterFly_7_or_31_nl
      & butterFly_7_and_374_nl);
  yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= STD_LOGIC_VECTOR'( and_1022_seb
      & butterFly_7_butterFly_7_or_95_rmff);
  and_dcpl_1165 <= NOT(mux_100_cse OR (fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(0))
      OR (fsm_output(7)) OR (NOT (fsm_output(3))));
  and_dcpl_1178 <= (fsm_output(4)) AND (NOT (fsm_output(2))) AND nor_1375_cse AND
      (NOT (fsm_output(6))) AND (fsm_output(7)) AND (fsm_output(5)) AND (fsm_output(3));
  or_tmp_4090 <= (NOT (fsm_output(3))) OR (NOT (fsm_output(0))) OR (fsm_output(6));
  and_2399_cse <= nor_2178_cse_1 AND and_2083_cse;
  and_dcpl_1206 <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_1210 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_1222 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_1241 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("10"));
  and_dcpl_1246 <= (fsm_output(4)) AND (NOT (fsm_output(2)));
  and_dcpl_1257 <= CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("01"));
  and_dcpl_1324 <= NOT((NOT (fsm_output(6))) OR (fsm_output(7)) OR (fsm_output(5))
      OR (fsm_output(3)));
  and_dcpl_1455 <= (fsm_output(4)) AND (NOT (fsm_output(0)));
  and_dcpl_1566 <= (NOT (fsm_output(6))) AND (NOT (fsm_output(7))) AND (fsm_output(5))
      AND (fsm_output(3));
  and_dcpl_1573 <= (NOT (fsm_output(1))) AND (fsm_output(2)) AND (fsm_output(4))
      AND (NOT (fsm_output(0)));
  and_dcpl_1596 <= and_dcpl_1246 AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("00"));
  and_dcpl_1633 <= (fsm_output(4)) AND (fsm_output(2)) AND and_1317_cse;
  nor_2367_nl <= NOT((NOT (fsm_output(7))) OR (fsm_output(1)));
  nor_2368_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(1))));
  mux_4244_nl <= MUX_s_1_2_2(nor_2367_nl, nor_2368_nl, fsm_output(5));
  and_2383_ssc <= mux_4244_nl AND (fsm_output(2)) AND (NOT (fsm_output(4))) AND (fsm_output(0))
      AND nor_1395_cse;
  mux_tmp_4267 <= MUX_s_1_2_2(nor_tmp_35, (fsm_output(6)), fsm_output(3));
  mux_tmp_4268 <= MUX_s_1_2_2((NOT (fsm_output(7))), (fsm_output(7)), fsm_output(6));
  or_tmp_4112 <= CONV_SL_1_1(fsm_output(7 DOWNTO 6)/=STD_LOGIC_VECTOR'("00"));
  or_tmp_4115 <= (fsm_output(4)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(7));
  or_tmp_4117 <= (NOT (fsm_output(2))) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  or_tmp_4118 <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (fsm_output(7));
  or_tmp_4121 <= (NOT (fsm_output(2))) OR (fsm_output(6)) OR (NOT (fsm_output(7)));
  or_tmp_4152 <= (fsm_output(5)) OR (fsm_output(1)) OR (fsm_output(3));
  mux_tmp_4334 <= MUX_s_1_2_2((fsm_output(7)), or_tmp_48, fsm_output(1));
  or_tmp_4164 <= (NOT (fsm_output(1))) OR (fsm_output(7)) OR (fsm_output(5));
  or_tmp_4177 <= (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(5));
  mux_tmp_4373 <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), fsm_output(5));
  mux_tmp_4374 <= MUX_s_1_2_2((NOT (fsm_output(4))), and_2083_cse, fsm_output(5));
  or_tmp_4199 <= (fsm_output(4)) OR and_2141_cse;
  mux_tmp_4396 <= MUX_s_1_2_2(or_tmp_4199, or_2272_cse, fsm_output(0));
  or_tmp_4208 <= (fsm_output(7)) OR and_2120_cse;
  nor_2338_nl <= NOT((fsm_output(7)) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(4))
      OR (NOT (fsm_output(2))));
  nor_2340_nl <= NOT((fsm_output(6)) OR (NOT (fsm_output(1))) OR (NOT (fsm_output(4)))
      OR (fsm_output(2)));
  mux_4240_nl <= MUX_s_1_2_2(nor_2307_cse, nor_2340_nl, fsm_output(7));
  mux_4241_nl <= MUX_s_1_2_2(nor_2338_nl, mux_4240_nl, fsm_output(5));
  and_2348_ssc <= mux_4241_nl AND (fsm_output(0)) AND (fsm_output(3));
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND mux_104_nl) = '1' ) THEN
        m_sva <= MUX_v_32_2_2(m_rsci_idat, (xx_rsc_10_0_i_qa_d(31 DOWNTO 0)), and_dcpl_77);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( core_wen = '1' ) THEN
        revArr_rsci_s_raddr_core_4 <= S1_OUTER_LOOP_for_acc_svs_4;
        revArr_rsci_s_raddr_core_3_0 <= S1_OUTER_LOOP_for_acc_svs_3_0;
        reg_tw_rsci_s_raddr_core_cse <= S34_OUTER_LOOP_for_tf_mul_cmp_z_oreg;
        reg_x_rsc_0_0_i_s_raddr_core_cse <= MUX_v_5_2_2((reg_S2_COPY_LOOP_for_i_5_0_1_reg
            & reg_S2_COPY_LOOP_for_i_5_0_2_reg), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
            & reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg), and_dcpl_934);
        reg_x_rsc_0_0_i_s_waddr_core_cse <= MUX_v_5_2_2((reg_S2_COPY_LOOP_for_i_5_0_1_reg
            & reg_S2_COPY_LOOP_for_i_5_0_2_reg), (reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
            & reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg), and_dcpl_935);
        reg_x_rsc_0_0_i_s_dout_core_cse <= MUX1HOT_v_32_33_2(S2_INNER_LOOP1_tf_sva,
            S2_INNER_LOOP1_tfh_sva, operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm,
            tmp_13_sva_4, tmp_16_sva_4, tmp_13_sva_5, tmp_13_sva_6, tmp_12_sva_2,
            tmp_16_sva_8, tmp_13_sva_7, m_sva, modulo_add_base_1_sva, tmp_12_sva_4,
            mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm, mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm,
            mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm, operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm,
            tmp_12_sva_5, tmp_12_sva_6, operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm,
            tmp_12_sva_7, tmp_1_sva_7, tmp_16_sva_22, tmp_16_sva_23, tmp_13_sva_2,
            tmp_10_sva_2, tmp_16_sva_26, tmp_10_sva_4, tmp_10_sva_5, tmp_10_sva_6,
            tmp_10_sva_7, tmp_16_sva_31, tmp_55_lpi_3_dfm, STD_LOGIC_VECTOR'( S1_OUTER_LOOP_for_and_62_nl
            & S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_nl & S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_1_nl
            & S1_OUTER_LOOP_for_and_63_nl & S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_3_nl
            & S1_OUTER_LOOP_for_and_64_nl & S1_OUTER_LOOP_for_and_65_nl & S1_OUTER_LOOP_for_and_66_nl
            & S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_7_nl & S1_OUTER_LOOP_for_and_67_nl
            & S1_OUTER_LOOP_for_and_68_nl & S1_OUTER_LOOP_for_and_69_nl & S1_OUTER_LOOP_for_and_70_nl
            & S1_OUTER_LOOP_for_and_71_nl & S1_OUTER_LOOP_for_and_72_nl & S1_OUTER_LOOP_for_and_73_nl
            & S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_15_nl & S1_OUTER_LOOP_for_and_74_nl
            & S1_OUTER_LOOP_for_and_75_nl & S1_OUTER_LOOP_for_and_76_nl & S1_OUTER_LOOP_for_and_77_nl
            & S1_OUTER_LOOP_for_and_78_nl & S1_OUTER_LOOP_for_and_79_nl & S1_OUTER_LOOP_for_and_80_nl
            & S1_OUTER_LOOP_for_and_81_nl & S1_OUTER_LOOP_for_and_82_nl & S1_OUTER_LOOP_for_and_83_nl
            & S1_OUTER_LOOP_for_and_84_nl & S1_OUTER_LOOP_for_and_85_nl & S1_OUTER_LOOP_for_and_86_nl
            & S1_OUTER_LOOP_for_and_87_nl & S1_OUTER_LOOP_for_and_88_nl & and_dcpl_935));
        S34_OUTER_LOOP_for_tf_mul_cmp_a <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
            S34_OUTER_LOOP_for_tf_mux_1_nl, not_10627_nl);
        S34_OUTER_LOOP_for_k_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), S34_OUTER_LOOP_for_k_mux_nl,
            not_nl);
        tmp_16_sva_22 <= MUX1HOT_v_32_7_2(x_rsc_22_0_i_s_din_mxwt, (yy_rsc_22_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_2_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_1_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_22_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_1_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_1_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_16_sva_23 <= MUX1HOT_v_32_7_2(x_rsc_23_0_i_s_din_mxwt, (yy_rsc_23_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_6_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_5_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_23_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_5_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_5_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_16_sva_26 <= MUX1HOT_v_32_7_2(x_rsc_26_0_i_s_din_mxwt, (yy_rsc_26_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_14_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_13_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_26_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_13_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_13_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_16_sva_31 <= MUX1HOT_v_32_7_2(x_rsc_31_0_i_s_din_mxwt, (yy_rsc_31_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_3_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_2_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_31_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_2_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_2_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_16_sva_4 <= MUX1HOT_v_32_7_2(x_rsc_4_0_i_s_din_mxwt, (yy_rsc_4_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_7_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_6_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_4_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_6_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_6_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_16_sva_8 <= MUX1HOT_v_32_7_2(x_rsc_8_0_i_s_din_mxwt, (yy_rsc_8_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_15_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_14_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_8_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_14_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_14_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_26_sva_10 <= MUX1HOT_v_32_10_2(x_rsc_10_0_i_s_din_mxwt, (yy_rsc_10_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_14_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_14_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_15_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_10_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_10_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_14_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_14_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_10_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112 & and_dcpl_1113 & and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1116 & and_dcpl_1109
            & and_dcpl_1110 & and_dcpl_77));
        tmp_26_sva_5 <= MUX1HOT_v_32_10_2(x_rsc_5_0_i_s_din_mxwt, (yy_rsc_5_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_3_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_3_0_i_qa_d(31 DOWNTO
            0)), (xx_rsc_1_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_5_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_5_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_3_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_3_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_5_0_i_qa_d(63 DOWNTO 32)),
            STD_LOGIC_VECTOR'( and_dcpl_1112 & and_dcpl_1113 & and_dcpl_1114 & and_dcpl_1105
            & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1116 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_26_sva_6 <= MUX1HOT_v_32_10_2(x_rsc_6_0_i_s_din_mxwt, (yy_rsc_6_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_7_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_7_0_i_qa_d(31 DOWNTO
            0)), (xx_rsc_5_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_6_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_6_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_7_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_7_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_6_0_i_qa_d(63 DOWNTO 32)),
            STD_LOGIC_VECTOR'( and_dcpl_1112 & and_dcpl_1113 & and_dcpl_1114 & and_dcpl_1105
            & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1116 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_1_sva_7 <= MUX1HOT_v_32_8_2(x_rsc_21_0_i_s_din_mxwt, (yy_rsc_21_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_29_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_29_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_30_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_21_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_29_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_29_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_1101 & and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1108 & and_dcpl_1109 & and_dcpl_1110));
        tmp_10_sva_2 <= MUX1HOT_v_32_7_2(x_rsc_25_0_i_s_din_mxwt, (yy_rsc_25_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_10_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_9_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_25_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_9_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_9_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_10_sva_4 <= MUX1HOT_v_32_7_2(x_rsc_27_0_i_s_din_mxwt, (yy_rsc_27_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_18_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_17_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_27_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_17_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_17_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_10_sva_5 <= MUX1HOT_v_32_7_2(x_rsc_28_0_i_s_din_mxwt, (yy_rsc_28_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_22_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_21_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_28_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_21_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_21_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_10_sva_6 <= MUX1HOT_v_32_7_2(x_rsc_29_0_i_s_din_mxwt, (yy_rsc_29_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_26_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_25_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_29_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_25_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_25_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_10_sva_7 <= MUX1HOT_v_32_7_2(x_rsc_30_0_i_s_din_mxwt, (yy_rsc_30_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_30_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_29_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_30_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_29_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_29_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_12_sva_2 <= MUX1HOT_v_32_7_2(x_rsc_7_0_i_s_din_mxwt, (yy_rsc_7_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_11_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_10_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_7_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_10_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_10_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_1108 & and_dcpl_1109
            & and_dcpl_1110));
        tmp_14_sva_1 <= MUX1HOT_v_32_9_2(x_rsc_12_0_i_s_din_mxwt, (yy_rsc_12_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_4_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_4_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_12_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_12_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_4_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_4_0_i_qa_d(31 DOWNTO
            0)), (xx_rsc_12_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112
            & and_dcpl_1113 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1116
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_14_sva_6 <= MUX1HOT_v_32_9_2(x_rsc_17_0_i_s_din_mxwt, (yy_rsc_17_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_24_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_24_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_17_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_17_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_24_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_24_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_17_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112
            & and_dcpl_1113 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1116
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_14_sva_7 <= MUX1HOT_v_32_9_2(x_rsc_18_0_i_s_din_mxwt, (yy_rsc_18_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_28_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_28_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_18_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_18_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_28_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_28_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_18_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112
            & and_dcpl_1113 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1116
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_15_sva_2 <= MUX1HOT_v_32_9_2(x_rsc_20_0_i_s_din_mxwt, (yy_rsc_20_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_8_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_8_0_i_qa_d(31 DOWNTO
            0)), (yy_rsc_20_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_20_0_i_qa_d(31 DOWNTO
            0)), (yy_rsc_8_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_8_0_i_qa_d(63 DOWNTO
            32)), (xx_rsc_20_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112
            & and_dcpl_1113 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1116
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_15_sva_6 <= MUX1HOT_v_32_5_2(x_rsc_24_0_i_s_din_mxwt, (yy_rsc_24_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_24_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_24_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_24_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112
            & and_1222_nl & and_1225_nl & and_1229_nl & and_1231_nl));
        tmp_21_sva_4 <= MUX1HOT_v_32_9_2(x_rsc_3_0_i_s_din_mxwt, (yy_rsc_3_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_17_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_19_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_3_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_3_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_19_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_19_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_3_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112
            & and_dcpl_1113 & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1116
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_22_sva_4 <= MUX1HOT_v_32_10_2(x_rsc_9_0_i_s_din_mxwt, (yy_rsc_9_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_19_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_19_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_17_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_9_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_9_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_19_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_19_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_9_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1112 & and_dcpl_1113 & and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1116 & and_dcpl_1109
            & and_dcpl_1110 & and_dcpl_77));
        reg_tmp_54_lpi_3_dfm_cse <= MUX1HOT_v_32_32_2(S2_INNER_LOOP1_tf_sva, S2_INNER_LOOP1_tfh_sva,
            operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm,
            tmp_21_sva_4, tmp_16_sva_4, tmp_26_sva_5, tmp_26_sva_6, tmp_12_sva_2,
            tmp_16_sva_8, tmp_22_sva_4, tmp_26_sva_10, modulo_add_base_1_sva, tmp_14_sva_1,
            mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm, mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm,
            mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm, operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm,
            tmp_14_sva_6, tmp_14_sva_7, operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm,
            tmp_15_sva_2, tmp_1_sva_7, tmp_16_sva_22, tmp_16_sva_23, tmp_15_sva_6,
            tmp_10_sva_2, tmp_16_sva_26, tmp_10_sva_4, tmp_10_sva_5, tmp_10_sva_6,
            tmp_10_sva_7, tmp_16_sva_31, STD_LOGIC_VECTOR'( S1_OUTER_LOOP_for_mux_25_nl
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_2_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_4_itm & S1_OUTER_LOOP_for_mux_26_nl
            & S1_OUTER_LOOP_for_mux_27_nl & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54
            & S1_OUTER_LOOP_for_mux_28_nl & S1_OUTER_LOOP_for_mux_29_nl & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56 & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_18_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_19_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_20_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_21_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_22_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_23_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_24_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_25_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_26_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_27_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_28_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_29_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_30_itm));
        tmp_26_sva <= MUX1HOT_v_32_8_2(x_rsc_0_0_i_s_din_mxwt, (xx_rsc_2_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_2_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_3_0_i_qa_d(31 DOWNTO
            0)), (yy_rsc_0_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_2_0_i_qa_d(63 DOWNTO
            32)), (xx_rsc_2_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_0_0_i_qa_d(63 DOWNTO
            32)), STD_LOGIC_VECTOR'( and_dcpl_1136 & and_dcpl_1114 & and_dcpl_1105
            & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_26_sva_1 <= MUX1HOT_v_32_8_2(x_rsc_1_0_i_s_din_mxwt, (xx_rsc_6_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_6_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_7_0_i_qa_d(31 DOWNTO
            0)), (yy_rsc_1_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_6_0_i_qa_d(63 DOWNTO
            32)), (xx_rsc_6_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_1_0_i_qa_d(63 DOWNTO
            32)), STD_LOGIC_VECTOR'( and_dcpl_1136 & and_dcpl_1114 & and_dcpl_1105
            & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_26_sva_26 <= MUX1HOT_v_32_7_2(x_rsc_26_0_i_s_din_mxwt, (xx_rsc_1_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_3_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_26_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_3_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_3_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_26_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_26_sva_27 <= MUX1HOT_v_32_7_2(x_rsc_27_0_i_s_din_mxwt, (xx_rsc_5_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_7_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_27_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_7_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_7_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_27_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_26_sva_29 <= MUX1HOT_v_32_7_2(x_rsc_29_0_i_s_din_mxwt, (xx_rsc_13_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_15_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_29_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_15_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_15_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_29_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_26_sva_8 <= MUX1HOT_v_32_8_2(x_rsc_8_0_i_s_din_mxwt, (xx_rsc_15_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_15_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_13_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_8_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_15_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_15_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_8_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136 & and_dcpl_1114 & and_dcpl_1105
            & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_14_sva <= MUX1HOT_v_32_7_2(x_rsc_11_0_i_s_din_mxwt, (xx_rsc_0_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_0_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_11_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_0_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_0_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_11_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_14_sva_2 <= MUX1HOT_v_32_7_2(x_rsc_13_0_i_s_din_mxwt, (xx_rsc_8_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_8_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_13_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_8_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_8_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_13_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_14_sva_3 <= MUX1HOT_v_32_7_2(x_rsc_14_0_i_s_din_mxwt, (xx_rsc_12_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_12_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_14_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_12_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_12_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_14_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_14_sva_4 <= MUX1HOT_v_32_7_2(x_rsc_15_0_i_s_din_mxwt, (xx_rsc_16_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_16_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_15_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_16_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_16_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_15_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_14_sva_5 <= MUX1HOT_v_32_7_2(x_rsc_16_0_i_s_din_mxwt, (xx_rsc_20_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_20_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_16_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_20_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_20_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_16_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_15_sva <= MUX1HOT_v_32_7_2(x_rsc_19_0_i_s_din_mxwt, (xx_rsc_0_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_0_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_19_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_0_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_0_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_19_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_15_sva_1 <= MUX1HOT_v_32_7_2(x_rsc_2_0_i_s_din_mxwt, (xx_rsc_4_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_4_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_2_0_i_qa_d(63 DOWNTO
            32)), (yy_rsc_4_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_4_0_i_qa_d(63 DOWNTO
            32)), (xx_rsc_2_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_15_sva_3 <= MUX1HOT_v_32_7_2(x_rsc_21_0_i_s_din_mxwt, (xx_rsc_12_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_12_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_21_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_12_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_12_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_21_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_15_sva_4 <= MUX1HOT_v_32_7_2(x_rsc_22_0_i_s_din_mxwt, (xx_rsc_16_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_16_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_22_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_16_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_16_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_22_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_15_sva_5 <= MUX1HOT_v_32_7_2(x_rsc_23_0_i_s_din_mxwt, (xx_rsc_20_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_20_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_23_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_20_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_20_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_23_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_15_sva_7 <= MUX1HOT_v_32_7_2(x_rsc_25_0_i_s_din_mxwt, (xx_rsc_28_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_28_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_25_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_28_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_28_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_25_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_21_sva_2 <= MUX1HOT_v_32_7_2(x_rsc_28_0_i_s_din_mxwt, (xx_rsc_9_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_11_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_28_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_11_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_11_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_28_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_21_sva_5 <= MUX1HOT_v_32_7_2(x_rsc_30_0_i_s_din_mxwt, (xx_rsc_21_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_23_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_30_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_23_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_23_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_30_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_21_sva_6 <= MUX1HOT_v_32_7_2(x_rsc_31_0_i_s_din_mxwt, (xx_rsc_25_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_27_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_31_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_27_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_27_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_31_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_21_sva_7 <= MUX1HOT_v_32_7_2(x_rsc_4_0_i_s_din_mxwt, (xx_rsc_29_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_31_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_4_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_31_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_31_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_4_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136
            & and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_22_sva_2 <= MUX1HOT_v_32_8_2(x_rsc_7_0_i_s_din_mxwt, (xx_rsc_11_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_11_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_9_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_7_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_11_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_11_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_7_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1136 & and_dcpl_1114 & and_dcpl_1105
            & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_55_lpi_3_dfm <= MUX1HOT_v_32_32_2(tmp_26_sva, tmp_26_sva_1, tmp_15_sva_1,
            tmp_21_sva_4, tmp_21_sva_7, tmp_26_sva_5, tmp_26_sva_6, tmp_22_sva_2,
            tmp_26_sva_8, tmp_22_sva_4, tmp_26_sva_10, tmp_14_sva, tmp_14_sva_1,
            tmp_14_sva_2, tmp_14_sva_3, tmp_14_sva_4, tmp_14_sva_5, tmp_14_sva_6,
            tmp_14_sva_7, tmp_15_sva, tmp_15_sva_2, tmp_15_sva_3, tmp_15_sva_4, tmp_15_sva_5,
            tmp_15_sva_6, tmp_15_sva_7, tmp_26_sva_26, tmp_26_sva_27, tmp_21_sva_2,
            tmp_26_sva_29, tmp_21_sva_5, tmp_21_sva_6, STD_LOGIC_VECTOR'( S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_1_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_82_nl & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_83_nl
            & S1_OUTER_LOOP_for_mux_30_nl & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58
            & S1_OUTER_LOOP_for_mux_31_nl & S1_OUTER_LOOP_for_mux_32_nl & S1_OUTER_LOOP_for_mux_33_nl
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_66 & S1_OUTER_LOOP_for_mux_34_nl
            & S1_OUTER_LOOP_for_mux_35_nl & S1_OUTER_LOOP_for_mux_36_nl & S1_OUTER_LOOP_for_mux_37_nl
            & S1_OUTER_LOOP_for_mux_38_nl & S1_OUTER_LOOP_for_mux_39_nl & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_45_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_84_nl & S1_OUTER_LOOP_for_mux_40_nl
            & S1_OUTER_LOOP_for_mux_41_nl & S1_OUTER_LOOP_for_mux_42_nl & S1_OUTER_LOOP_for_mux_43_nl
            & S1_OUTER_LOOP_for_mux_44_nl & S1_OUTER_LOOP_for_mux_45_nl & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_53_itm
            & S1_OUTER_LOOP_for_mux_46_nl & S1_OUTER_LOOP_for_mux_47_nl & S1_OUTER_LOOP_for_mux_48_nl
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_57_itm & S1_OUTER_LOOP_for_mux_49_nl
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_59_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_60_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_61_itm));
        S2_OUTER_LOOP_c_2_sva <= NOT(mux_4091_nl AND (fsm_output(4)) AND and_2893_cse
            AND (NOT (fsm_output(6))) AND (fsm_output(3)));
        tmp_12_sva_4 <= MUX1HOT_v_32_6_2((xx_rsc_19_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_18_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_12_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_18_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_18_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_12_0_i_qa_d(31
            DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_12_sva_5 <= MUX1HOT_v_32_6_2((xx_rsc_23_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_22_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_17_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_22_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_22_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_17_0_i_qa_d(31
            DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_12_sva_6 <= MUX1HOT_v_32_6_2((xx_rsc_27_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_26_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_18_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_26_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_26_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_18_0_i_qa_d(31
            DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_12_sva_7 <= MUX1HOT_v_32_6_2((xx_rsc_31_0_i_qa_d(63 DOWNTO 32)), (yy_rsc_30_0_i_qa_d(63
            DOWNTO 32)), (yy_rsc_20_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_30_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_30_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_20_0_i_qa_d(31
            DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1103 & and_dcpl_1105 & and_dcpl_93
            & and_dcpl_1109 & and_dcpl_1110 & and_dcpl_77));
        tmp_13_sva_2 <= MUX1HOT_v_32_7_2((xx_rsc_10_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_10_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_11_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_24_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_10_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_10_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_24_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_13_sva_4 <= MUX1HOT_v_32_7_2((xx_rsc_18_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_18_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_19_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_3_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_18_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_18_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_3_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_13_sva_5 <= MUX1HOT_v_32_7_2((xx_rsc_22_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_22_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_23_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_5_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_22_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_22_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_5_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_13_sva_6 <= MUX1HOT_v_32_7_2((xx_rsc_26_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_26_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_27_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_6_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_26_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_26_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_6_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_13_sva_7 <= MUX1HOT_v_32_7_2((xx_rsc_30_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_30_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_31_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_9_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_30_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_30_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_9_0_i_qa_d(31 DOWNTO 0)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110
            & and_dcpl_77));
        tmp_22_sva_5 <= MUX1HOT_v_32_6_2((xx_rsc_23_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_23_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_21_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_10_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_23_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_23_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1114 & and_dcpl_1105 & and_dcpl_1115
            & and_dcpl_93 & and_dcpl_1109 & and_dcpl_1110));
        tmp_22_sva_6 <= MUX1HOT_v_32_5_2((xx_rsc_27_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_27_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_25_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_27_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_27_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1109 & and_dcpl_1110));
        tmp_22_sva_7 <= MUX1HOT_v_32_5_2((xx_rsc_31_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_31_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_29_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_31_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_31_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_1114
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1109 & and_dcpl_1110));
        mult_3_res_sva <= acc_1_nl(32 DOWNTO 1);
        reg_mult_3_res_lpi_4_dfm_cse <= MUX_v_32_2_2(z_out_5, mult_3_res_sva, z_out_17_32);
        reg_mult_2_res_lpi_4_dfm_cse <= MUX_v_32_2_2(z_out_6, mult_3_res_sva, z_out_17_32);
        modulo_sub_3_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_3_sva_1(30
            DOWNTO 0))), z_out_7, modulo_sub_base_3_sva_1(31));
        mult_1_res_sva <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm)
            - UNSIGNED(mult_z_mul_cmp_z(31 DOWNTO 0)), 32));
        reg_mult_1_res_lpi_4_dfm_cse <= MUX_v_32_2_2(z_out_5, mult_1_res_sva, z_out_19_32);
        modulo_sub_2_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_2_sva_1(30
            DOWNTO 0))), z_out_8, modulo_sub_base_2_sva_1(31));
        reg_mult_res_lpi_4_dfm_cse <= MUX_v_32_2_2(z_out_6, mult_3_res_sva, z_out_19_32);
        modulo_sub_1_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_1_sva_1(30
            DOWNTO 0))), z_out_9, modulo_sub_base_1_sva_1(31));
        modulo_sub_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_sva_1(30
            DOWNTO 0))), z_out_10, modulo_sub_base_sva_1(31));
        modulo_sub_7_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_7_sva_1(30
            DOWNTO 0))), z_out_11, modulo_sub_base_7_sva_1(31));
        modulo_sub_6_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_6_sva_1(30
            DOWNTO 0))), z_out_7, modulo_sub_base_6_sva_1(31));
        modulo_sub_5_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_5_sva_1(30
            DOWNTO 0))), z_out_13, modulo_sub_base_5_sva_1(31));
        modulo_sub_4_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_4_sva_1(30
            DOWNTO 0))), z_out_10, modulo_sub_base_4_sva_1(31));
        modulo_sub_11_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_11_sva_1(30
            DOWNTO 0))), z_out_8, modulo_sub_base_11_sva_1(31));
        modulo_sub_10_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_10_sva_1(30
            DOWNTO 0))), z_out_9, modulo_sub_base_10_sva_1(31));
        modulo_sub_9_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_9_sva_1(30
            DOWNTO 0))), z_out_9, modulo_sub_base_9_sva_1(31));
        modulo_sub_8_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_8_sva_1(30
            DOWNTO 0))), z_out_10, modulo_sub_base_8_sva_1(31));
        S34_OUTER_LOOP_for_tf_h_sva <= tw_h_rsci_s_din_mxwt;
        tmp_36_lpi_3_dfm <= MUX1HOT_v_32_32_2(tmp_26_sva, tmp_26_sva_1, tmp_15_sva_1,
            tmp_21_sva_4, tmp_21_sva_7, tmp_26_sva_5, tmp_26_sva_6, tmp_22_sva_2,
            tmp_26_sva_8, tmp_22_sva_4, tmp_26_sva_10, tmp_14_sva, tmp_14_sva_1,
            tmp_14_sva_2, tmp_14_sva_3, tmp_14_sva_4, tmp_14_sva_5, tmp_14_sva_6,
            tmp_14_sva_7, tmp_15_sva, tmp_15_sva_2, tmp_15_sva_3, tmp_15_sva_4, tmp_15_sva_5,
            tmp_15_sva_6, tmp_15_sva_7, tmp_26_sva_26, tmp_26_sva_27, tmp_21_sva_2,
            tmp_26_sva_29, tmp_21_sva_5, tmp_21_sva_6, STD_LOGIC_VECTOR'( S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_nl & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_1_nl
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_66
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_15_nl
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm
            & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm & S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm
            & S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm));
        S34_OUTER_LOOP_for_tf_sva <= tw_rsci_s_din_mxwt;
        modulo_sub_15_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_15_sva_1(30
            DOWNTO 0))), z_out_11, modulo_sub_base_15_sva_1(31));
        modulo_sub_14_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_14_sva_1(30
            DOWNTO 0))), z_out_7, modulo_sub_base_14_sva_1(31));
        modulo_sub_13_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_13_sva_1(30
            DOWNTO 0))), z_out_13, modulo_sub_base_13_sva_1(31));
        modulo_sub_12_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_12_sva_1(30
            DOWNTO 0))), z_out_14, modulo_sub_base_12_sva_1(31));
        modulo_sub_19_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_19_sva_1(30
            DOWNTO 0))), z_out_11, modulo_sub_base_19_sva_1(31));
        reg_modulo_sub_18_qr_lpi_4_dfm_cse <= MUX_v_32_2_2(('0' & (z_out_12(30 DOWNTO
            0))), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_sub_18_qif_acc_nl),
            32)), z_out_12(31));
        modulo_sub_17_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_17_sva_1(30
            DOWNTO 0))), z_out_13, modulo_sub_base_17_sva_1(31));
        modulo_sub_16_qr_lpi_4_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_16_sva_1(30
            DOWNTO 0))), z_out_14, modulo_sub_base_16_sva_1(31));
        modulo_sub_23_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_23_sva_1(30
            DOWNTO 0))), z_out_9, modulo_sub_base_23_sva_1(31));
        modulo_sub_21_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_21_sva_1(30
            DOWNTO 0))), z_out_8, modulo_sub_base_21_sva_1(31));
        modulo_sub_20_qr_lpi_3_dfm <= MUX_v_32_2_2(('0' & (modulo_sub_base_20_sva_1(30
            DOWNTO 0))), z_out_14, modulo_sub_base_20_sva_1(31));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_twiddle_rsci_oswt_cse <= '0';
        reg_revArr_rsci_oswt_cse <= '0';
        reg_tw_rsci_oswt_cse <= '0';
        reg_xx_rsc_0_0_cgo_cse <= '0';
        reg_xx_rsc_1_0_cgo_cse <= '0';
        reg_xx_rsc_2_0_cgo_cse <= '0';
        reg_xx_rsc_3_0_cgo_cse <= '0';
        reg_xx_rsc_4_0_cgo_cse <= '0';
        reg_xx_rsc_5_0_cgo_cse <= '0';
        reg_xx_rsc_6_0_cgo_cse <= '0';
        reg_xx_rsc_7_0_cgo_cse <= '0';
        reg_xx_rsc_8_0_cgo_cse <= '0';
        reg_xx_rsc_9_0_cgo_cse <= '0';
        reg_xx_rsc_10_0_cgo_cse <= '0';
        reg_xx_rsc_11_0_cgo_cse <= '0';
        reg_xx_rsc_12_0_cgo_cse <= '0';
        reg_xx_rsc_13_0_cgo_cse <= '0';
        reg_xx_rsc_14_0_cgo_cse <= '0';
        reg_xx_rsc_15_0_cgo_cse <= '0';
        reg_xx_rsc_16_0_cgo_cse <= '0';
        reg_xx_rsc_17_0_cgo_cse <= '0';
        reg_xx_rsc_18_0_cgo_cse <= '0';
        reg_xx_rsc_19_0_cgo_cse <= '0';
        reg_xx_rsc_20_0_cgo_cse <= '0';
        reg_xx_rsc_21_0_cgo_cse <= '0';
        reg_xx_rsc_22_0_cgo_cse <= '0';
        reg_xx_rsc_23_0_cgo_cse <= '0';
        reg_xx_rsc_24_0_cgo_cse <= '0';
        reg_xx_rsc_25_0_cgo_cse <= '0';
        reg_xx_rsc_26_0_cgo_cse <= '0';
        reg_xx_rsc_27_0_cgo_cse <= '0';
        reg_xx_rsc_28_0_cgo_cse <= '0';
        reg_xx_rsc_29_0_cgo_cse <= '0';
        reg_xx_rsc_30_0_cgo_cse <= '0';
        reg_xx_rsc_31_0_cgo_cse <= '0';
        reg_yy_rsc_0_0_cgo_cse <= '0';
        reg_yy_rsc_1_0_cgo_cse <= '0';
        reg_yy_rsc_2_0_cgo_cse <= '0';
        reg_yy_rsc_3_0_cgo_cse <= '0';
        reg_yy_rsc_4_0_cgo_cse <= '0';
        reg_yy_rsc_5_0_cgo_cse <= '0';
        reg_yy_rsc_6_0_cgo_cse <= '0';
        reg_yy_rsc_7_0_cgo_cse <= '0';
        reg_yy_rsc_8_0_cgo_cse <= '0';
        reg_yy_rsc_9_0_cgo_cse <= '0';
        reg_yy_rsc_10_0_cgo_cse <= '0';
        reg_yy_rsc_11_0_cgo_cse <= '0';
        reg_yy_rsc_12_0_cgo_cse <= '0';
        reg_yy_rsc_13_0_cgo_cse <= '0';
        reg_yy_rsc_14_0_cgo_cse <= '0';
        reg_yy_rsc_15_0_cgo_cse <= '0';
        reg_yy_rsc_16_0_cgo_cse <= '0';
        reg_yy_rsc_17_0_cgo_cse <= '0';
        reg_yy_rsc_18_0_cgo_cse <= '0';
        reg_yy_rsc_19_0_cgo_cse <= '0';
        reg_yy_rsc_20_0_cgo_cse <= '0';
        reg_yy_rsc_21_0_cgo_cse <= '0';
        reg_yy_rsc_22_0_cgo_cse <= '0';
        reg_yy_rsc_23_0_cgo_cse <= '0';
        reg_yy_rsc_24_0_cgo_cse <= '0';
        reg_yy_rsc_25_0_cgo_cse <= '0';
        reg_yy_rsc_26_0_cgo_cse <= '0';
        reg_yy_rsc_27_0_cgo_cse <= '0';
        reg_yy_rsc_28_0_cgo_cse <= '0';
        reg_yy_rsc_29_0_cgo_cse <= '0';
        reg_yy_rsc_30_0_cgo_cse <= '0';
        reg_yy_rsc_31_0_cgo_cse <= '0';
        reg_x_rsc_0_0_i_oswt_cse <= '0';
        reg_x_rsc_0_0_i_oswt_1_cse <= '0';
        reg_x_rsc_1_0_i_oswt_cse <= '0';
        reg_x_rsc_1_0_i_oswt_1_cse <= '0';
        reg_x_rsc_2_0_i_oswt_cse <= '0';
        reg_x_rsc_2_0_i_oswt_1_cse <= '0';
        reg_x_rsc_3_0_i_oswt_cse <= '0';
        reg_x_rsc_3_0_i_oswt_1_cse <= '0';
        reg_x_rsc_4_0_i_oswt_cse <= '0';
        reg_x_rsc_4_0_i_oswt_1_cse <= '0';
        reg_x_rsc_5_0_i_oswt_cse <= '0';
        reg_x_rsc_5_0_i_oswt_1_cse <= '0';
        reg_x_rsc_6_0_i_oswt_cse <= '0';
        reg_x_rsc_6_0_i_oswt_1_cse <= '0';
        reg_x_rsc_7_0_i_oswt_cse <= '0';
        reg_x_rsc_7_0_i_oswt_1_cse <= '0';
        reg_x_rsc_8_0_i_oswt_cse <= '0';
        reg_x_rsc_8_0_i_oswt_1_cse <= '0';
        reg_x_rsc_9_0_i_oswt_cse <= '0';
        reg_x_rsc_9_0_i_oswt_1_cse <= '0';
        reg_x_rsc_10_0_i_oswt_cse <= '0';
        reg_x_rsc_10_0_i_oswt_1_cse <= '0';
        reg_x_rsc_11_0_i_oswt_cse <= '0';
        reg_x_rsc_11_0_i_oswt_1_cse <= '0';
        reg_x_rsc_12_0_i_oswt_cse <= '0';
        reg_x_rsc_12_0_i_oswt_1_cse <= '0';
        reg_x_rsc_13_0_i_oswt_cse <= '0';
        reg_x_rsc_13_0_i_oswt_1_cse <= '0';
        reg_x_rsc_14_0_i_oswt_cse <= '0';
        reg_x_rsc_14_0_i_oswt_1_cse <= '0';
        reg_x_rsc_15_0_i_oswt_cse <= '0';
        reg_x_rsc_15_0_i_oswt_1_cse <= '0';
        reg_x_rsc_16_0_i_oswt_cse <= '0';
        reg_x_rsc_16_0_i_oswt_1_cse <= '0';
        reg_x_rsc_17_0_i_oswt_cse <= '0';
        reg_x_rsc_17_0_i_oswt_1_cse <= '0';
        reg_x_rsc_18_0_i_oswt_cse <= '0';
        reg_x_rsc_18_0_i_oswt_1_cse <= '0';
        reg_x_rsc_19_0_i_oswt_cse <= '0';
        reg_x_rsc_19_0_i_oswt_1_cse <= '0';
        reg_x_rsc_20_0_i_oswt_cse <= '0';
        reg_x_rsc_20_0_i_oswt_1_cse <= '0';
        reg_x_rsc_21_0_i_oswt_cse <= '0';
        reg_x_rsc_21_0_i_oswt_1_cse <= '0';
        reg_x_rsc_22_0_i_oswt_cse <= '0';
        reg_x_rsc_22_0_i_oswt_1_cse <= '0';
        reg_x_rsc_23_0_i_oswt_cse <= '0';
        reg_x_rsc_23_0_i_oswt_1_cse <= '0';
        reg_x_rsc_24_0_i_oswt_cse <= '0';
        reg_x_rsc_24_0_i_oswt_1_cse <= '0';
        reg_x_rsc_25_0_i_oswt_cse <= '0';
        reg_x_rsc_25_0_i_oswt_1_cse <= '0';
        reg_x_rsc_26_0_i_oswt_cse <= '0';
        reg_x_rsc_26_0_i_oswt_1_cse <= '0';
        reg_x_rsc_27_0_i_oswt_cse <= '0';
        reg_x_rsc_27_0_i_oswt_1_cse <= '0';
        reg_x_rsc_28_0_i_oswt_cse <= '0';
        reg_x_rsc_28_0_i_oswt_1_cse <= '0';
        reg_x_rsc_29_0_i_oswt_cse <= '0';
        reg_x_rsc_29_0_i_oswt_1_cse <= '0';
        reg_x_rsc_30_0_i_oswt_cse <= '0';
        reg_x_rsc_30_0_i_oswt_1_cse <= '0';
        reg_x_rsc_31_0_i_oswt_cse <= '0';
        reg_x_rsc_31_0_i_oswt_1_cse <= '0';
        reg_x_rsc_triosy_31_0_obj_iswt0_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        reg_ensig_cgo_1_cse <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_9_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_19_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_23_itm <= '0';
        reg_modulo_add_3_slc_32_svs_st_cse <= '0';
        reg_modulo_add_2_slc_32_svs_st_cse <= '0';
        reg_modulo_add_1_slc_32_svs_st_cse <= '0';
        reg_modulo_add_7_slc_32_svs_st_cse <= '0';
        reg_modulo_add_6_slc_32_svs_st_cse <= '0';
        reg_modulo_add_5_slc_32_svs_st_cse <= '0';
        reg_modulo_add_11_slc_32_svs_st_cse <= '0';
        modulo_add_13_slc_32_svs_st <= '0';
      ELSIF ( core_wen = '1' ) THEN
        reg_twiddle_rsci_oswt_cse <= mux_111_rmff;
        reg_revArr_rsci_oswt_cse <= and_dcpl_88;
        reg_tw_rsci_oswt_cse <= and_dcpl_93;
        reg_xx_rsc_0_0_cgo_cse <= NOT mux_138_itm;
        reg_xx_rsc_1_0_cgo_cse <= mux_191_rmff;
        reg_xx_rsc_2_0_cgo_cse <= mux_241_rmff;
        reg_xx_rsc_3_0_cgo_cse <= mux_293_rmff;
        reg_xx_rsc_4_0_cgo_cse <= NOT mux_357_itm;
        reg_xx_rsc_5_0_cgo_cse <= mux_408_rmff;
        reg_xx_rsc_6_0_cgo_cse <= mux_455_rmff;
        reg_xx_rsc_7_0_cgo_cse <= mux_504_rmff;
        reg_xx_rsc_8_0_cgo_cse <= NOT mux_566_itm;
        reg_xx_rsc_9_0_cgo_cse <= mux_614_rmff;
        reg_xx_rsc_10_0_cgo_cse <= mux_661_rmff;
        reg_xx_rsc_11_0_cgo_cse <= mux_710_rmff;
        reg_xx_rsc_12_0_cgo_cse <= NOT mux_772_itm;
        reg_xx_rsc_13_0_cgo_cse <= mux_820_rmff;
        reg_xx_rsc_14_0_cgo_cse <= mux_867_rmff;
        reg_xx_rsc_15_0_cgo_cse <= mux_916_rmff;
        reg_xx_rsc_16_0_cgo_cse <= NOT mux_979_itm;
        reg_xx_rsc_17_0_cgo_cse <= mux_1030_rmff;
        reg_xx_rsc_18_0_cgo_cse <= mux_1080_rmff;
        reg_xx_rsc_19_0_cgo_cse <= mux_1132_rmff;
        reg_xx_rsc_20_0_cgo_cse <= NOT mux_1196_itm;
        reg_xx_rsc_21_0_cgo_cse <= mux_1248_rmff;
        reg_xx_rsc_22_0_cgo_cse <= mux_1298_rmff;
        reg_xx_rsc_23_0_cgo_cse <= mux_1350_rmff;
        reg_xx_rsc_24_0_cgo_cse <= NOT mux_1414_itm;
        reg_xx_rsc_25_0_cgo_cse <= mux_1465_rmff;
        reg_xx_rsc_26_0_cgo_cse <= mux_1515_rmff;
        reg_xx_rsc_27_0_cgo_cse <= mux_1567_rmff;
        reg_xx_rsc_28_0_cgo_cse <= NOT mux_1631_itm;
        reg_xx_rsc_29_0_cgo_cse <= mux_1682_rmff;
        reg_xx_rsc_30_0_cgo_cse <= mux_1732_rmff;
        reg_xx_rsc_31_0_cgo_cse <= mux_1781_rmff;
        reg_yy_rsc_0_0_cgo_cse <= NOT mux_1843_itm;
        reg_yy_rsc_1_0_cgo_cse <= NOT mux_1902_itm;
        reg_yy_rsc_2_0_cgo_cse <= NOT mux_1950_itm;
        reg_yy_rsc_3_0_cgo_cse <= NOT mux_2010_itm;
        reg_yy_rsc_4_0_cgo_cse <= NOT mux_2075_itm;
        reg_yy_rsc_5_0_cgo_cse <= NOT mux_2130_itm;
        reg_yy_rsc_6_0_cgo_cse <= NOT mux_2175_itm;
        reg_yy_rsc_7_0_cgo_cse <= NOT mux_2233_itm;
        reg_yy_rsc_8_0_cgo_cse <= NOT mux_2295_itm;
        reg_yy_rsc_9_0_cgo_cse <= NOT mux_2350_itm;
        reg_yy_rsc_10_0_cgo_cse <= NOT mux_2395_itm;
        reg_yy_rsc_11_0_cgo_cse <= NOT mux_2453_itm;
        reg_yy_rsc_12_0_cgo_cse <= NOT mux_2515_itm;
        reg_yy_rsc_13_0_cgo_cse <= NOT mux_2570_itm;
        reg_yy_rsc_14_0_cgo_cse <= NOT mux_2615_itm;
        reg_yy_rsc_15_0_cgo_cse <= NOT mux_2673_itm;
        reg_yy_rsc_16_0_cgo_cse <= NOT mux_2735_itm;
        reg_yy_rsc_17_0_cgo_cse <= NOT mux_2790_itm;
        reg_yy_rsc_18_0_cgo_cse <= NOT mux_2835_itm;
        reg_yy_rsc_19_0_cgo_cse <= NOT mux_2893_itm;
        reg_yy_rsc_20_0_cgo_cse <= NOT mux_2955_itm;
        reg_yy_rsc_21_0_cgo_cse <= NOT mux_3010_itm;
        reg_yy_rsc_22_0_cgo_cse <= NOT mux_3055_itm;
        reg_yy_rsc_23_0_cgo_cse <= NOT mux_3113_itm;
        reg_yy_rsc_24_0_cgo_cse <= NOT mux_3175_itm;
        reg_yy_rsc_25_0_cgo_cse <= NOT mux_3230_itm;
        reg_yy_rsc_26_0_cgo_cse <= NOT mux_3275_itm;
        reg_yy_rsc_27_0_cgo_cse <= NOT mux_3333_itm;
        reg_yy_rsc_28_0_cgo_cse <= NOT mux_3395_itm;
        reg_yy_rsc_29_0_cgo_cse <= NOT mux_3450_itm;
        reg_yy_rsc_30_0_cgo_cse <= NOT mux_3495_itm;
        reg_yy_rsc_31_0_cgo_cse <= NOT mux_3553_itm;
        reg_x_rsc_0_0_i_oswt_cse <= mux_3592_nl AND and_dcpl_927;
        reg_x_rsc_0_0_i_oswt_1_cse <= (NOT mux_3593_nl) AND and_dcpl_932;
        reg_x_rsc_1_0_i_oswt_cse <= mux_3594_nl AND and_dcpl_927;
        reg_x_rsc_1_0_i_oswt_1_cse <= (NOT mux_3595_nl) AND and_dcpl_932;
        reg_x_rsc_2_0_i_oswt_cse <= mux_3596_nl AND and_dcpl_927;
        reg_x_rsc_2_0_i_oswt_1_cse <= (NOT mux_3597_nl) AND and_dcpl_932;
        reg_x_rsc_3_0_i_oswt_cse <= mux_3598_nl AND and_dcpl_927;
        reg_x_rsc_3_0_i_oswt_1_cse <= (NOT mux_3599_nl) AND and_dcpl_932;
        reg_x_rsc_4_0_i_oswt_cse <= mux_3600_nl AND and_dcpl_927;
        reg_x_rsc_4_0_i_oswt_1_cse <= (NOT mux_3601_nl) AND and_dcpl_932;
        reg_x_rsc_5_0_i_oswt_cse <= mux_3602_nl AND and_dcpl_927;
        reg_x_rsc_5_0_i_oswt_1_cse <= (NOT mux_3603_nl) AND and_dcpl_932;
        reg_x_rsc_6_0_i_oswt_cse <= mux_3604_nl AND and_dcpl_927;
        reg_x_rsc_6_0_i_oswt_1_cse <= (NOT mux_3605_nl) AND and_dcpl_932;
        reg_x_rsc_7_0_i_oswt_cse <= mux_3606_nl AND and_dcpl_927;
        reg_x_rsc_7_0_i_oswt_1_cse <= (NOT mux_3607_nl) AND and_dcpl_932;
        reg_x_rsc_8_0_i_oswt_cse <= mux_3608_nl AND and_dcpl_927;
        reg_x_rsc_8_0_i_oswt_1_cse <= (NOT mux_3609_nl) AND and_dcpl_932;
        reg_x_rsc_9_0_i_oswt_cse <= mux_3610_nl AND and_dcpl_927;
        reg_x_rsc_9_0_i_oswt_1_cse <= (NOT mux_3611_nl) AND and_dcpl_932;
        reg_x_rsc_10_0_i_oswt_cse <= mux_3612_nl AND and_dcpl_927;
        reg_x_rsc_10_0_i_oswt_1_cse <= (NOT mux_3613_nl) AND and_dcpl_932;
        reg_x_rsc_11_0_i_oswt_cse <= mux_3614_nl AND and_dcpl_927;
        reg_x_rsc_11_0_i_oswt_1_cse <= (NOT mux_3615_nl) AND and_dcpl_932;
        reg_x_rsc_12_0_i_oswt_cse <= mux_3616_nl AND and_dcpl_927;
        reg_x_rsc_12_0_i_oswt_1_cse <= (NOT mux_3617_nl) AND and_dcpl_932;
        reg_x_rsc_13_0_i_oswt_cse <= mux_3618_nl AND and_dcpl_927;
        reg_x_rsc_13_0_i_oswt_1_cse <= (NOT mux_3619_nl) AND and_dcpl_932;
        reg_x_rsc_14_0_i_oswt_cse <= mux_3620_nl AND and_dcpl_927;
        reg_x_rsc_14_0_i_oswt_1_cse <= (NOT mux_3621_nl) AND and_dcpl_932;
        reg_x_rsc_15_0_i_oswt_cse <= mux_3622_nl AND and_dcpl_927;
        reg_x_rsc_15_0_i_oswt_1_cse <= (NOT mux_3623_nl) AND and_dcpl_932;
        reg_x_rsc_16_0_i_oswt_cse <= mux_3624_nl AND and_dcpl_927;
        reg_x_rsc_16_0_i_oswt_1_cse <= (NOT mux_3625_nl) AND and_dcpl_932;
        reg_x_rsc_17_0_i_oswt_cse <= mux_3626_nl AND and_dcpl_927;
        reg_x_rsc_17_0_i_oswt_1_cse <= (NOT mux_3627_nl) AND and_dcpl_932;
        reg_x_rsc_18_0_i_oswt_cse <= mux_3628_nl AND and_dcpl_927;
        reg_x_rsc_18_0_i_oswt_1_cse <= (NOT mux_3629_nl) AND and_dcpl_932;
        reg_x_rsc_19_0_i_oswt_cse <= mux_3630_nl AND and_dcpl_927;
        reg_x_rsc_19_0_i_oswt_1_cse <= (NOT mux_3631_nl) AND and_dcpl_932;
        reg_x_rsc_20_0_i_oswt_cse <= mux_3632_nl AND and_dcpl_927;
        reg_x_rsc_20_0_i_oswt_1_cse <= (NOT mux_3633_nl) AND and_dcpl_932;
        reg_x_rsc_21_0_i_oswt_cse <= mux_3634_nl AND and_dcpl_927;
        reg_x_rsc_21_0_i_oswt_1_cse <= (NOT mux_3635_nl) AND and_dcpl_932;
        reg_x_rsc_22_0_i_oswt_cse <= mux_3636_nl AND and_dcpl_927;
        reg_x_rsc_22_0_i_oswt_1_cse <= (NOT mux_3637_nl) AND and_dcpl_932;
        reg_x_rsc_23_0_i_oswt_cse <= mux_3638_nl AND and_dcpl_927;
        reg_x_rsc_23_0_i_oswt_1_cse <= (NOT mux_3639_nl) AND and_dcpl_932;
        reg_x_rsc_24_0_i_oswt_cse <= mux_3640_nl AND and_dcpl_927;
        reg_x_rsc_24_0_i_oswt_1_cse <= (NOT mux_3641_nl) AND and_dcpl_932;
        reg_x_rsc_25_0_i_oswt_cse <= mux_3642_nl AND and_dcpl_927;
        reg_x_rsc_25_0_i_oswt_1_cse <= (NOT mux_3643_nl) AND and_dcpl_932;
        reg_x_rsc_26_0_i_oswt_cse <= mux_3644_nl AND and_dcpl_927;
        reg_x_rsc_26_0_i_oswt_1_cse <= (NOT mux_3645_nl) AND and_dcpl_932;
        reg_x_rsc_27_0_i_oswt_cse <= mux_3646_nl AND and_dcpl_927;
        reg_x_rsc_27_0_i_oswt_1_cse <= (NOT mux_3647_nl) AND and_dcpl_932;
        reg_x_rsc_28_0_i_oswt_cse <= mux_3648_nl AND and_dcpl_927;
        reg_x_rsc_28_0_i_oswt_1_cse <= (NOT mux_3649_nl) AND and_dcpl_932;
        reg_x_rsc_29_0_i_oswt_cse <= mux_3650_nl AND and_dcpl_927;
        reg_x_rsc_29_0_i_oswt_1_cse <= (NOT mux_3651_nl) AND and_dcpl_932;
        reg_x_rsc_30_0_i_oswt_cse <= mux_3652_nl AND and_dcpl_927;
        reg_x_rsc_30_0_i_oswt_1_cse <= (NOT mux_3653_nl) AND and_dcpl_932;
        reg_x_rsc_31_0_i_oswt_cse <= mux_3654_nl AND and_dcpl_927;
        reg_x_rsc_31_0_i_oswt_1_cse <= mux_3655_nl AND and_dcpl_932;
        reg_x_rsc_triosy_31_0_obj_iswt0_cse <= nor_tmp_3 AND (NOT (fsm_output(2)))
            AND and_dcpl_1000 AND and_2881_cse AND (fsm_output(7)) AND (z_out(5));
        reg_ensig_cgo_cse <= and_1109_rmff;
        reg_ensig_cgo_1_cse <= NOT mux_3669_itm;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_9_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_9_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_8_itm_mx0w1, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_9_nl,
            STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_93 & and_dcpl_77));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_19_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_19_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_11_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_19_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1096 & and_dcpl_93 & and_dcpl_77));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_23_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_23_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_17_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_23_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1096 & and_dcpl_93 & and_dcpl_77));
        reg_modulo_add_3_slc_32_svs_st_cse <= acc_15_nl(33);
        reg_modulo_add_2_slc_32_svs_st_cse <= acc_17_nl(33);
        reg_modulo_add_1_slc_32_svs_st_cse <= acc_19_nl(33);
        reg_modulo_add_7_slc_32_svs_st_cse <= acc_20_nl(33);
        reg_modulo_add_6_slc_32_svs_st_cse <= acc_21_nl(33);
        reg_modulo_add_5_slc_32_svs_st_cse <= acc_18_nl(33);
        reg_modulo_add_11_slc_32_svs_st_cse <= acc_22_nl(33);
        modulo_add_13_slc_32_svs_st <= modulo_add_13_acc_1_nl(32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND ((NOT (S1_OUTER_LOOP_k_5_0_sva_2(5))) OR (S2_INNER_LOOP1_r_4_0_sva_2(4))
          OR operator_20_true_8_slc_operator_20_true_8_acc_14_itm)) = '1' ) THEN
        S34_OUTER_LOOP_for_k_slc_S34_OUTER_LOOP_for_k_sva_19_5_4_0_1 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
            (S1_OUTER_LOOP_for_p_sva_1(9 DOWNTO 5)), and_1112_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg <= '0';
      ELSIF ( ((NOT mux_4278_nl) AND core_wen) = '1' ) THEN
        reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg <= S2_COPY_LOOP_p_asn_S2_COPY_LOOP_p_5_0_sva_4_0_S1_OUTER_LOOP_k_and_rgt(4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( ((NOT mux_4293_nl) AND core_wen) = '1' ) THEN
        reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg <= S2_COPY_LOOP_p_asn_S2_COPY_LOOP_p_5_0_sva_4_0_S1_OUTER_LOOP_k_and_rgt(3
            DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S2_COPY_LOOP_for_i_5_0_sva_1_5 <= '0';
      ELSIF ( (mux_4303_nl AND core_wen) = '1' ) THEN
        S2_COPY_LOOP_for_i_5_0_sva_1_5 <= S2_COPY_LOOP_for_i_mux1h_2_rgt(5);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_S2_COPY_LOOP_for_i_5_0_1_reg <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (mux_4318_nl AND core_wen) = '1' ) THEN
        reg_S2_COPY_LOOP_for_i_5_0_1_reg <= S2_COPY_LOOP_for_i_mux1h_2_rgt(4 DOWNTO
            3);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_S2_COPY_LOOP_for_i_5_0_2_reg <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( ((NOT mux_4334_nl) AND core_wen) = '1' ) THEN
        reg_S2_COPY_LOOP_for_i_5_0_2_reg <= S2_COPY_LOOP_for_i_mux1h_2_rgt(2 DOWNTO
            0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_p_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000");
      ELSIF ( (core_wen AND (and_dcpl_1082 OR S1_OUTER_LOOP_for_p_sva_1_mx0c1 OR
          and_dcpl_1084)) = '1' ) THEN
        S1_OUTER_LOOP_for_p_sva_1 <= MUX_v_20_2_2(z_out_26, (STD_LOGIC_VECTOR'( "00000")
            & S2_INNER_LOOP1_S2_INNER_LOOP1_and_nl), S1_OUTER_LOOP_for_p_sva_1_mx0c1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( operator_20_true_1_and_cse = '1' ) THEN
        operator_20_true_1_slc_operator_20_true_1_acc_14_itm <= z_out_16_14;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_33_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_35_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_36_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_37_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_39_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_40_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_41_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_42_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_43_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_44_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_47_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_49_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_51_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_55_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58_itm <= '0';
      ELSIF ( operator_20_true_1_and_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_33_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_35_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_36_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_37_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_39_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_40_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_41_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_42_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_43_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_44_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_47_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_49_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_51_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_55_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm_mx0w0;
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_acc_svs_4 <= '0';
      ELSIF ( ((NOT mux_4361_nl) AND core_wen) = '1' ) THEN
        S1_OUTER_LOOP_for_acc_svs_4 <= S34_OUTER_LOOP_for_a_and_rgt(4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_acc_svs_3_0 <= STD_LOGIC_VECTOR'( "0000");
      ELSIF ( (mux_4373_nl AND core_wen) = '1' ) THEN
        S1_OUTER_LOOP_for_acc_svs_3_0 <= S34_OUTER_LOOP_for_a_and_rgt(3 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_1_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_60_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_61_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_1_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_1_itm <= MUX1HOT_s_1_3_2(S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_nor_itm_mx0w0,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_9_itm_mx0w1, nor_2152_cse, STD_LOGIC_VECTOR'(
            and_dcpl_1091 & and_dcpl_93 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_60_itm <= MUX1HOT_s_1_3_2(S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_29_itm_mx0w0,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_4_itm_mx0w1, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_60_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1091 & and_dcpl_93 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_61_itm <= MUX1HOT_s_1_3_2(and_1344_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_5_itm_mx0w1, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_61_cse,
            STD_LOGIC_VECTOR'( and_dcpl_1091 & and_dcpl_93 & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_nor_25_itm <= '0';
        S1_OUTER_LOOP_for_nor_26_itm <= '0';
        S1_OUTER_LOOP_for_nor_39_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_6_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_2_cse = '1' ) THEN
        S1_OUTER_LOOP_for_nor_25_itm <= MUX1HOT_s_1_3_2(S34_OUTER_LOOP_for_a_nor_itm_mx0w0,
            S34_OUTER_LOOP_for_a_nor_1_itm_mx0w1, S6_OUTER_LOOP_for_nor_25_nl, STD_LOGIC_VECTOR'(
            and_dcpl_1091 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_nor_26_itm <= MUX1HOT_s_1_3_2(S34_OUTER_LOOP_for_a_nor_1_itm_mx0w1,
            S34_OUTER_LOOP_for_a_nor_14_itm_mx0w1, S6_OUTER_LOOP_for_nor_26_nl, STD_LOGIC_VECTOR'(
            and_dcpl_1091 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_nor_39_itm <= MUX1HOT_s_1_3_2(S34_OUTER_LOOP_for_a_nor_14_itm_mx0w1,
            S34_OUTER_LOOP_for_a_nor_itm_mx0w0, S6_OUTER_LOOP_for_nor_39_nl, STD_LOGIC_VECTOR'(
            and_dcpl_1091 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_6_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_6_itm_mx0w0,
            and_1329_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_6_nl, STD_LOGIC_VECTOR'(
            and_dcpl_1091 & and_dcpl_1092 & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_nor_28_itm <= '0';
        S1_OUTER_LOOP_for_nor_32_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_5_cse = '1' ) THEN
        S1_OUTER_LOOP_for_nor_28_itm <= MUX_s_1_2_2(S34_OUTER_LOOP_for_a_nor_3_nl,
            S6_OUTER_LOOP_for_nor_28_nl, and_dcpl_1084);
        S1_OUTER_LOOP_for_nor_32_itm <= MUX_s_1_2_2(S34_OUTER_LOOP_for_a_nor_7_nl,
            S6_OUTER_LOOP_for_nor_32_nl, and_dcpl_1084);
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_itm <= MUX_s_1_2_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_nor_itm_mx0w1,
            S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_nor_nl, and_dcpl_1084);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_45_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_53_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_57_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_16_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_45_itm <= MUX1HOT_s_1_4_2(and_1532_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_5_itm_mx0w1, S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_25_itm_mx0w2,
            S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_45_nl, STD_LOGIC_VECTOR'( and_dcpl_1091
            & and_dcpl_1088 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_53_itm <= MUX1HOT_s_1_4_2(and_1447_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_8_itm_mx0w1, S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_27_itm_mx0w2,
            S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_53_nl, STD_LOGIC_VECTOR'( and_dcpl_1091
            & and_dcpl_1088 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_57_itm <= MUX1HOT_s_1_4_2(and_1403_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_9_itm_mx0w1, and_1366_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_57_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1091 & and_dcpl_1088 & and_dcpl_1092 & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_59_itm <= '0';
      ELSIF ( (core_wen AND (and_dcpl_1091 OR and_dcpl_88 OR and_dcpl_1092 OR and_dcpl_1084))
          = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_59_itm <= MUX1HOT_s_1_4_2(and_1373_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_nor_itm_mx0w1, and_1350_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_59_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1091 & and_dcpl_88 & and_dcpl_1092 & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_nor_itm <= '0';
        S1_OUTER_LOOP_for_nor_1_itm <= '0';
        S1_OUTER_LOOP_for_nor_3_itm <= '0';
        S1_OUTER_LOOP_for_nor_7_itm <= '0';
        S1_OUTER_LOOP_for_nor_14_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_34_cse = '1' ) THEN
        S1_OUTER_LOOP_for_nor_itm <= MUX_s_1_2_2(S2_COPY_LOOP_for_nor_nl, S6_OUTER_LOOP_for_nor_nl,
            and_dcpl_1084);
        S1_OUTER_LOOP_for_nor_1_itm <= MUX_s_1_2_2(S2_COPY_LOOP_for_nor_1_nl, S6_OUTER_LOOP_for_nor_1_nl,
            and_dcpl_1084);
        S1_OUTER_LOOP_for_nor_3_itm <= MUX_s_1_2_2(S2_COPY_LOOP_for_nor_3_nl, S6_OUTER_LOOP_for_nor_3_nl,
            and_dcpl_1084);
        S1_OUTER_LOOP_for_nor_7_itm <= MUX_s_1_2_2(S2_COPY_LOOP_for_nor_7_nl, S6_OUTER_LOOP_for_nor_7_nl,
            and_dcpl_1084);
        S1_OUTER_LOOP_for_nor_14_itm <= MUX_s_1_2_2(S2_COPY_LOOP_for_nor_14_nl, S6_OUTER_LOOP_for_nor_14_nl,
            and_dcpl_1084);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_39_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_10_itm_mx0w0,
            butterFly_7_f1_butterFly_7_f1_nor_nl, and_1532_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_10_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & not_tmp_1436 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_12_itm_mx0w0,
            butterFly_7_f1_butterFly_7_f1_and_4_nl, and_1403_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_12_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & not_tmp_1436 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_13_itm_mx0w0,
            butterFly_7_f1_butterFly_7_f1_and_5_nl, and_1373_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_13_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & not_tmp_1436 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_14_itm_mx0w0,
            and_1380_cse, S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_29_itm_mx0w0,
            and_1919_cse, STD_LOGIC_VECTOR'( and_dcpl_1095 & not_tmp_1436 & and_dcpl_1092
            & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_18_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_20_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_21_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_24_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_27_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_28_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_29_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_44_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_18_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_18_itm_mx0w0,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_10_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_18_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_20_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_20_itm_mx0w0,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_13_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_20_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_21_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_21_itm_mx0w0,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_14_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_21_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_24_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_24_itm_mx0w0,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_18_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_24_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_27_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_27_itm_mx0w2,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_20_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_27_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_28_itm <= MUX1HOT_s_1_3_2(and_1366_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_21_itm_mx0w0, and_1740_cse, STD_LOGIC_VECTOR'(
            and_dcpl_1095 & and_dcpl_1092 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_29_itm <= MUX1HOT_s_1_3_2(and_1350_cse,
            and_1435_cse, and_1721_cse, STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_1092
            & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_22_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_25_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_26_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_30_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_47_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_22_itm <= MUX1HOT_s_1_3_2(and_1435_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_16_itm_mx0w1, and_1827_cse, STD_LOGIC_VECTOR'(
            and_dcpl_1095 & and_dcpl_93 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_25_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_25_itm_mx0w2,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_19_itm_mx0w1, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_25_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1095 & and_dcpl_93 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_26_itm <= MUX1HOT_s_1_3_2(and_1391_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_2_itm_mx0w1, and_1773_cse, STD_LOGIC_VECTOR'(
            and_dcpl_1095 & and_dcpl_93 & and_dcpl_1084));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_30_itm <= MUX1HOT_s_1_3_2(and_1329_cse,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_23_itm_mx0w1, and_1692_cse, STD_LOGIC_VECTOR'(
            and_dcpl_1095 & and_dcpl_93 & and_dcpl_1084));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_2_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_4_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_55_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_2_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_2_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_12_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_2_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1096 & and_dcpl_1092 & and_dcpl_77));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_4_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_4_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_24_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_4_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1096 & and_dcpl_1092 & and_dcpl_77));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm <= '0';
      ELSIF ( (core_wen AND (and_dcpl_934 OR and_dcpl_88 OR and_dcpl_1092 OR and_dcpl_77))
          = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_5_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_6_itm_mx0w0, and_1391_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_5_nl,
            STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_88 & and_dcpl_1092 & and_dcpl_77));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_8_itm <= '0';
      ELSIF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1092 OR and_dcpl_77)) = '1'
          ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_8_itm <= MUX1HOT_s_1_3_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_8_itm_mx0w1,
            S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_6_itm_mx0w0, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_8_nl,
            STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_1092 & and_dcpl_77));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm <= '0';
      ELSIF ( (core_wen AND (and_dcpl_1096 OR not_tmp_1436 OR and_dcpl_1092 OR and_dcpl_77))
          = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_11_itm_mx0w0,
            butterFly_7_f1_butterFly_7_f1_and_2_nl, and_1447_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_11_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1096 & not_tmp_1436 & and_dcpl_1092 & and_dcpl_77));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm <= '0';
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm <= '0';
      ELSIF ( S1_OUTER_LOOP_for_and_60_cse = '1' ) THEN
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_16_itm_mx0w1,
            butterFly_4_f1_butterFly_4_f1_nor_cse, and_1344_cse, S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_16_nl,
            STD_LOGIC_VECTOR'( and_dcpl_1096 & and_dcpl_1097 & and_dcpl_1092 & and_dcpl_77));
        S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm <= MUX1HOT_s_1_4_2(S2_COPY_LOOP_for_S2_COPY_LOOP_for_and_17_itm_mx0w0,
            butterFly_4_f1_butterFly_4_f1_and_2_nl, S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_nor_itm_mx0w0,
            S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_17_nl, STD_LOGIC_VECTOR'( and_dcpl_1096
            & and_dcpl_1097 & and_dcpl_1092 & and_dcpl_77));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR modulo_add_base_1_sva_mx0c3
          OR modulo_add_base_1_sva_mx0c4 OR and_dcpl_479 OR and_dcpl_556 OR and_dcpl_540
          OR and_dcpl_1105 OR modulo_add_base_1_sva_mx0c9 OR and_dcpl_102 OR and_dcpl_184
          OR and_dcpl_171 OR and_dcpl_1115 OR modulo_add_base_1_sva_mx0c14 OR and_dcpl_459
          OR and_dcpl_552 OR and_dcpl_534 OR modulo_add_base_1_sva_mx0c18 OR and_dcpl_1108
          OR and_dcpl_1109 OR modulo_add_base_1_sva_mx0c21 OR and_dcpl_129 OR and_dcpl_191
          OR and_dcpl_179 OR and_dcpl_1110 OR modulo_add_base_1_sva_mx0c26 OR and_dcpl_480
          OR and_dcpl_557 OR and_dcpl_541 OR modulo_add_base_1_sva_mx0c30 OR and_dcpl_131
          OR and_dcpl_192 OR and_dcpl_180)) = '1' ) THEN
        modulo_add_base_1_sva <= MUX1HOT_v_32_34_2(x_rsc_11_0_i_s_din_mxwt, (yy_rsc_11_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_1_0_i_qa_d(31 DOWNTO 0)), (mult_z_mul_cmp_z(31 DOWNTO
            0)), modulo_add_base_3_sva_mx0w4, modulo_add_base_2_sva_mx0w5, modulo_add_base_1_sva_mx0w6,
            modulo_add_base_sva_mx0w7, (yy_rsc_1_0_i_qa_d(31 DOWNTO 0)), modulo_add_base_7_sva_mx0w9,
            modulo_add_base_6_sva_mx0w10, modulo_add_base_5_sva_mx0w11, modulo_add_base_4_sva_mx0w12,
            (xx_rsc_2_0_i_qa_d(31 DOWNTO 0)), modulo_add_base_11_sva_mx0w14, modulo_add_base_10_sva_mx0w15,
            modulo_add_base_9_sva_mx0w16, modulo_add_base_8_sva_mx0w17, mult_12_z_mul_cmp_z,
            (xx_rsc_11_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_1_0_i_qa_d(63 DOWNTO 32)),
            modulo_add_base_15_sva_mx0w21, modulo_add_base_14_sva_mx0w22, modulo_add_base_13_sva_mx0w23,
            modulo_add_base_12_sva_mx0w24, (xx_rsc_1_0_i_qa_d(63 DOWNTO 32)), modulo_add_base_19_sva_mx0w26,
            modulo_add_base_18_sva_mx0w27, modulo_add_base_17_sva_mx0w28, modulo_add_base_16_sva_mx0w29,
            modulo_add_base_23_sva_mx0w30, modulo_add_base_22_sva_mx0w31, modulo_add_base_21_sva_mx0w32,
            modulo_add_base_20_sva_mx0w33, STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_1101
            & and_dcpl_1114 & modulo_add_base_1_sva_mx0c3 & modulo_add_base_1_sva_mx0c4
            & and_dcpl_479 & and_dcpl_556 & and_dcpl_540 & and_dcpl_1105 & modulo_add_base_1_sva_mx0c9
            & and_dcpl_102 & and_dcpl_184 & and_dcpl_171 & and_dcpl_1115 & modulo_add_base_1_sva_mx0c14
            & and_dcpl_459 & and_dcpl_552 & and_dcpl_534 & modulo_add_base_1_sva_mx0c18
            & and_dcpl_1108 & and_dcpl_1109 & modulo_add_base_1_sva_mx0c21 & and_dcpl_129
            & and_dcpl_191 & and_dcpl_179 & and_dcpl_1110 & modulo_add_base_1_sva_mx0c26
            & and_dcpl_480 & and_dcpl_557 & and_dcpl_541 & modulo_add_base_1_sva_mx0c30
            & and_dcpl_131 & and_dcpl_192 & and_dcpl_180));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3
          OR not_tmp_1349 OR and_dcpl_1105 OR and_dcpl_1115 OR mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c7
          OR and_dcpl_1108 OR and_dcpl_1109 OR and_dcpl_1110)) = '1' ) THEN
        mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm <= MUX1HOT_v_32_11_2(x_rsc_13_0_i_s_din_mxwt,
            (yy_rsc_13_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_5_0_i_qa_d(31 DOWNTO 0)),
            (mult_z_mul_cmp_z(51 DOWNTO 20)), (mult_z_mul_cmp_z(31 DOWNTO 0)), (yy_rsc_5_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_6_0_i_qa_d(31 DOWNTO 0)), mult_12_z_mul_cmp_z, (xx_rsc_13_0_i_qa_d(31
            DOWNTO 0)), (yy_rsc_5_0_i_qa_d(63 DOWNTO 32)), (xx_rsc_5_0_i_qa_d(63
            DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_1101 & and_dcpl_1114
            & mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3 & not_tmp_1349 & and_dcpl_1105
            & and_dcpl_1115 & mult_10_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c7 & and_dcpl_1108
            & and_dcpl_1109 & and_dcpl_1110));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3
          OR and_dcpl_1105 OR and_dcpl_1115 OR and_dcpl_1108 OR and_dcpl_1109 OR
          and_dcpl_1110)) = '1' ) THEN
        mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm <= MUX1HOT_v_32_9_2(x_rsc_14_0_i_s_din_mxwt,
            (yy_rsc_14_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_9_0_i_qa_d(31 DOWNTO 0)),
            (mult_z_mul_cmp_z(31 DOWNTO 0)), (yy_rsc_9_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_10_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_14_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_9_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_9_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1114 & mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1108 & and_dcpl_1109 & and_dcpl_1110));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3
          OR and_dcpl_1105 OR and_dcpl_1115 OR and_dcpl_1108 OR and_dcpl_1109 OR
          and_dcpl_1110)) = '1' ) THEN
        mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm <= MUX1HOT_v_32_9_2(x_rsc_15_0_i_s_din_mxwt,
            (yy_rsc_15_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_13_0_i_qa_d(31 DOWNTO 0)),
            (mult_z_mul_cmp_z(31 DOWNTO 0)), (yy_rsc_13_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_14_0_i_qa_d(31
            DOWNTO 0)), (xx_rsc_15_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_13_0_i_qa_d(63
            DOWNTO 32)), (xx_rsc_13_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934
            & and_dcpl_1101 & and_dcpl_1114 & mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm_mx0c3
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1108 & and_dcpl_1109 & and_dcpl_1110));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm_mx0c3
          OR and_dcpl_1105 OR and_dcpl_1115 OR and_dcpl_1108 OR and_dcpl_1109 OR
          and_dcpl_1110)) = '1' ) THEN
        operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm <=
            MUX1HOT_v_32_9_2(x_rsc_16_0_i_s_din_mxwt, (yy_rsc_16_0_i_qa_d(31 DOWNTO
            0)), (xx_rsc_17_0_i_qa_d(31 DOWNTO 0)), (mult_z_mul_cmp_z(51 DOWNTO 20)),
            (yy_rsc_17_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_18_0_i_qa_d(31 DOWNTO 0)),
            (xx_rsc_16_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_17_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_17_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934 &
            and_dcpl_1101 & and_dcpl_1114 & operator_96_false_10_operator_96_false_10_slc_mult_10_t_mul_51_20_itm_mx0c3
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1108 & and_dcpl_1109 & and_dcpl_1110));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm_mx0c3
          OR and_dcpl_1105 OR and_dcpl_1115 OR and_dcpl_1108 OR and_dcpl_1109 OR
          and_dcpl_1110)) = '1' ) THEN
        operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm <=
            MUX1HOT_v_32_9_2(x_rsc_19_0_i_s_din_mxwt, (yy_rsc_19_0_i_qa_d(31 DOWNTO
            0)), (xx_rsc_21_0_i_qa_d(31 DOWNTO 0)), (mult_z_mul_cmp_z(51 DOWNTO 20)),
            (yy_rsc_21_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_22_0_i_qa_d(31 DOWNTO 0)),
            (xx_rsc_19_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_21_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_21_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934 &
            and_dcpl_1101 & and_dcpl_1114 & operator_96_false_16_operator_96_false_16_slc_mult_16_t_mul_51_20_itm_mx0c3
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1108 & and_dcpl_1109 & and_dcpl_1110));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (and_dcpl_934 OR and_dcpl_1101 OR and_dcpl_1114 OR operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm_mx0c3
          OR and_dcpl_1105 OR and_dcpl_1115 OR and_dcpl_1108 OR and_dcpl_1109 OR
          and_dcpl_1110)) = '1' ) THEN
        operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm <=
            MUX1HOT_v_32_9_2(x_rsc_2_0_i_s_din_mxwt, (yy_rsc_2_0_i_qa_d(31 DOWNTO
            0)), (xx_rsc_25_0_i_qa_d(31 DOWNTO 0)), (mult_z_mul_cmp_z(51 DOWNTO 20)),
            (yy_rsc_25_0_i_qa_d(31 DOWNTO 0)), (xx_rsc_26_0_i_qa_d(31 DOWNTO 0)),
            (xx_rsc_2_0_i_qa_d(31 DOWNTO 0)), (yy_rsc_25_0_i_qa_d(63 DOWNTO 32)),
            (xx_rsc_25_0_i_qa_d(63 DOWNTO 32)), STD_LOGIC_VECTOR'( and_dcpl_934 &
            and_dcpl_1101 & and_dcpl_1114 & operator_96_false_17_operator_96_false_17_slc_mult_17_t_mul_51_20_itm_mx0c3
            & and_dcpl_1105 & and_dcpl_1115 & and_dcpl_1108 & and_dcpl_1109 & and_dcpl_1110));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( S2_INNER_LOOP1_tf_and_1_cse = '1' ) THEN
        S2_INNER_LOOP1_tf_sva <= MUX1HOT_v_32_4_2(x_rsc_0_0_i_s_din_mxwt, (yy_rsc_0_0_i_qa_d(31
            DOWNTO 0)), twiddle_rsci_qb_d_mxwt, (xx_rsc_0_0_i_qa_d(31 DOWNTO 0)),
            STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_1101 & not_tmp_1520 & and_dcpl_1108));
        S2_INNER_LOOP1_tfh_sva <= MUX1HOT_v_32_4_2(x_rsc_1_0_i_s_din_mxwt, (yy_rsc_1_0_i_qa_d(31
            DOWNTO 0)), twiddle_h_rsci_qb_d_mxwt, (xx_rsc_1_0_i_qa_d(31 DOWNTO 0)),
            STD_LOGIC_VECTOR'( and_dcpl_934 & and_dcpl_1101 & not_tmp_1520 & and_dcpl_1108));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_drf_revArr_ptr_1_smx_9_0_reg <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (mux_4391_nl AND core_wen) = '1' ) THEN
        reg_drf_revArr_ptr_1_smx_9_0_reg <= S2_COPY_LOOP_for_S2_COPY_LOOP_for_mux_6_rgt(4
            DOWNTO 3);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_drf_revArr_ptr_1_smx_9_0_1_reg <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (mux_4397_nl AND core_wen) = '1' ) THEN
        reg_drf_revArr_ptr_1_smx_9_0_1_reg <= S2_COPY_LOOP_for_S2_COPY_LOOP_for_mux_6_rgt(2
            DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S2_OUTER_LOOP_c_1_sva <= '0';
      ELSIF ( (core_wen AND (((NOT mux_tmp_3812) AND and_dcpl_1085 AND and_dcpl_79)
          OR S2_OUTER_LOOP_c_1_sva_mx0c1 OR S2_OUTER_LOOP_c_1_sva_mx0c2)) = '1' )
          THEN
        S2_OUTER_LOOP_c_1_sva <= (S2_OUTER_LOOP_c_1_sva OR (S2_INNER_LOOP1_r_4_0_sva_2(4)))
            AND (S2_OUTER_LOOP_c_1_sva_mx0c1 OR S2_OUTER_LOOP_c_1_sva_mx0c2);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_4404_nl AND core_wen) = '1' ) THEN
        operator_33_true_return_2_3_0_sva_3 <= z_out_3(3);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (mux_4410_nl AND core_wen) = '1' ) THEN
        operator_33_true_return_2_3_0_sva_2_0 <= z_out_3(2 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly_f1_and_cse = '1' ) THEN
        tmp_lpi_4_dfm <= tmp_lpi_4_dfm_mx0w0;
        tmp_2_lpi_4_dfm <= tmp_2_lpi_4_dfm_mx0w0;
        tmp_4_lpi_4_dfm <= tmp_4_lpi_4_dfm_mx0w0;
        tmp_6_lpi_4_dfm <= tmp_6_lpi_4_dfm_mx0w0;
        tmp_1_lpi_4_dfm <= tmp_1_lpi_4_dfm_mx0w0;
        tmp_3_lpi_4_dfm <= tmp_3_lpi_4_dfm_mx0w0;
        tmp_5_lpi_4_dfm <= tmp_5_lpi_4_dfm_mx0w0;
        tmp_7_lpi_4_dfm <= tmp_7_lpi_4_dfm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly_4_f1_and_cse = '1' ) THEN
        tmp_28_lpi_4_dfm <= tmp_2_lpi_4_dfm_mx0w0;
        tmp_30_lpi_4_dfm <= tmp_4_lpi_4_dfm_mx0w0;
        tmp_32_lpi_4_dfm <= tmp_lpi_4_dfm_mx0w0;
        tmp_34_lpi_4_dfm <= tmp_6_lpi_4_dfm_mx0w0;
        tmp_29_lpi_4_dfm <= tmp_1_lpi_4_dfm_mx0w0;
        tmp_31_lpi_4_dfm <= tmp_3_lpi_4_dfm_mx0w0;
        tmp_33_lpi_4_dfm <= tmp_5_lpi_4_dfm_mx0w0;
        tmp_35_lpi_4_dfm <= tmp_7_lpi_4_dfm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly_8_f1_and_cse = '1' ) THEN
        tmp_8_lpi_3_dfm <= tmp_lpi_4_dfm_mx0w0;
        tmp_10_lpi_3_dfm <= tmp_2_lpi_4_dfm_mx0w0;
        tmp_12_lpi_3_dfm <= tmp_4_lpi_4_dfm_mx0w0;
        tmp_14_lpi_3_dfm <= tmp_6_lpi_4_dfm_mx0w0;
        tmp_9_lpi_3_dfm <= tmp_5_lpi_4_dfm_mx0w0;
        tmp_11_lpi_3_dfm <= tmp_1_lpi_4_dfm_mx0w0;
        tmp_13_lpi_3_dfm <= tmp_3_lpi_4_dfm_mx0w0;
        tmp_15_lpi_3_dfm <= tmp_7_lpi_4_dfm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( operator_20_true_8_and_cse = '1' ) THEN
        operator_20_true_8_slc_operator_20_true_8_acc_14_itm <= z_out_16_14;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm <= '0';
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm <= '0';
      ELSIF ( operator_20_true_8_and_cse = '1' ) THEN
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_2_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_4_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_5_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_6_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_8_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_9_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_10_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_11_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_12_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_13_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_16_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_17_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_18_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_19_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_20_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_21_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_23_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_24_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_25_itm_mx0w0;
        S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm <= S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_27_itm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly_12_f1_and_cse = '1' ) THEN
        tmp_38_lpi_4_dfm <= tmp_2_lpi_4_dfm_mx0w0;
        tmp_40_lpi_4_dfm <= tmp_4_lpi_4_dfm_mx0w0;
        tmp_42_lpi_4_dfm <= tmp_lpi_4_dfm_mx0w0;
        tmp_44_lpi_4_dfm <= tmp_6_lpi_4_dfm_mx0w0;
        tmp_39_lpi_4_dfm <= tmp_1_lpi_4_dfm_mx0w0;
        tmp_41_lpi_4_dfm <= tmp_3_lpi_4_dfm_mx0w0;
        tmp_43_lpi_4_dfm <= tmp_5_lpi_4_dfm_mx0w0;
        tmp_45_lpi_4_dfm <= tmp_7_lpi_4_dfm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly_16_f1_and_cse = '1' ) THEN
        tmp_17_lpi_4_dfm <= tmp_2_lpi_4_dfm_mx0w0;
        tmp_19_lpi_4_dfm <= tmp_4_lpi_4_dfm_mx0w0;
        tmp_21_lpi_4_dfm <= tmp_lpi_4_dfm_mx0w0;
        tmp_23_lpi_4_dfm <= tmp_6_lpi_4_dfm_mx0w0;
        tmp_18_lpi_4_dfm <= tmp_1_lpi_4_dfm_mx0w0;
        tmp_20_lpi_4_dfm <= tmp_3_lpi_4_dfm_mx0w0;
        tmp_22_lpi_4_dfm <= tmp_5_lpi_4_dfm_mx0w0;
        tmp_24_lpi_4_dfm <= tmp_7_lpi_4_dfm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly_20_f1_and_cse = '1' ) THEN
        tmp_46_lpi_3_dfm <= tmp_2_lpi_4_dfm_mx0w0;
        tmp_48_lpi_3_dfm <= tmp_4_lpi_4_dfm_mx0w0;
        tmp_50_lpi_3_dfm <= tmp_lpi_4_dfm_mx0w0;
        tmp_52_lpi_3_dfm <= tmp_6_lpi_4_dfm_mx0w0;
        tmp_47_lpi_3_dfm <= tmp_1_lpi_4_dfm_mx0w0;
        tmp_49_lpi_3_dfm <= tmp_3_lpi_4_dfm_mx0w0;
        tmp_51_lpi_3_dfm <= tmp_5_lpi_4_dfm_mx0w0;
        tmp_53_lpi_3_dfm <= tmp_7_lpi_4_dfm_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( operator_20_true_15_and_cse = '1' ) THEN
        operator_20_true_15_slc_operator_20_true_15_acc_14_itm <= z_out_16_14;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_33_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_35_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_36_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_37_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_39_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_40_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_41_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_42_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_43_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_44_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_47_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_48_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_49_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_50_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_51_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_52_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_54_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_55_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_56_itm <= '0';
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_58_itm <= '0';
      ELSIF ( operator_20_true_15_and_cse = '1' ) THEN
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_33_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("00011"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_35_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("00101"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_36_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("00110"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_37_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("00111"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_39_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01001"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_40_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01010"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_41_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01011"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_42_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01100"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_43_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01101"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_44_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01110"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_47_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10001"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_48_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10010"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_49_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10011"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_50_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10100"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_51_itm <= (S6_OUTER_LOOP_for_acc_tmp(4))
            AND (S6_OUTER_LOOP_for_acc_tmp(2)) AND (S6_OUTER_LOOP_for_acc_tmp(0))
            AND S6_OUTER_LOOP_for_nor_44_cse;
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_52_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10110"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_54_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11000"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_55_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11001"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_56_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11010"));
        S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_58_itm <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11100"));
      END IF;
    END IF;
  END PROCESS;
  nor_2174_nl <= NOT(CONV_SL_1_1(fsm_output(6 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000000")));
  or_285_nl <= (fsm_output(6)) OR and_1306_cse;
  mux_102_nl <= MUX_s_1_2_2((fsm_output(6)), or_285_nl, fsm_output(5));
  mux_101_nl <= MUX_s_1_2_2((fsm_output(6)), or_4376_cse, fsm_output(5));
  mux_103_nl <= MUX_s_1_2_2(mux_102_nl, mux_101_nl, fsm_output(3));
  mux_104_nl <= MUX_s_1_2_2(nor_2174_nl, mux_103_nl, fsm_output(7));
  nor_1463_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR (S1_OUTER_LOOP_for_acc_svs_3_0(2))
      OR (NOT (fsm_output(1))));
  nor_1464_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3592_nl <= MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output(0));
  mux_3593_nl <= MUX_s_1_2_2(or_309_cse, or_dcpl_180, fsm_output(0));
  S1_OUTER_LOOP_for_and_62_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_itm AND
      (NOT and_dcpl_935);
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_nl <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))
      AND S1_OUTER_LOOP_for_nor_itm AND (NOT and_dcpl_935);
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_1_nl <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1))
      AND S1_OUTER_LOOP_for_nor_1_itm AND (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_63_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_2_itm AND
      (NOT and_dcpl_935);
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_3_nl <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      AND S1_OUTER_LOOP_for_nor_3_itm AND (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_64_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_4_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_65_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_66_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_6_itm AND
      (NOT and_dcpl_935);
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_7_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND S1_OUTER_LOOP_for_nor_7_itm AND (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_67_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_8_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_68_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_9_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_69_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_10_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_70_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_11_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_71_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_12_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_72_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_13_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_73_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_14_itm AND
      (NOT and_dcpl_935);
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_15_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND S1_OUTER_LOOP_for_nor_14_itm AND (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_74_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_16_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_75_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_17_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_76_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_18_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_77_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_19_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_78_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_20_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_79_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_21_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_80_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_22_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_81_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_23_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_82_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_24_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_83_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_25_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_84_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_26_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_85_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_27_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_86_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_28_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_87_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_29_itm AND
      (NOT and_dcpl_935);
  S1_OUTER_LOOP_for_and_88_nl <= S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_30_itm AND
      (NOT and_dcpl_935);
  nor_1462_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3594_nl <= MUX_s_1_2_2(nor_2144_cse, nor_1462_nl, fsm_output(0));
  mux_3595_nl <= MUX_s_1_2_2(or_387_cse, or_dcpl_182, fsm_output(0));
  nor_1459_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR (S1_OUTER_LOOP_for_acc_svs_3_0(2))
      OR (NOT (fsm_output(1))));
  nor_1460_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3596_nl <= MUX_s_1_2_2(nor_1459_nl, nor_1460_nl, fsm_output(0));
  mux_3597_nl <= MUX_s_1_2_2(or_445_cse, or_dcpl_184, fsm_output(0));
  nor_1457_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR (S1_OUTER_LOOP_for_acc_svs_3_0(2))
      OR (NOT (fsm_output(1))));
  nor_1458_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3598_nl <= MUX_s_1_2_2(nor_1457_nl, nor_1458_nl, fsm_output(0));
  mux_3599_nl <= MUX_s_1_2_2(or_501_cse, or_dcpl_185, fsm_output(0));
  nor_1455_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR not_tmp_1278);
  nor_1456_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3600_nl <= MUX_s_1_2_2(nor_1455_nl, nor_1456_nl, fsm_output(0));
  mux_3601_nl <= MUX_s_1_2_2(or_549_cse, or_dcpl_188, fsm_output(0));
  nor_1453_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR not_tmp_1278);
  nor_1454_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3602_nl <= MUX_s_1_2_2(nor_1453_nl, nor_1454_nl, fsm_output(0));
  mux_3603_nl <= MUX_s_1_2_2(or_618_cse, or_dcpl_189, fsm_output(0));
  nor_1451_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR not_tmp_1278);
  nor_1452_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3604_nl <= MUX_s_1_2_2(nor_1451_nl, nor_1452_nl, fsm_output(0));
  mux_3605_nl <= MUX_s_1_2_2(or_682_cse, or_dcpl_191, fsm_output(0));
  nor_1449_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR S1_OUTER_LOOP_for_acc_svs_4 OR not_tmp_1278);
  nor_1450_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3606_nl <= MUX_s_1_2_2(nor_1449_nl, nor_1450_nl, fsm_output(0));
  mux_3607_nl <= MUX_s_1_2_2(or_735_cse, or_dcpl_192, fsm_output(0));
  nor_1447_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR S1_OUTER_LOOP_for_acc_svs_4
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1448_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3608_nl <= MUX_s_1_2_2(nor_1447_nl, nor_1448_nl, fsm_output(0));
  mux_3609_nl <= MUX_s_1_2_2(or_789_cse, or_dcpl_194, fsm_output(0));
  nor_1446_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3610_nl <= MUX_s_1_2_2(nor_2032_cse, nor_1446_nl, fsm_output(0));
  mux_3611_nl <= MUX_s_1_2_2(or_856_cse, or_dcpl_196, fsm_output(0));
  nor_1443_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR S1_OUTER_LOOP_for_acc_svs_4
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1444_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3612_nl <= MUX_s_1_2_2(nor_1443_nl, nor_1444_nl, fsm_output(0));
  mux_3613_nl <= MUX_s_1_2_2(or_908_cse, or_dcpl_197, fsm_output(0));
  nor_1441_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR S1_OUTER_LOOP_for_acc_svs_4
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1442_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3614_nl <= MUX_s_1_2_2(nor_1441_nl, nor_1442_nl, fsm_output(0));
  mux_3615_nl <= MUX_s_1_2_2(or_955_cse, or_dcpl_198, fsm_output(0));
  nor_1439_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR S1_OUTER_LOOP_for_acc_svs_4
      OR not_tmp_1278);
  nor_1440_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3616_nl <= MUX_s_1_2_2(nor_1439_nl, nor_1440_nl, fsm_output(0));
  mux_3617_nl <= MUX_s_1_2_2(or_1006_cse, or_dcpl_199, fsm_output(0));
  nor_1437_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR S1_OUTER_LOOP_for_acc_svs_4
      OR not_tmp_1278);
  nor_1438_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3618_nl <= MUX_s_1_2_2(nor_1437_nl, nor_1438_nl, fsm_output(0));
  mux_3619_nl <= MUX_s_1_2_2(or_1073_cse, or_dcpl_200, fsm_output(0));
  nor_1435_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR S1_OUTER_LOOP_for_acc_svs_4
      OR not_tmp_1278);
  nor_1436_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3620_nl <= MUX_s_1_2_2(nor_1435_nl, nor_1436_nl, fsm_output(0));
  mux_3621_nl <= MUX_s_1_2_2(or_1130_cse, or_dcpl_201, fsm_output(0));
  nor_1433_nl <= NOT((NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) AND (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND (S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND (NOT S1_OUTER_LOOP_for_acc_svs_4)))
      OR not_tmp_1278);
  nor_1434_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3622_nl <= MUX_s_1_2_2(nor_1433_nl, nor_1434_nl, fsm_output(0));
  mux_3623_nl <= MUX_s_1_2_2(nand_449_cse, or_dcpl_202, fsm_output(0));
  nor_1431_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1432_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3624_nl <= MUX_s_1_2_2(nor_1431_nl, nor_1432_nl, fsm_output(0));
  or_1283_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3625_nl <= MUX_s_1_2_2(or_1283_nl, or_dcpl_205, fsm_output(0));
  nor_1430_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3626_nl <= MUX_s_1_2_2(nor_1930_cse, nor_1430_nl, fsm_output(0));
  or_1340_nl <= (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3627_nl <= MUX_s_1_2_2(or_1340_nl, or_dcpl_206, fsm_output(0));
  nor_1427_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1428_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3628_nl <= MUX_s_1_2_2(nor_1427_nl, nor_1428_nl, fsm_output(0));
  or_1393_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3629_nl <= MUX_s_1_2_2(or_1393_nl, or_dcpl_208, fsm_output(0));
  nor_1425_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1426_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3630_nl <= MUX_s_1_2_2(nor_1425_nl, nor_1426_nl, fsm_output(0));
  or_1445_nl <= (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3631_nl <= MUX_s_1_2_2(or_1445_nl, or_dcpl_209, fsm_output(0));
  nor_1423_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_1311);
  nor_1424_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3632_nl <= MUX_s_1_2_2(nor_1423_nl, nor_1424_nl, fsm_output(0));
  or_1510_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_551;
  mux_3633_nl <= MUX_s_1_2_2(or_1510_nl, or_dcpl_212, fsm_output(0));
  nor_1421_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_1311);
  nor_1422_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3634_nl <= MUX_s_1_2_2(nor_1421_nl, nor_1422_nl, fsm_output(0));
  or_1578_nl <= (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_551;
  mux_3635_nl <= MUX_s_1_2_2(or_1578_nl, or_dcpl_213, fsm_output(0));
  nor_1419_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_1311);
  nor_1420_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3636_nl <= MUX_s_1_2_2(nor_1419_nl, nor_1420_nl, fsm_output(0));
  or_1638_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_551;
  mux_3637_nl <= MUX_s_1_2_2(or_1638_nl, or_dcpl_215, fsm_output(0));
  nor_1417_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_1311);
  nor_1418_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3638_nl <= MUX_s_1_2_2(nor_1417_nl, nor_1418_nl, fsm_output(0));
  or_1697_nl <= (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(3)) OR not_tmp_551;
  mux_3639_nl <= MUX_s_1_2_2(or_1697_nl, or_dcpl_216, fsm_output(0));
  nor_1415_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1416_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3640_nl <= MUX_s_1_2_2(nor_1415_nl, nor_1416_nl, fsm_output(0));
  or_1758_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3641_nl <= MUX_s_1_2_2(or_1758_nl, or_dcpl_217, fsm_output(0));
  nor_1413_nl <= NOT((NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1414_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3642_nl <= MUX_s_1_2_2(nor_1413_nl, nor_1414_nl, fsm_output(0));
  or_1814_nl <= (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(0))) OR (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3643_nl <= MUX_s_1_2_2(or_1814_nl, or_dcpl_218, fsm_output(0));
  nor_1411_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2)) OR (NOT (fsm_output(1))));
  nor_1412_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3644_nl <= MUX_s_1_2_2(nor_1411_nl, nor_1412_nl, fsm_output(0));
  or_1867_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(1)))
      OR (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(3))) OR (NOT S1_OUTER_LOOP_for_acc_svs_4)
      OR (S1_OUTER_LOOP_for_acc_svs_3_0(2));
  mux_3645_nl <= MUX_s_1_2_2(or_1867_nl, or_dcpl_219, fsm_output(0));
  and_2133_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) AND (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND (S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4 AND
      (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(2))) AND (fsm_output(1));
  nor_1410_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (fsm_output(1)));
  mux_3646_nl <= MUX_s_1_2_2(and_2133_nl, nor_1410_nl, fsm_output(0));
  nand_378_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) AND (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND (S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4 AND
      (NOT (S1_OUTER_LOOP_for_acc_svs_3_0(2))));
  mux_3647_nl <= MUX_s_1_2_2(nand_378_nl, or_dcpl_220, fsm_output(0));
  nor_1407_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR not_tmp_1328);
  nor_1408_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3648_nl <= MUX_s_1_2_2(nor_1407_nl, nor_1408_nl, fsm_output(0));
  or_1988_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))
      OR nand_517_cse;
  mux_3649_nl <= MUX_s_1_2_2(or_1988_nl, or_dcpl_221, fsm_output(0));
  nor_1405_nl <= NOT(CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR not_tmp_1328);
  nor_1406_nl <= NOT((NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0))) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3650_nl <= MUX_s_1_2_2(nor_1405_nl, nor_1406_nl, fsm_output(0));
  or_2042_nl <= CONV_SL_1_1(S1_OUTER_LOOP_for_acc_svs_3_0(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("01"))
      OR nand_517_cse;
  mux_3651_nl <= MUX_s_1_2_2(or_2042_nl, or_dcpl_222, fsm_output(0));
  nor_1403_nl <= NOT((S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR (NOT((S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND (S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4 AND
      (S1_OUTER_LOOP_for_acc_svs_3_0(2)) AND (fsm_output(1)))));
  nor_1404_nl <= NOT((reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)))
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))) OR (NOT reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg)
      OR (NOT (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2))) OR (fsm_output(1)));
  mux_3652_nl <= MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output(0));
  or_2091_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) OR nand_351_cse;
  mux_3653_nl <= MUX_s_1_2_2(or_2091_nl, or_dcpl_223, fsm_output(0));
  and_1324_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0)) AND (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND (S1_OUTER_LOOP_for_acc_svs_3_0(3)) AND S1_OUTER_LOOP_for_acc_svs_4 AND
      (S1_OUTER_LOOP_for_acc_svs_3_0(2)) AND (fsm_output(1));
  and_1325_nl <= (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)) AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3)) AND reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      AND (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) AND (NOT (fsm_output(1)));
  mux_3654_nl <= MUX_s_1_2_2(and_1324_nl, and_1325_nl, fsm_output(0));
  mux_3655_nl <= MUX_s_1_2_2(and_1713_cse, and_1692_cse, fsm_output(0));
  S34_OUTER_LOOP_for_tf_mux_1_nl <= MUX_v_5_2_2((reg_S2_COPY_LOOP_for_i_5_0_1_reg
      & reg_S2_COPY_LOOP_for_i_5_0_2_reg), (S1_OUTER_LOOP_k_5_0_sva_2(4 DOWNTO 0)),
      and_dcpl_1010);
  not_10627_nl <= NOT and_dcpl_1008;
  S34_OUTER_LOOP_for_k_mux_nl <= MUX_v_5_2_2((S1_OUTER_LOOP_for_p_sva_1(4 DOWNTO
      0)), (S1_OUTER_LOOP_k_5_0_sva_2(4 DOWNTO 0)), and_dcpl_1010);
  not_nl <= NOT and_dcpl_1008;
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_9_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_19_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_23_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND butterFly_4_f1_butterFly_4_f1_nor_cse;
  mux_3909_nl <= MUX_s_1_2_2((NOT (fsm_output(1))), (fsm_output(1)), fsm_output(5));
  and_1287_nl <= (fsm_output(3)) AND mux_3909_nl;
  mux_3910_nl <= MUX_s_1_2_2(and_1287_nl, nor_1311_cse, fsm_output(7));
  and_1222_nl <= mux_3910_nl AND and_dcpl_925 AND and_dcpl_1000;
  nor_1309_nl <= NOT((fsm_output(0)) OR (fsm_output(2)) OR (NOT (fsm_output(4))));
  nor_1310_nl <= NOT((NOT (fsm_output(0))) OR (fsm_output(2)) OR (fsm_output(4)));
  mux_3911_nl <= MUX_s_1_2_2(nor_1309_nl, nor_1310_nl, fsm_output(6));
  and_1286_nl <= (fsm_output(6)) AND (fsm_output(0)) AND (fsm_output(2)) AND (NOT
      (fsm_output(4)));
  mux_3912_nl <= MUX_s_1_2_2(mux_3911_nl, and_1286_nl, fsm_output(5));
  and_1225_nl <= mux_3912_nl AND (fsm_output(1)) AND (NOT (fsm_output(3))) AND (NOT
      (fsm_output(7)));
  nor_1307_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(0)));
  mux_3913_nl <= MUX_s_1_2_2(nor_1307_nl, nor_1308_cse, fsm_output(3));
  and_1229_nl <= mux_3913_nl AND (fsm_output(4)) AND nor_2178_cse_1 AND CONV_SL_1_1(fsm_output(7
      DOWNTO 6)=STD_LOGIC_VECTOR'("01"));
  and_1285_nl <= (fsm_output(5)) AND (fsm_output(2)) AND (fsm_output(1)) AND (fsm_output(4));
  nor_1306_nl <= NOT((fsm_output(5)) OR (fsm_output(2)) OR (fsm_output(1)) OR (fsm_output(4)));
  mux_3914_nl <= MUX_s_1_2_2(and_1285_nl, nor_1306_nl, fsm_output(3));
  and_1231_nl <= mux_3914_nl AND and_dcpl_1000 AND (fsm_output(7));
  S1_OUTER_LOOP_for_mux_25_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_nor_itm,
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_59_itm, and_dcpl_1165);
  S1_OUTER_LOOP_for_mux_26_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm,
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_45_itm, and_dcpl_1165);
  S1_OUTER_LOOP_for_mux_27_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_6_itm,
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_5_itm, and_dcpl_1165);
  S1_OUTER_LOOP_for_mux_28_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_8_itm,
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_53_itm, and_dcpl_1165);
  S1_OUTER_LOOP_for_mux_29_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_9_itm,
      S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_57_itm, and_dcpl_1165);
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_82_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0))
      AND S1_OUTER_LOOP_for_nor_25_itm;
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_83_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND S1_OUTER_LOOP_for_nor_26_itm;
  S1_OUTER_LOOP_for_mux_30_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_33_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_33_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_31_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_35_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_35_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_32_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_36_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_36_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_33_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_37_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_37_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_34_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_39_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_39_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_35_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_40_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_40_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_36_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_41_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_41_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_37_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_42_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_42_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_38_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_43_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_43_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_39_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_44_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_44_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_84_nl <= S1_OUTER_LOOP_for_acc_svs_4 AND
      S1_OUTER_LOOP_for_nor_39_itm;
  S1_OUTER_LOOP_for_mux_40_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_47_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_47_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_41_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_48_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_48_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_42_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_49_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_49_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_43_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_50_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_50_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_44_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_51_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_51_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_45_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_52_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_52_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_46_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_54_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_54_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_47_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_55_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_55_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_48_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_56_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_56_itm, and_dcpl_1178);
  S1_OUTER_LOOP_for_mux_49_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_S1_OUTER_LOOP_for_and_58_itm,
      S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_58_itm, and_dcpl_1178);
  mux_4091_nl <= MUX_s_1_2_2(and_1274_cse, nor_2412_cse, fsm_output(7));
  and_2897_nl <= (fsm_output(7)) AND (fsm_output(5)) AND (fsm_output(3)) AND (fsm_output(1))
      AND (fsm_output(2)) AND (NOT (fsm_output(0))) AND (NOT (fsm_output(6)));
  nor_2426_nl <= NOT((NOT (fsm_output(1))) OR (fsm_output(2)) OR (fsm_output(0))
      OR (NOT (fsm_output(6))));
  nor_2427_nl <= NOT((NOT (fsm_output(1))) OR (NOT (fsm_output(2))) OR (fsm_output(0))
      OR (fsm_output(6)));
  mux_4416_nl <= MUX_s_1_2_2(nor_2426_nl, nor_2427_nl, fsm_output(3));
  or_4856_nl <= (fsm_output(0)) OR (fsm_output(6));
  nand_573_nl <= NOT((fsm_output(0)) AND (fsm_output(6)));
  mux_4417_nl <= MUX_s_1_2_2(or_4856_nl, nand_573_nl, fsm_output(2));
  nor_2428_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(1)) OR mux_4417_nl);
  mux_4415_nl <= MUX_s_1_2_2(mux_4416_nl, nor_2428_nl, fsm_output(5));
  nor_2429_nl <= NOT((fsm_output(5)) OR (fsm_output(3)) OR (NOT (fsm_output(1)))
      OR (NOT (fsm_output(2))) OR (fsm_output(0)) OR (fsm_output(6)));
  mux_4414_nl <= MUX_s_1_2_2(mux_4415_nl, nor_2429_nl, fsm_output(7));
  mux_4413_nl <= MUX_s_1_2_2(and_2897_nl, mux_4414_nl, fsm_output(4));
  or_4857_nl <= (fsm_output(3)) OR (fsm_output(0)) OR (NOT (fsm_output(6)));
  mux_4419_nl <= MUX_s_1_2_2(or_4857_nl, or_tmp_4090, fsm_output(4));
  nor_2430_nl <= NOT((fsm_output(2)) OR (fsm_output(7)) OR (NOT (fsm_output(5)))
      OR mux_4419_nl);
  nand_574_nl <= NOT((fsm_output(3)) AND (fsm_output(0)) AND (fsm_output(6)));
  mux_4422_nl <= MUX_s_1_2_2(nand_574_nl, or_tmp_4090, fsm_output(4));
  nand_575_nl <= NOT((fsm_output(4)) AND (fsm_output(3)) AND (NOT (fsm_output(0)))
      AND (fsm_output(6)));
  mux_4421_nl <= MUX_s_1_2_2(mux_4422_nl, nand_575_nl, fsm_output(5));
  or_4858_nl <= (NOT (fsm_output(4))) OR (fsm_output(3)) OR (NOT (fsm_output(0)))
      OR (fsm_output(6));
  or_4859_nl <= (fsm_output(4)) OR (NOT (fsm_output(3))) OR (NOT (fsm_output(0)))
      OR (fsm_output(6));
  mux_4423_nl <= MUX_s_1_2_2(or_4858_nl, or_4859_nl, fsm_output(5));
  mux_4420_nl <= MUX_s_1_2_2(mux_4421_nl, mux_4423_nl, fsm_output(7));
  and_2898_nl <= (fsm_output(2)) AND (NOT mux_4420_nl);
  mux_4418_nl <= MUX_s_1_2_2(nor_2430_nl, and_2898_nl, fsm_output(1));
  or_4860_nl <= (NOT (fsm_output(5))) OR (fsm_output(6)) OR (fsm_output(3)) OR (NOT
      (fsm_output(0))) OR (fsm_output(7));
  or_4861_nl <= (fsm_output(5)) OR (NOT (fsm_output(6))) OR (fsm_output(3)) OR (NOT
      (fsm_output(0))) OR (fsm_output(7));
  mux_4425_nl <= MUX_s_1_2_2(or_4860_nl, or_4861_nl, fsm_output(4));
  nor_2431_nl <= NOT((fsm_output(1)) OR mux_4425_nl);
  nor_2432_nl <= NOT((NOT (fsm_output(5))) OR (fsm_output(6)) OR (NOT((fsm_output(3))
      AND (fsm_output(0)) AND (fsm_output(7)))));
  nor_2433_nl <= NOT((fsm_output(6)) OR (fsm_output(3)) OR (NOT((fsm_output(0)) AND
      (fsm_output(7)))));
  nor_2434_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(3))) OR (fsm_output(0))
      OR (fsm_output(7)));
  mux_4428_nl <= MUX_s_1_2_2(nor_2433_nl, nor_2434_nl, fsm_output(5));
  mux_4427_nl <= MUX_s_1_2_2(nor_2432_nl, mux_4428_nl, fsm_output(4));
  nor_2435_nl <= NOT((NOT (fsm_output(4))) OR (NOT (fsm_output(5))) OR (fsm_output(6))
      OR (fsm_output(3)) OR (NOT (fsm_output(0))) OR (fsm_output(7)));
  mux_4426_nl <= MUX_s_1_2_2(mux_4427_nl, nor_2435_nl, fsm_output(1));
  mux_4424_nl <= MUX_s_1_2_2(nor_2431_nl, mux_4426_nl, fsm_output(2));
  mult_3_res_mux1h_2_nl <= MUX1HOT_v_32_3_2(mult_16_z_slc_mult_z_mul_cmp_z_31_0_itm,
      modulo_add_base_1_sva, mult_17_z_slc_mult_z_mul_cmp_z_31_0_itm, STD_LOGIC_VECTOR'(
      mux_4413_nl & mux_4418_nl & mux_4424_nl));
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_res_mux1h_2_nl & '1')
      + UNSIGNED((NOT (mult_z_mul_cmp_z(31 DOWNTO 0))) & '1'), 33));
  and_2918_nl <= (fsm_output(4)) AND (NOT (fsm_output(2))) AND (fsm_output(1)) AND
      (NOT (fsm_output(0))) AND (NOT (fsm_output(6))) AND (fsm_output(7)) AND and_dcpl_103;
  modulo_add_3_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT modulo_add_base_3_sva_mx0w4),
      (NOT modulo_add_base_sva_mx0w7), (NOT modulo_add_base_20_sva_mx0w33), STD_LOGIC_VECTOR'(
      (NOT (fsm_output(1))) & (fsm_output(0)) & and_2918_nl));
  acc_15_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_3_mux1h_3_nl
      & '1'), 33), 34), 34));
  and_2925_nl <= (NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR (NOT
      (fsm_output(0))))) AND and_dcpl_1222 AND (NOT (fsm_output(5))) AND (NOT (fsm_output(3)));
  modulo_add_2_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT modulo_add_base_2_sva_mx0w5),
      (NOT modulo_add_base_12_sva_mx0w24), (NOT modulo_add_base_16_sva_mx0w29), STD_LOGIC_VECTOR'(
      (fsm_output(5)) & and_2925_nl & (fsm_output(3))));
  acc_17_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_2_mux1h_3_nl
      & '1'), 33), 34), 34));
  and_2929_nl <= (NOT (fsm_output(4))) AND (NOT (fsm_output(2))) AND and_dcpl_1241
      AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("00")) AND and_dcpl_103;
  and_2930_nl <= and_dcpl_1246 AND and_dcpl_1241 AND (fsm_output(6)) AND (NOT (fsm_output(7)))
      AND (NOT (fsm_output(5))) AND (NOT (fsm_output(3)));
  and_2931_nl <= and_dcpl_1596 AND and_dcpl_1222 AND (NOT (fsm_output(5))) AND (fsm_output(3));
  and_2932_nl <= and_dcpl_1596 AND and_dcpl_1222 AND and_dcpl_103;
  modulo_add_1_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_1_sva_mx0w6),
      (NOT modulo_add_base_10_sva_mx0w15), (NOT modulo_add_base_18_sva_mx0w27), (NOT
      modulo_add_base_22_sva_mx0w31), STD_LOGIC_VECTOR'( and_2929_nl & and_2930_nl
      & and_2931_nl & and_2932_nl));
  acc_19_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_1_mux1h_3_nl
      & '1'), 33), 34), 34));
  modulo_add_7_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT modulo_add_base_7_sva_mx0w9),
      (NOT modulo_add_base_15_sva_mx0w21), (NOT modulo_add_base_23_sva_mx0w30), STD_LOGIC_VECTOR'(
      and_2913_cse & (fsm_output(6)) & (fsm_output(7))));
  acc_20_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_7_mux1h_3_nl
      & '1'), 33), 34), 34));
  and_2934_nl <= and_dcpl_1246 AND (fsm_output(1)) AND (NOT (fsm_output(0))) AND
      (NOT (fsm_output(6))) AND (NOT (fsm_output(7))) AND and_2881_cse;
  and_2935_nl <= and_dcpl_1246 AND and_1317_cse AND and_dcpl_1210 AND nor_1711_cse;
  and_2936_nl <= and_dcpl_1633 AND and_dcpl_1210 AND and_2881_cse;
  and_2937_nl <= and_dcpl_1633 AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("10"))
      AND nor_1711_cse;
  modulo_add_6_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_6_sva_mx0w10),
      (NOT modulo_add_base_9_sva_mx0w16), (NOT modulo_add_base_14_sva_mx0w22), (NOT
      modulo_add_base_19_sva_mx0w26), STD_LOGIC_VECTOR'( and_2934_nl & and_2935_nl
      & and_2936_nl & and_2937_nl));
  acc_21_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_6_mux1h_3_nl
      & '1'), 33), 34), 34));
  and_2926_nl <= (fsm_output(1)) AND (NOT (fsm_output(2))) AND (fsm_output(4)) AND
      (fsm_output(0)) AND and_dcpl_1566;
  and_2927_nl <= and_dcpl_1573 AND and_dcpl_1566;
  and_2928_nl <= and_dcpl_1573 AND CONV_SL_1_1(fsm_output(7 DOWNTO 6)=STD_LOGIC_VECTOR'("01"))
      AND nor_1711_cse;
  modulo_add_5_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT modulo_add_base_5_sva_mx0w11),
      (NOT modulo_add_base_4_sva_mx0w12), (NOT modulo_add_base_8_sva_mx0w17), STD_LOGIC_VECTOR'(
      and_2926_nl & and_2927_nl & and_2928_nl));
  acc_18_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_5_mux1h_3_nl
      & '1'), 33), 34), 34));
  and_2938_nl <= nor_2178_cse_1 AND (fsm_output(4)) AND (fsm_output(0)) AND (fsm_output(6))
      AND (NOT (fsm_output(7))) AND (NOT (fsm_output(5))) AND (NOT (fsm_output(3)));
  modulo_add_11_mux1h_3_nl <= MUX1HOT_v_32_3_2((NOT modulo_add_base_11_sva_mx0w14),
      (NOT modulo_add_base_17_sva_mx0w28), (NOT modulo_add_base_21_sva_mx0w32), STD_LOGIC_VECTOR'(
      and_2938_nl & (fsm_output(3)) & (fsm_output(5))));
  acc_22_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_11_mux1h_3_nl
      & '1'), 33), 34), 34));
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(0))
      AND S1_OUTER_LOOP_for_nor_39_itm;
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_1_nl <= (S1_OUTER_LOOP_for_acc_svs_3_0(1))
      AND S1_OUTER_LOOP_for_nor_25_itm;
  S34_OUTER_LOOP_for_a_S34_OUTER_LOOP_for_a_and_15_nl <= S1_OUTER_LOOP_for_acc_svs_4
      AND S1_OUTER_LOOP_for_nor_26_itm;
  modulo_add_13_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & m_sva)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT modulo_add_base_13_sva_mx0w23),
      32), 33) + UNSIGNED'( "000000000000000000000000000000001"), 33));
  modulo_sub_18_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (z_out_12(30
      DOWNTO 0))) + UNSIGNED(m_sva), 32));
  and_1112_nl <= and_dcpl_447 AND and_dcpl_108;
  mux_4274_nl <= MUX_s_1_2_2(nor_tmp_35, mux_tmp_4268, or_2194_cse);
  mux_4273_nl <= MUX_s_1_2_2(mux_tmp_4268, nor_tmp_35, and_2893_cse);
  mux_4275_nl <= MUX_s_1_2_2(mux_4274_nl, mux_4273_nl, fsm_output(3));
  mux_4276_nl <= MUX_s_1_2_2(mux_4275_nl, mux_tmp_4267, fsm_output(4));
  mux_4271_nl <= MUX_s_1_2_2(mux_tmp_4268, nor_tmp_35, fsm_output(2));
  mux_4272_nl <= MUX_s_1_2_2(mux_4271_nl, mux_tmp_4267, fsm_output(4));
  mux_4277_nl <= MUX_s_1_2_2(mux_4276_nl, mux_4272_nl, fsm_output(1));
  mux_4266_nl <= MUX_s_1_2_2((fsm_output(6)), nor_tmp_35, fsm_output(2));
  and_2894_nl <= or_4854_cse AND (fsm_output(7));
  mux_4267_nl <= MUX_s_1_2_2(mux_4266_nl, and_2894_nl, fsm_output(4));
  mux_nl <= MUX_s_1_2_2((fsm_output(6)), nor_tmp_35, or_2194_cse);
  mux_4264_nl <= MUX_s_1_2_2((fsm_output(6)), mux_nl, fsm_output(3));
  and_2895_nl <= ((NOT((NOT (fsm_output(3))) OR (fsm_output(0)))) OR (fsm_output(2))
      OR (fsm_output(6))) AND (fsm_output(7));
  mux_4265_nl <= MUX_s_1_2_2(mux_4264_nl, and_2895_nl, fsm_output(4));
  mux_4268_nl <= MUX_s_1_2_2(mux_4267_nl, mux_4265_nl, fsm_output(1));
  mux_4278_nl <= MUX_s_1_2_2(mux_4277_nl, mux_4268_nl, fsm_output(5));
  mux_4290_nl <= MUX_s_1_2_2(or_tmp_4112, or_338_cse, fsm_output(2));
  or_4766_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00")) OR mux_4290_nl;
  or_4764_nl <= (fsm_output(4)) OR (NOT (fsm_output(2))) OR (fsm_output(6)) OR (NOT
      (fsm_output(7)));
  mux_4288_nl <= MUX_s_1_2_2(or_tmp_4118, or_tmp_4121, fsm_output(4));
  mux_4289_nl <= MUX_s_1_2_2(or_4764_nl, mux_4288_nl, fsm_output(3));
  mux_4291_nl <= MUX_s_1_2_2(or_4766_nl, mux_4289_nl, fsm_output(0));
  or_4762_nl <= (fsm_output(4)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(6)))
      OR (fsm_output(7));
  mux_4286_nl <= MUX_s_1_2_2(or_tmp_4117, or_tmp_4121, fsm_output(4));
  or_4761_nl <= (fsm_output(3)) OR mux_4286_nl;
  mux_4287_nl <= MUX_s_1_2_2(or_4762_nl, or_4761_nl, fsm_output(0));
  mux_4292_nl <= MUX_s_1_2_2(mux_4291_nl, mux_4287_nl, fsm_output(5));
  mux_4283_nl <= MUX_s_1_2_2(or_tmp_4118, or_tmp_4117, fsm_output(4));
  or_4758_nl <= (fsm_output(3)) OR mux_4283_nl;
  mux_4284_nl <= MUX_s_1_2_2(or_tmp_4115, or_4758_nl, fsm_output(0));
  or_4755_nl <= (fsm_output(3)) OR (fsm_output(4)) OR (NOT (fsm_output(2))) OR (fsm_output(6))
      OR (fsm_output(7));
  or_4753_nl <= (fsm_output(2)) OR (NOT (fsm_output(6))) OR (fsm_output(7));
  mux_4279_nl <= MUX_s_1_2_2(or_338_cse, or_tmp_4112, fsm_output(2));
  mux_4280_nl <= MUX_s_1_2_2(or_4753_nl, mux_4279_nl, fsm_output(4));
  mux_4281_nl <= MUX_s_1_2_2(or_tmp_4115, mux_4280_nl, fsm_output(3));
  mux_4282_nl <= MUX_s_1_2_2(or_4755_nl, mux_4281_nl, fsm_output(0));
  mux_4285_nl <= MUX_s_1_2_2(mux_4284_nl, mux_4282_nl, fsm_output(5));
  mux_4293_nl <= MUX_s_1_2_2(mux_4292_nl, mux_4285_nl, fsm_output(1));
  mux_4299_nl <= MUX_s_1_2_2((NOT or_4342_cse), or_4342_cse, fsm_output(5));
  mux_4300_nl <= MUX_s_1_2_2(nand_569_cse, mux_4299_nl, fsm_output(3));
  mux_4301_nl <= MUX_s_1_2_2(mux_4300_nl, nand_570_cse, fsm_output(4));
  mux_4297_nl <= MUX_s_1_2_2(or_4342_cse, nand_531_cse, fsm_output(5));
  nand_562_nl <= NOT((fsm_output(5)) AND nand_536_cse);
  mux_4298_nl <= MUX_s_1_2_2(mux_4297_nl, nand_562_nl, fsm_output(3));
  or_4853_nl <= (fsm_output(4)) OR mux_4298_nl;
  mux_4302_nl <= MUX_s_1_2_2(mux_4301_nl, or_4853_nl, fsm_output(6));
  nor_2423_nl <= NOT((fsm_output(3)) OR (fsm_output(5)) OR and_1317_cse OR (NOT (fsm_output(2))));
  mux_4294_nl <= MUX_s_1_2_2(nand_536_cse, or_4769_cse, fsm_output(0));
  or_4768_nl <= nor_2186_cse OR (fsm_output(2));
  mux_4295_nl <= MUX_s_1_2_2((NOT mux_4294_nl), or_4768_nl, fsm_output(5));
  and_2866_nl <= (fsm_output(3)) AND mux_4295_nl;
  mux_4296_nl <= MUX_s_1_2_2(nor_2423_nl, and_2866_nl, fsm_output(4));
  nor_2422_nl <= NOT((fsm_output(6)) OR mux_4296_nl);
  mux_4303_nl <= MUX_s_1_2_2(mux_4302_nl, nor_2422_nl, fsm_output(7));
  mux_4313_nl <= MUX_s_1_2_2(nor_2178_cse_1, and_2141_cse, fsm_output(0));
  mux_4314_nl <= MUX_s_1_2_2(mux_4313_nl, (NOT or_4342_cse), fsm_output(3));
  mux_4312_nl <= MUX_s_1_2_2((NOT and_2141_cse), or_4342_cse, fsm_output(3));
  mux_4315_nl <= MUX_s_1_2_2(mux_4314_nl, mux_4312_nl, fsm_output(5));
  mux_4316_nl <= MUX_s_1_2_2(mux_4315_nl, nand_570_cse, fsm_output(4));
  or_4782_nl <= CONV_SL_1_1(fsm_output(3 DOWNTO 0)/=STD_LOGIC_VECTOR'("0000"));
  mux_4411_nl <= MUX_s_1_2_2(and_2141_cse, (NOT or_4769_cse), fsm_output(0));
  mux_4309_nl <= MUX_s_1_2_2(mux_4411_nl, and_2141_cse, fsm_output(3));
  mux_4310_nl <= MUX_s_1_2_2(or_4782_nl, mux_4309_nl, fsm_output(5));
  mux_4311_nl <= MUX_s_1_2_2(mux_4310_nl, or_4781_cse, fsm_output(4));
  mux_4317_nl <= MUX_s_1_2_2(mux_4316_nl, mux_4311_nl, fsm_output(6));
  mux_4307_nl <= MUX_s_1_2_2((NOT (fsm_output(2))), or_4769_cse, fsm_output(0));
  nor_2421_nl <= NOT((fsm_output(5)) OR (fsm_output(3)) OR mux_4307_nl);
  mux_4305_nl <= MUX_s_1_2_2(and_2141_cse, (NOT or_4769_cse), fsm_output(0));
  and_2889_nl <= (fsm_output(3)) AND mux_4305_nl;
  or_4776_nl <= CONV_SL_1_1(fsm_output(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("01"));
  mux_4304_nl <= MUX_s_1_2_2(and_2141_cse, or_4776_nl, fsm_output(3));
  mux_4306_nl <= MUX_s_1_2_2(and_2889_nl, mux_4304_nl, fsm_output(5));
  mux_4308_nl <= MUX_s_1_2_2(nor_2421_nl, mux_4306_nl, fsm_output(4));
  nor_2420_nl <= NOT((fsm_output(6)) OR mux_4308_nl);
  mux_4318_nl <= MUX_s_1_2_2(mux_4317_nl, nor_2420_nl, fsm_output(7));
  or_4796_nl <= (fsm_output(2)) OR (fsm_output(5)) OR (fsm_output(1));
  or_4795_nl <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR (NOT (fsm_output(3)));
  or_4793_nl <= (NOT (fsm_output(1))) OR (fsm_output(3));
  mux_4329_nl <= MUX_s_1_2_2(or_4793_nl, or_4797_cse, fsm_output(5));
  mux_4330_nl <= MUX_s_1_2_2(or_4795_nl, mux_4329_nl, fsm_output(2));
  mux_4331_nl <= MUX_s_1_2_2(or_4796_nl, mux_4330_nl, fsm_output(0));
  mux_4328_nl <= MUX_s_1_2_2(or_tmp_4152, (NOT nor_tmp_31), fsm_output(2));
  or_4792_nl <= (fsm_output(0)) OR mux_4328_nl;
  mux_4332_nl <= MUX_s_1_2_2(mux_4331_nl, or_4792_nl, fsm_output(4));
  or_4790_nl <= (NOT (fsm_output(5))) OR (fsm_output(1)) OR (fsm_output(3));
  mux_4325_nl <= MUX_s_1_2_2(or_tmp_4152, or_4790_nl, fsm_output(2));
  mux_4326_nl <= MUX_s_1_2_2(nand_569_cse, mux_4325_nl, fsm_output(0));
  or_4789_nl <= (NOT (fsm_output(2))) OR (fsm_output(5)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3));
  mux_4327_nl <= MUX_s_1_2_2(mux_4326_nl, or_4789_nl, fsm_output(4));
  mux_4333_nl <= MUX_s_1_2_2(mux_4332_nl, mux_4327_nl, fsm_output(6));
  or_4787_nl <= (NOT (fsm_output(0))) OR (fsm_output(5)) OR (NOT (fsm_output(1)))
      OR (fsm_output(3));
  or_4786_nl <= (fsm_output(1)) OR (NOT (fsm_output(3)));
  mux_4321_nl <= MUX_s_1_2_2(or_4786_nl, or_4797_cse, fsm_output(5));
  mux_4322_nl <= MUX_s_1_2_2((NOT nor_tmp_31), mux_4321_nl, fsm_output(2));
  mux_4319_nl <= MUX_s_1_2_2(nand_568_cse, or_4797_cse, fsm_output(5));
  mux_4320_nl <= MUX_s_1_2_2((NOT nor_tmp_31), mux_4319_nl, fsm_output(2));
  mux_4323_nl <= MUX_s_1_2_2(mux_4322_nl, mux_4320_nl, fsm_output(0));
  mux_4324_nl <= MUX_s_1_2_2(or_4787_nl, mux_4323_nl, fsm_output(4));
  or_4788_nl <= (fsm_output(6)) OR mux_4324_nl;
  mux_4334_nl <= MUX_s_1_2_2(mux_4333_nl, or_4788_nl, fsm_output(7));
  or_290_nl <= (fsm_output(6)) OR (NOT (fsm_output(2))) OR (NOT (fsm_output(1)))
      OR (fsm_output(4));
  or_289_nl <= (NOT (fsm_output(6))) OR (NOT (fsm_output(2))) OR (fsm_output(1))
      OR (fsm_output(4));
  mux_105_nl <= MUX_s_1_2_2(or_290_nl, or_289_nl, fsm_output(5));
  or_4683_nl <= (fsm_output(3)) OR mux_105_nl;
  or_4684_nl <= (NOT (fsm_output(3))) OR (NOT (fsm_output(5))) OR (fsm_output(6))
      OR (fsm_output(2)) OR (NOT nor_tmp_3);
  mux_106_nl <= MUX_s_1_2_2(or_4683_nl, or_4684_nl, fsm_output(7));
  nor_2209_nl <= NOT(mux_106_nl OR (fsm_output(0)));
  S2_INNER_LOOP1_S2_INNER_LOOP1_and_nl <= MUX_v_15_2_2(STD_LOGIC_VECTOR'("000000000000000"),
      (S1_OUTER_LOOP_for_p_sva_1(19 DOWNTO 5)), nor_2209_nl);
  mux_4357_nl <= MUX_s_1_2_2(or_tmp_48, or_4805_cse, fsm_output(0));
  mux_4355_nl <= MUX_s_1_2_2(or_4162_cse, or_tmp_48, fsm_output(1));
  mux_4356_nl <= MUX_s_1_2_2(mux_tmp_4334, mux_4355_nl, fsm_output(0));
  mux_4358_nl <= MUX_s_1_2_2(mux_4357_nl, mux_4356_nl, fsm_output(3));
  mux_4353_nl <= MUX_s_1_2_2(or_tmp_48, (fsm_output(7)), fsm_output(1));
  mux_4354_nl <= MUX_s_1_2_2(or_tmp_4164, mux_4353_nl, fsm_output(3));
  mux_4359_nl <= MUX_s_1_2_2((NOT mux_4358_nl), mux_4354_nl, fsm_output(6));
  and_2885_nl <= ((NOT (fsm_output(1))) OR (fsm_output(7))) AND (fsm_output(5));
  mux_4348_nl <= MUX_s_1_2_2((NOT (fsm_output(5))), (fsm_output(5)), fsm_output(7));
  mux_4349_nl <= MUX_s_1_2_2(and_2112_cse, mux_4348_nl, fsm_output(1));
  mux_4350_nl <= MUX_s_1_2_2(and_2885_nl, mux_4349_nl, fsm_output(0));
  mux_4351_nl <= MUX_s_1_2_2(mux_4350_nl, or_tmp_4164, fsm_output(3));
  mux_4346_nl <= MUX_s_1_2_2(or_tmp_48, (fsm_output(7)), fsm_output(0));
  mux_4345_nl <= MUX_s_1_2_2(or_tmp_48, (fsm_output(7)), and_1317_cse);
  mux_4347_nl <= MUX_s_1_2_2(mux_4346_nl, mux_4345_nl, fsm_output(3));
  mux_4352_nl <= MUX_s_1_2_2((NOT mux_4351_nl), mux_4347_nl, fsm_output(6));
  mux_4360_nl <= MUX_s_1_2_2(mux_4359_nl, mux_4352_nl, fsm_output(2));
  nor_2417_nl <= NOT((fsm_output(0)) OR (fsm_output(1)) OR (fsm_output(7)) OR (fsm_output(5)));
  mux_4342_nl <= MUX_s_1_2_2(nor_2417_nl, and_2112_cse, fsm_output(3));
  mux_4340_nl <= MUX_s_1_2_2((fsm_output(7)), or_4162_cse, or_3894_cse);
  mux_4341_nl <= MUX_s_1_2_2((fsm_output(7)), mux_4340_nl, fsm_output(3));
  mux_4343_nl <= MUX_s_1_2_2(mux_4342_nl, mux_4341_nl, fsm_output(6));
  nor_2418_nl <= NOT((fsm_output(1)) OR (NOT and_2112_cse));
  mux_4337_nl <= MUX_s_1_2_2(nor_2418_nl, and_2112_cse, fsm_output(0));
  mux_4338_nl <= MUX_s_1_2_2(mux_4337_nl, mux_tmp_4334, fsm_output(3));
  mux_4335_nl <= MUX_s_1_2_2((fsm_output(7)), or_4162_cse, or_4797_cse);
  mux_4339_nl <= MUX_s_1_2_2(mux_4338_nl, mux_4335_nl, fsm_output(6));
  mux_4344_nl <= MUX_s_1_2_2(mux_4343_nl, mux_4339_nl, fsm_output(2));
  mux_4361_nl <= MUX_s_1_2_2(mux_4360_nl, mux_4344_nl, fsm_output(4));
  nor_2410_nl <= NOT((fsm_output(2)) OR (NOT (fsm_output(6))) OR (NOT (fsm_output(1)))
      OR (fsm_output(5)));
  mux_4369_nl <= MUX_s_1_2_2(and_1274_cse, (NOT or_tmp_4177), fsm_output(2));
  mux_4370_nl <= MUX_s_1_2_2(nor_2410_nl, mux_4369_nl, fsm_output(3));
  mux_4366_nl <= MUX_s_1_2_2(nor_2411_cse, (fsm_output(5)), fsm_output(6));
  mux_4367_nl <= MUX_s_1_2_2((NOT or_tmp_4177), mux_4366_nl, fsm_output(2));
  mux_4365_nl <= MUX_s_1_2_2(nor_2412_cse, and_1274_cse, fsm_output(6));
  mux_4368_nl <= MUX_s_1_2_2(mux_4367_nl, mux_4365_nl, fsm_output(3));
  mux_4371_nl <= MUX_s_1_2_2(mux_4370_nl, mux_4368_nl, fsm_output(0));
  nor_2413_nl <= NOT((NOT (fsm_output(3))) OR (fsm_output(2)) OR (NOT (fsm_output(6)))
      OR (fsm_output(1)) OR (fsm_output(5)));
  nor_2414_nl <= NOT((fsm_output(3)) OR (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(1))
      OR (fsm_output(5)));
  mux_4364_nl <= MUX_s_1_2_2(nor_2413_nl, nor_2414_nl, fsm_output(0));
  mux_4372_nl <= MUX_s_1_2_2(mux_4371_nl, mux_4364_nl, fsm_output(4));
  or_4810_nl <= (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(1)) OR (NOT (fsm_output(5)));
  or_4808_nl <= (fsm_output(2)) OR (fsm_output(6)) OR (fsm_output(1)) OR (fsm_output(5));
  mux_4362_nl <= MUX_s_1_2_2(or_4810_nl, or_4808_nl, fsm_output(3));
  nor_2415_nl <= NOT((fsm_output(0)) OR mux_4362_nl);
  nor_2416_nl <= NOT((fsm_output(0)) OR (fsm_output(3)) OR (NOT (fsm_output(2)))
      OR (fsm_output(6)) OR (NOT and_1274_cse));
  mux_4363_nl <= MUX_s_1_2_2(nor_2415_nl, nor_2416_nl, fsm_output(4));
  mux_4373_nl <= MUX_s_1_2_2(mux_4372_nl, mux_4363_nl, fsm_output(7));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_60_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11110"));
  S6_OUTER_LOOP_for_nor_25_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(4 DOWNTO
      1)/=STD_LOGIC_VECTOR'("0000")));
  S6_OUTER_LOOP_for_nor_26_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(4)) OR (S6_OUTER_LOOP_for_acc_tmp(3))
      OR (S6_OUTER_LOOP_for_acc_tmp(2)) OR (S6_OUTER_LOOP_for_acc_tmp(0)));
  S6_OUTER_LOOP_for_nor_39_nl <= NOT(CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp(3 DOWNTO
      0)/=STD_LOGIC_VECTOR'("0000")));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_6_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("111"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("00"));
  S34_OUTER_LOOP_for_a_nor_3_nl <= NOT((S34_OUTER_LOOP_for_a_acc_2_tmp(4)) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(3))
      OR (S34_OUTER_LOOP_for_a_acc_2_tmp(1)) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(0)));
  S6_OUTER_LOOP_for_nor_28_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(4)) OR (S6_OUTER_LOOP_for_acc_tmp(3))
      OR (S6_OUTER_LOOP_for_acc_tmp(1)) OR (S6_OUTER_LOOP_for_acc_tmp(0)));
  S34_OUTER_LOOP_for_a_nor_7_nl <= NOT((S34_OUTER_LOOP_for_a_acc_2_tmp(4)) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(2))
      OR (S34_OUTER_LOOP_for_a_acc_2_tmp(1)) OR (S34_OUTER_LOOP_for_a_acc_2_tmp(0)));
  S6_OUTER_LOOP_for_nor_32_nl <= NOT((S6_OUTER_LOOP_for_acc_tmp(4)) OR (S6_OUTER_LOOP_for_acc_tmp(2))
      OR (S6_OUTER_LOOP_for_acc_tmp(1)) OR (S6_OUTER_LOOP_for_acc_tmp(0)));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_nor_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_45_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("01111"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_53_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("10111"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_57_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11011"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_59_nl <= CONV_SL_1_1(S6_OUTER_LOOP_for_acc_tmp=STD_LOGIC_VECTOR'("11101"));
  S2_COPY_LOOP_for_nor_nl <= NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3
      DOWNTO 1)/=STD_LOGIC_VECTOR'("000")));
  S6_OUTER_LOOP_for_nor_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  S2_COPY_LOOP_for_nor_1_nl <= NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)));
  S6_OUTER_LOOP_for_nor_1_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)));
  S2_COPY_LOOP_for_nor_3_nl <= NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(3))
      OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(1)) OR (reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(0)));
  S6_OUTER_LOOP_for_nor_3_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  S2_COPY_LOOP_for_nor_7_nl <= NOT(reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg OR CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg(2
      DOWNTO 0)/=STD_LOGIC_VECTOR'("000")));
  S6_OUTER_LOOP_for_nor_7_nl <= NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  S2_COPY_LOOP_for_nor_14_nl <= NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg/=STD_LOGIC_VECTOR'("0000")));
  S6_OUTER_LOOP_for_nor_14_nl <= NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg/=STD_LOGIC_VECTOR'("000")));
  butterFly_7_f1_butterFly_7_f1_nor_nl <= NOT(CONV_SL_1_1(operator_20_true_28_acc_tmp/=STD_LOGIC_VECTOR'("000")));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_10_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))));
  butterFly_7_f1_butterFly_7_f1_and_4_nl <= CONV_SL_1_1(operator_20_true_28_acc_tmp=STD_LOGIC_VECTOR'("101"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_12_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))
      AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1))));
  butterFly_7_f1_butterFly_7_f1_and_5_nl <= CONV_SL_1_1(operator_20_true_28_acc_tmp=STD_LOGIC_VECTOR'("110"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_13_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_18_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_20_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))
      AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_21_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)=STD_LOGIC_VECTOR'("11"))
      AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_24_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND S6_OUTER_LOOP_for_nor_22_cse;
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_27_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("100"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_25_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg=STD_LOGIC_VECTOR'("11"))
      AND CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("010"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_2_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_4_nl <= (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_5_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (NOT(CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_1_reg/=STD_LOGIC_VECTOR'("00"))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_8_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
  butterFly_7_f1_butterFly_7_f1_and_2_nl <= CONV_SL_1_1(operator_20_true_28_acc_tmp=STD_LOGIC_VECTOR'("011"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_11_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(1 DOWNTO 0)/=STD_LOGIC_VECTOR'("00"))));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_16_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0)) AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      OR CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg(2 DOWNTO 1)/=STD_LOGIC_VECTOR'("00"))));
  butterFly_4_f1_butterFly_4_f1_and_2_nl <= CONV_SL_1_1(reg_S2_COPY_LOOP_for_i_5_0_2_reg=STD_LOGIC_VECTOR'("011"));
  S6_OUTER_LOOP_for_S6_OUTER_LOOP_for_and_17_nl <= (reg_S2_COPY_LOOP_for_i_5_0_1_reg(1))
      AND (reg_S2_COPY_LOOP_for_i_5_0_2_reg(1)) AND (NOT((reg_S2_COPY_LOOP_for_i_5_0_1_reg(0))
      OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(2)) OR (reg_S2_COPY_LOOP_for_i_5_0_2_reg(0))));
  or_4824_nl <= (fsm_output(5)) OR and_2083_cse;
  mux_4387_nl <= MUX_s_1_2_2(or_4824_nl, (fsm_output(4)), fsm_output(1));
  nor_2402_nl <= NOT(nor_1308_cse OR (fsm_output(4)));
  mux_4386_nl <= MUX_s_1_2_2(nor_2402_nl, mux_tmp_4374, fsm_output(1));
  mux_4388_nl <= MUX_s_1_2_2((NOT mux_4387_nl), mux_4386_nl, fsm_output(3));
  mux_4385_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), and_2881_cse);
  mux_4389_nl <= MUX_s_1_2_2(mux_4388_nl, mux_4385_nl, fsm_output(2));
  mux_4382_nl <= MUX_s_1_2_2((NOT and_2083_cse), (fsm_output(4)), or_4805_cse);
  mux_4383_nl <= MUX_s_1_2_2(mux_4382_nl, mux_tmp_4373, fsm_output(3));
  or_4821_nl <= (fsm_output(0)) OR (fsm_output(4));
  mux_4380_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), or_4821_nl, fsm_output(5));
  mux_4381_nl <= MUX_s_1_2_2(mux_tmp_4373, mux_4380_nl, fsm_output(1));
  mux_4384_nl <= MUX_s_1_2_2(mux_4383_nl, mux_4381_nl, fsm_output(2));
  mux_4390_nl <= MUX_s_1_2_2((NOT mux_4389_nl), mux_4384_nl, fsm_output(6));
  mux_4377_nl <= MUX_s_1_2_2(mux_tmp_4374, mux_tmp_4373, fsm_output(1));
  and_2882_nl <= ((fsm_output(1)) OR (fsm_output(5)) OR (fsm_output(0))) AND (fsm_output(4));
  mux_4378_nl <= MUX_s_1_2_2(mux_4377_nl, and_2882_nl, fsm_output(3));
  mux_4374_nl <= MUX_s_1_2_2((NOT (fsm_output(4))), (fsm_output(4)), or_4818_cse);
  mux_4379_nl <= MUX_s_1_2_2(mux_4378_nl, mux_4374_nl, fsm_output(2));
  nor_2403_nl <= NOT((fsm_output(6)) OR mux_4379_nl);
  mux_4391_nl <= MUX_s_1_2_2(mux_4390_nl, nor_2403_nl, fsm_output(7));
  nor_2404_nl <= NOT((NOT (fsm_output(3))) OR (NOT (fsm_output(7))) OR (fsm_output(4))
      OR (fsm_output(1)));
  nor_2405_nl <= NOT((fsm_output(7)) OR (NOT (fsm_output(4))) OR (fsm_output(1)));
  nor_2406_nl <= NOT((fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(1)));
  mux_4393_nl <= MUX_s_1_2_2(nor_2405_nl, nor_2406_nl, fsm_output(3));
  mux_4394_nl <= MUX_s_1_2_2(nor_2404_nl, mux_4393_nl, fsm_output(0));
  or_4831_nl <= (NOT (fsm_output(7))) OR (fsm_output(4)) OR (fsm_output(1));
  or_4830_nl <= (fsm_output(7)) OR (fsm_output(4)) OR (NOT (fsm_output(1)));
  mux_4392_nl <= MUX_s_1_2_2(or_4831_nl, or_4830_nl, fsm_output(3));
  nor_2407_nl <= NOT((fsm_output(0)) OR mux_4392_nl);
  mux_4395_nl <= MUX_s_1_2_2(mux_4394_nl, nor_2407_nl, fsm_output(5));
  nor_2408_nl <= NOT((fsm_output(5)) OR (fsm_output(0)) OR (fsm_output(3)) OR (fsm_output(7))
      OR (fsm_output(4)) OR (NOT (fsm_output(1))));
  mux_4396_nl <= MUX_s_1_2_2(mux_4395_nl, nor_2408_nl, fsm_output(6));
  nor_2409_nl <= NOT((NOT (fsm_output(6))) OR (NOT (fsm_output(5))) OR (NOT (fsm_output(0)))
      OR (fsm_output(7)) OR (fsm_output(4)) OR (NOT (fsm_output(1))));
  mux_4397_nl <= MUX_s_1_2_2(mux_4396_nl, nor_2409_nl, fsm_output(2));
  and_2879_nl <= (fsm_output(3)) AND (fsm_output(0));
  mux_4401_nl <= MUX_s_1_2_2((fsm_output(4)), or_tmp_4199, and_2879_nl);
  or_4842_nl <= (fsm_output(3)) OR mux_tmp_4396;
  mux_4402_nl <= MUX_s_1_2_2((NOT mux_4401_nl), or_4842_nl, fsm_output(7));
  mux_4400_nl <= MUX_s_1_2_2((fsm_output(4)), or_tmp_4199, fsm_output(0));
  or_4841_nl <= (fsm_output(7)) OR (fsm_output(3)) OR mux_4400_nl;
  mux_4403_nl <= MUX_s_1_2_2(mux_4402_nl, or_4841_nl, fsm_output(5));
  mux_4399_nl <= MUX_s_1_2_2((fsm_output(4)), mux_tmp_4396, fsm_output(3));
  or_4839_nl <= (NOT (fsm_output(5))) OR (fsm_output(7)) OR (NOT mux_4399_nl);
  mux_4404_nl <= MUX_s_1_2_2(mux_4403_nl, or_4839_nl, fsm_output(6));
  and_2875_nl <= (fsm_output(7)) AND (CONV_SL_1_1(fsm_output(2 DOWNTO 0)/=STD_LOGIC_VECTOR'("101")));
  mux_4408_nl <= MUX_s_1_2_2(and_2875_nl, or_tmp_4208, fsm_output(3));
  and_2877_nl <= (fsm_output(3)) AND (fsm_output(7)) AND (fsm_output(1)) AND (fsm_output(2));
  mux_4409_nl <= MUX_s_1_2_2((NOT mux_4408_nl), and_2877_nl, fsm_output(4));
  or_4849_nl <= (fsm_output(6)) OR mux_4409_nl;
  or_4846_nl <= CONV_SL_1_1(fsm_output(4 DOWNTO 3)/=STD_LOGIC_VECTOR'("00"));
  mux_4406_nl <= MUX_s_1_2_2(or_tmp_4208, (fsm_output(7)), or_4846_nl);
  or_4845_nl <= (NOT (fsm_output(3))) OR (fsm_output(7)) OR (NOT(or_3894_cse AND
      (fsm_output(2))));
  mux_4405_nl <= MUX_s_1_2_2(or_4845_nl, (fsm_output(7)), fsm_output(4));
  mux_4407_nl <= MUX_s_1_2_2(mux_4406_nl, mux_4405_nl, fsm_output(6));
  mux_4410_nl <= MUX_s_1_2_2(or_4849_nl, mux_4407_nl, fsm_output(5));
  S5_COPY_LOOP_for_mux_3_nl <= MUX_s_1_2_2(S1_OUTER_LOOP_for_acc_svs_4, reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg,
      and_2348_ssc);
  S5_COPY_LOOP_for_mux_4_nl <= MUX_v_4_2_2(S1_OUTER_LOOP_for_acc_svs_3_0, reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg,
      and_2348_ssc);
  z_out <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(S5_COPY_LOOP_for_mux_3_nl
      & S5_COPY_LOOP_for_mux_4_nl), 5), 6) + UNSIGNED'( "000001"), 6));
  mult_3_if_or_4_nl <= (nor_2178_cse_1 AND and_dcpl_1085 AND nor_1346_cse AND and_dcpl_103)
      OR (and_dcpl_1206 AND and_2083_cse AND nor_1346_cse AND and_2881_cse) OR (and_2399_cse
      AND and_dcpl_1210 AND nor_1711_cse) OR (and_dcpl_1206 AND and_dcpl_82 AND and_dcpl_1210
      AND and_dcpl_103) OR (nor_2178_cse_1 AND and_dcpl_82 AND and_dcpl_1222 AND
      nor_1711_cse) OR (and_2399_cse AND and_dcpl_1222 AND and_dcpl_460) OR (and_2399_cse
      AND and_dcpl_1222 AND and_dcpl_103);
  mult_3_if_mux_1_nl <= MUX_v_32_2_2(mult_3_res_sva, mult_1_res_sva, mult_3_if_or_4_nl);
  acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_if_mux_1_nl & '1') +
      UNSIGNED((NOT m_sva) & '1'), 33));
  z_out_5 <= acc_2_nl(32 DOWNTO 1);
  acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_res_sva & '1') + UNSIGNED((NOT
      m_sva) & '1'), 33));
  z_out_6 <= acc_3_nl(32 DOWNTO 1);
  and_2906_nl <= (fsm_output(1)) AND (NOT (fsm_output(2))) AND (fsm_output(4)) AND
      (NOT (fsm_output(0))) AND nor_1346_cse AND and_2881_cse;
  and_2907_nl <= (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(4)) AND (fsm_output(0))
      AND (fsm_output(6)) AND (NOT (fsm_output(7))) AND and_2881_cse;
  modulo_sub_3_qif_mux1h_2_nl <= MUX1HOT_v_31_3_2((modulo_sub_base_3_sva_1(30 DOWNTO
      0)), (modulo_sub_base_6_sva_1(30 DOWNTO 0)), (modulo_sub_base_14_sva_1(30 DOWNTO
      0)), STD_LOGIC_VECTOR'( (NOT (fsm_output(4))) & and_2906_nl & and_2907_nl));
  z_out_7 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_3_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  nor_2436_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (NOT and_dcpl_1257) OR
      (fsm_output(6)) OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  and_2908_nl <= (fsm_output(4)) AND (NOT (fsm_output(2))) AND and_dcpl_1257 AND
      (fsm_output(6)) AND (NOT (fsm_output(7))) AND (NOT (fsm_output(5))) AND (NOT
      (fsm_output(3)));
  modulo_sub_2_qif_mux1h_2_nl <= MUX1HOT_v_31_3_2((modulo_sub_base_2_sva_1(30 DOWNTO
      0)), (modulo_sub_base_11_sva_1(30 DOWNTO 0)), (modulo_sub_base_21_sva_1(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( nor_2436_nl & and_2908_nl & (fsm_output(7))));
  z_out_8 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_2_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  nor_2437_nl <= NOT((NOT and_dcpl_1206) OR (fsm_output(4)) OR (fsm_output(0)) OR
      (fsm_output(6)) OR (fsm_output(7)) OR (NOT (fsm_output(5))) OR (fsm_output(3)));
  and_2909_nl <= and_dcpl_1206 AND (fsm_output(4)) AND (NOT (fsm_output(0))) AND
      and_dcpl_1324;
  and_2910_nl <= and_dcpl_1206 AND (fsm_output(4)) AND (fsm_output(0)) AND and_dcpl_1324;
  and_2911_nl <= CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("10101111"));
  modulo_sub_1_qif_mux1h_2_nl <= MUX1HOT_v_31_4_2((modulo_sub_base_1_sva_1(30 DOWNTO
      0)), (modulo_sub_base_10_sva_1(30 DOWNTO 0)), (modulo_sub_base_9_sva_1(30 DOWNTO
      0)), (modulo_sub_base_23_sva_1(30 DOWNTO 0)), STD_LOGIC_VECTOR'( nor_2437_nl
      & and_2909_nl & and_2910_nl & and_2911_nl));
  z_out_9 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_1_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  and_2912_nl <= and_dcpl_925 AND CONV_SL_1_1(fsm_output(1 DOWNTO 0)=STD_LOGIC_VECTOR'("11"))
      AND nor_1346_cse AND (fsm_output(5)) AND (NOT (fsm_output(3)));
  modulo_sub_qif_mux1h_2_nl <= MUX1HOT_v_31_3_2((modulo_sub_base_sva_1(30 DOWNTO
      0)), (modulo_sub_base_4_sva_1(30 DOWNTO 0)), (modulo_sub_base_8_sva_1(30 DOWNTO
      0)), STD_LOGIC_VECTOR'( and_2912_nl & (fsm_output(3)) & (NOT (fsm_output(5)))));
  z_out_10 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  and_2913_cse <= nor_2178_cse_1 AND (fsm_output(4)) AND (fsm_output(0)) AND (NOT
      (fsm_output(6))) AND (NOT (fsm_output(7))) AND and_2881_cse;
  and_2914_nl <= (fsm_output(1)) AND (fsm_output(2)) AND (fsm_output(4)) AND (NOT
      (fsm_output(0))) AND (fsm_output(6)) AND (NOT (fsm_output(7))) AND and_2881_cse;
  modulo_sub_7_qif_mux1h_2_nl <= MUX1HOT_v_31_3_2((modulo_sub_base_7_sva_1(30 DOWNTO
      0)), (modulo_sub_base_15_sva_1(30 DOWNTO 0)), (modulo_sub_base_19_sva_1(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( and_2913_cse & and_2914_nl & (fsm_output(7))));
  z_out_11 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_7_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  and_2915_nl <= (fsm_output(4)) AND (NOT (fsm_output(2))) AND nor_1375_cse AND (NOT
      (fsm_output(6))) AND (fsm_output(7)) AND (fsm_output(5)) AND (NOT (fsm_output(3)));
  butterFly_18_mux_2_nl <= MUX_v_32_2_2(tmp_21_lpi_4_dfm, tmp_50_lpi_3_dfm, and_2915_nl);
  acc_9_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(butterFly_18_mux_2_nl & '1')
      + UNSIGNED((NOT reg_mult_3_res_lpi_4_dfm_cse) & '1'), 33));
  z_out_12 <= acc_9_nl(32 DOWNTO 1);
  and_2916_nl <= nor_2178_cse_1 AND (fsm_output(4)) AND (fsm_output(0)) AND (NOT
      (fsm_output(6))) AND (fsm_output(7)) AND (NOT (fsm_output(5))) AND (fsm_output(3));
  modulo_sub_5_qif_mux1h_2_nl <= MUX1HOT_v_31_3_2((modulo_sub_base_5_sva_1(30 DOWNTO
      0)), (modulo_sub_base_13_sva_1(30 DOWNTO 0)), (modulo_sub_base_17_sva_1(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(5)) & (NOT (fsm_output(3))) & and_2916_nl));
  z_out_13 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_5_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  nor_2438_nl <= NOT((fsm_output(4)) OR (fsm_output(2)) OR (fsm_output(1)) OR (NOT
      (fsm_output(0))) OR (NOT and_dcpl_1222) OR (fsm_output(5)) OR (fsm_output(3)));
  and_2917_nl <= (fsm_output(4)) AND (NOT (fsm_output(2))) AND (fsm_output(1)) AND
      (NOT (fsm_output(0))) AND and_dcpl_1222 AND (fsm_output(5)) AND (NOT (fsm_output(3)));
  modulo_sub_12_qif_mux1h_2_nl <= MUX1HOT_v_31_3_2((modulo_sub_base_12_sva_1(30 DOWNTO
      0)), (modulo_sub_base_16_sva_1(30 DOWNTO 0)), (modulo_sub_base_20_sva_1(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( nor_2438_nl & (fsm_output(3)) & and_2917_nl));
  z_out_14 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_12_qif_mux1h_2_nl)
      + UNSIGNED(m_sva), 32));
  operator_20_true_15_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_26(19
      DOWNTO 5)) + UNSIGNED'( "111111111111111"), 15));
  z_out_16_14 <= operator_20_true_15_acc_nl(14);
  acc_14_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_3_res_sva & '1')
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT m_sva) & '1'), 33), 34), 34));
  z_out_17_32 <= acc_14_nl(33);
  mult_1_if_or_2_nl <= (and_dcpl_1206 AND and_dcpl_82 AND nor_1346_cse AND and_dcpl_103)
      OR (nor_2178_cse_1 AND and_dcpl_1455 AND nor_1346_cse AND and_2881_cse) OR
      (and_dcpl_1206 AND and_dcpl_1455 AND and_dcpl_1210 AND nor_1711_cse) OR (CONV_SL_1_1(fsm_output(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("10")) AND and_2083_cse AND and_dcpl_1210 AND and_2881_cse)
      OR (and_2141_cse AND and_dcpl_1455 AND and_dcpl_1222 AND nor_1711_cse) OR (and_2141_cse
      AND and_dcpl_82 AND and_dcpl_1222 AND and_2881_cse);
  mult_1_if_mult_1_if_mux_1_nl <= MUX_v_32_2_2(mult_1_res_sva, mult_3_res_sva, mult_1_if_or_2_nl);
  acc_16_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_1_if_mult_1_if_mux_1_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT m_sva) & '1'), 33), 34),
      34));
  z_out_19_32 <= acc_16_nl(33);
  and_2939_nl <= CONV_SL_1_1(fsm_output=STD_LOGIC_VECTOR'("10110110"));
  S34_OUTER_LOOP_for_mux_3_nl <= MUX_v_5_2_2((reg_S2_COPY_LOOP_p_5_0_sva_4_0_reg
      & reg_S2_COPY_LOOP_p_5_0_sva_4_0_1_reg), (reg_S2_COPY_LOOP_for_i_5_0_1_reg
      & reg_S2_COPY_LOOP_for_i_5_0_2_reg), and_2939_nl);
  z_out_26 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED((S1_OUTER_LOOP_for_p_sva_1(14
      DOWNTO 0)) & S34_OUTER_LOOP_for_mux_3_nl) + UNSIGNED'( "00000000000000000001"),
      20));
END v14;

-- ------------------------------------------------------------------
--  Design Unit:    hybrid
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_DPRAM_RBW_DUAL_pkg.ALL;


ENTITY hybrid IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    x_rsc_0_0_s_tdone : IN STD_LOGIC;
    x_rsc_0_0_tr_write_done : IN STD_LOGIC;
    x_rsc_0_0_RREADY : IN STD_LOGIC;
    x_rsc_0_0_RVALID : OUT STD_LOGIC;
    x_rsc_0_0_RUSER : OUT STD_LOGIC;
    x_rsc_0_0_RLAST : OUT STD_LOGIC;
    x_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_RID : OUT STD_LOGIC;
    x_rsc_0_0_ARREADY : OUT STD_LOGIC;
    x_rsc_0_0_ARVALID : IN STD_LOGIC;
    x_rsc_0_0_ARUSER : IN STD_LOGIC;
    x_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_ARLOCK : IN STD_LOGIC;
    x_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_0_0_ARID : IN STD_LOGIC;
    x_rsc_0_0_BREADY : IN STD_LOGIC;
    x_rsc_0_0_BVALID : OUT STD_LOGIC;
    x_rsc_0_0_BUSER : OUT STD_LOGIC;
    x_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_BID : OUT STD_LOGIC;
    x_rsc_0_0_WREADY : OUT STD_LOGIC;
    x_rsc_0_0_WVALID : IN STD_LOGIC;
    x_rsc_0_0_WUSER : IN STD_LOGIC;
    x_rsc_0_0_WLAST : IN STD_LOGIC;
    x_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_0_0_AWREADY : OUT STD_LOGIC;
    x_rsc_0_0_AWVALID : IN STD_LOGIC;
    x_rsc_0_0_AWUSER : IN STD_LOGIC;
    x_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_0_0_AWLOCK : IN STD_LOGIC;
    x_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_0_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    x_rsc_1_0_s_tdone : IN STD_LOGIC;
    x_rsc_1_0_tr_write_done : IN STD_LOGIC;
    x_rsc_1_0_RREADY : IN STD_LOGIC;
    x_rsc_1_0_RVALID : OUT STD_LOGIC;
    x_rsc_1_0_RUSER : OUT STD_LOGIC;
    x_rsc_1_0_RLAST : OUT STD_LOGIC;
    x_rsc_1_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_RID : OUT STD_LOGIC;
    x_rsc_1_0_ARREADY : OUT STD_LOGIC;
    x_rsc_1_0_ARVALID : IN STD_LOGIC;
    x_rsc_1_0_ARUSER : IN STD_LOGIC;
    x_rsc_1_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_ARLOCK : IN STD_LOGIC;
    x_rsc_1_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_1_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_1_0_ARID : IN STD_LOGIC;
    x_rsc_1_0_BREADY : IN STD_LOGIC;
    x_rsc_1_0_BVALID : OUT STD_LOGIC;
    x_rsc_1_0_BUSER : OUT STD_LOGIC;
    x_rsc_1_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_BID : OUT STD_LOGIC;
    x_rsc_1_0_WREADY : OUT STD_LOGIC;
    x_rsc_1_0_WVALID : IN STD_LOGIC;
    x_rsc_1_0_WUSER : IN STD_LOGIC;
    x_rsc_1_0_WLAST : IN STD_LOGIC;
    x_rsc_1_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_1_0_AWREADY : OUT STD_LOGIC;
    x_rsc_1_0_AWVALID : IN STD_LOGIC;
    x_rsc_1_0_AWUSER : IN STD_LOGIC;
    x_rsc_1_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_1_0_AWLOCK : IN STD_LOGIC;
    x_rsc_1_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_1_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_1_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_1_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_1_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    x_rsc_2_0_s_tdone : IN STD_LOGIC;
    x_rsc_2_0_tr_write_done : IN STD_LOGIC;
    x_rsc_2_0_RREADY : IN STD_LOGIC;
    x_rsc_2_0_RVALID : OUT STD_LOGIC;
    x_rsc_2_0_RUSER : OUT STD_LOGIC;
    x_rsc_2_0_RLAST : OUT STD_LOGIC;
    x_rsc_2_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_RID : OUT STD_LOGIC;
    x_rsc_2_0_ARREADY : OUT STD_LOGIC;
    x_rsc_2_0_ARVALID : IN STD_LOGIC;
    x_rsc_2_0_ARUSER : IN STD_LOGIC;
    x_rsc_2_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_ARLOCK : IN STD_LOGIC;
    x_rsc_2_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_2_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_2_0_ARID : IN STD_LOGIC;
    x_rsc_2_0_BREADY : IN STD_LOGIC;
    x_rsc_2_0_BVALID : OUT STD_LOGIC;
    x_rsc_2_0_BUSER : OUT STD_LOGIC;
    x_rsc_2_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_BID : OUT STD_LOGIC;
    x_rsc_2_0_WREADY : OUT STD_LOGIC;
    x_rsc_2_0_WVALID : IN STD_LOGIC;
    x_rsc_2_0_WUSER : IN STD_LOGIC;
    x_rsc_2_0_WLAST : IN STD_LOGIC;
    x_rsc_2_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_2_0_AWREADY : OUT STD_LOGIC;
    x_rsc_2_0_AWVALID : IN STD_LOGIC;
    x_rsc_2_0_AWUSER : IN STD_LOGIC;
    x_rsc_2_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_2_0_AWLOCK : IN STD_LOGIC;
    x_rsc_2_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_2_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_2_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_2_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_2_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_2_0_lz : OUT STD_LOGIC;
    x_rsc_3_0_s_tdone : IN STD_LOGIC;
    x_rsc_3_0_tr_write_done : IN STD_LOGIC;
    x_rsc_3_0_RREADY : IN STD_LOGIC;
    x_rsc_3_0_RVALID : OUT STD_LOGIC;
    x_rsc_3_0_RUSER : OUT STD_LOGIC;
    x_rsc_3_0_RLAST : OUT STD_LOGIC;
    x_rsc_3_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_RID : OUT STD_LOGIC;
    x_rsc_3_0_ARREADY : OUT STD_LOGIC;
    x_rsc_3_0_ARVALID : IN STD_LOGIC;
    x_rsc_3_0_ARUSER : IN STD_LOGIC;
    x_rsc_3_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_ARLOCK : IN STD_LOGIC;
    x_rsc_3_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_3_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_3_0_ARID : IN STD_LOGIC;
    x_rsc_3_0_BREADY : IN STD_LOGIC;
    x_rsc_3_0_BVALID : OUT STD_LOGIC;
    x_rsc_3_0_BUSER : OUT STD_LOGIC;
    x_rsc_3_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_BID : OUT STD_LOGIC;
    x_rsc_3_0_WREADY : OUT STD_LOGIC;
    x_rsc_3_0_WVALID : IN STD_LOGIC;
    x_rsc_3_0_WUSER : IN STD_LOGIC;
    x_rsc_3_0_WLAST : IN STD_LOGIC;
    x_rsc_3_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_3_0_AWREADY : OUT STD_LOGIC;
    x_rsc_3_0_AWVALID : IN STD_LOGIC;
    x_rsc_3_0_AWUSER : IN STD_LOGIC;
    x_rsc_3_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_3_0_AWLOCK : IN STD_LOGIC;
    x_rsc_3_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_3_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_3_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_3_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_3_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_3_0_lz : OUT STD_LOGIC;
    x_rsc_4_0_s_tdone : IN STD_LOGIC;
    x_rsc_4_0_tr_write_done : IN STD_LOGIC;
    x_rsc_4_0_RREADY : IN STD_LOGIC;
    x_rsc_4_0_RVALID : OUT STD_LOGIC;
    x_rsc_4_0_RUSER : OUT STD_LOGIC;
    x_rsc_4_0_RLAST : OUT STD_LOGIC;
    x_rsc_4_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_RID : OUT STD_LOGIC;
    x_rsc_4_0_ARREADY : OUT STD_LOGIC;
    x_rsc_4_0_ARVALID : IN STD_LOGIC;
    x_rsc_4_0_ARUSER : IN STD_LOGIC;
    x_rsc_4_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_ARLOCK : IN STD_LOGIC;
    x_rsc_4_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_4_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_4_0_ARID : IN STD_LOGIC;
    x_rsc_4_0_BREADY : IN STD_LOGIC;
    x_rsc_4_0_BVALID : OUT STD_LOGIC;
    x_rsc_4_0_BUSER : OUT STD_LOGIC;
    x_rsc_4_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_BID : OUT STD_LOGIC;
    x_rsc_4_0_WREADY : OUT STD_LOGIC;
    x_rsc_4_0_WVALID : IN STD_LOGIC;
    x_rsc_4_0_WUSER : IN STD_LOGIC;
    x_rsc_4_0_WLAST : IN STD_LOGIC;
    x_rsc_4_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_4_0_AWREADY : OUT STD_LOGIC;
    x_rsc_4_0_AWVALID : IN STD_LOGIC;
    x_rsc_4_0_AWUSER : IN STD_LOGIC;
    x_rsc_4_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_4_0_AWLOCK : IN STD_LOGIC;
    x_rsc_4_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_4_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_4_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_4_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_4_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_4_0_lz : OUT STD_LOGIC;
    x_rsc_5_0_s_tdone : IN STD_LOGIC;
    x_rsc_5_0_tr_write_done : IN STD_LOGIC;
    x_rsc_5_0_RREADY : IN STD_LOGIC;
    x_rsc_5_0_RVALID : OUT STD_LOGIC;
    x_rsc_5_0_RUSER : OUT STD_LOGIC;
    x_rsc_5_0_RLAST : OUT STD_LOGIC;
    x_rsc_5_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_RID : OUT STD_LOGIC;
    x_rsc_5_0_ARREADY : OUT STD_LOGIC;
    x_rsc_5_0_ARVALID : IN STD_LOGIC;
    x_rsc_5_0_ARUSER : IN STD_LOGIC;
    x_rsc_5_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_ARLOCK : IN STD_LOGIC;
    x_rsc_5_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_5_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_5_0_ARID : IN STD_LOGIC;
    x_rsc_5_0_BREADY : IN STD_LOGIC;
    x_rsc_5_0_BVALID : OUT STD_LOGIC;
    x_rsc_5_0_BUSER : OUT STD_LOGIC;
    x_rsc_5_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_BID : OUT STD_LOGIC;
    x_rsc_5_0_WREADY : OUT STD_LOGIC;
    x_rsc_5_0_WVALID : IN STD_LOGIC;
    x_rsc_5_0_WUSER : IN STD_LOGIC;
    x_rsc_5_0_WLAST : IN STD_LOGIC;
    x_rsc_5_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_5_0_AWREADY : OUT STD_LOGIC;
    x_rsc_5_0_AWVALID : IN STD_LOGIC;
    x_rsc_5_0_AWUSER : IN STD_LOGIC;
    x_rsc_5_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_5_0_AWLOCK : IN STD_LOGIC;
    x_rsc_5_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_5_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_5_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_5_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_5_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_5_0_lz : OUT STD_LOGIC;
    x_rsc_6_0_s_tdone : IN STD_LOGIC;
    x_rsc_6_0_tr_write_done : IN STD_LOGIC;
    x_rsc_6_0_RREADY : IN STD_LOGIC;
    x_rsc_6_0_RVALID : OUT STD_LOGIC;
    x_rsc_6_0_RUSER : OUT STD_LOGIC;
    x_rsc_6_0_RLAST : OUT STD_LOGIC;
    x_rsc_6_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_RID : OUT STD_LOGIC;
    x_rsc_6_0_ARREADY : OUT STD_LOGIC;
    x_rsc_6_0_ARVALID : IN STD_LOGIC;
    x_rsc_6_0_ARUSER : IN STD_LOGIC;
    x_rsc_6_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_ARLOCK : IN STD_LOGIC;
    x_rsc_6_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_6_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_6_0_ARID : IN STD_LOGIC;
    x_rsc_6_0_BREADY : IN STD_LOGIC;
    x_rsc_6_0_BVALID : OUT STD_LOGIC;
    x_rsc_6_0_BUSER : OUT STD_LOGIC;
    x_rsc_6_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_BID : OUT STD_LOGIC;
    x_rsc_6_0_WREADY : OUT STD_LOGIC;
    x_rsc_6_0_WVALID : IN STD_LOGIC;
    x_rsc_6_0_WUSER : IN STD_LOGIC;
    x_rsc_6_0_WLAST : IN STD_LOGIC;
    x_rsc_6_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_6_0_AWREADY : OUT STD_LOGIC;
    x_rsc_6_0_AWVALID : IN STD_LOGIC;
    x_rsc_6_0_AWUSER : IN STD_LOGIC;
    x_rsc_6_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_6_0_AWLOCK : IN STD_LOGIC;
    x_rsc_6_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_6_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_6_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_6_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_6_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_6_0_lz : OUT STD_LOGIC;
    x_rsc_7_0_s_tdone : IN STD_LOGIC;
    x_rsc_7_0_tr_write_done : IN STD_LOGIC;
    x_rsc_7_0_RREADY : IN STD_LOGIC;
    x_rsc_7_0_RVALID : OUT STD_LOGIC;
    x_rsc_7_0_RUSER : OUT STD_LOGIC;
    x_rsc_7_0_RLAST : OUT STD_LOGIC;
    x_rsc_7_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_RID : OUT STD_LOGIC;
    x_rsc_7_0_ARREADY : OUT STD_LOGIC;
    x_rsc_7_0_ARVALID : IN STD_LOGIC;
    x_rsc_7_0_ARUSER : IN STD_LOGIC;
    x_rsc_7_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_ARLOCK : IN STD_LOGIC;
    x_rsc_7_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_7_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_7_0_ARID : IN STD_LOGIC;
    x_rsc_7_0_BREADY : IN STD_LOGIC;
    x_rsc_7_0_BVALID : OUT STD_LOGIC;
    x_rsc_7_0_BUSER : OUT STD_LOGIC;
    x_rsc_7_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_BID : OUT STD_LOGIC;
    x_rsc_7_0_WREADY : OUT STD_LOGIC;
    x_rsc_7_0_WVALID : IN STD_LOGIC;
    x_rsc_7_0_WUSER : IN STD_LOGIC;
    x_rsc_7_0_WLAST : IN STD_LOGIC;
    x_rsc_7_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_7_0_AWREADY : OUT STD_LOGIC;
    x_rsc_7_0_AWVALID : IN STD_LOGIC;
    x_rsc_7_0_AWUSER : IN STD_LOGIC;
    x_rsc_7_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_7_0_AWLOCK : IN STD_LOGIC;
    x_rsc_7_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_7_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_7_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_7_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_7_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_7_0_lz : OUT STD_LOGIC;
    x_rsc_8_0_s_tdone : IN STD_LOGIC;
    x_rsc_8_0_tr_write_done : IN STD_LOGIC;
    x_rsc_8_0_RREADY : IN STD_LOGIC;
    x_rsc_8_0_RVALID : OUT STD_LOGIC;
    x_rsc_8_0_RUSER : OUT STD_LOGIC;
    x_rsc_8_0_RLAST : OUT STD_LOGIC;
    x_rsc_8_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_RID : OUT STD_LOGIC;
    x_rsc_8_0_ARREADY : OUT STD_LOGIC;
    x_rsc_8_0_ARVALID : IN STD_LOGIC;
    x_rsc_8_0_ARUSER : IN STD_LOGIC;
    x_rsc_8_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_ARLOCK : IN STD_LOGIC;
    x_rsc_8_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_8_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_8_0_ARID : IN STD_LOGIC;
    x_rsc_8_0_BREADY : IN STD_LOGIC;
    x_rsc_8_0_BVALID : OUT STD_LOGIC;
    x_rsc_8_0_BUSER : OUT STD_LOGIC;
    x_rsc_8_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_BID : OUT STD_LOGIC;
    x_rsc_8_0_WREADY : OUT STD_LOGIC;
    x_rsc_8_0_WVALID : IN STD_LOGIC;
    x_rsc_8_0_WUSER : IN STD_LOGIC;
    x_rsc_8_0_WLAST : IN STD_LOGIC;
    x_rsc_8_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_8_0_AWREADY : OUT STD_LOGIC;
    x_rsc_8_0_AWVALID : IN STD_LOGIC;
    x_rsc_8_0_AWUSER : IN STD_LOGIC;
    x_rsc_8_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_8_0_AWLOCK : IN STD_LOGIC;
    x_rsc_8_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_8_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_8_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_8_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_8_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_8_0_lz : OUT STD_LOGIC;
    x_rsc_9_0_s_tdone : IN STD_LOGIC;
    x_rsc_9_0_tr_write_done : IN STD_LOGIC;
    x_rsc_9_0_RREADY : IN STD_LOGIC;
    x_rsc_9_0_RVALID : OUT STD_LOGIC;
    x_rsc_9_0_RUSER : OUT STD_LOGIC;
    x_rsc_9_0_RLAST : OUT STD_LOGIC;
    x_rsc_9_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_RID : OUT STD_LOGIC;
    x_rsc_9_0_ARREADY : OUT STD_LOGIC;
    x_rsc_9_0_ARVALID : IN STD_LOGIC;
    x_rsc_9_0_ARUSER : IN STD_LOGIC;
    x_rsc_9_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_ARLOCK : IN STD_LOGIC;
    x_rsc_9_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_9_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_9_0_ARID : IN STD_LOGIC;
    x_rsc_9_0_BREADY : IN STD_LOGIC;
    x_rsc_9_0_BVALID : OUT STD_LOGIC;
    x_rsc_9_0_BUSER : OUT STD_LOGIC;
    x_rsc_9_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_BID : OUT STD_LOGIC;
    x_rsc_9_0_WREADY : OUT STD_LOGIC;
    x_rsc_9_0_WVALID : IN STD_LOGIC;
    x_rsc_9_0_WUSER : IN STD_LOGIC;
    x_rsc_9_0_WLAST : IN STD_LOGIC;
    x_rsc_9_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_9_0_AWREADY : OUT STD_LOGIC;
    x_rsc_9_0_AWVALID : IN STD_LOGIC;
    x_rsc_9_0_AWUSER : IN STD_LOGIC;
    x_rsc_9_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_9_0_AWLOCK : IN STD_LOGIC;
    x_rsc_9_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_9_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_9_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_9_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_9_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_9_0_lz : OUT STD_LOGIC;
    x_rsc_10_0_s_tdone : IN STD_LOGIC;
    x_rsc_10_0_tr_write_done : IN STD_LOGIC;
    x_rsc_10_0_RREADY : IN STD_LOGIC;
    x_rsc_10_0_RVALID : OUT STD_LOGIC;
    x_rsc_10_0_RUSER : OUT STD_LOGIC;
    x_rsc_10_0_RLAST : OUT STD_LOGIC;
    x_rsc_10_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_RID : OUT STD_LOGIC;
    x_rsc_10_0_ARREADY : OUT STD_LOGIC;
    x_rsc_10_0_ARVALID : IN STD_LOGIC;
    x_rsc_10_0_ARUSER : IN STD_LOGIC;
    x_rsc_10_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_ARLOCK : IN STD_LOGIC;
    x_rsc_10_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_10_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_10_0_ARID : IN STD_LOGIC;
    x_rsc_10_0_BREADY : IN STD_LOGIC;
    x_rsc_10_0_BVALID : OUT STD_LOGIC;
    x_rsc_10_0_BUSER : OUT STD_LOGIC;
    x_rsc_10_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_BID : OUT STD_LOGIC;
    x_rsc_10_0_WREADY : OUT STD_LOGIC;
    x_rsc_10_0_WVALID : IN STD_LOGIC;
    x_rsc_10_0_WUSER : IN STD_LOGIC;
    x_rsc_10_0_WLAST : IN STD_LOGIC;
    x_rsc_10_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_10_0_AWREADY : OUT STD_LOGIC;
    x_rsc_10_0_AWVALID : IN STD_LOGIC;
    x_rsc_10_0_AWUSER : IN STD_LOGIC;
    x_rsc_10_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_10_0_AWLOCK : IN STD_LOGIC;
    x_rsc_10_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_10_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_10_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_10_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_10_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_10_0_lz : OUT STD_LOGIC;
    x_rsc_11_0_s_tdone : IN STD_LOGIC;
    x_rsc_11_0_tr_write_done : IN STD_LOGIC;
    x_rsc_11_0_RREADY : IN STD_LOGIC;
    x_rsc_11_0_RVALID : OUT STD_LOGIC;
    x_rsc_11_0_RUSER : OUT STD_LOGIC;
    x_rsc_11_0_RLAST : OUT STD_LOGIC;
    x_rsc_11_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_RID : OUT STD_LOGIC;
    x_rsc_11_0_ARREADY : OUT STD_LOGIC;
    x_rsc_11_0_ARVALID : IN STD_LOGIC;
    x_rsc_11_0_ARUSER : IN STD_LOGIC;
    x_rsc_11_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_ARLOCK : IN STD_LOGIC;
    x_rsc_11_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_11_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_11_0_ARID : IN STD_LOGIC;
    x_rsc_11_0_BREADY : IN STD_LOGIC;
    x_rsc_11_0_BVALID : OUT STD_LOGIC;
    x_rsc_11_0_BUSER : OUT STD_LOGIC;
    x_rsc_11_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_BID : OUT STD_LOGIC;
    x_rsc_11_0_WREADY : OUT STD_LOGIC;
    x_rsc_11_0_WVALID : IN STD_LOGIC;
    x_rsc_11_0_WUSER : IN STD_LOGIC;
    x_rsc_11_0_WLAST : IN STD_LOGIC;
    x_rsc_11_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_11_0_AWREADY : OUT STD_LOGIC;
    x_rsc_11_0_AWVALID : IN STD_LOGIC;
    x_rsc_11_0_AWUSER : IN STD_LOGIC;
    x_rsc_11_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_11_0_AWLOCK : IN STD_LOGIC;
    x_rsc_11_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_11_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_11_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_11_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_11_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_11_0_lz : OUT STD_LOGIC;
    x_rsc_12_0_s_tdone : IN STD_LOGIC;
    x_rsc_12_0_tr_write_done : IN STD_LOGIC;
    x_rsc_12_0_RREADY : IN STD_LOGIC;
    x_rsc_12_0_RVALID : OUT STD_LOGIC;
    x_rsc_12_0_RUSER : OUT STD_LOGIC;
    x_rsc_12_0_RLAST : OUT STD_LOGIC;
    x_rsc_12_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_RID : OUT STD_LOGIC;
    x_rsc_12_0_ARREADY : OUT STD_LOGIC;
    x_rsc_12_0_ARVALID : IN STD_LOGIC;
    x_rsc_12_0_ARUSER : IN STD_LOGIC;
    x_rsc_12_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_ARLOCK : IN STD_LOGIC;
    x_rsc_12_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_12_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_12_0_ARID : IN STD_LOGIC;
    x_rsc_12_0_BREADY : IN STD_LOGIC;
    x_rsc_12_0_BVALID : OUT STD_LOGIC;
    x_rsc_12_0_BUSER : OUT STD_LOGIC;
    x_rsc_12_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_BID : OUT STD_LOGIC;
    x_rsc_12_0_WREADY : OUT STD_LOGIC;
    x_rsc_12_0_WVALID : IN STD_LOGIC;
    x_rsc_12_0_WUSER : IN STD_LOGIC;
    x_rsc_12_0_WLAST : IN STD_LOGIC;
    x_rsc_12_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_12_0_AWREADY : OUT STD_LOGIC;
    x_rsc_12_0_AWVALID : IN STD_LOGIC;
    x_rsc_12_0_AWUSER : IN STD_LOGIC;
    x_rsc_12_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_12_0_AWLOCK : IN STD_LOGIC;
    x_rsc_12_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_12_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_12_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_12_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_12_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_12_0_lz : OUT STD_LOGIC;
    x_rsc_13_0_s_tdone : IN STD_LOGIC;
    x_rsc_13_0_tr_write_done : IN STD_LOGIC;
    x_rsc_13_0_RREADY : IN STD_LOGIC;
    x_rsc_13_0_RVALID : OUT STD_LOGIC;
    x_rsc_13_0_RUSER : OUT STD_LOGIC;
    x_rsc_13_0_RLAST : OUT STD_LOGIC;
    x_rsc_13_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_RID : OUT STD_LOGIC;
    x_rsc_13_0_ARREADY : OUT STD_LOGIC;
    x_rsc_13_0_ARVALID : IN STD_LOGIC;
    x_rsc_13_0_ARUSER : IN STD_LOGIC;
    x_rsc_13_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_ARLOCK : IN STD_LOGIC;
    x_rsc_13_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_13_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_13_0_ARID : IN STD_LOGIC;
    x_rsc_13_0_BREADY : IN STD_LOGIC;
    x_rsc_13_0_BVALID : OUT STD_LOGIC;
    x_rsc_13_0_BUSER : OUT STD_LOGIC;
    x_rsc_13_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_BID : OUT STD_LOGIC;
    x_rsc_13_0_WREADY : OUT STD_LOGIC;
    x_rsc_13_0_WVALID : IN STD_LOGIC;
    x_rsc_13_0_WUSER : IN STD_LOGIC;
    x_rsc_13_0_WLAST : IN STD_LOGIC;
    x_rsc_13_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_13_0_AWREADY : OUT STD_LOGIC;
    x_rsc_13_0_AWVALID : IN STD_LOGIC;
    x_rsc_13_0_AWUSER : IN STD_LOGIC;
    x_rsc_13_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_13_0_AWLOCK : IN STD_LOGIC;
    x_rsc_13_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_13_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_13_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_13_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_13_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_13_0_lz : OUT STD_LOGIC;
    x_rsc_14_0_s_tdone : IN STD_LOGIC;
    x_rsc_14_0_tr_write_done : IN STD_LOGIC;
    x_rsc_14_0_RREADY : IN STD_LOGIC;
    x_rsc_14_0_RVALID : OUT STD_LOGIC;
    x_rsc_14_0_RUSER : OUT STD_LOGIC;
    x_rsc_14_0_RLAST : OUT STD_LOGIC;
    x_rsc_14_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_RID : OUT STD_LOGIC;
    x_rsc_14_0_ARREADY : OUT STD_LOGIC;
    x_rsc_14_0_ARVALID : IN STD_LOGIC;
    x_rsc_14_0_ARUSER : IN STD_LOGIC;
    x_rsc_14_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_ARLOCK : IN STD_LOGIC;
    x_rsc_14_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_14_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_14_0_ARID : IN STD_LOGIC;
    x_rsc_14_0_BREADY : IN STD_LOGIC;
    x_rsc_14_0_BVALID : OUT STD_LOGIC;
    x_rsc_14_0_BUSER : OUT STD_LOGIC;
    x_rsc_14_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_BID : OUT STD_LOGIC;
    x_rsc_14_0_WREADY : OUT STD_LOGIC;
    x_rsc_14_0_WVALID : IN STD_LOGIC;
    x_rsc_14_0_WUSER : IN STD_LOGIC;
    x_rsc_14_0_WLAST : IN STD_LOGIC;
    x_rsc_14_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_14_0_AWREADY : OUT STD_LOGIC;
    x_rsc_14_0_AWVALID : IN STD_LOGIC;
    x_rsc_14_0_AWUSER : IN STD_LOGIC;
    x_rsc_14_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_14_0_AWLOCK : IN STD_LOGIC;
    x_rsc_14_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_14_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_14_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_14_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_14_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_14_0_lz : OUT STD_LOGIC;
    x_rsc_15_0_s_tdone : IN STD_LOGIC;
    x_rsc_15_0_tr_write_done : IN STD_LOGIC;
    x_rsc_15_0_RREADY : IN STD_LOGIC;
    x_rsc_15_0_RVALID : OUT STD_LOGIC;
    x_rsc_15_0_RUSER : OUT STD_LOGIC;
    x_rsc_15_0_RLAST : OUT STD_LOGIC;
    x_rsc_15_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_RID : OUT STD_LOGIC;
    x_rsc_15_0_ARREADY : OUT STD_LOGIC;
    x_rsc_15_0_ARVALID : IN STD_LOGIC;
    x_rsc_15_0_ARUSER : IN STD_LOGIC;
    x_rsc_15_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_ARLOCK : IN STD_LOGIC;
    x_rsc_15_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_15_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_15_0_ARID : IN STD_LOGIC;
    x_rsc_15_0_BREADY : IN STD_LOGIC;
    x_rsc_15_0_BVALID : OUT STD_LOGIC;
    x_rsc_15_0_BUSER : OUT STD_LOGIC;
    x_rsc_15_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_BID : OUT STD_LOGIC;
    x_rsc_15_0_WREADY : OUT STD_LOGIC;
    x_rsc_15_0_WVALID : IN STD_LOGIC;
    x_rsc_15_0_WUSER : IN STD_LOGIC;
    x_rsc_15_0_WLAST : IN STD_LOGIC;
    x_rsc_15_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_15_0_AWREADY : OUT STD_LOGIC;
    x_rsc_15_0_AWVALID : IN STD_LOGIC;
    x_rsc_15_0_AWUSER : IN STD_LOGIC;
    x_rsc_15_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_15_0_AWLOCK : IN STD_LOGIC;
    x_rsc_15_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_15_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_15_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_15_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_15_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_15_0_lz : OUT STD_LOGIC;
    x_rsc_16_0_s_tdone : IN STD_LOGIC;
    x_rsc_16_0_tr_write_done : IN STD_LOGIC;
    x_rsc_16_0_RREADY : IN STD_LOGIC;
    x_rsc_16_0_RVALID : OUT STD_LOGIC;
    x_rsc_16_0_RUSER : OUT STD_LOGIC;
    x_rsc_16_0_RLAST : OUT STD_LOGIC;
    x_rsc_16_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_RID : OUT STD_LOGIC;
    x_rsc_16_0_ARREADY : OUT STD_LOGIC;
    x_rsc_16_0_ARVALID : IN STD_LOGIC;
    x_rsc_16_0_ARUSER : IN STD_LOGIC;
    x_rsc_16_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_ARLOCK : IN STD_LOGIC;
    x_rsc_16_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_16_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_16_0_ARID : IN STD_LOGIC;
    x_rsc_16_0_BREADY : IN STD_LOGIC;
    x_rsc_16_0_BVALID : OUT STD_LOGIC;
    x_rsc_16_0_BUSER : OUT STD_LOGIC;
    x_rsc_16_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_BID : OUT STD_LOGIC;
    x_rsc_16_0_WREADY : OUT STD_LOGIC;
    x_rsc_16_0_WVALID : IN STD_LOGIC;
    x_rsc_16_0_WUSER : IN STD_LOGIC;
    x_rsc_16_0_WLAST : IN STD_LOGIC;
    x_rsc_16_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_16_0_AWREADY : OUT STD_LOGIC;
    x_rsc_16_0_AWVALID : IN STD_LOGIC;
    x_rsc_16_0_AWUSER : IN STD_LOGIC;
    x_rsc_16_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_16_0_AWLOCK : IN STD_LOGIC;
    x_rsc_16_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_16_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_16_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_16_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_16_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_16_0_lz : OUT STD_LOGIC;
    x_rsc_17_0_s_tdone : IN STD_LOGIC;
    x_rsc_17_0_tr_write_done : IN STD_LOGIC;
    x_rsc_17_0_RREADY : IN STD_LOGIC;
    x_rsc_17_0_RVALID : OUT STD_LOGIC;
    x_rsc_17_0_RUSER : OUT STD_LOGIC;
    x_rsc_17_0_RLAST : OUT STD_LOGIC;
    x_rsc_17_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_RID : OUT STD_LOGIC;
    x_rsc_17_0_ARREADY : OUT STD_LOGIC;
    x_rsc_17_0_ARVALID : IN STD_LOGIC;
    x_rsc_17_0_ARUSER : IN STD_LOGIC;
    x_rsc_17_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_ARLOCK : IN STD_LOGIC;
    x_rsc_17_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_17_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_17_0_ARID : IN STD_LOGIC;
    x_rsc_17_0_BREADY : IN STD_LOGIC;
    x_rsc_17_0_BVALID : OUT STD_LOGIC;
    x_rsc_17_0_BUSER : OUT STD_LOGIC;
    x_rsc_17_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_BID : OUT STD_LOGIC;
    x_rsc_17_0_WREADY : OUT STD_LOGIC;
    x_rsc_17_0_WVALID : IN STD_LOGIC;
    x_rsc_17_0_WUSER : IN STD_LOGIC;
    x_rsc_17_0_WLAST : IN STD_LOGIC;
    x_rsc_17_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_17_0_AWREADY : OUT STD_LOGIC;
    x_rsc_17_0_AWVALID : IN STD_LOGIC;
    x_rsc_17_0_AWUSER : IN STD_LOGIC;
    x_rsc_17_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_17_0_AWLOCK : IN STD_LOGIC;
    x_rsc_17_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_17_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_17_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_17_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_17_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_17_0_lz : OUT STD_LOGIC;
    x_rsc_18_0_s_tdone : IN STD_LOGIC;
    x_rsc_18_0_tr_write_done : IN STD_LOGIC;
    x_rsc_18_0_RREADY : IN STD_LOGIC;
    x_rsc_18_0_RVALID : OUT STD_LOGIC;
    x_rsc_18_0_RUSER : OUT STD_LOGIC;
    x_rsc_18_0_RLAST : OUT STD_LOGIC;
    x_rsc_18_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_RID : OUT STD_LOGIC;
    x_rsc_18_0_ARREADY : OUT STD_LOGIC;
    x_rsc_18_0_ARVALID : IN STD_LOGIC;
    x_rsc_18_0_ARUSER : IN STD_LOGIC;
    x_rsc_18_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_ARLOCK : IN STD_LOGIC;
    x_rsc_18_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_18_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_18_0_ARID : IN STD_LOGIC;
    x_rsc_18_0_BREADY : IN STD_LOGIC;
    x_rsc_18_0_BVALID : OUT STD_LOGIC;
    x_rsc_18_0_BUSER : OUT STD_LOGIC;
    x_rsc_18_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_BID : OUT STD_LOGIC;
    x_rsc_18_0_WREADY : OUT STD_LOGIC;
    x_rsc_18_0_WVALID : IN STD_LOGIC;
    x_rsc_18_0_WUSER : IN STD_LOGIC;
    x_rsc_18_0_WLAST : IN STD_LOGIC;
    x_rsc_18_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_18_0_AWREADY : OUT STD_LOGIC;
    x_rsc_18_0_AWVALID : IN STD_LOGIC;
    x_rsc_18_0_AWUSER : IN STD_LOGIC;
    x_rsc_18_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_18_0_AWLOCK : IN STD_LOGIC;
    x_rsc_18_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_18_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_18_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_18_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_18_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_18_0_lz : OUT STD_LOGIC;
    x_rsc_19_0_s_tdone : IN STD_LOGIC;
    x_rsc_19_0_tr_write_done : IN STD_LOGIC;
    x_rsc_19_0_RREADY : IN STD_LOGIC;
    x_rsc_19_0_RVALID : OUT STD_LOGIC;
    x_rsc_19_0_RUSER : OUT STD_LOGIC;
    x_rsc_19_0_RLAST : OUT STD_LOGIC;
    x_rsc_19_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_RID : OUT STD_LOGIC;
    x_rsc_19_0_ARREADY : OUT STD_LOGIC;
    x_rsc_19_0_ARVALID : IN STD_LOGIC;
    x_rsc_19_0_ARUSER : IN STD_LOGIC;
    x_rsc_19_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_ARLOCK : IN STD_LOGIC;
    x_rsc_19_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_19_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_19_0_ARID : IN STD_LOGIC;
    x_rsc_19_0_BREADY : IN STD_LOGIC;
    x_rsc_19_0_BVALID : OUT STD_LOGIC;
    x_rsc_19_0_BUSER : OUT STD_LOGIC;
    x_rsc_19_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_BID : OUT STD_LOGIC;
    x_rsc_19_0_WREADY : OUT STD_LOGIC;
    x_rsc_19_0_WVALID : IN STD_LOGIC;
    x_rsc_19_0_WUSER : IN STD_LOGIC;
    x_rsc_19_0_WLAST : IN STD_LOGIC;
    x_rsc_19_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_19_0_AWREADY : OUT STD_LOGIC;
    x_rsc_19_0_AWVALID : IN STD_LOGIC;
    x_rsc_19_0_AWUSER : IN STD_LOGIC;
    x_rsc_19_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_19_0_AWLOCK : IN STD_LOGIC;
    x_rsc_19_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_19_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_19_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_19_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_19_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_19_0_lz : OUT STD_LOGIC;
    x_rsc_20_0_s_tdone : IN STD_LOGIC;
    x_rsc_20_0_tr_write_done : IN STD_LOGIC;
    x_rsc_20_0_RREADY : IN STD_LOGIC;
    x_rsc_20_0_RVALID : OUT STD_LOGIC;
    x_rsc_20_0_RUSER : OUT STD_LOGIC;
    x_rsc_20_0_RLAST : OUT STD_LOGIC;
    x_rsc_20_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_RID : OUT STD_LOGIC;
    x_rsc_20_0_ARREADY : OUT STD_LOGIC;
    x_rsc_20_0_ARVALID : IN STD_LOGIC;
    x_rsc_20_0_ARUSER : IN STD_LOGIC;
    x_rsc_20_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_ARLOCK : IN STD_LOGIC;
    x_rsc_20_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_20_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_20_0_ARID : IN STD_LOGIC;
    x_rsc_20_0_BREADY : IN STD_LOGIC;
    x_rsc_20_0_BVALID : OUT STD_LOGIC;
    x_rsc_20_0_BUSER : OUT STD_LOGIC;
    x_rsc_20_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_BID : OUT STD_LOGIC;
    x_rsc_20_0_WREADY : OUT STD_LOGIC;
    x_rsc_20_0_WVALID : IN STD_LOGIC;
    x_rsc_20_0_WUSER : IN STD_LOGIC;
    x_rsc_20_0_WLAST : IN STD_LOGIC;
    x_rsc_20_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_20_0_AWREADY : OUT STD_LOGIC;
    x_rsc_20_0_AWVALID : IN STD_LOGIC;
    x_rsc_20_0_AWUSER : IN STD_LOGIC;
    x_rsc_20_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_20_0_AWLOCK : IN STD_LOGIC;
    x_rsc_20_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_20_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_20_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_20_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_20_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_20_0_lz : OUT STD_LOGIC;
    x_rsc_21_0_s_tdone : IN STD_LOGIC;
    x_rsc_21_0_tr_write_done : IN STD_LOGIC;
    x_rsc_21_0_RREADY : IN STD_LOGIC;
    x_rsc_21_0_RVALID : OUT STD_LOGIC;
    x_rsc_21_0_RUSER : OUT STD_LOGIC;
    x_rsc_21_0_RLAST : OUT STD_LOGIC;
    x_rsc_21_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_RID : OUT STD_LOGIC;
    x_rsc_21_0_ARREADY : OUT STD_LOGIC;
    x_rsc_21_0_ARVALID : IN STD_LOGIC;
    x_rsc_21_0_ARUSER : IN STD_LOGIC;
    x_rsc_21_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_ARLOCK : IN STD_LOGIC;
    x_rsc_21_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_21_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_21_0_ARID : IN STD_LOGIC;
    x_rsc_21_0_BREADY : IN STD_LOGIC;
    x_rsc_21_0_BVALID : OUT STD_LOGIC;
    x_rsc_21_0_BUSER : OUT STD_LOGIC;
    x_rsc_21_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_BID : OUT STD_LOGIC;
    x_rsc_21_0_WREADY : OUT STD_LOGIC;
    x_rsc_21_0_WVALID : IN STD_LOGIC;
    x_rsc_21_0_WUSER : IN STD_LOGIC;
    x_rsc_21_0_WLAST : IN STD_LOGIC;
    x_rsc_21_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_21_0_AWREADY : OUT STD_LOGIC;
    x_rsc_21_0_AWVALID : IN STD_LOGIC;
    x_rsc_21_0_AWUSER : IN STD_LOGIC;
    x_rsc_21_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_21_0_AWLOCK : IN STD_LOGIC;
    x_rsc_21_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_21_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_21_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_21_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_21_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_21_0_lz : OUT STD_LOGIC;
    x_rsc_22_0_s_tdone : IN STD_LOGIC;
    x_rsc_22_0_tr_write_done : IN STD_LOGIC;
    x_rsc_22_0_RREADY : IN STD_LOGIC;
    x_rsc_22_0_RVALID : OUT STD_LOGIC;
    x_rsc_22_0_RUSER : OUT STD_LOGIC;
    x_rsc_22_0_RLAST : OUT STD_LOGIC;
    x_rsc_22_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_RID : OUT STD_LOGIC;
    x_rsc_22_0_ARREADY : OUT STD_LOGIC;
    x_rsc_22_0_ARVALID : IN STD_LOGIC;
    x_rsc_22_0_ARUSER : IN STD_LOGIC;
    x_rsc_22_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_ARLOCK : IN STD_LOGIC;
    x_rsc_22_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_22_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_22_0_ARID : IN STD_LOGIC;
    x_rsc_22_0_BREADY : IN STD_LOGIC;
    x_rsc_22_0_BVALID : OUT STD_LOGIC;
    x_rsc_22_0_BUSER : OUT STD_LOGIC;
    x_rsc_22_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_BID : OUT STD_LOGIC;
    x_rsc_22_0_WREADY : OUT STD_LOGIC;
    x_rsc_22_0_WVALID : IN STD_LOGIC;
    x_rsc_22_0_WUSER : IN STD_LOGIC;
    x_rsc_22_0_WLAST : IN STD_LOGIC;
    x_rsc_22_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_22_0_AWREADY : OUT STD_LOGIC;
    x_rsc_22_0_AWVALID : IN STD_LOGIC;
    x_rsc_22_0_AWUSER : IN STD_LOGIC;
    x_rsc_22_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_22_0_AWLOCK : IN STD_LOGIC;
    x_rsc_22_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_22_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_22_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_22_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_22_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_22_0_lz : OUT STD_LOGIC;
    x_rsc_23_0_s_tdone : IN STD_LOGIC;
    x_rsc_23_0_tr_write_done : IN STD_LOGIC;
    x_rsc_23_0_RREADY : IN STD_LOGIC;
    x_rsc_23_0_RVALID : OUT STD_LOGIC;
    x_rsc_23_0_RUSER : OUT STD_LOGIC;
    x_rsc_23_0_RLAST : OUT STD_LOGIC;
    x_rsc_23_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_RID : OUT STD_LOGIC;
    x_rsc_23_0_ARREADY : OUT STD_LOGIC;
    x_rsc_23_0_ARVALID : IN STD_LOGIC;
    x_rsc_23_0_ARUSER : IN STD_LOGIC;
    x_rsc_23_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_ARLOCK : IN STD_LOGIC;
    x_rsc_23_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_23_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_23_0_ARID : IN STD_LOGIC;
    x_rsc_23_0_BREADY : IN STD_LOGIC;
    x_rsc_23_0_BVALID : OUT STD_LOGIC;
    x_rsc_23_0_BUSER : OUT STD_LOGIC;
    x_rsc_23_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_BID : OUT STD_LOGIC;
    x_rsc_23_0_WREADY : OUT STD_LOGIC;
    x_rsc_23_0_WVALID : IN STD_LOGIC;
    x_rsc_23_0_WUSER : IN STD_LOGIC;
    x_rsc_23_0_WLAST : IN STD_LOGIC;
    x_rsc_23_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_23_0_AWREADY : OUT STD_LOGIC;
    x_rsc_23_0_AWVALID : IN STD_LOGIC;
    x_rsc_23_0_AWUSER : IN STD_LOGIC;
    x_rsc_23_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_23_0_AWLOCK : IN STD_LOGIC;
    x_rsc_23_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_23_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_23_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_23_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_23_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_23_0_lz : OUT STD_LOGIC;
    x_rsc_24_0_s_tdone : IN STD_LOGIC;
    x_rsc_24_0_tr_write_done : IN STD_LOGIC;
    x_rsc_24_0_RREADY : IN STD_LOGIC;
    x_rsc_24_0_RVALID : OUT STD_LOGIC;
    x_rsc_24_0_RUSER : OUT STD_LOGIC;
    x_rsc_24_0_RLAST : OUT STD_LOGIC;
    x_rsc_24_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_RID : OUT STD_LOGIC;
    x_rsc_24_0_ARREADY : OUT STD_LOGIC;
    x_rsc_24_0_ARVALID : IN STD_LOGIC;
    x_rsc_24_0_ARUSER : IN STD_LOGIC;
    x_rsc_24_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_ARLOCK : IN STD_LOGIC;
    x_rsc_24_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_24_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_24_0_ARID : IN STD_LOGIC;
    x_rsc_24_0_BREADY : IN STD_LOGIC;
    x_rsc_24_0_BVALID : OUT STD_LOGIC;
    x_rsc_24_0_BUSER : OUT STD_LOGIC;
    x_rsc_24_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_BID : OUT STD_LOGIC;
    x_rsc_24_0_WREADY : OUT STD_LOGIC;
    x_rsc_24_0_WVALID : IN STD_LOGIC;
    x_rsc_24_0_WUSER : IN STD_LOGIC;
    x_rsc_24_0_WLAST : IN STD_LOGIC;
    x_rsc_24_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_24_0_AWREADY : OUT STD_LOGIC;
    x_rsc_24_0_AWVALID : IN STD_LOGIC;
    x_rsc_24_0_AWUSER : IN STD_LOGIC;
    x_rsc_24_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_24_0_AWLOCK : IN STD_LOGIC;
    x_rsc_24_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_24_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_24_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_24_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_24_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_24_0_lz : OUT STD_LOGIC;
    x_rsc_25_0_s_tdone : IN STD_LOGIC;
    x_rsc_25_0_tr_write_done : IN STD_LOGIC;
    x_rsc_25_0_RREADY : IN STD_LOGIC;
    x_rsc_25_0_RVALID : OUT STD_LOGIC;
    x_rsc_25_0_RUSER : OUT STD_LOGIC;
    x_rsc_25_0_RLAST : OUT STD_LOGIC;
    x_rsc_25_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_RID : OUT STD_LOGIC;
    x_rsc_25_0_ARREADY : OUT STD_LOGIC;
    x_rsc_25_0_ARVALID : IN STD_LOGIC;
    x_rsc_25_0_ARUSER : IN STD_LOGIC;
    x_rsc_25_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_ARLOCK : IN STD_LOGIC;
    x_rsc_25_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_25_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_25_0_ARID : IN STD_LOGIC;
    x_rsc_25_0_BREADY : IN STD_LOGIC;
    x_rsc_25_0_BVALID : OUT STD_LOGIC;
    x_rsc_25_0_BUSER : OUT STD_LOGIC;
    x_rsc_25_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_BID : OUT STD_LOGIC;
    x_rsc_25_0_WREADY : OUT STD_LOGIC;
    x_rsc_25_0_WVALID : IN STD_LOGIC;
    x_rsc_25_0_WUSER : IN STD_LOGIC;
    x_rsc_25_0_WLAST : IN STD_LOGIC;
    x_rsc_25_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_25_0_AWREADY : OUT STD_LOGIC;
    x_rsc_25_0_AWVALID : IN STD_LOGIC;
    x_rsc_25_0_AWUSER : IN STD_LOGIC;
    x_rsc_25_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_25_0_AWLOCK : IN STD_LOGIC;
    x_rsc_25_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_25_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_25_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_25_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_25_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_25_0_lz : OUT STD_LOGIC;
    x_rsc_26_0_s_tdone : IN STD_LOGIC;
    x_rsc_26_0_tr_write_done : IN STD_LOGIC;
    x_rsc_26_0_RREADY : IN STD_LOGIC;
    x_rsc_26_0_RVALID : OUT STD_LOGIC;
    x_rsc_26_0_RUSER : OUT STD_LOGIC;
    x_rsc_26_0_RLAST : OUT STD_LOGIC;
    x_rsc_26_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_RID : OUT STD_LOGIC;
    x_rsc_26_0_ARREADY : OUT STD_LOGIC;
    x_rsc_26_0_ARVALID : IN STD_LOGIC;
    x_rsc_26_0_ARUSER : IN STD_LOGIC;
    x_rsc_26_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_ARLOCK : IN STD_LOGIC;
    x_rsc_26_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_26_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_26_0_ARID : IN STD_LOGIC;
    x_rsc_26_0_BREADY : IN STD_LOGIC;
    x_rsc_26_0_BVALID : OUT STD_LOGIC;
    x_rsc_26_0_BUSER : OUT STD_LOGIC;
    x_rsc_26_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_BID : OUT STD_LOGIC;
    x_rsc_26_0_WREADY : OUT STD_LOGIC;
    x_rsc_26_0_WVALID : IN STD_LOGIC;
    x_rsc_26_0_WUSER : IN STD_LOGIC;
    x_rsc_26_0_WLAST : IN STD_LOGIC;
    x_rsc_26_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_26_0_AWREADY : OUT STD_LOGIC;
    x_rsc_26_0_AWVALID : IN STD_LOGIC;
    x_rsc_26_0_AWUSER : IN STD_LOGIC;
    x_rsc_26_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_26_0_AWLOCK : IN STD_LOGIC;
    x_rsc_26_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_26_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_26_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_26_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_26_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_26_0_lz : OUT STD_LOGIC;
    x_rsc_27_0_s_tdone : IN STD_LOGIC;
    x_rsc_27_0_tr_write_done : IN STD_LOGIC;
    x_rsc_27_0_RREADY : IN STD_LOGIC;
    x_rsc_27_0_RVALID : OUT STD_LOGIC;
    x_rsc_27_0_RUSER : OUT STD_LOGIC;
    x_rsc_27_0_RLAST : OUT STD_LOGIC;
    x_rsc_27_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_RID : OUT STD_LOGIC;
    x_rsc_27_0_ARREADY : OUT STD_LOGIC;
    x_rsc_27_0_ARVALID : IN STD_LOGIC;
    x_rsc_27_0_ARUSER : IN STD_LOGIC;
    x_rsc_27_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_ARLOCK : IN STD_LOGIC;
    x_rsc_27_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_27_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_27_0_ARID : IN STD_LOGIC;
    x_rsc_27_0_BREADY : IN STD_LOGIC;
    x_rsc_27_0_BVALID : OUT STD_LOGIC;
    x_rsc_27_0_BUSER : OUT STD_LOGIC;
    x_rsc_27_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_BID : OUT STD_LOGIC;
    x_rsc_27_0_WREADY : OUT STD_LOGIC;
    x_rsc_27_0_WVALID : IN STD_LOGIC;
    x_rsc_27_0_WUSER : IN STD_LOGIC;
    x_rsc_27_0_WLAST : IN STD_LOGIC;
    x_rsc_27_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_27_0_AWREADY : OUT STD_LOGIC;
    x_rsc_27_0_AWVALID : IN STD_LOGIC;
    x_rsc_27_0_AWUSER : IN STD_LOGIC;
    x_rsc_27_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_27_0_AWLOCK : IN STD_LOGIC;
    x_rsc_27_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_27_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_27_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_27_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_27_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_27_0_lz : OUT STD_LOGIC;
    x_rsc_28_0_s_tdone : IN STD_LOGIC;
    x_rsc_28_0_tr_write_done : IN STD_LOGIC;
    x_rsc_28_0_RREADY : IN STD_LOGIC;
    x_rsc_28_0_RVALID : OUT STD_LOGIC;
    x_rsc_28_0_RUSER : OUT STD_LOGIC;
    x_rsc_28_0_RLAST : OUT STD_LOGIC;
    x_rsc_28_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_RID : OUT STD_LOGIC;
    x_rsc_28_0_ARREADY : OUT STD_LOGIC;
    x_rsc_28_0_ARVALID : IN STD_LOGIC;
    x_rsc_28_0_ARUSER : IN STD_LOGIC;
    x_rsc_28_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_ARLOCK : IN STD_LOGIC;
    x_rsc_28_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_28_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_28_0_ARID : IN STD_LOGIC;
    x_rsc_28_0_BREADY : IN STD_LOGIC;
    x_rsc_28_0_BVALID : OUT STD_LOGIC;
    x_rsc_28_0_BUSER : OUT STD_LOGIC;
    x_rsc_28_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_BID : OUT STD_LOGIC;
    x_rsc_28_0_WREADY : OUT STD_LOGIC;
    x_rsc_28_0_WVALID : IN STD_LOGIC;
    x_rsc_28_0_WUSER : IN STD_LOGIC;
    x_rsc_28_0_WLAST : IN STD_LOGIC;
    x_rsc_28_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_28_0_AWREADY : OUT STD_LOGIC;
    x_rsc_28_0_AWVALID : IN STD_LOGIC;
    x_rsc_28_0_AWUSER : IN STD_LOGIC;
    x_rsc_28_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_28_0_AWLOCK : IN STD_LOGIC;
    x_rsc_28_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_28_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_28_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_28_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_28_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_28_0_lz : OUT STD_LOGIC;
    x_rsc_29_0_s_tdone : IN STD_LOGIC;
    x_rsc_29_0_tr_write_done : IN STD_LOGIC;
    x_rsc_29_0_RREADY : IN STD_LOGIC;
    x_rsc_29_0_RVALID : OUT STD_LOGIC;
    x_rsc_29_0_RUSER : OUT STD_LOGIC;
    x_rsc_29_0_RLAST : OUT STD_LOGIC;
    x_rsc_29_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_RID : OUT STD_LOGIC;
    x_rsc_29_0_ARREADY : OUT STD_LOGIC;
    x_rsc_29_0_ARVALID : IN STD_LOGIC;
    x_rsc_29_0_ARUSER : IN STD_LOGIC;
    x_rsc_29_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_ARLOCK : IN STD_LOGIC;
    x_rsc_29_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_29_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_29_0_ARID : IN STD_LOGIC;
    x_rsc_29_0_BREADY : IN STD_LOGIC;
    x_rsc_29_0_BVALID : OUT STD_LOGIC;
    x_rsc_29_0_BUSER : OUT STD_LOGIC;
    x_rsc_29_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_BID : OUT STD_LOGIC;
    x_rsc_29_0_WREADY : OUT STD_LOGIC;
    x_rsc_29_0_WVALID : IN STD_LOGIC;
    x_rsc_29_0_WUSER : IN STD_LOGIC;
    x_rsc_29_0_WLAST : IN STD_LOGIC;
    x_rsc_29_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_29_0_AWREADY : OUT STD_LOGIC;
    x_rsc_29_0_AWVALID : IN STD_LOGIC;
    x_rsc_29_0_AWUSER : IN STD_LOGIC;
    x_rsc_29_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_29_0_AWLOCK : IN STD_LOGIC;
    x_rsc_29_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_29_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_29_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_29_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_29_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_29_0_lz : OUT STD_LOGIC;
    x_rsc_30_0_s_tdone : IN STD_LOGIC;
    x_rsc_30_0_tr_write_done : IN STD_LOGIC;
    x_rsc_30_0_RREADY : IN STD_LOGIC;
    x_rsc_30_0_RVALID : OUT STD_LOGIC;
    x_rsc_30_0_RUSER : OUT STD_LOGIC;
    x_rsc_30_0_RLAST : OUT STD_LOGIC;
    x_rsc_30_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_RID : OUT STD_LOGIC;
    x_rsc_30_0_ARREADY : OUT STD_LOGIC;
    x_rsc_30_0_ARVALID : IN STD_LOGIC;
    x_rsc_30_0_ARUSER : IN STD_LOGIC;
    x_rsc_30_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_ARLOCK : IN STD_LOGIC;
    x_rsc_30_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_30_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_30_0_ARID : IN STD_LOGIC;
    x_rsc_30_0_BREADY : IN STD_LOGIC;
    x_rsc_30_0_BVALID : OUT STD_LOGIC;
    x_rsc_30_0_BUSER : OUT STD_LOGIC;
    x_rsc_30_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_BID : OUT STD_LOGIC;
    x_rsc_30_0_WREADY : OUT STD_LOGIC;
    x_rsc_30_0_WVALID : IN STD_LOGIC;
    x_rsc_30_0_WUSER : IN STD_LOGIC;
    x_rsc_30_0_WLAST : IN STD_LOGIC;
    x_rsc_30_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_30_0_AWREADY : OUT STD_LOGIC;
    x_rsc_30_0_AWVALID : IN STD_LOGIC;
    x_rsc_30_0_AWUSER : IN STD_LOGIC;
    x_rsc_30_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_30_0_AWLOCK : IN STD_LOGIC;
    x_rsc_30_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_30_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_30_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_30_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_30_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_30_0_lz : OUT STD_LOGIC;
    x_rsc_31_0_s_tdone : IN STD_LOGIC;
    x_rsc_31_0_tr_write_done : IN STD_LOGIC;
    x_rsc_31_0_RREADY : IN STD_LOGIC;
    x_rsc_31_0_RVALID : OUT STD_LOGIC;
    x_rsc_31_0_RUSER : OUT STD_LOGIC;
    x_rsc_31_0_RLAST : OUT STD_LOGIC;
    x_rsc_31_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_RID : OUT STD_LOGIC;
    x_rsc_31_0_ARREADY : OUT STD_LOGIC;
    x_rsc_31_0_ARVALID : IN STD_LOGIC;
    x_rsc_31_0_ARUSER : IN STD_LOGIC;
    x_rsc_31_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_ARLOCK : IN STD_LOGIC;
    x_rsc_31_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_31_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_31_0_ARID : IN STD_LOGIC;
    x_rsc_31_0_BREADY : IN STD_LOGIC;
    x_rsc_31_0_BVALID : OUT STD_LOGIC;
    x_rsc_31_0_BUSER : OUT STD_LOGIC;
    x_rsc_31_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_BID : OUT STD_LOGIC;
    x_rsc_31_0_WREADY : OUT STD_LOGIC;
    x_rsc_31_0_WVALID : IN STD_LOGIC;
    x_rsc_31_0_WUSER : IN STD_LOGIC;
    x_rsc_31_0_WLAST : IN STD_LOGIC;
    x_rsc_31_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    x_rsc_31_0_AWREADY : OUT STD_LOGIC;
    x_rsc_31_0_AWVALID : IN STD_LOGIC;
    x_rsc_31_0_AWUSER : IN STD_LOGIC;
    x_rsc_31_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    x_rsc_31_0_AWLOCK : IN STD_LOGIC;
    x_rsc_31_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    x_rsc_31_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    x_rsc_31_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    x_rsc_31_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    x_rsc_31_0_AWID : IN STD_LOGIC;
    x_rsc_triosy_31_0_lz : OUT STD_LOGIC;
    m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    m_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_rsc_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_h_rsc_adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
    twiddle_h_rsc_qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_triosy_lz : OUT STD_LOGIC;
    revArr_rsc_s_tdone : IN STD_LOGIC;
    revArr_rsc_tr_write_done : IN STD_LOGIC;
    revArr_rsc_RREADY : IN STD_LOGIC;
    revArr_rsc_RVALID : OUT STD_LOGIC;
    revArr_rsc_RUSER : OUT STD_LOGIC;
    revArr_rsc_RLAST : OUT STD_LOGIC;
    revArr_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    revArr_rsc_RID : OUT STD_LOGIC;
    revArr_rsc_ARREADY : OUT STD_LOGIC;
    revArr_rsc_ARVALID : IN STD_LOGIC;
    revArr_rsc_ARUSER : IN STD_LOGIC;
    revArr_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_ARLOCK : IN STD_LOGIC;
    revArr_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    revArr_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    revArr_rsc_ARID : IN STD_LOGIC;
    revArr_rsc_BREADY : IN STD_LOGIC;
    revArr_rsc_BVALID : OUT STD_LOGIC;
    revArr_rsc_BUSER : OUT STD_LOGIC;
    revArr_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_BID : OUT STD_LOGIC;
    revArr_rsc_WREADY : OUT STD_LOGIC;
    revArr_rsc_WVALID : IN STD_LOGIC;
    revArr_rsc_WUSER : IN STD_LOGIC;
    revArr_rsc_WLAST : IN STD_LOGIC;
    revArr_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    revArr_rsc_AWREADY : OUT STD_LOGIC;
    revArr_rsc_AWVALID : IN STD_LOGIC;
    revArr_rsc_AWUSER : IN STD_LOGIC;
    revArr_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    revArr_rsc_AWLOCK : IN STD_LOGIC;
    revArr_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    revArr_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    revArr_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    revArr_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    revArr_rsc_AWID : IN STD_LOGIC;
    revArr_rsc_triosy_lz : OUT STD_LOGIC;
    tw_rsc_s_tdone : IN STD_LOGIC;
    tw_rsc_tr_write_done : IN STD_LOGIC;
    tw_rsc_RREADY : IN STD_LOGIC;
    tw_rsc_RVALID : OUT STD_LOGIC;
    tw_rsc_RUSER : OUT STD_LOGIC;
    tw_rsc_RLAST : OUT STD_LOGIC;
    tw_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_rsc_RID : OUT STD_LOGIC;
    tw_rsc_ARREADY : OUT STD_LOGIC;
    tw_rsc_ARVALID : IN STD_LOGIC;
    tw_rsc_ARUSER : IN STD_LOGIC;
    tw_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_ARLOCK : IN STD_LOGIC;
    tw_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_rsc_ARID : IN STD_LOGIC;
    tw_rsc_BREADY : IN STD_LOGIC;
    tw_rsc_BVALID : OUT STD_LOGIC;
    tw_rsc_BUSER : OUT STD_LOGIC;
    tw_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_BID : OUT STD_LOGIC;
    tw_rsc_WREADY : OUT STD_LOGIC;
    tw_rsc_WVALID : IN STD_LOGIC;
    tw_rsc_WUSER : IN STD_LOGIC;
    tw_rsc_WLAST : IN STD_LOGIC;
    tw_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_rsc_AWREADY : OUT STD_LOGIC;
    tw_rsc_AWVALID : IN STD_LOGIC;
    tw_rsc_AWUSER : IN STD_LOGIC;
    tw_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_rsc_AWLOCK : IN STD_LOGIC;
    tw_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_rsc_AWID : IN STD_LOGIC;
    tw_rsc_triosy_lz : OUT STD_LOGIC;
    tw_h_rsc_s_tdone : IN STD_LOGIC;
    tw_h_rsc_tr_write_done : IN STD_LOGIC;
    tw_h_rsc_RREADY : IN STD_LOGIC;
    tw_h_rsc_RVALID : OUT STD_LOGIC;
    tw_h_rsc_RUSER : OUT STD_LOGIC;
    tw_h_rsc_RLAST : OUT STD_LOGIC;
    tw_h_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_h_rsc_RID : OUT STD_LOGIC;
    tw_h_rsc_ARREADY : OUT STD_LOGIC;
    tw_h_rsc_ARVALID : IN STD_LOGIC;
    tw_h_rsc_ARUSER : IN STD_LOGIC;
    tw_h_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_ARLOCK : IN STD_LOGIC;
    tw_h_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_h_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_h_rsc_ARID : IN STD_LOGIC;
    tw_h_rsc_BREADY : IN STD_LOGIC;
    tw_h_rsc_BVALID : OUT STD_LOGIC;
    tw_h_rsc_BUSER : OUT STD_LOGIC;
    tw_h_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_BID : OUT STD_LOGIC;
    tw_h_rsc_WREADY : OUT STD_LOGIC;
    tw_h_rsc_WVALID : IN STD_LOGIC;
    tw_h_rsc_WUSER : IN STD_LOGIC;
    tw_h_rsc_WLAST : IN STD_LOGIC;
    tw_h_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    tw_h_rsc_AWREADY : OUT STD_LOGIC;
    tw_h_rsc_AWVALID : IN STD_LOGIC;
    tw_h_rsc_AWUSER : IN STD_LOGIC;
    tw_h_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    tw_h_rsc_AWLOCK : IN STD_LOGIC;
    tw_h_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    tw_h_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    tw_h_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    tw_h_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    tw_h_rsc_AWID : IN STD_LOGIC;
    tw_h_rsc_triosy_lz : OUT STD_LOGIC
  );
END hybrid;

ARCHITECTURE v14 OF hybrid IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsci_adrb_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsci_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL twiddle_h_rsci_adrb_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_h_rsci_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xx_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_2_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_2_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_3_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_3_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_4_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_4_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_5_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_5_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_6_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_6_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_7_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_7_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_8_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_8_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_9_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_9_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_10_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_10_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_11_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_11_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_12_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_12_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_13_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_13_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_14_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_14_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_15_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_15_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_16_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_16_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_17_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_17_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_18_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_18_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_19_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_19_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_20_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_20_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_21_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_21_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_22_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_22_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_23_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_23_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_24_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_24_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_25_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_25_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_26_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_26_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_27_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_27_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_28_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_28_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_29_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_29_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_30_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_30_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_31_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_clka_en_d : STD_LOGIC;
  SIGNAL xx_rsc_31_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_2_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_2_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_3_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_3_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_4_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_4_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_5_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_5_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_6_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_6_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_7_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_7_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_8_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_8_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_9_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_9_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_10_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_10_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_11_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_11_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_12_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_12_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_13_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_13_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_14_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_14_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_15_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_15_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_16_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_16_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_17_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_17_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_18_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_18_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_19_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_19_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_20_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_20_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_21_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_21_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_22_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_22_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_23_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_23_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_24_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_24_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_25_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_25_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_26_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_26_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_27_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_27_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_28_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_28_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_29_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_29_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_30_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_30_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_31_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_clka_en_d : STD_LOGIC;
  SIGNAL yy_rsc_31_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL S34_OUTER_LOOP_for_tf_mul_cmp_a : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL S34_OUTER_LOOP_for_tf_mul_cmp_b : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_0_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_0_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_0_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_web : STD_LOGIC;
  SIGNAL xx_rsc_0_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_0_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_0_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_1_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_1_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_1_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_web : STD_LOGIC;
  SIGNAL xx_rsc_1_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_1_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_1_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_2_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_2_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_2_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_web : STD_LOGIC;
  SIGNAL xx_rsc_2_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_2_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_2_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_3_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_3_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_3_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_web : STD_LOGIC;
  SIGNAL xx_rsc_3_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_3_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_3_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_4_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_4_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_4_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_web : STD_LOGIC;
  SIGNAL xx_rsc_4_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_4_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_4_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_5_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_5_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_5_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_web : STD_LOGIC;
  SIGNAL xx_rsc_5_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_5_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_5_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_6_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_6_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_6_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_web : STD_LOGIC;
  SIGNAL xx_rsc_6_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_6_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_6_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_7_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_7_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_7_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_web : STD_LOGIC;
  SIGNAL xx_rsc_7_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_7_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_7_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_8_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_8_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_8_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_web : STD_LOGIC;
  SIGNAL xx_rsc_8_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_8_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_8_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_9_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_9_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_9_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_web : STD_LOGIC;
  SIGNAL xx_rsc_9_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_9_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_9_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_10_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_10_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_10_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_web : STD_LOGIC;
  SIGNAL xx_rsc_10_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_10_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_10_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_11_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_11_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_11_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_web : STD_LOGIC;
  SIGNAL xx_rsc_11_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_11_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_11_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_12_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_12_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_12_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_web : STD_LOGIC;
  SIGNAL xx_rsc_12_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_12_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_12_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_13_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_13_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_13_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_web : STD_LOGIC;
  SIGNAL xx_rsc_13_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_13_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_13_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_14_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_14_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_14_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_web : STD_LOGIC;
  SIGNAL xx_rsc_14_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_14_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_14_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_15_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_15_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_15_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_web : STD_LOGIC;
  SIGNAL xx_rsc_15_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_15_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_15_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_16_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_16_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_16_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_web : STD_LOGIC;
  SIGNAL xx_rsc_16_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_16_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_16_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_17_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_17_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_17_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_web : STD_LOGIC;
  SIGNAL xx_rsc_17_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_17_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_17_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_18_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_18_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_18_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_web : STD_LOGIC;
  SIGNAL xx_rsc_18_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_18_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_18_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_19_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_19_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_19_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_web : STD_LOGIC;
  SIGNAL xx_rsc_19_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_19_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_19_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_20_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_20_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_20_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_web : STD_LOGIC;
  SIGNAL xx_rsc_20_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_20_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_20_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_21_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_21_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_21_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_web : STD_LOGIC;
  SIGNAL xx_rsc_21_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_21_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_21_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_22_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_22_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_22_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_web : STD_LOGIC;
  SIGNAL xx_rsc_22_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_22_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_22_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_23_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_23_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_23_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_web : STD_LOGIC;
  SIGNAL xx_rsc_23_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_23_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_23_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_24_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_24_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_24_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_web : STD_LOGIC;
  SIGNAL xx_rsc_24_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_24_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_24_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_25_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_25_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_25_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_web : STD_LOGIC;
  SIGNAL xx_rsc_25_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_25_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_25_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_26_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_26_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_26_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_web : STD_LOGIC;
  SIGNAL xx_rsc_26_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_26_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_26_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_27_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_27_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_27_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_web : STD_LOGIC;
  SIGNAL xx_rsc_27_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_27_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_27_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_28_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_28_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_28_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_web : STD_LOGIC;
  SIGNAL xx_rsc_28_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_28_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_28_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_29_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_29_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_29_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_web : STD_LOGIC;
  SIGNAL xx_rsc_29_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_29_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_29_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_30_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_30_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_30_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_web : STD_LOGIC;
  SIGNAL xx_rsc_30_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_30_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_30_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_31_0_clkb_en : STD_LOGIC;
  SIGNAL xx_rsc_31_0_clka_en : STD_LOGIC;
  SIGNAL xx_rsc_31_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_web : STD_LOGIC;
  SIGNAL xx_rsc_31_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_31_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_wea : STD_LOGIC;
  SIGNAL xx_rsc_31_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_0_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_0_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_0_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_web : STD_LOGIC;
  SIGNAL yy_rsc_0_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_0_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_0_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_1_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_1_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_1_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_web : STD_LOGIC;
  SIGNAL yy_rsc_1_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_1_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_1_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_2_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_2_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_2_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_web : STD_LOGIC;
  SIGNAL yy_rsc_2_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_2_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_2_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_3_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_3_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_3_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_web : STD_LOGIC;
  SIGNAL yy_rsc_3_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_3_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_3_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_4_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_4_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_4_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_web : STD_LOGIC;
  SIGNAL yy_rsc_4_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_4_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_4_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_5_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_5_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_5_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_web : STD_LOGIC;
  SIGNAL yy_rsc_5_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_5_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_5_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_6_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_6_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_6_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_web : STD_LOGIC;
  SIGNAL yy_rsc_6_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_6_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_6_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_7_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_7_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_7_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_web : STD_LOGIC;
  SIGNAL yy_rsc_7_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_7_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_7_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_8_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_8_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_8_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_web : STD_LOGIC;
  SIGNAL yy_rsc_8_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_8_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_8_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_9_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_9_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_9_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_web : STD_LOGIC;
  SIGNAL yy_rsc_9_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_9_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_9_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_10_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_10_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_10_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_web : STD_LOGIC;
  SIGNAL yy_rsc_10_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_10_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_10_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_11_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_11_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_11_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_web : STD_LOGIC;
  SIGNAL yy_rsc_11_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_11_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_11_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_12_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_12_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_12_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_web : STD_LOGIC;
  SIGNAL yy_rsc_12_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_12_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_12_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_13_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_13_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_13_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_web : STD_LOGIC;
  SIGNAL yy_rsc_13_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_13_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_13_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_14_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_14_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_14_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_web : STD_LOGIC;
  SIGNAL yy_rsc_14_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_14_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_14_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_15_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_15_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_15_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_web : STD_LOGIC;
  SIGNAL yy_rsc_15_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_15_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_15_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_16_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_16_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_16_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_web : STD_LOGIC;
  SIGNAL yy_rsc_16_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_16_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_16_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_17_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_17_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_17_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_web : STD_LOGIC;
  SIGNAL yy_rsc_17_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_17_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_17_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_18_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_18_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_18_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_web : STD_LOGIC;
  SIGNAL yy_rsc_18_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_18_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_18_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_19_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_19_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_19_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_web : STD_LOGIC;
  SIGNAL yy_rsc_19_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_19_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_19_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_20_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_20_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_20_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_web : STD_LOGIC;
  SIGNAL yy_rsc_20_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_20_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_20_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_21_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_21_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_21_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_web : STD_LOGIC;
  SIGNAL yy_rsc_21_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_21_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_21_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_22_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_22_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_22_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_web : STD_LOGIC;
  SIGNAL yy_rsc_22_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_22_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_22_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_23_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_23_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_23_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_web : STD_LOGIC;
  SIGNAL yy_rsc_23_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_23_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_23_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_24_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_24_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_24_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_web : STD_LOGIC;
  SIGNAL yy_rsc_24_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_24_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_24_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_25_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_25_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_25_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_web : STD_LOGIC;
  SIGNAL yy_rsc_25_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_25_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_25_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_26_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_26_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_26_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_web : STD_LOGIC;
  SIGNAL yy_rsc_26_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_26_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_26_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_27_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_27_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_27_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_web : STD_LOGIC;
  SIGNAL yy_rsc_27_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_27_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_27_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_28_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_28_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_28_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_web : STD_LOGIC;
  SIGNAL yy_rsc_28_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_28_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_28_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_29_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_29_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_29_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_web : STD_LOGIC;
  SIGNAL yy_rsc_29_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_29_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_29_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_30_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_30_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_30_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_web : STD_LOGIC;
  SIGNAL yy_rsc_30_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_30_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_30_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_31_0_clkb_en : STD_LOGIC;
  SIGNAL yy_rsc_31_0_clka_en : STD_LOGIC;
  SIGNAL yy_rsc_31_0_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_web : STD_LOGIC;
  SIGNAL yy_rsc_31_0_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_31_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_wea : STD_LOGIC;
  SIGNAL yy_rsc_31_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_da_d_iff : STD_LOGIC_VECTOR (63 DOWNTO 0);

  SIGNAL xx_rsc_0_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_0_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_0_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_1_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_1_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_1_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_2_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_2_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_2_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_3_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_3_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_3_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_4_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_4_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_4_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_5_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_5_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_5_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_6_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_6_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_6_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_7_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_7_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_7_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_8_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_8_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_8_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_9_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_9_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_9_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_10_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_10_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_10_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_11_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_11_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_11_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_12_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_12_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_12_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_13_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_13_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_13_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_14_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_14_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_14_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_15_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_15_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_15_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_16_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_16_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_16_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_17_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_17_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_17_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_18_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_18_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_18_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_19_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_19_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_19_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_20_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_20_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_20_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_21_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_21_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_21_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_22_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_22_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_22_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_23_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_23_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_23_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_24_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_24_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_24_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_25_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_25_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_25_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_26_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_26_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_26_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_27_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_27_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_27_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_28_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_28_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_28_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_29_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_29_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_29_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_30_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_30_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_30_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL xx_rsc_31_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_31_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_31_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_0_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_0_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_0_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_1_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_1_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_1_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_2_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_2_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_2_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_3_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_3_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_3_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_4_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_4_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_4_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_5_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_5_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_5_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_6_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_6_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_6_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_7_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_7_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_7_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_8_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_8_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_8_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_9_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_9_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_9_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_10_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_10_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_10_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_11_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_11_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_11_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_12_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_12_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_12_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_13_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_13_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_13_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_14_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_14_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_14_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_15_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_15_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_15_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_16_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_16_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_16_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_17_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_17_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_17_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_18_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_18_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_18_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_19_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_19_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_19_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_20_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_20_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_20_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_21_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_21_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_21_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_22_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_22_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_22_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_23_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_23_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_23_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_24_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_24_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_24_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_25_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_25_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_25_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_26_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_26_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_26_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_27_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_27_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_27_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_28_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_28_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_28_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_29_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_29_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_29_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_30_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_30_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_30_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yy_rsc_31_0_comp_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_31_0_comp_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_31_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_comp_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_3_5_32_32_32_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_rsci_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsci_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsci_adrb_d_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_rsci_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_4_5_32_32_32_32_1_gen
    PORT(
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adrb_d : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
      qb_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      readB_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL twiddle_h_rsci_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsci_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_h_rsci_adrb_d_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL twiddle_h_rsci_qb_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_1_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_2_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_3_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_4_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_5_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_6_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_7_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_8_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_9_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_10_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_11_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_12_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_13_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_14_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_15_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_16_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_17_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_18_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_19_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_20_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_21_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_22_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_23_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_24_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_25_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_26_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_27_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_28_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_39_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_29_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_40_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_30_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_41_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL xx_rsc_31_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_42_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_0_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_43_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_1_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_44_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_2_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_45_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_3_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_46_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_4_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_47_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_5_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_6_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_7_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_8_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_9_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_52_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_10_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_53_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_11_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_54_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_12_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_55_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_13_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_56_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_14_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_57_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_15_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_58_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_16_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_59_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_17_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_60_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_18_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_61_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_19_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_62_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_20_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_63_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_21_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_64_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_22_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_65_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_23_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_66_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_24_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_67_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_25_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_68_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_26_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_69_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_27_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_70_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_28_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_71_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_29_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_72_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_30_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_73_5_32_32_32_32_1_gen
    PORT(
      clkb_en : OUT STD_LOGIC;
      clka_en : OUT STD_LOGIC;
      qb : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      web : OUT STD_LOGIC;
      db : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adrb : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      clka : IN STD_LOGIC;
      clka_en_d : IN STD_LOGIC;
      clkb_en_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      wea_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC_VECTOR (1 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL yy_rsc_31_0_i_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_db : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_adrb : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_adra : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_adra_d_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_da_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_qa_d_1 : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_wea_d_1 : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 : STD_LOGIC_VECTOR (1 DOWNTO
      0);

  COMPONENT hybrid_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      x_rsc_0_0_s_tdone : IN STD_LOGIC;
      x_rsc_0_0_tr_write_done : IN STD_LOGIC;
      x_rsc_0_0_RREADY : IN STD_LOGIC;
      x_rsc_0_0_RVALID : OUT STD_LOGIC;
      x_rsc_0_0_RUSER : OUT STD_LOGIC;
      x_rsc_0_0_RLAST : OUT STD_LOGIC;
      x_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_RID : OUT STD_LOGIC;
      x_rsc_0_0_ARREADY : OUT STD_LOGIC;
      x_rsc_0_0_ARVALID : IN STD_LOGIC;
      x_rsc_0_0_ARUSER : IN STD_LOGIC;
      x_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_ARLOCK : IN STD_LOGIC;
      x_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_0_0_ARID : IN STD_LOGIC;
      x_rsc_0_0_BREADY : IN STD_LOGIC;
      x_rsc_0_0_BVALID : OUT STD_LOGIC;
      x_rsc_0_0_BUSER : OUT STD_LOGIC;
      x_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_BID : OUT STD_LOGIC;
      x_rsc_0_0_WREADY : OUT STD_LOGIC;
      x_rsc_0_0_WVALID : IN STD_LOGIC;
      x_rsc_0_0_WUSER : IN STD_LOGIC;
      x_rsc_0_0_WLAST : IN STD_LOGIC;
      x_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_0_0_AWREADY : OUT STD_LOGIC;
      x_rsc_0_0_AWVALID : IN STD_LOGIC;
      x_rsc_0_0_AWUSER : IN STD_LOGIC;
      x_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_0_0_AWLOCK : IN STD_LOGIC;
      x_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_0_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      x_rsc_1_0_s_tdone : IN STD_LOGIC;
      x_rsc_1_0_tr_write_done : IN STD_LOGIC;
      x_rsc_1_0_RREADY : IN STD_LOGIC;
      x_rsc_1_0_RVALID : OUT STD_LOGIC;
      x_rsc_1_0_RUSER : OUT STD_LOGIC;
      x_rsc_1_0_RLAST : OUT STD_LOGIC;
      x_rsc_1_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_RID : OUT STD_LOGIC;
      x_rsc_1_0_ARREADY : OUT STD_LOGIC;
      x_rsc_1_0_ARVALID : IN STD_LOGIC;
      x_rsc_1_0_ARUSER : IN STD_LOGIC;
      x_rsc_1_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_ARLOCK : IN STD_LOGIC;
      x_rsc_1_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_1_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_1_0_ARID : IN STD_LOGIC;
      x_rsc_1_0_BREADY : IN STD_LOGIC;
      x_rsc_1_0_BVALID : OUT STD_LOGIC;
      x_rsc_1_0_BUSER : OUT STD_LOGIC;
      x_rsc_1_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_BID : OUT STD_LOGIC;
      x_rsc_1_0_WREADY : OUT STD_LOGIC;
      x_rsc_1_0_WVALID : IN STD_LOGIC;
      x_rsc_1_0_WUSER : IN STD_LOGIC;
      x_rsc_1_0_WLAST : IN STD_LOGIC;
      x_rsc_1_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_1_0_AWREADY : OUT STD_LOGIC;
      x_rsc_1_0_AWVALID : IN STD_LOGIC;
      x_rsc_1_0_AWUSER : IN STD_LOGIC;
      x_rsc_1_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_1_0_AWLOCK : IN STD_LOGIC;
      x_rsc_1_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_1_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_1_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_1_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_1_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      x_rsc_2_0_s_tdone : IN STD_LOGIC;
      x_rsc_2_0_tr_write_done : IN STD_LOGIC;
      x_rsc_2_0_RREADY : IN STD_LOGIC;
      x_rsc_2_0_RVALID : OUT STD_LOGIC;
      x_rsc_2_0_RUSER : OUT STD_LOGIC;
      x_rsc_2_0_RLAST : OUT STD_LOGIC;
      x_rsc_2_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_RID : OUT STD_LOGIC;
      x_rsc_2_0_ARREADY : OUT STD_LOGIC;
      x_rsc_2_0_ARVALID : IN STD_LOGIC;
      x_rsc_2_0_ARUSER : IN STD_LOGIC;
      x_rsc_2_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_ARLOCK : IN STD_LOGIC;
      x_rsc_2_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_2_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_2_0_ARID : IN STD_LOGIC;
      x_rsc_2_0_BREADY : IN STD_LOGIC;
      x_rsc_2_0_BVALID : OUT STD_LOGIC;
      x_rsc_2_0_BUSER : OUT STD_LOGIC;
      x_rsc_2_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_BID : OUT STD_LOGIC;
      x_rsc_2_0_WREADY : OUT STD_LOGIC;
      x_rsc_2_0_WVALID : IN STD_LOGIC;
      x_rsc_2_0_WUSER : IN STD_LOGIC;
      x_rsc_2_0_WLAST : IN STD_LOGIC;
      x_rsc_2_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_2_0_AWREADY : OUT STD_LOGIC;
      x_rsc_2_0_AWVALID : IN STD_LOGIC;
      x_rsc_2_0_AWUSER : IN STD_LOGIC;
      x_rsc_2_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_2_0_AWLOCK : IN STD_LOGIC;
      x_rsc_2_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_2_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_2_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_2_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_2_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_2_0_lz : OUT STD_LOGIC;
      x_rsc_3_0_s_tdone : IN STD_LOGIC;
      x_rsc_3_0_tr_write_done : IN STD_LOGIC;
      x_rsc_3_0_RREADY : IN STD_LOGIC;
      x_rsc_3_0_RVALID : OUT STD_LOGIC;
      x_rsc_3_0_RUSER : OUT STD_LOGIC;
      x_rsc_3_0_RLAST : OUT STD_LOGIC;
      x_rsc_3_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_RID : OUT STD_LOGIC;
      x_rsc_3_0_ARREADY : OUT STD_LOGIC;
      x_rsc_3_0_ARVALID : IN STD_LOGIC;
      x_rsc_3_0_ARUSER : IN STD_LOGIC;
      x_rsc_3_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_ARLOCK : IN STD_LOGIC;
      x_rsc_3_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_3_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_3_0_ARID : IN STD_LOGIC;
      x_rsc_3_0_BREADY : IN STD_LOGIC;
      x_rsc_3_0_BVALID : OUT STD_LOGIC;
      x_rsc_3_0_BUSER : OUT STD_LOGIC;
      x_rsc_3_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_BID : OUT STD_LOGIC;
      x_rsc_3_0_WREADY : OUT STD_LOGIC;
      x_rsc_3_0_WVALID : IN STD_LOGIC;
      x_rsc_3_0_WUSER : IN STD_LOGIC;
      x_rsc_3_0_WLAST : IN STD_LOGIC;
      x_rsc_3_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_3_0_AWREADY : OUT STD_LOGIC;
      x_rsc_3_0_AWVALID : IN STD_LOGIC;
      x_rsc_3_0_AWUSER : IN STD_LOGIC;
      x_rsc_3_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_3_0_AWLOCK : IN STD_LOGIC;
      x_rsc_3_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_3_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_3_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_3_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_3_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_3_0_lz : OUT STD_LOGIC;
      x_rsc_4_0_s_tdone : IN STD_LOGIC;
      x_rsc_4_0_tr_write_done : IN STD_LOGIC;
      x_rsc_4_0_RREADY : IN STD_LOGIC;
      x_rsc_4_0_RVALID : OUT STD_LOGIC;
      x_rsc_4_0_RUSER : OUT STD_LOGIC;
      x_rsc_4_0_RLAST : OUT STD_LOGIC;
      x_rsc_4_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_RID : OUT STD_LOGIC;
      x_rsc_4_0_ARREADY : OUT STD_LOGIC;
      x_rsc_4_0_ARVALID : IN STD_LOGIC;
      x_rsc_4_0_ARUSER : IN STD_LOGIC;
      x_rsc_4_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_ARLOCK : IN STD_LOGIC;
      x_rsc_4_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_4_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_4_0_ARID : IN STD_LOGIC;
      x_rsc_4_0_BREADY : IN STD_LOGIC;
      x_rsc_4_0_BVALID : OUT STD_LOGIC;
      x_rsc_4_0_BUSER : OUT STD_LOGIC;
      x_rsc_4_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_BID : OUT STD_LOGIC;
      x_rsc_4_0_WREADY : OUT STD_LOGIC;
      x_rsc_4_0_WVALID : IN STD_LOGIC;
      x_rsc_4_0_WUSER : IN STD_LOGIC;
      x_rsc_4_0_WLAST : IN STD_LOGIC;
      x_rsc_4_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_4_0_AWREADY : OUT STD_LOGIC;
      x_rsc_4_0_AWVALID : IN STD_LOGIC;
      x_rsc_4_0_AWUSER : IN STD_LOGIC;
      x_rsc_4_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_4_0_AWLOCK : IN STD_LOGIC;
      x_rsc_4_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_4_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_4_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_4_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_4_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_4_0_lz : OUT STD_LOGIC;
      x_rsc_5_0_s_tdone : IN STD_LOGIC;
      x_rsc_5_0_tr_write_done : IN STD_LOGIC;
      x_rsc_5_0_RREADY : IN STD_LOGIC;
      x_rsc_5_0_RVALID : OUT STD_LOGIC;
      x_rsc_5_0_RUSER : OUT STD_LOGIC;
      x_rsc_5_0_RLAST : OUT STD_LOGIC;
      x_rsc_5_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_RID : OUT STD_LOGIC;
      x_rsc_5_0_ARREADY : OUT STD_LOGIC;
      x_rsc_5_0_ARVALID : IN STD_LOGIC;
      x_rsc_5_0_ARUSER : IN STD_LOGIC;
      x_rsc_5_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_ARLOCK : IN STD_LOGIC;
      x_rsc_5_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_5_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_5_0_ARID : IN STD_LOGIC;
      x_rsc_5_0_BREADY : IN STD_LOGIC;
      x_rsc_5_0_BVALID : OUT STD_LOGIC;
      x_rsc_5_0_BUSER : OUT STD_LOGIC;
      x_rsc_5_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_BID : OUT STD_LOGIC;
      x_rsc_5_0_WREADY : OUT STD_LOGIC;
      x_rsc_5_0_WVALID : IN STD_LOGIC;
      x_rsc_5_0_WUSER : IN STD_LOGIC;
      x_rsc_5_0_WLAST : IN STD_LOGIC;
      x_rsc_5_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_5_0_AWREADY : OUT STD_LOGIC;
      x_rsc_5_0_AWVALID : IN STD_LOGIC;
      x_rsc_5_0_AWUSER : IN STD_LOGIC;
      x_rsc_5_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_5_0_AWLOCK : IN STD_LOGIC;
      x_rsc_5_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_5_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_5_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_5_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_5_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_5_0_lz : OUT STD_LOGIC;
      x_rsc_6_0_s_tdone : IN STD_LOGIC;
      x_rsc_6_0_tr_write_done : IN STD_LOGIC;
      x_rsc_6_0_RREADY : IN STD_LOGIC;
      x_rsc_6_0_RVALID : OUT STD_LOGIC;
      x_rsc_6_0_RUSER : OUT STD_LOGIC;
      x_rsc_6_0_RLAST : OUT STD_LOGIC;
      x_rsc_6_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_RID : OUT STD_LOGIC;
      x_rsc_6_0_ARREADY : OUT STD_LOGIC;
      x_rsc_6_0_ARVALID : IN STD_LOGIC;
      x_rsc_6_0_ARUSER : IN STD_LOGIC;
      x_rsc_6_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_ARLOCK : IN STD_LOGIC;
      x_rsc_6_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_6_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_6_0_ARID : IN STD_LOGIC;
      x_rsc_6_0_BREADY : IN STD_LOGIC;
      x_rsc_6_0_BVALID : OUT STD_LOGIC;
      x_rsc_6_0_BUSER : OUT STD_LOGIC;
      x_rsc_6_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_BID : OUT STD_LOGIC;
      x_rsc_6_0_WREADY : OUT STD_LOGIC;
      x_rsc_6_0_WVALID : IN STD_LOGIC;
      x_rsc_6_0_WUSER : IN STD_LOGIC;
      x_rsc_6_0_WLAST : IN STD_LOGIC;
      x_rsc_6_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_6_0_AWREADY : OUT STD_LOGIC;
      x_rsc_6_0_AWVALID : IN STD_LOGIC;
      x_rsc_6_0_AWUSER : IN STD_LOGIC;
      x_rsc_6_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_6_0_AWLOCK : IN STD_LOGIC;
      x_rsc_6_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_6_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_6_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_6_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_6_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_6_0_lz : OUT STD_LOGIC;
      x_rsc_7_0_s_tdone : IN STD_LOGIC;
      x_rsc_7_0_tr_write_done : IN STD_LOGIC;
      x_rsc_7_0_RREADY : IN STD_LOGIC;
      x_rsc_7_0_RVALID : OUT STD_LOGIC;
      x_rsc_7_0_RUSER : OUT STD_LOGIC;
      x_rsc_7_0_RLAST : OUT STD_LOGIC;
      x_rsc_7_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_RID : OUT STD_LOGIC;
      x_rsc_7_0_ARREADY : OUT STD_LOGIC;
      x_rsc_7_0_ARVALID : IN STD_LOGIC;
      x_rsc_7_0_ARUSER : IN STD_LOGIC;
      x_rsc_7_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_ARLOCK : IN STD_LOGIC;
      x_rsc_7_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_7_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_7_0_ARID : IN STD_LOGIC;
      x_rsc_7_0_BREADY : IN STD_LOGIC;
      x_rsc_7_0_BVALID : OUT STD_LOGIC;
      x_rsc_7_0_BUSER : OUT STD_LOGIC;
      x_rsc_7_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_BID : OUT STD_LOGIC;
      x_rsc_7_0_WREADY : OUT STD_LOGIC;
      x_rsc_7_0_WVALID : IN STD_LOGIC;
      x_rsc_7_0_WUSER : IN STD_LOGIC;
      x_rsc_7_0_WLAST : IN STD_LOGIC;
      x_rsc_7_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_7_0_AWREADY : OUT STD_LOGIC;
      x_rsc_7_0_AWVALID : IN STD_LOGIC;
      x_rsc_7_0_AWUSER : IN STD_LOGIC;
      x_rsc_7_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_7_0_AWLOCK : IN STD_LOGIC;
      x_rsc_7_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_7_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_7_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_7_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_7_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_7_0_lz : OUT STD_LOGIC;
      x_rsc_8_0_s_tdone : IN STD_LOGIC;
      x_rsc_8_0_tr_write_done : IN STD_LOGIC;
      x_rsc_8_0_RREADY : IN STD_LOGIC;
      x_rsc_8_0_RVALID : OUT STD_LOGIC;
      x_rsc_8_0_RUSER : OUT STD_LOGIC;
      x_rsc_8_0_RLAST : OUT STD_LOGIC;
      x_rsc_8_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_RID : OUT STD_LOGIC;
      x_rsc_8_0_ARREADY : OUT STD_LOGIC;
      x_rsc_8_0_ARVALID : IN STD_LOGIC;
      x_rsc_8_0_ARUSER : IN STD_LOGIC;
      x_rsc_8_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_ARLOCK : IN STD_LOGIC;
      x_rsc_8_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_8_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_8_0_ARID : IN STD_LOGIC;
      x_rsc_8_0_BREADY : IN STD_LOGIC;
      x_rsc_8_0_BVALID : OUT STD_LOGIC;
      x_rsc_8_0_BUSER : OUT STD_LOGIC;
      x_rsc_8_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_BID : OUT STD_LOGIC;
      x_rsc_8_0_WREADY : OUT STD_LOGIC;
      x_rsc_8_0_WVALID : IN STD_LOGIC;
      x_rsc_8_0_WUSER : IN STD_LOGIC;
      x_rsc_8_0_WLAST : IN STD_LOGIC;
      x_rsc_8_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_8_0_AWREADY : OUT STD_LOGIC;
      x_rsc_8_0_AWVALID : IN STD_LOGIC;
      x_rsc_8_0_AWUSER : IN STD_LOGIC;
      x_rsc_8_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_8_0_AWLOCK : IN STD_LOGIC;
      x_rsc_8_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_8_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_8_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_8_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_8_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_8_0_lz : OUT STD_LOGIC;
      x_rsc_9_0_s_tdone : IN STD_LOGIC;
      x_rsc_9_0_tr_write_done : IN STD_LOGIC;
      x_rsc_9_0_RREADY : IN STD_LOGIC;
      x_rsc_9_0_RVALID : OUT STD_LOGIC;
      x_rsc_9_0_RUSER : OUT STD_LOGIC;
      x_rsc_9_0_RLAST : OUT STD_LOGIC;
      x_rsc_9_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_RID : OUT STD_LOGIC;
      x_rsc_9_0_ARREADY : OUT STD_LOGIC;
      x_rsc_9_0_ARVALID : IN STD_LOGIC;
      x_rsc_9_0_ARUSER : IN STD_LOGIC;
      x_rsc_9_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_ARLOCK : IN STD_LOGIC;
      x_rsc_9_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_9_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_9_0_ARID : IN STD_LOGIC;
      x_rsc_9_0_BREADY : IN STD_LOGIC;
      x_rsc_9_0_BVALID : OUT STD_LOGIC;
      x_rsc_9_0_BUSER : OUT STD_LOGIC;
      x_rsc_9_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_BID : OUT STD_LOGIC;
      x_rsc_9_0_WREADY : OUT STD_LOGIC;
      x_rsc_9_0_WVALID : IN STD_LOGIC;
      x_rsc_9_0_WUSER : IN STD_LOGIC;
      x_rsc_9_0_WLAST : IN STD_LOGIC;
      x_rsc_9_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_9_0_AWREADY : OUT STD_LOGIC;
      x_rsc_9_0_AWVALID : IN STD_LOGIC;
      x_rsc_9_0_AWUSER : IN STD_LOGIC;
      x_rsc_9_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_9_0_AWLOCK : IN STD_LOGIC;
      x_rsc_9_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_9_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_9_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_9_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_9_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_9_0_lz : OUT STD_LOGIC;
      x_rsc_10_0_s_tdone : IN STD_LOGIC;
      x_rsc_10_0_tr_write_done : IN STD_LOGIC;
      x_rsc_10_0_RREADY : IN STD_LOGIC;
      x_rsc_10_0_RVALID : OUT STD_LOGIC;
      x_rsc_10_0_RUSER : OUT STD_LOGIC;
      x_rsc_10_0_RLAST : OUT STD_LOGIC;
      x_rsc_10_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_RID : OUT STD_LOGIC;
      x_rsc_10_0_ARREADY : OUT STD_LOGIC;
      x_rsc_10_0_ARVALID : IN STD_LOGIC;
      x_rsc_10_0_ARUSER : IN STD_LOGIC;
      x_rsc_10_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_ARLOCK : IN STD_LOGIC;
      x_rsc_10_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_10_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_10_0_ARID : IN STD_LOGIC;
      x_rsc_10_0_BREADY : IN STD_LOGIC;
      x_rsc_10_0_BVALID : OUT STD_LOGIC;
      x_rsc_10_0_BUSER : OUT STD_LOGIC;
      x_rsc_10_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_BID : OUT STD_LOGIC;
      x_rsc_10_0_WREADY : OUT STD_LOGIC;
      x_rsc_10_0_WVALID : IN STD_LOGIC;
      x_rsc_10_0_WUSER : IN STD_LOGIC;
      x_rsc_10_0_WLAST : IN STD_LOGIC;
      x_rsc_10_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_10_0_AWREADY : OUT STD_LOGIC;
      x_rsc_10_0_AWVALID : IN STD_LOGIC;
      x_rsc_10_0_AWUSER : IN STD_LOGIC;
      x_rsc_10_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_10_0_AWLOCK : IN STD_LOGIC;
      x_rsc_10_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_10_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_10_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_10_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_10_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_10_0_lz : OUT STD_LOGIC;
      x_rsc_11_0_s_tdone : IN STD_LOGIC;
      x_rsc_11_0_tr_write_done : IN STD_LOGIC;
      x_rsc_11_0_RREADY : IN STD_LOGIC;
      x_rsc_11_0_RVALID : OUT STD_LOGIC;
      x_rsc_11_0_RUSER : OUT STD_LOGIC;
      x_rsc_11_0_RLAST : OUT STD_LOGIC;
      x_rsc_11_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_RID : OUT STD_LOGIC;
      x_rsc_11_0_ARREADY : OUT STD_LOGIC;
      x_rsc_11_0_ARVALID : IN STD_LOGIC;
      x_rsc_11_0_ARUSER : IN STD_LOGIC;
      x_rsc_11_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_ARLOCK : IN STD_LOGIC;
      x_rsc_11_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_11_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_11_0_ARID : IN STD_LOGIC;
      x_rsc_11_0_BREADY : IN STD_LOGIC;
      x_rsc_11_0_BVALID : OUT STD_LOGIC;
      x_rsc_11_0_BUSER : OUT STD_LOGIC;
      x_rsc_11_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_BID : OUT STD_LOGIC;
      x_rsc_11_0_WREADY : OUT STD_LOGIC;
      x_rsc_11_0_WVALID : IN STD_LOGIC;
      x_rsc_11_0_WUSER : IN STD_LOGIC;
      x_rsc_11_0_WLAST : IN STD_LOGIC;
      x_rsc_11_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_11_0_AWREADY : OUT STD_LOGIC;
      x_rsc_11_0_AWVALID : IN STD_LOGIC;
      x_rsc_11_0_AWUSER : IN STD_LOGIC;
      x_rsc_11_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_11_0_AWLOCK : IN STD_LOGIC;
      x_rsc_11_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_11_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_11_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_11_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_11_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_11_0_lz : OUT STD_LOGIC;
      x_rsc_12_0_s_tdone : IN STD_LOGIC;
      x_rsc_12_0_tr_write_done : IN STD_LOGIC;
      x_rsc_12_0_RREADY : IN STD_LOGIC;
      x_rsc_12_0_RVALID : OUT STD_LOGIC;
      x_rsc_12_0_RUSER : OUT STD_LOGIC;
      x_rsc_12_0_RLAST : OUT STD_LOGIC;
      x_rsc_12_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_RID : OUT STD_LOGIC;
      x_rsc_12_0_ARREADY : OUT STD_LOGIC;
      x_rsc_12_0_ARVALID : IN STD_LOGIC;
      x_rsc_12_0_ARUSER : IN STD_LOGIC;
      x_rsc_12_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_ARLOCK : IN STD_LOGIC;
      x_rsc_12_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_12_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_12_0_ARID : IN STD_LOGIC;
      x_rsc_12_0_BREADY : IN STD_LOGIC;
      x_rsc_12_0_BVALID : OUT STD_LOGIC;
      x_rsc_12_0_BUSER : OUT STD_LOGIC;
      x_rsc_12_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_BID : OUT STD_LOGIC;
      x_rsc_12_0_WREADY : OUT STD_LOGIC;
      x_rsc_12_0_WVALID : IN STD_LOGIC;
      x_rsc_12_0_WUSER : IN STD_LOGIC;
      x_rsc_12_0_WLAST : IN STD_LOGIC;
      x_rsc_12_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_12_0_AWREADY : OUT STD_LOGIC;
      x_rsc_12_0_AWVALID : IN STD_LOGIC;
      x_rsc_12_0_AWUSER : IN STD_LOGIC;
      x_rsc_12_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_12_0_AWLOCK : IN STD_LOGIC;
      x_rsc_12_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_12_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_12_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_12_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_12_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_12_0_lz : OUT STD_LOGIC;
      x_rsc_13_0_s_tdone : IN STD_LOGIC;
      x_rsc_13_0_tr_write_done : IN STD_LOGIC;
      x_rsc_13_0_RREADY : IN STD_LOGIC;
      x_rsc_13_0_RVALID : OUT STD_LOGIC;
      x_rsc_13_0_RUSER : OUT STD_LOGIC;
      x_rsc_13_0_RLAST : OUT STD_LOGIC;
      x_rsc_13_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_RID : OUT STD_LOGIC;
      x_rsc_13_0_ARREADY : OUT STD_LOGIC;
      x_rsc_13_0_ARVALID : IN STD_LOGIC;
      x_rsc_13_0_ARUSER : IN STD_LOGIC;
      x_rsc_13_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_ARLOCK : IN STD_LOGIC;
      x_rsc_13_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_13_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_13_0_ARID : IN STD_LOGIC;
      x_rsc_13_0_BREADY : IN STD_LOGIC;
      x_rsc_13_0_BVALID : OUT STD_LOGIC;
      x_rsc_13_0_BUSER : OUT STD_LOGIC;
      x_rsc_13_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_BID : OUT STD_LOGIC;
      x_rsc_13_0_WREADY : OUT STD_LOGIC;
      x_rsc_13_0_WVALID : IN STD_LOGIC;
      x_rsc_13_0_WUSER : IN STD_LOGIC;
      x_rsc_13_0_WLAST : IN STD_LOGIC;
      x_rsc_13_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_13_0_AWREADY : OUT STD_LOGIC;
      x_rsc_13_0_AWVALID : IN STD_LOGIC;
      x_rsc_13_0_AWUSER : IN STD_LOGIC;
      x_rsc_13_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_13_0_AWLOCK : IN STD_LOGIC;
      x_rsc_13_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_13_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_13_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_13_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_13_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_13_0_lz : OUT STD_LOGIC;
      x_rsc_14_0_s_tdone : IN STD_LOGIC;
      x_rsc_14_0_tr_write_done : IN STD_LOGIC;
      x_rsc_14_0_RREADY : IN STD_LOGIC;
      x_rsc_14_0_RVALID : OUT STD_LOGIC;
      x_rsc_14_0_RUSER : OUT STD_LOGIC;
      x_rsc_14_0_RLAST : OUT STD_LOGIC;
      x_rsc_14_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_RID : OUT STD_LOGIC;
      x_rsc_14_0_ARREADY : OUT STD_LOGIC;
      x_rsc_14_0_ARVALID : IN STD_LOGIC;
      x_rsc_14_0_ARUSER : IN STD_LOGIC;
      x_rsc_14_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_ARLOCK : IN STD_LOGIC;
      x_rsc_14_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_14_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_14_0_ARID : IN STD_LOGIC;
      x_rsc_14_0_BREADY : IN STD_LOGIC;
      x_rsc_14_0_BVALID : OUT STD_LOGIC;
      x_rsc_14_0_BUSER : OUT STD_LOGIC;
      x_rsc_14_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_BID : OUT STD_LOGIC;
      x_rsc_14_0_WREADY : OUT STD_LOGIC;
      x_rsc_14_0_WVALID : IN STD_LOGIC;
      x_rsc_14_0_WUSER : IN STD_LOGIC;
      x_rsc_14_0_WLAST : IN STD_LOGIC;
      x_rsc_14_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_14_0_AWREADY : OUT STD_LOGIC;
      x_rsc_14_0_AWVALID : IN STD_LOGIC;
      x_rsc_14_0_AWUSER : IN STD_LOGIC;
      x_rsc_14_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_14_0_AWLOCK : IN STD_LOGIC;
      x_rsc_14_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_14_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_14_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_14_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_14_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_14_0_lz : OUT STD_LOGIC;
      x_rsc_15_0_s_tdone : IN STD_LOGIC;
      x_rsc_15_0_tr_write_done : IN STD_LOGIC;
      x_rsc_15_0_RREADY : IN STD_LOGIC;
      x_rsc_15_0_RVALID : OUT STD_LOGIC;
      x_rsc_15_0_RUSER : OUT STD_LOGIC;
      x_rsc_15_0_RLAST : OUT STD_LOGIC;
      x_rsc_15_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_RID : OUT STD_LOGIC;
      x_rsc_15_0_ARREADY : OUT STD_LOGIC;
      x_rsc_15_0_ARVALID : IN STD_LOGIC;
      x_rsc_15_0_ARUSER : IN STD_LOGIC;
      x_rsc_15_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_ARLOCK : IN STD_LOGIC;
      x_rsc_15_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_15_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_15_0_ARID : IN STD_LOGIC;
      x_rsc_15_0_BREADY : IN STD_LOGIC;
      x_rsc_15_0_BVALID : OUT STD_LOGIC;
      x_rsc_15_0_BUSER : OUT STD_LOGIC;
      x_rsc_15_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_BID : OUT STD_LOGIC;
      x_rsc_15_0_WREADY : OUT STD_LOGIC;
      x_rsc_15_0_WVALID : IN STD_LOGIC;
      x_rsc_15_0_WUSER : IN STD_LOGIC;
      x_rsc_15_0_WLAST : IN STD_LOGIC;
      x_rsc_15_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_15_0_AWREADY : OUT STD_LOGIC;
      x_rsc_15_0_AWVALID : IN STD_LOGIC;
      x_rsc_15_0_AWUSER : IN STD_LOGIC;
      x_rsc_15_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_15_0_AWLOCK : IN STD_LOGIC;
      x_rsc_15_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_15_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_15_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_15_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_15_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_15_0_lz : OUT STD_LOGIC;
      x_rsc_16_0_s_tdone : IN STD_LOGIC;
      x_rsc_16_0_tr_write_done : IN STD_LOGIC;
      x_rsc_16_0_RREADY : IN STD_LOGIC;
      x_rsc_16_0_RVALID : OUT STD_LOGIC;
      x_rsc_16_0_RUSER : OUT STD_LOGIC;
      x_rsc_16_0_RLAST : OUT STD_LOGIC;
      x_rsc_16_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_RID : OUT STD_LOGIC;
      x_rsc_16_0_ARREADY : OUT STD_LOGIC;
      x_rsc_16_0_ARVALID : IN STD_LOGIC;
      x_rsc_16_0_ARUSER : IN STD_LOGIC;
      x_rsc_16_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_ARLOCK : IN STD_LOGIC;
      x_rsc_16_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_16_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_16_0_ARID : IN STD_LOGIC;
      x_rsc_16_0_BREADY : IN STD_LOGIC;
      x_rsc_16_0_BVALID : OUT STD_LOGIC;
      x_rsc_16_0_BUSER : OUT STD_LOGIC;
      x_rsc_16_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_BID : OUT STD_LOGIC;
      x_rsc_16_0_WREADY : OUT STD_LOGIC;
      x_rsc_16_0_WVALID : IN STD_LOGIC;
      x_rsc_16_0_WUSER : IN STD_LOGIC;
      x_rsc_16_0_WLAST : IN STD_LOGIC;
      x_rsc_16_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_16_0_AWREADY : OUT STD_LOGIC;
      x_rsc_16_0_AWVALID : IN STD_LOGIC;
      x_rsc_16_0_AWUSER : IN STD_LOGIC;
      x_rsc_16_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_16_0_AWLOCK : IN STD_LOGIC;
      x_rsc_16_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_16_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_16_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_16_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_16_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_16_0_lz : OUT STD_LOGIC;
      x_rsc_17_0_s_tdone : IN STD_LOGIC;
      x_rsc_17_0_tr_write_done : IN STD_LOGIC;
      x_rsc_17_0_RREADY : IN STD_LOGIC;
      x_rsc_17_0_RVALID : OUT STD_LOGIC;
      x_rsc_17_0_RUSER : OUT STD_LOGIC;
      x_rsc_17_0_RLAST : OUT STD_LOGIC;
      x_rsc_17_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_RID : OUT STD_LOGIC;
      x_rsc_17_0_ARREADY : OUT STD_LOGIC;
      x_rsc_17_0_ARVALID : IN STD_LOGIC;
      x_rsc_17_0_ARUSER : IN STD_LOGIC;
      x_rsc_17_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_ARLOCK : IN STD_LOGIC;
      x_rsc_17_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_17_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_17_0_ARID : IN STD_LOGIC;
      x_rsc_17_0_BREADY : IN STD_LOGIC;
      x_rsc_17_0_BVALID : OUT STD_LOGIC;
      x_rsc_17_0_BUSER : OUT STD_LOGIC;
      x_rsc_17_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_BID : OUT STD_LOGIC;
      x_rsc_17_0_WREADY : OUT STD_LOGIC;
      x_rsc_17_0_WVALID : IN STD_LOGIC;
      x_rsc_17_0_WUSER : IN STD_LOGIC;
      x_rsc_17_0_WLAST : IN STD_LOGIC;
      x_rsc_17_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_17_0_AWREADY : OUT STD_LOGIC;
      x_rsc_17_0_AWVALID : IN STD_LOGIC;
      x_rsc_17_0_AWUSER : IN STD_LOGIC;
      x_rsc_17_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_17_0_AWLOCK : IN STD_LOGIC;
      x_rsc_17_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_17_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_17_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_17_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_17_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_17_0_lz : OUT STD_LOGIC;
      x_rsc_18_0_s_tdone : IN STD_LOGIC;
      x_rsc_18_0_tr_write_done : IN STD_LOGIC;
      x_rsc_18_0_RREADY : IN STD_LOGIC;
      x_rsc_18_0_RVALID : OUT STD_LOGIC;
      x_rsc_18_0_RUSER : OUT STD_LOGIC;
      x_rsc_18_0_RLAST : OUT STD_LOGIC;
      x_rsc_18_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_RID : OUT STD_LOGIC;
      x_rsc_18_0_ARREADY : OUT STD_LOGIC;
      x_rsc_18_0_ARVALID : IN STD_LOGIC;
      x_rsc_18_0_ARUSER : IN STD_LOGIC;
      x_rsc_18_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_ARLOCK : IN STD_LOGIC;
      x_rsc_18_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_18_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_18_0_ARID : IN STD_LOGIC;
      x_rsc_18_0_BREADY : IN STD_LOGIC;
      x_rsc_18_0_BVALID : OUT STD_LOGIC;
      x_rsc_18_0_BUSER : OUT STD_LOGIC;
      x_rsc_18_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_BID : OUT STD_LOGIC;
      x_rsc_18_0_WREADY : OUT STD_LOGIC;
      x_rsc_18_0_WVALID : IN STD_LOGIC;
      x_rsc_18_0_WUSER : IN STD_LOGIC;
      x_rsc_18_0_WLAST : IN STD_LOGIC;
      x_rsc_18_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_18_0_AWREADY : OUT STD_LOGIC;
      x_rsc_18_0_AWVALID : IN STD_LOGIC;
      x_rsc_18_0_AWUSER : IN STD_LOGIC;
      x_rsc_18_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_18_0_AWLOCK : IN STD_LOGIC;
      x_rsc_18_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_18_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_18_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_18_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_18_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_18_0_lz : OUT STD_LOGIC;
      x_rsc_19_0_s_tdone : IN STD_LOGIC;
      x_rsc_19_0_tr_write_done : IN STD_LOGIC;
      x_rsc_19_0_RREADY : IN STD_LOGIC;
      x_rsc_19_0_RVALID : OUT STD_LOGIC;
      x_rsc_19_0_RUSER : OUT STD_LOGIC;
      x_rsc_19_0_RLAST : OUT STD_LOGIC;
      x_rsc_19_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_RID : OUT STD_LOGIC;
      x_rsc_19_0_ARREADY : OUT STD_LOGIC;
      x_rsc_19_0_ARVALID : IN STD_LOGIC;
      x_rsc_19_0_ARUSER : IN STD_LOGIC;
      x_rsc_19_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_ARLOCK : IN STD_LOGIC;
      x_rsc_19_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_19_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_19_0_ARID : IN STD_LOGIC;
      x_rsc_19_0_BREADY : IN STD_LOGIC;
      x_rsc_19_0_BVALID : OUT STD_LOGIC;
      x_rsc_19_0_BUSER : OUT STD_LOGIC;
      x_rsc_19_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_BID : OUT STD_LOGIC;
      x_rsc_19_0_WREADY : OUT STD_LOGIC;
      x_rsc_19_0_WVALID : IN STD_LOGIC;
      x_rsc_19_0_WUSER : IN STD_LOGIC;
      x_rsc_19_0_WLAST : IN STD_LOGIC;
      x_rsc_19_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_19_0_AWREADY : OUT STD_LOGIC;
      x_rsc_19_0_AWVALID : IN STD_LOGIC;
      x_rsc_19_0_AWUSER : IN STD_LOGIC;
      x_rsc_19_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_19_0_AWLOCK : IN STD_LOGIC;
      x_rsc_19_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_19_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_19_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_19_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_19_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_19_0_lz : OUT STD_LOGIC;
      x_rsc_20_0_s_tdone : IN STD_LOGIC;
      x_rsc_20_0_tr_write_done : IN STD_LOGIC;
      x_rsc_20_0_RREADY : IN STD_LOGIC;
      x_rsc_20_0_RVALID : OUT STD_LOGIC;
      x_rsc_20_0_RUSER : OUT STD_LOGIC;
      x_rsc_20_0_RLAST : OUT STD_LOGIC;
      x_rsc_20_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_RID : OUT STD_LOGIC;
      x_rsc_20_0_ARREADY : OUT STD_LOGIC;
      x_rsc_20_0_ARVALID : IN STD_LOGIC;
      x_rsc_20_0_ARUSER : IN STD_LOGIC;
      x_rsc_20_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_ARLOCK : IN STD_LOGIC;
      x_rsc_20_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_20_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_20_0_ARID : IN STD_LOGIC;
      x_rsc_20_0_BREADY : IN STD_LOGIC;
      x_rsc_20_0_BVALID : OUT STD_LOGIC;
      x_rsc_20_0_BUSER : OUT STD_LOGIC;
      x_rsc_20_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_BID : OUT STD_LOGIC;
      x_rsc_20_0_WREADY : OUT STD_LOGIC;
      x_rsc_20_0_WVALID : IN STD_LOGIC;
      x_rsc_20_0_WUSER : IN STD_LOGIC;
      x_rsc_20_0_WLAST : IN STD_LOGIC;
      x_rsc_20_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_20_0_AWREADY : OUT STD_LOGIC;
      x_rsc_20_0_AWVALID : IN STD_LOGIC;
      x_rsc_20_0_AWUSER : IN STD_LOGIC;
      x_rsc_20_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_20_0_AWLOCK : IN STD_LOGIC;
      x_rsc_20_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_20_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_20_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_20_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_20_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_20_0_lz : OUT STD_LOGIC;
      x_rsc_21_0_s_tdone : IN STD_LOGIC;
      x_rsc_21_0_tr_write_done : IN STD_LOGIC;
      x_rsc_21_0_RREADY : IN STD_LOGIC;
      x_rsc_21_0_RVALID : OUT STD_LOGIC;
      x_rsc_21_0_RUSER : OUT STD_LOGIC;
      x_rsc_21_0_RLAST : OUT STD_LOGIC;
      x_rsc_21_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_RID : OUT STD_LOGIC;
      x_rsc_21_0_ARREADY : OUT STD_LOGIC;
      x_rsc_21_0_ARVALID : IN STD_LOGIC;
      x_rsc_21_0_ARUSER : IN STD_LOGIC;
      x_rsc_21_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_ARLOCK : IN STD_LOGIC;
      x_rsc_21_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_21_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_21_0_ARID : IN STD_LOGIC;
      x_rsc_21_0_BREADY : IN STD_LOGIC;
      x_rsc_21_0_BVALID : OUT STD_LOGIC;
      x_rsc_21_0_BUSER : OUT STD_LOGIC;
      x_rsc_21_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_BID : OUT STD_LOGIC;
      x_rsc_21_0_WREADY : OUT STD_LOGIC;
      x_rsc_21_0_WVALID : IN STD_LOGIC;
      x_rsc_21_0_WUSER : IN STD_LOGIC;
      x_rsc_21_0_WLAST : IN STD_LOGIC;
      x_rsc_21_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_21_0_AWREADY : OUT STD_LOGIC;
      x_rsc_21_0_AWVALID : IN STD_LOGIC;
      x_rsc_21_0_AWUSER : IN STD_LOGIC;
      x_rsc_21_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_21_0_AWLOCK : IN STD_LOGIC;
      x_rsc_21_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_21_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_21_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_21_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_21_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_21_0_lz : OUT STD_LOGIC;
      x_rsc_22_0_s_tdone : IN STD_LOGIC;
      x_rsc_22_0_tr_write_done : IN STD_LOGIC;
      x_rsc_22_0_RREADY : IN STD_LOGIC;
      x_rsc_22_0_RVALID : OUT STD_LOGIC;
      x_rsc_22_0_RUSER : OUT STD_LOGIC;
      x_rsc_22_0_RLAST : OUT STD_LOGIC;
      x_rsc_22_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_RID : OUT STD_LOGIC;
      x_rsc_22_0_ARREADY : OUT STD_LOGIC;
      x_rsc_22_0_ARVALID : IN STD_LOGIC;
      x_rsc_22_0_ARUSER : IN STD_LOGIC;
      x_rsc_22_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_ARLOCK : IN STD_LOGIC;
      x_rsc_22_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_22_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_22_0_ARID : IN STD_LOGIC;
      x_rsc_22_0_BREADY : IN STD_LOGIC;
      x_rsc_22_0_BVALID : OUT STD_LOGIC;
      x_rsc_22_0_BUSER : OUT STD_LOGIC;
      x_rsc_22_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_BID : OUT STD_LOGIC;
      x_rsc_22_0_WREADY : OUT STD_LOGIC;
      x_rsc_22_0_WVALID : IN STD_LOGIC;
      x_rsc_22_0_WUSER : IN STD_LOGIC;
      x_rsc_22_0_WLAST : IN STD_LOGIC;
      x_rsc_22_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_22_0_AWREADY : OUT STD_LOGIC;
      x_rsc_22_0_AWVALID : IN STD_LOGIC;
      x_rsc_22_0_AWUSER : IN STD_LOGIC;
      x_rsc_22_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_22_0_AWLOCK : IN STD_LOGIC;
      x_rsc_22_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_22_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_22_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_22_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_22_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_22_0_lz : OUT STD_LOGIC;
      x_rsc_23_0_s_tdone : IN STD_LOGIC;
      x_rsc_23_0_tr_write_done : IN STD_LOGIC;
      x_rsc_23_0_RREADY : IN STD_LOGIC;
      x_rsc_23_0_RVALID : OUT STD_LOGIC;
      x_rsc_23_0_RUSER : OUT STD_LOGIC;
      x_rsc_23_0_RLAST : OUT STD_LOGIC;
      x_rsc_23_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_RID : OUT STD_LOGIC;
      x_rsc_23_0_ARREADY : OUT STD_LOGIC;
      x_rsc_23_0_ARVALID : IN STD_LOGIC;
      x_rsc_23_0_ARUSER : IN STD_LOGIC;
      x_rsc_23_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_ARLOCK : IN STD_LOGIC;
      x_rsc_23_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_23_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_23_0_ARID : IN STD_LOGIC;
      x_rsc_23_0_BREADY : IN STD_LOGIC;
      x_rsc_23_0_BVALID : OUT STD_LOGIC;
      x_rsc_23_0_BUSER : OUT STD_LOGIC;
      x_rsc_23_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_BID : OUT STD_LOGIC;
      x_rsc_23_0_WREADY : OUT STD_LOGIC;
      x_rsc_23_0_WVALID : IN STD_LOGIC;
      x_rsc_23_0_WUSER : IN STD_LOGIC;
      x_rsc_23_0_WLAST : IN STD_LOGIC;
      x_rsc_23_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_23_0_AWREADY : OUT STD_LOGIC;
      x_rsc_23_0_AWVALID : IN STD_LOGIC;
      x_rsc_23_0_AWUSER : IN STD_LOGIC;
      x_rsc_23_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_23_0_AWLOCK : IN STD_LOGIC;
      x_rsc_23_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_23_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_23_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_23_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_23_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_23_0_lz : OUT STD_LOGIC;
      x_rsc_24_0_s_tdone : IN STD_LOGIC;
      x_rsc_24_0_tr_write_done : IN STD_LOGIC;
      x_rsc_24_0_RREADY : IN STD_LOGIC;
      x_rsc_24_0_RVALID : OUT STD_LOGIC;
      x_rsc_24_0_RUSER : OUT STD_LOGIC;
      x_rsc_24_0_RLAST : OUT STD_LOGIC;
      x_rsc_24_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_RID : OUT STD_LOGIC;
      x_rsc_24_0_ARREADY : OUT STD_LOGIC;
      x_rsc_24_0_ARVALID : IN STD_LOGIC;
      x_rsc_24_0_ARUSER : IN STD_LOGIC;
      x_rsc_24_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_ARLOCK : IN STD_LOGIC;
      x_rsc_24_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_24_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_24_0_ARID : IN STD_LOGIC;
      x_rsc_24_0_BREADY : IN STD_LOGIC;
      x_rsc_24_0_BVALID : OUT STD_LOGIC;
      x_rsc_24_0_BUSER : OUT STD_LOGIC;
      x_rsc_24_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_BID : OUT STD_LOGIC;
      x_rsc_24_0_WREADY : OUT STD_LOGIC;
      x_rsc_24_0_WVALID : IN STD_LOGIC;
      x_rsc_24_0_WUSER : IN STD_LOGIC;
      x_rsc_24_0_WLAST : IN STD_LOGIC;
      x_rsc_24_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_24_0_AWREADY : OUT STD_LOGIC;
      x_rsc_24_0_AWVALID : IN STD_LOGIC;
      x_rsc_24_0_AWUSER : IN STD_LOGIC;
      x_rsc_24_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_24_0_AWLOCK : IN STD_LOGIC;
      x_rsc_24_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_24_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_24_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_24_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_24_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_24_0_lz : OUT STD_LOGIC;
      x_rsc_25_0_s_tdone : IN STD_LOGIC;
      x_rsc_25_0_tr_write_done : IN STD_LOGIC;
      x_rsc_25_0_RREADY : IN STD_LOGIC;
      x_rsc_25_0_RVALID : OUT STD_LOGIC;
      x_rsc_25_0_RUSER : OUT STD_LOGIC;
      x_rsc_25_0_RLAST : OUT STD_LOGIC;
      x_rsc_25_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_RID : OUT STD_LOGIC;
      x_rsc_25_0_ARREADY : OUT STD_LOGIC;
      x_rsc_25_0_ARVALID : IN STD_LOGIC;
      x_rsc_25_0_ARUSER : IN STD_LOGIC;
      x_rsc_25_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_ARLOCK : IN STD_LOGIC;
      x_rsc_25_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_25_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_25_0_ARID : IN STD_LOGIC;
      x_rsc_25_0_BREADY : IN STD_LOGIC;
      x_rsc_25_0_BVALID : OUT STD_LOGIC;
      x_rsc_25_0_BUSER : OUT STD_LOGIC;
      x_rsc_25_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_BID : OUT STD_LOGIC;
      x_rsc_25_0_WREADY : OUT STD_LOGIC;
      x_rsc_25_0_WVALID : IN STD_LOGIC;
      x_rsc_25_0_WUSER : IN STD_LOGIC;
      x_rsc_25_0_WLAST : IN STD_LOGIC;
      x_rsc_25_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_25_0_AWREADY : OUT STD_LOGIC;
      x_rsc_25_0_AWVALID : IN STD_LOGIC;
      x_rsc_25_0_AWUSER : IN STD_LOGIC;
      x_rsc_25_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_25_0_AWLOCK : IN STD_LOGIC;
      x_rsc_25_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_25_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_25_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_25_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_25_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_25_0_lz : OUT STD_LOGIC;
      x_rsc_26_0_s_tdone : IN STD_LOGIC;
      x_rsc_26_0_tr_write_done : IN STD_LOGIC;
      x_rsc_26_0_RREADY : IN STD_LOGIC;
      x_rsc_26_0_RVALID : OUT STD_LOGIC;
      x_rsc_26_0_RUSER : OUT STD_LOGIC;
      x_rsc_26_0_RLAST : OUT STD_LOGIC;
      x_rsc_26_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_RID : OUT STD_LOGIC;
      x_rsc_26_0_ARREADY : OUT STD_LOGIC;
      x_rsc_26_0_ARVALID : IN STD_LOGIC;
      x_rsc_26_0_ARUSER : IN STD_LOGIC;
      x_rsc_26_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_ARLOCK : IN STD_LOGIC;
      x_rsc_26_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_26_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_26_0_ARID : IN STD_LOGIC;
      x_rsc_26_0_BREADY : IN STD_LOGIC;
      x_rsc_26_0_BVALID : OUT STD_LOGIC;
      x_rsc_26_0_BUSER : OUT STD_LOGIC;
      x_rsc_26_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_BID : OUT STD_LOGIC;
      x_rsc_26_0_WREADY : OUT STD_LOGIC;
      x_rsc_26_0_WVALID : IN STD_LOGIC;
      x_rsc_26_0_WUSER : IN STD_LOGIC;
      x_rsc_26_0_WLAST : IN STD_LOGIC;
      x_rsc_26_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_26_0_AWREADY : OUT STD_LOGIC;
      x_rsc_26_0_AWVALID : IN STD_LOGIC;
      x_rsc_26_0_AWUSER : IN STD_LOGIC;
      x_rsc_26_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_26_0_AWLOCK : IN STD_LOGIC;
      x_rsc_26_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_26_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_26_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_26_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_26_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_26_0_lz : OUT STD_LOGIC;
      x_rsc_27_0_s_tdone : IN STD_LOGIC;
      x_rsc_27_0_tr_write_done : IN STD_LOGIC;
      x_rsc_27_0_RREADY : IN STD_LOGIC;
      x_rsc_27_0_RVALID : OUT STD_LOGIC;
      x_rsc_27_0_RUSER : OUT STD_LOGIC;
      x_rsc_27_0_RLAST : OUT STD_LOGIC;
      x_rsc_27_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_RID : OUT STD_LOGIC;
      x_rsc_27_0_ARREADY : OUT STD_LOGIC;
      x_rsc_27_0_ARVALID : IN STD_LOGIC;
      x_rsc_27_0_ARUSER : IN STD_LOGIC;
      x_rsc_27_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_ARLOCK : IN STD_LOGIC;
      x_rsc_27_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_27_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_27_0_ARID : IN STD_LOGIC;
      x_rsc_27_0_BREADY : IN STD_LOGIC;
      x_rsc_27_0_BVALID : OUT STD_LOGIC;
      x_rsc_27_0_BUSER : OUT STD_LOGIC;
      x_rsc_27_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_BID : OUT STD_LOGIC;
      x_rsc_27_0_WREADY : OUT STD_LOGIC;
      x_rsc_27_0_WVALID : IN STD_LOGIC;
      x_rsc_27_0_WUSER : IN STD_LOGIC;
      x_rsc_27_0_WLAST : IN STD_LOGIC;
      x_rsc_27_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_27_0_AWREADY : OUT STD_LOGIC;
      x_rsc_27_0_AWVALID : IN STD_LOGIC;
      x_rsc_27_0_AWUSER : IN STD_LOGIC;
      x_rsc_27_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_27_0_AWLOCK : IN STD_LOGIC;
      x_rsc_27_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_27_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_27_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_27_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_27_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_27_0_lz : OUT STD_LOGIC;
      x_rsc_28_0_s_tdone : IN STD_LOGIC;
      x_rsc_28_0_tr_write_done : IN STD_LOGIC;
      x_rsc_28_0_RREADY : IN STD_LOGIC;
      x_rsc_28_0_RVALID : OUT STD_LOGIC;
      x_rsc_28_0_RUSER : OUT STD_LOGIC;
      x_rsc_28_0_RLAST : OUT STD_LOGIC;
      x_rsc_28_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_RID : OUT STD_LOGIC;
      x_rsc_28_0_ARREADY : OUT STD_LOGIC;
      x_rsc_28_0_ARVALID : IN STD_LOGIC;
      x_rsc_28_0_ARUSER : IN STD_LOGIC;
      x_rsc_28_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_ARLOCK : IN STD_LOGIC;
      x_rsc_28_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_28_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_28_0_ARID : IN STD_LOGIC;
      x_rsc_28_0_BREADY : IN STD_LOGIC;
      x_rsc_28_0_BVALID : OUT STD_LOGIC;
      x_rsc_28_0_BUSER : OUT STD_LOGIC;
      x_rsc_28_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_BID : OUT STD_LOGIC;
      x_rsc_28_0_WREADY : OUT STD_LOGIC;
      x_rsc_28_0_WVALID : IN STD_LOGIC;
      x_rsc_28_0_WUSER : IN STD_LOGIC;
      x_rsc_28_0_WLAST : IN STD_LOGIC;
      x_rsc_28_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_28_0_AWREADY : OUT STD_LOGIC;
      x_rsc_28_0_AWVALID : IN STD_LOGIC;
      x_rsc_28_0_AWUSER : IN STD_LOGIC;
      x_rsc_28_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_28_0_AWLOCK : IN STD_LOGIC;
      x_rsc_28_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_28_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_28_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_28_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_28_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_28_0_lz : OUT STD_LOGIC;
      x_rsc_29_0_s_tdone : IN STD_LOGIC;
      x_rsc_29_0_tr_write_done : IN STD_LOGIC;
      x_rsc_29_0_RREADY : IN STD_LOGIC;
      x_rsc_29_0_RVALID : OUT STD_LOGIC;
      x_rsc_29_0_RUSER : OUT STD_LOGIC;
      x_rsc_29_0_RLAST : OUT STD_LOGIC;
      x_rsc_29_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_RID : OUT STD_LOGIC;
      x_rsc_29_0_ARREADY : OUT STD_LOGIC;
      x_rsc_29_0_ARVALID : IN STD_LOGIC;
      x_rsc_29_0_ARUSER : IN STD_LOGIC;
      x_rsc_29_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_ARLOCK : IN STD_LOGIC;
      x_rsc_29_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_29_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_29_0_ARID : IN STD_LOGIC;
      x_rsc_29_0_BREADY : IN STD_LOGIC;
      x_rsc_29_0_BVALID : OUT STD_LOGIC;
      x_rsc_29_0_BUSER : OUT STD_LOGIC;
      x_rsc_29_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_BID : OUT STD_LOGIC;
      x_rsc_29_0_WREADY : OUT STD_LOGIC;
      x_rsc_29_0_WVALID : IN STD_LOGIC;
      x_rsc_29_0_WUSER : IN STD_LOGIC;
      x_rsc_29_0_WLAST : IN STD_LOGIC;
      x_rsc_29_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_29_0_AWREADY : OUT STD_LOGIC;
      x_rsc_29_0_AWVALID : IN STD_LOGIC;
      x_rsc_29_0_AWUSER : IN STD_LOGIC;
      x_rsc_29_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_29_0_AWLOCK : IN STD_LOGIC;
      x_rsc_29_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_29_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_29_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_29_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_29_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_29_0_lz : OUT STD_LOGIC;
      x_rsc_30_0_s_tdone : IN STD_LOGIC;
      x_rsc_30_0_tr_write_done : IN STD_LOGIC;
      x_rsc_30_0_RREADY : IN STD_LOGIC;
      x_rsc_30_0_RVALID : OUT STD_LOGIC;
      x_rsc_30_0_RUSER : OUT STD_LOGIC;
      x_rsc_30_0_RLAST : OUT STD_LOGIC;
      x_rsc_30_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_RID : OUT STD_LOGIC;
      x_rsc_30_0_ARREADY : OUT STD_LOGIC;
      x_rsc_30_0_ARVALID : IN STD_LOGIC;
      x_rsc_30_0_ARUSER : IN STD_LOGIC;
      x_rsc_30_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_ARLOCK : IN STD_LOGIC;
      x_rsc_30_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_30_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_30_0_ARID : IN STD_LOGIC;
      x_rsc_30_0_BREADY : IN STD_LOGIC;
      x_rsc_30_0_BVALID : OUT STD_LOGIC;
      x_rsc_30_0_BUSER : OUT STD_LOGIC;
      x_rsc_30_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_BID : OUT STD_LOGIC;
      x_rsc_30_0_WREADY : OUT STD_LOGIC;
      x_rsc_30_0_WVALID : IN STD_LOGIC;
      x_rsc_30_0_WUSER : IN STD_LOGIC;
      x_rsc_30_0_WLAST : IN STD_LOGIC;
      x_rsc_30_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_30_0_AWREADY : OUT STD_LOGIC;
      x_rsc_30_0_AWVALID : IN STD_LOGIC;
      x_rsc_30_0_AWUSER : IN STD_LOGIC;
      x_rsc_30_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_30_0_AWLOCK : IN STD_LOGIC;
      x_rsc_30_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_30_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_30_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_30_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_30_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_30_0_lz : OUT STD_LOGIC;
      x_rsc_31_0_s_tdone : IN STD_LOGIC;
      x_rsc_31_0_tr_write_done : IN STD_LOGIC;
      x_rsc_31_0_RREADY : IN STD_LOGIC;
      x_rsc_31_0_RVALID : OUT STD_LOGIC;
      x_rsc_31_0_RUSER : OUT STD_LOGIC;
      x_rsc_31_0_RLAST : OUT STD_LOGIC;
      x_rsc_31_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_RID : OUT STD_LOGIC;
      x_rsc_31_0_ARREADY : OUT STD_LOGIC;
      x_rsc_31_0_ARVALID : IN STD_LOGIC;
      x_rsc_31_0_ARUSER : IN STD_LOGIC;
      x_rsc_31_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_ARLOCK : IN STD_LOGIC;
      x_rsc_31_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_31_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_31_0_ARID : IN STD_LOGIC;
      x_rsc_31_0_BREADY : IN STD_LOGIC;
      x_rsc_31_0_BVALID : OUT STD_LOGIC;
      x_rsc_31_0_BUSER : OUT STD_LOGIC;
      x_rsc_31_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_BID : OUT STD_LOGIC;
      x_rsc_31_0_WREADY : OUT STD_LOGIC;
      x_rsc_31_0_WVALID : IN STD_LOGIC;
      x_rsc_31_0_WUSER : IN STD_LOGIC;
      x_rsc_31_0_WLAST : IN STD_LOGIC;
      x_rsc_31_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      x_rsc_31_0_AWREADY : OUT STD_LOGIC;
      x_rsc_31_0_AWVALID : IN STD_LOGIC;
      x_rsc_31_0_AWUSER : IN STD_LOGIC;
      x_rsc_31_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      x_rsc_31_0_AWLOCK : IN STD_LOGIC;
      x_rsc_31_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      x_rsc_31_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      x_rsc_31_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      x_rsc_31_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      x_rsc_31_0_AWID : IN STD_LOGIC;
      x_rsc_triosy_31_0_lz : OUT STD_LOGIC;
      m_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      m_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_h_rsc_triosy_lz : OUT STD_LOGIC;
      revArr_rsc_s_tdone : IN STD_LOGIC;
      revArr_rsc_tr_write_done : IN STD_LOGIC;
      revArr_rsc_RREADY : IN STD_LOGIC;
      revArr_rsc_RVALID : OUT STD_LOGIC;
      revArr_rsc_RUSER : OUT STD_LOGIC;
      revArr_rsc_RLAST : OUT STD_LOGIC;
      revArr_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      revArr_rsc_RID : OUT STD_LOGIC;
      revArr_rsc_ARREADY : OUT STD_LOGIC;
      revArr_rsc_ARVALID : IN STD_LOGIC;
      revArr_rsc_ARUSER : IN STD_LOGIC;
      revArr_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_ARLOCK : IN STD_LOGIC;
      revArr_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      revArr_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      revArr_rsc_ARID : IN STD_LOGIC;
      revArr_rsc_BREADY : IN STD_LOGIC;
      revArr_rsc_BVALID : OUT STD_LOGIC;
      revArr_rsc_BUSER : OUT STD_LOGIC;
      revArr_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_BID : OUT STD_LOGIC;
      revArr_rsc_WREADY : OUT STD_LOGIC;
      revArr_rsc_WVALID : IN STD_LOGIC;
      revArr_rsc_WUSER : IN STD_LOGIC;
      revArr_rsc_WLAST : IN STD_LOGIC;
      revArr_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      revArr_rsc_AWREADY : OUT STD_LOGIC;
      revArr_rsc_AWVALID : IN STD_LOGIC;
      revArr_rsc_AWUSER : IN STD_LOGIC;
      revArr_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      revArr_rsc_AWLOCK : IN STD_LOGIC;
      revArr_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      revArr_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      revArr_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      revArr_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      revArr_rsc_AWID : IN STD_LOGIC;
      revArr_rsc_triosy_lz : OUT STD_LOGIC;
      tw_rsc_s_tdone : IN STD_LOGIC;
      tw_rsc_tr_write_done : IN STD_LOGIC;
      tw_rsc_RREADY : IN STD_LOGIC;
      tw_rsc_RVALID : OUT STD_LOGIC;
      tw_rsc_RUSER : OUT STD_LOGIC;
      tw_rsc_RLAST : OUT STD_LOGIC;
      tw_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_rsc_RID : OUT STD_LOGIC;
      tw_rsc_ARREADY : OUT STD_LOGIC;
      tw_rsc_ARVALID : IN STD_LOGIC;
      tw_rsc_ARUSER : IN STD_LOGIC;
      tw_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_ARLOCK : IN STD_LOGIC;
      tw_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_rsc_ARID : IN STD_LOGIC;
      tw_rsc_BREADY : IN STD_LOGIC;
      tw_rsc_BVALID : OUT STD_LOGIC;
      tw_rsc_BUSER : OUT STD_LOGIC;
      tw_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_BID : OUT STD_LOGIC;
      tw_rsc_WREADY : OUT STD_LOGIC;
      tw_rsc_WVALID : IN STD_LOGIC;
      tw_rsc_WUSER : IN STD_LOGIC;
      tw_rsc_WLAST : IN STD_LOGIC;
      tw_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_rsc_AWREADY : OUT STD_LOGIC;
      tw_rsc_AWVALID : IN STD_LOGIC;
      tw_rsc_AWUSER : IN STD_LOGIC;
      tw_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_rsc_AWLOCK : IN STD_LOGIC;
      tw_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_rsc_AWID : IN STD_LOGIC;
      tw_rsc_triosy_lz : OUT STD_LOGIC;
      tw_h_rsc_s_tdone : IN STD_LOGIC;
      tw_h_rsc_tr_write_done : IN STD_LOGIC;
      tw_h_rsc_RREADY : IN STD_LOGIC;
      tw_h_rsc_RVALID : OUT STD_LOGIC;
      tw_h_rsc_RUSER : OUT STD_LOGIC;
      tw_h_rsc_RLAST : OUT STD_LOGIC;
      tw_h_rsc_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_h_rsc_RID : OUT STD_LOGIC;
      tw_h_rsc_ARREADY : OUT STD_LOGIC;
      tw_h_rsc_ARVALID : IN STD_LOGIC;
      tw_h_rsc_ARUSER : IN STD_LOGIC;
      tw_h_rsc_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_ARLOCK : IN STD_LOGIC;
      tw_h_rsc_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_h_rsc_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_h_rsc_ARID : IN STD_LOGIC;
      tw_h_rsc_BREADY : IN STD_LOGIC;
      tw_h_rsc_BVALID : OUT STD_LOGIC;
      tw_h_rsc_BUSER : OUT STD_LOGIC;
      tw_h_rsc_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_BID : OUT STD_LOGIC;
      tw_h_rsc_WREADY : OUT STD_LOGIC;
      tw_h_rsc_WVALID : IN STD_LOGIC;
      tw_h_rsc_WUSER : IN STD_LOGIC;
      tw_h_rsc_WLAST : IN STD_LOGIC;
      tw_h_rsc_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      tw_h_rsc_AWREADY : OUT STD_LOGIC;
      tw_h_rsc_AWVALID : IN STD_LOGIC;
      tw_h_rsc_AWUSER : IN STD_LOGIC;
      tw_h_rsc_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      tw_h_rsc_AWLOCK : IN STD_LOGIC;
      tw_h_rsc_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      tw_h_rsc_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      tw_h_rsc_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      tw_h_rsc_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      tw_h_rsc_AWID : IN STD_LOGIC;
      tw_h_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      twiddle_h_rsci_adrb_d : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      twiddle_h_rsci_qb_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xx_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_1_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_2_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_2_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_2_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_3_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_3_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_3_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_4_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_4_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_4_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_5_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_5_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_5_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_6_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_6_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_6_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_7_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_7_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_7_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_8_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_8_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_8_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_9_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_9_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_9_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_10_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_10_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_10_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_11_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_11_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_11_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_12_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_12_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_12_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_13_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_13_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_13_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_14_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_14_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_14_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_15_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_15_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_15_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_16_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_16_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_16_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_17_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_17_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_17_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_18_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_18_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_18_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_19_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_19_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_19_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_20_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_20_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_20_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_21_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_21_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_21_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_22_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_22_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_22_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_23_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_23_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_23_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_24_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_24_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_24_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_25_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_25_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_25_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_26_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_26_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_26_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_27_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_27_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_27_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_28_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_28_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_28_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_29_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_29_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_29_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_30_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_30_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_30_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_31_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
      xx_rsc_31_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_31_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_0_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_0_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_0_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_1_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_1_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_1_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_2_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_2_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_2_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_2_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_3_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_3_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_3_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_3_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_4_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_4_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_4_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_4_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_5_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_5_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_5_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_5_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_6_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_6_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_6_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_6_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_7_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_7_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_7_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_7_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_8_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_8_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_8_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_8_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_9_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_9_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_9_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_9_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_10_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_10_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_10_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_10_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_11_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_11_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_11_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_11_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_12_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_12_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_12_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_12_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_13_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_13_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_13_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_13_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_14_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_14_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_14_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_14_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_15_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_15_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_15_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_15_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_16_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_16_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_16_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_16_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_17_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_17_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_17_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_17_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_18_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_18_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_18_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_18_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_19_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_19_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_19_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_19_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_20_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_20_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_20_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_20_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_21_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_21_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_21_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_21_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_22_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_22_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_22_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_22_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_23_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_23_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_23_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_23_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_24_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_24_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_24_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_24_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_25_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_25_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_25_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_25_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_26_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_26_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_26_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_26_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_27_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_27_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_27_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_27_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_28_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_28_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_28_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_28_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_29_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_29_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_29_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_29_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_30_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_30_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_30_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_30_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_31_0_i_adra_d : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      yy_rsc_31_0_i_clka_en_d : OUT STD_LOGIC;
      yy_rsc_31_0_i_qa_d : IN STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_31_0_i_wea_d : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : OUT STD_LOGIC_VECTOR (1 DOWNTO
          0);
      S34_OUTER_LOOP_for_tf_mul_cmp_a : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
      S34_OUTER_LOOP_for_tf_mul_cmp_b : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      S34_OUTER_LOOP_for_tf_mul_cmp_z : IN STD_LOGIC_VECTOR (9 DOWNTO 0);
      xx_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_1_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_2_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      xx_rsc_3_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_1_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_2_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0);
      yy_rsc_3_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL hybrid_core_inst_x_rsc_0_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_0_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_1_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_2_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_3_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_4_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_5_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_6_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_7_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_8_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_9_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_10_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_11_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_12_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_13_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_14_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_15_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_16_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_17_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_18_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_19_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_20_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_21_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_22_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_23_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_24_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_25_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_26_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_27_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_28_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_29_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_30_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_x_rsc_31_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_m_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_revArr_rsc_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_rsc_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL hybrid_core_inst_tw_h_rsc_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL hybrid_core_inst_twiddle_rsci_adrb_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_inst_twiddle_rsci_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_twiddle_h_rsci_adrb_d : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL hybrid_core_inst_twiddle_h_rsci_qb_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_2_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_2_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_2_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_3_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_3_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_3_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_4_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_4_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_4_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_5_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_5_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_5_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_6_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_6_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_6_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_7_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_7_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_7_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_8_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_8_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_8_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_9_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_9_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_9_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_10_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_10_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_10_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_11_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_11_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_11_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_12_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_12_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_12_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_13_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_13_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_13_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_14_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_14_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_14_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_15_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_15_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_15_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_16_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_16_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_16_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_17_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_17_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_17_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_18_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_18_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_18_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_19_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_19_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_19_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_20_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_20_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_20_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_21_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_21_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_21_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_22_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_22_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_22_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_23_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_23_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_23_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_24_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_24_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_24_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_25_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_25_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_25_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_26_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_26_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_26_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_27_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_27_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_27_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_28_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_28_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_28_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_29_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_29_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_29_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_30_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_30_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_30_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_31_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_31_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_31_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_0_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_1_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_2_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_2_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_2_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_3_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_3_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_3_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_4_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_4_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_4_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_5_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_5_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_5_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_6_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_6_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_6_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_7_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_7_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_7_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_8_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_8_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_8_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_9_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_9_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_9_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_10_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_10_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_10_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_11_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_11_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_11_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_12_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_12_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_12_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_13_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_13_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_13_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_14_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_14_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_14_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_15_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_15_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_15_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_16_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_16_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_16_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_17_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_17_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_17_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_18_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_18_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_18_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_19_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_19_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_19_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_20_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_20_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_20_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_21_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_21_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_21_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_22_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_22_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_22_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_23_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_23_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_23_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_24_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_24_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_24_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_25_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_25_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_25_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_26_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_26_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_26_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_27_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_27_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_27_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_28_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_28_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_28_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_29_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_29_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_29_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_30_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_30_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_30_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_31_0_i_adra_d : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_31_0_i_qa_d : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_31_0_i_wea_d : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_a : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  SIGNAL hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_b : STD_LOGIC_VECTOR (9 DOWNTO
      0);
  SIGNAL hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z : STD_LOGIC_VECTOR (9 DOWNTO
      0);
  SIGNAL hybrid_core_inst_xx_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_1_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_2_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_xx_rsc_3_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_1_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_2_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);
  SIGNAL hybrid_core_inst_yy_rsc_3_0_i_da_d_pff : STD_LOGIC_VECTOR (63 DOWNTO 0);

BEGIN
  xx_rsc_0_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_0_0_comp_adra,
      adrb => xx_rsc_0_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_0_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_0_0_clkb_en,
      da => xx_rsc_0_0_comp_da,
      db => xx_rsc_0_0_comp_db,
      qa => xx_rsc_0_0_comp_qa,
      qb => xx_rsc_0_0_comp_qb,
      wea => xx_rsc_0_0_wea,
      web => xx_rsc_0_0_web
    );
  xx_rsc_0_0_comp_adra <= xx_rsc_0_0_adra;
  xx_rsc_0_0_comp_adrb <= xx_rsc_0_0_adrb;
  xx_rsc_0_0_comp_da <= xx_rsc_0_0_da;
  xx_rsc_0_0_comp_db <= xx_rsc_0_0_db;
  xx_rsc_0_0_qa <= xx_rsc_0_0_comp_qa;
  xx_rsc_0_0_qb <= xx_rsc_0_0_comp_qb;

  xx_rsc_1_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_1_0_comp_adra,
      adrb => xx_rsc_1_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_1_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_1_0_clkb_en,
      da => xx_rsc_1_0_comp_da,
      db => xx_rsc_1_0_comp_db,
      qa => xx_rsc_1_0_comp_qa,
      qb => xx_rsc_1_0_comp_qb,
      wea => xx_rsc_1_0_wea,
      web => xx_rsc_1_0_web
    );
  xx_rsc_1_0_comp_adra <= xx_rsc_1_0_adra;
  xx_rsc_1_0_comp_adrb <= xx_rsc_1_0_adrb;
  xx_rsc_1_0_comp_da <= xx_rsc_1_0_da;
  xx_rsc_1_0_comp_db <= xx_rsc_1_0_db;
  xx_rsc_1_0_qa <= xx_rsc_1_0_comp_qa;
  xx_rsc_1_0_qb <= xx_rsc_1_0_comp_qb;

  xx_rsc_2_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_2_0_comp_adra,
      adrb => xx_rsc_2_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_2_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_2_0_clkb_en,
      da => xx_rsc_2_0_comp_da,
      db => xx_rsc_2_0_comp_db,
      qa => xx_rsc_2_0_comp_qa,
      qb => xx_rsc_2_0_comp_qb,
      wea => xx_rsc_2_0_wea,
      web => xx_rsc_2_0_web
    );
  xx_rsc_2_0_comp_adra <= xx_rsc_2_0_adra;
  xx_rsc_2_0_comp_adrb <= xx_rsc_2_0_adrb;
  xx_rsc_2_0_comp_da <= xx_rsc_2_0_da;
  xx_rsc_2_0_comp_db <= xx_rsc_2_0_db;
  xx_rsc_2_0_qa <= xx_rsc_2_0_comp_qa;
  xx_rsc_2_0_qb <= xx_rsc_2_0_comp_qb;

  xx_rsc_3_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_3_0_comp_adra,
      adrb => xx_rsc_3_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_3_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_3_0_clkb_en,
      da => xx_rsc_3_0_comp_da,
      db => xx_rsc_3_0_comp_db,
      qa => xx_rsc_3_0_comp_qa,
      qb => xx_rsc_3_0_comp_qb,
      wea => xx_rsc_3_0_wea,
      web => xx_rsc_3_0_web
    );
  xx_rsc_3_0_comp_adra <= xx_rsc_3_0_adra;
  xx_rsc_3_0_comp_adrb <= xx_rsc_3_0_adrb;
  xx_rsc_3_0_comp_da <= xx_rsc_3_0_da;
  xx_rsc_3_0_comp_db <= xx_rsc_3_0_db;
  xx_rsc_3_0_qa <= xx_rsc_3_0_comp_qa;
  xx_rsc_3_0_qb <= xx_rsc_3_0_comp_qb;

  xx_rsc_4_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_4_0_comp_adra,
      adrb => xx_rsc_4_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_4_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_4_0_clkb_en,
      da => xx_rsc_4_0_comp_da,
      db => xx_rsc_4_0_comp_db,
      qa => xx_rsc_4_0_comp_qa,
      qb => xx_rsc_4_0_comp_qb,
      wea => xx_rsc_4_0_wea,
      web => xx_rsc_4_0_web
    );
  xx_rsc_4_0_comp_adra <= xx_rsc_4_0_adra;
  xx_rsc_4_0_comp_adrb <= xx_rsc_4_0_adrb;
  xx_rsc_4_0_comp_da <= xx_rsc_4_0_da;
  xx_rsc_4_0_comp_db <= xx_rsc_4_0_db;
  xx_rsc_4_0_qa <= xx_rsc_4_0_comp_qa;
  xx_rsc_4_0_qb <= xx_rsc_4_0_comp_qb;

  xx_rsc_5_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_5_0_comp_adra,
      adrb => xx_rsc_5_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_5_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_5_0_clkb_en,
      da => xx_rsc_5_0_comp_da,
      db => xx_rsc_5_0_comp_db,
      qa => xx_rsc_5_0_comp_qa,
      qb => xx_rsc_5_0_comp_qb,
      wea => xx_rsc_5_0_wea,
      web => xx_rsc_5_0_web
    );
  xx_rsc_5_0_comp_adra <= xx_rsc_5_0_adra;
  xx_rsc_5_0_comp_adrb <= xx_rsc_5_0_adrb;
  xx_rsc_5_0_comp_da <= xx_rsc_5_0_da;
  xx_rsc_5_0_comp_db <= xx_rsc_5_0_db;
  xx_rsc_5_0_qa <= xx_rsc_5_0_comp_qa;
  xx_rsc_5_0_qb <= xx_rsc_5_0_comp_qb;

  xx_rsc_6_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_6_0_comp_adra,
      adrb => xx_rsc_6_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_6_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_6_0_clkb_en,
      da => xx_rsc_6_0_comp_da,
      db => xx_rsc_6_0_comp_db,
      qa => xx_rsc_6_0_comp_qa,
      qb => xx_rsc_6_0_comp_qb,
      wea => xx_rsc_6_0_wea,
      web => xx_rsc_6_0_web
    );
  xx_rsc_6_0_comp_adra <= xx_rsc_6_0_adra;
  xx_rsc_6_0_comp_adrb <= xx_rsc_6_0_adrb;
  xx_rsc_6_0_comp_da <= xx_rsc_6_0_da;
  xx_rsc_6_0_comp_db <= xx_rsc_6_0_db;
  xx_rsc_6_0_qa <= xx_rsc_6_0_comp_qa;
  xx_rsc_6_0_qb <= xx_rsc_6_0_comp_qb;

  xx_rsc_7_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_7_0_comp_adra,
      adrb => xx_rsc_7_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_7_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_7_0_clkb_en,
      da => xx_rsc_7_0_comp_da,
      db => xx_rsc_7_0_comp_db,
      qa => xx_rsc_7_0_comp_qa,
      qb => xx_rsc_7_0_comp_qb,
      wea => xx_rsc_7_0_wea,
      web => xx_rsc_7_0_web
    );
  xx_rsc_7_0_comp_adra <= xx_rsc_7_0_adra;
  xx_rsc_7_0_comp_adrb <= xx_rsc_7_0_adrb;
  xx_rsc_7_0_comp_da <= xx_rsc_7_0_da;
  xx_rsc_7_0_comp_db <= xx_rsc_7_0_db;
  xx_rsc_7_0_qa <= xx_rsc_7_0_comp_qa;
  xx_rsc_7_0_qb <= xx_rsc_7_0_comp_qb;

  xx_rsc_8_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_8_0_comp_adra,
      adrb => xx_rsc_8_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_8_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_8_0_clkb_en,
      da => xx_rsc_8_0_comp_da,
      db => xx_rsc_8_0_comp_db,
      qa => xx_rsc_8_0_comp_qa,
      qb => xx_rsc_8_0_comp_qb,
      wea => xx_rsc_8_0_wea,
      web => xx_rsc_8_0_web
    );
  xx_rsc_8_0_comp_adra <= xx_rsc_8_0_adra;
  xx_rsc_8_0_comp_adrb <= xx_rsc_8_0_adrb;
  xx_rsc_8_0_comp_da <= xx_rsc_8_0_da;
  xx_rsc_8_0_comp_db <= xx_rsc_8_0_db;
  xx_rsc_8_0_qa <= xx_rsc_8_0_comp_qa;
  xx_rsc_8_0_qb <= xx_rsc_8_0_comp_qb;

  xx_rsc_9_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_9_0_comp_adra,
      adrb => xx_rsc_9_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_9_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_9_0_clkb_en,
      da => xx_rsc_9_0_comp_da,
      db => xx_rsc_9_0_comp_db,
      qa => xx_rsc_9_0_comp_qa,
      qb => xx_rsc_9_0_comp_qb,
      wea => xx_rsc_9_0_wea,
      web => xx_rsc_9_0_web
    );
  xx_rsc_9_0_comp_adra <= xx_rsc_9_0_adra;
  xx_rsc_9_0_comp_adrb <= xx_rsc_9_0_adrb;
  xx_rsc_9_0_comp_da <= xx_rsc_9_0_da;
  xx_rsc_9_0_comp_db <= xx_rsc_9_0_db;
  xx_rsc_9_0_qa <= xx_rsc_9_0_comp_qa;
  xx_rsc_9_0_qb <= xx_rsc_9_0_comp_qb;

  xx_rsc_10_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_10_0_comp_adra,
      adrb => xx_rsc_10_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_10_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_10_0_clkb_en,
      da => xx_rsc_10_0_comp_da,
      db => xx_rsc_10_0_comp_db,
      qa => xx_rsc_10_0_comp_qa,
      qb => xx_rsc_10_0_comp_qb,
      wea => xx_rsc_10_0_wea,
      web => xx_rsc_10_0_web
    );
  xx_rsc_10_0_comp_adra <= xx_rsc_10_0_adra;
  xx_rsc_10_0_comp_adrb <= xx_rsc_10_0_adrb;
  xx_rsc_10_0_comp_da <= xx_rsc_10_0_da;
  xx_rsc_10_0_comp_db <= xx_rsc_10_0_db;
  xx_rsc_10_0_qa <= xx_rsc_10_0_comp_qa;
  xx_rsc_10_0_qb <= xx_rsc_10_0_comp_qb;

  xx_rsc_11_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_11_0_comp_adra,
      adrb => xx_rsc_11_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_11_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_11_0_clkb_en,
      da => xx_rsc_11_0_comp_da,
      db => xx_rsc_11_0_comp_db,
      qa => xx_rsc_11_0_comp_qa,
      qb => xx_rsc_11_0_comp_qb,
      wea => xx_rsc_11_0_wea,
      web => xx_rsc_11_0_web
    );
  xx_rsc_11_0_comp_adra <= xx_rsc_11_0_adra;
  xx_rsc_11_0_comp_adrb <= xx_rsc_11_0_adrb;
  xx_rsc_11_0_comp_da <= xx_rsc_11_0_da;
  xx_rsc_11_0_comp_db <= xx_rsc_11_0_db;
  xx_rsc_11_0_qa <= xx_rsc_11_0_comp_qa;
  xx_rsc_11_0_qb <= xx_rsc_11_0_comp_qb;

  xx_rsc_12_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_12_0_comp_adra,
      adrb => xx_rsc_12_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_12_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_12_0_clkb_en,
      da => xx_rsc_12_0_comp_da,
      db => xx_rsc_12_0_comp_db,
      qa => xx_rsc_12_0_comp_qa,
      qb => xx_rsc_12_0_comp_qb,
      wea => xx_rsc_12_0_wea,
      web => xx_rsc_12_0_web
    );
  xx_rsc_12_0_comp_adra <= xx_rsc_12_0_adra;
  xx_rsc_12_0_comp_adrb <= xx_rsc_12_0_adrb;
  xx_rsc_12_0_comp_da <= xx_rsc_12_0_da;
  xx_rsc_12_0_comp_db <= xx_rsc_12_0_db;
  xx_rsc_12_0_qa <= xx_rsc_12_0_comp_qa;
  xx_rsc_12_0_qb <= xx_rsc_12_0_comp_qb;

  xx_rsc_13_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_13_0_comp_adra,
      adrb => xx_rsc_13_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_13_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_13_0_clkb_en,
      da => xx_rsc_13_0_comp_da,
      db => xx_rsc_13_0_comp_db,
      qa => xx_rsc_13_0_comp_qa,
      qb => xx_rsc_13_0_comp_qb,
      wea => xx_rsc_13_0_wea,
      web => xx_rsc_13_0_web
    );
  xx_rsc_13_0_comp_adra <= xx_rsc_13_0_adra;
  xx_rsc_13_0_comp_adrb <= xx_rsc_13_0_adrb;
  xx_rsc_13_0_comp_da <= xx_rsc_13_0_da;
  xx_rsc_13_0_comp_db <= xx_rsc_13_0_db;
  xx_rsc_13_0_qa <= xx_rsc_13_0_comp_qa;
  xx_rsc_13_0_qb <= xx_rsc_13_0_comp_qb;

  xx_rsc_14_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_14_0_comp_adra,
      adrb => xx_rsc_14_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_14_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_14_0_clkb_en,
      da => xx_rsc_14_0_comp_da,
      db => xx_rsc_14_0_comp_db,
      qa => xx_rsc_14_0_comp_qa,
      qb => xx_rsc_14_0_comp_qb,
      wea => xx_rsc_14_0_wea,
      web => xx_rsc_14_0_web
    );
  xx_rsc_14_0_comp_adra <= xx_rsc_14_0_adra;
  xx_rsc_14_0_comp_adrb <= xx_rsc_14_0_adrb;
  xx_rsc_14_0_comp_da <= xx_rsc_14_0_da;
  xx_rsc_14_0_comp_db <= xx_rsc_14_0_db;
  xx_rsc_14_0_qa <= xx_rsc_14_0_comp_qa;
  xx_rsc_14_0_qb <= xx_rsc_14_0_comp_qb;

  xx_rsc_15_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_15_0_comp_adra,
      adrb => xx_rsc_15_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_15_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_15_0_clkb_en,
      da => xx_rsc_15_0_comp_da,
      db => xx_rsc_15_0_comp_db,
      qa => xx_rsc_15_0_comp_qa,
      qb => xx_rsc_15_0_comp_qb,
      wea => xx_rsc_15_0_wea,
      web => xx_rsc_15_0_web
    );
  xx_rsc_15_0_comp_adra <= xx_rsc_15_0_adra;
  xx_rsc_15_0_comp_adrb <= xx_rsc_15_0_adrb;
  xx_rsc_15_0_comp_da <= xx_rsc_15_0_da;
  xx_rsc_15_0_comp_db <= xx_rsc_15_0_db;
  xx_rsc_15_0_qa <= xx_rsc_15_0_comp_qa;
  xx_rsc_15_0_qb <= xx_rsc_15_0_comp_qb;

  xx_rsc_16_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_16_0_comp_adra,
      adrb => xx_rsc_16_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_16_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_16_0_clkb_en,
      da => xx_rsc_16_0_comp_da,
      db => xx_rsc_16_0_comp_db,
      qa => xx_rsc_16_0_comp_qa,
      qb => xx_rsc_16_0_comp_qb,
      wea => xx_rsc_16_0_wea,
      web => xx_rsc_16_0_web
    );
  xx_rsc_16_0_comp_adra <= xx_rsc_16_0_adra;
  xx_rsc_16_0_comp_adrb <= xx_rsc_16_0_adrb;
  xx_rsc_16_0_comp_da <= xx_rsc_16_0_da;
  xx_rsc_16_0_comp_db <= xx_rsc_16_0_db;
  xx_rsc_16_0_qa <= xx_rsc_16_0_comp_qa;
  xx_rsc_16_0_qb <= xx_rsc_16_0_comp_qb;

  xx_rsc_17_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_17_0_comp_adra,
      adrb => xx_rsc_17_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_17_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_17_0_clkb_en,
      da => xx_rsc_17_0_comp_da,
      db => xx_rsc_17_0_comp_db,
      qa => xx_rsc_17_0_comp_qa,
      qb => xx_rsc_17_0_comp_qb,
      wea => xx_rsc_17_0_wea,
      web => xx_rsc_17_0_web
    );
  xx_rsc_17_0_comp_adra <= xx_rsc_17_0_adra;
  xx_rsc_17_0_comp_adrb <= xx_rsc_17_0_adrb;
  xx_rsc_17_0_comp_da <= xx_rsc_17_0_da;
  xx_rsc_17_0_comp_db <= xx_rsc_17_0_db;
  xx_rsc_17_0_qa <= xx_rsc_17_0_comp_qa;
  xx_rsc_17_0_qb <= xx_rsc_17_0_comp_qb;

  xx_rsc_18_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_18_0_comp_adra,
      adrb => xx_rsc_18_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_18_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_18_0_clkb_en,
      da => xx_rsc_18_0_comp_da,
      db => xx_rsc_18_0_comp_db,
      qa => xx_rsc_18_0_comp_qa,
      qb => xx_rsc_18_0_comp_qb,
      wea => xx_rsc_18_0_wea,
      web => xx_rsc_18_0_web
    );
  xx_rsc_18_0_comp_adra <= xx_rsc_18_0_adra;
  xx_rsc_18_0_comp_adrb <= xx_rsc_18_0_adrb;
  xx_rsc_18_0_comp_da <= xx_rsc_18_0_da;
  xx_rsc_18_0_comp_db <= xx_rsc_18_0_db;
  xx_rsc_18_0_qa <= xx_rsc_18_0_comp_qa;
  xx_rsc_18_0_qb <= xx_rsc_18_0_comp_qb;

  xx_rsc_19_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_19_0_comp_adra,
      adrb => xx_rsc_19_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_19_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_19_0_clkb_en,
      da => xx_rsc_19_0_comp_da,
      db => xx_rsc_19_0_comp_db,
      qa => xx_rsc_19_0_comp_qa,
      qb => xx_rsc_19_0_comp_qb,
      wea => xx_rsc_19_0_wea,
      web => xx_rsc_19_0_web
    );
  xx_rsc_19_0_comp_adra <= xx_rsc_19_0_adra;
  xx_rsc_19_0_comp_adrb <= xx_rsc_19_0_adrb;
  xx_rsc_19_0_comp_da <= xx_rsc_19_0_da;
  xx_rsc_19_0_comp_db <= xx_rsc_19_0_db;
  xx_rsc_19_0_qa <= xx_rsc_19_0_comp_qa;
  xx_rsc_19_0_qb <= xx_rsc_19_0_comp_qb;

  xx_rsc_20_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_20_0_comp_adra,
      adrb => xx_rsc_20_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_20_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_20_0_clkb_en,
      da => xx_rsc_20_0_comp_da,
      db => xx_rsc_20_0_comp_db,
      qa => xx_rsc_20_0_comp_qa,
      qb => xx_rsc_20_0_comp_qb,
      wea => xx_rsc_20_0_wea,
      web => xx_rsc_20_0_web
    );
  xx_rsc_20_0_comp_adra <= xx_rsc_20_0_adra;
  xx_rsc_20_0_comp_adrb <= xx_rsc_20_0_adrb;
  xx_rsc_20_0_comp_da <= xx_rsc_20_0_da;
  xx_rsc_20_0_comp_db <= xx_rsc_20_0_db;
  xx_rsc_20_0_qa <= xx_rsc_20_0_comp_qa;
  xx_rsc_20_0_qb <= xx_rsc_20_0_comp_qb;

  xx_rsc_21_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_21_0_comp_adra,
      adrb => xx_rsc_21_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_21_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_21_0_clkb_en,
      da => xx_rsc_21_0_comp_da,
      db => xx_rsc_21_0_comp_db,
      qa => xx_rsc_21_0_comp_qa,
      qb => xx_rsc_21_0_comp_qb,
      wea => xx_rsc_21_0_wea,
      web => xx_rsc_21_0_web
    );
  xx_rsc_21_0_comp_adra <= xx_rsc_21_0_adra;
  xx_rsc_21_0_comp_adrb <= xx_rsc_21_0_adrb;
  xx_rsc_21_0_comp_da <= xx_rsc_21_0_da;
  xx_rsc_21_0_comp_db <= xx_rsc_21_0_db;
  xx_rsc_21_0_qa <= xx_rsc_21_0_comp_qa;
  xx_rsc_21_0_qb <= xx_rsc_21_0_comp_qb;

  xx_rsc_22_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_22_0_comp_adra,
      adrb => xx_rsc_22_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_22_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_22_0_clkb_en,
      da => xx_rsc_22_0_comp_da,
      db => xx_rsc_22_0_comp_db,
      qa => xx_rsc_22_0_comp_qa,
      qb => xx_rsc_22_0_comp_qb,
      wea => xx_rsc_22_0_wea,
      web => xx_rsc_22_0_web
    );
  xx_rsc_22_0_comp_adra <= xx_rsc_22_0_adra;
  xx_rsc_22_0_comp_adrb <= xx_rsc_22_0_adrb;
  xx_rsc_22_0_comp_da <= xx_rsc_22_0_da;
  xx_rsc_22_0_comp_db <= xx_rsc_22_0_db;
  xx_rsc_22_0_qa <= xx_rsc_22_0_comp_qa;
  xx_rsc_22_0_qb <= xx_rsc_22_0_comp_qb;

  xx_rsc_23_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_23_0_comp_adra,
      adrb => xx_rsc_23_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_23_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_23_0_clkb_en,
      da => xx_rsc_23_0_comp_da,
      db => xx_rsc_23_0_comp_db,
      qa => xx_rsc_23_0_comp_qa,
      qb => xx_rsc_23_0_comp_qb,
      wea => xx_rsc_23_0_wea,
      web => xx_rsc_23_0_web
    );
  xx_rsc_23_0_comp_adra <= xx_rsc_23_0_adra;
  xx_rsc_23_0_comp_adrb <= xx_rsc_23_0_adrb;
  xx_rsc_23_0_comp_da <= xx_rsc_23_0_da;
  xx_rsc_23_0_comp_db <= xx_rsc_23_0_db;
  xx_rsc_23_0_qa <= xx_rsc_23_0_comp_qa;
  xx_rsc_23_0_qb <= xx_rsc_23_0_comp_qb;

  xx_rsc_24_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_24_0_comp_adra,
      adrb => xx_rsc_24_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_24_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_24_0_clkb_en,
      da => xx_rsc_24_0_comp_da,
      db => xx_rsc_24_0_comp_db,
      qa => xx_rsc_24_0_comp_qa,
      qb => xx_rsc_24_0_comp_qb,
      wea => xx_rsc_24_0_wea,
      web => xx_rsc_24_0_web
    );
  xx_rsc_24_0_comp_adra <= xx_rsc_24_0_adra;
  xx_rsc_24_0_comp_adrb <= xx_rsc_24_0_adrb;
  xx_rsc_24_0_comp_da <= xx_rsc_24_0_da;
  xx_rsc_24_0_comp_db <= xx_rsc_24_0_db;
  xx_rsc_24_0_qa <= xx_rsc_24_0_comp_qa;
  xx_rsc_24_0_qb <= xx_rsc_24_0_comp_qb;

  xx_rsc_25_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_25_0_comp_adra,
      adrb => xx_rsc_25_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_25_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_25_0_clkb_en,
      da => xx_rsc_25_0_comp_da,
      db => xx_rsc_25_0_comp_db,
      qa => xx_rsc_25_0_comp_qa,
      qb => xx_rsc_25_0_comp_qb,
      wea => xx_rsc_25_0_wea,
      web => xx_rsc_25_0_web
    );
  xx_rsc_25_0_comp_adra <= xx_rsc_25_0_adra;
  xx_rsc_25_0_comp_adrb <= xx_rsc_25_0_adrb;
  xx_rsc_25_0_comp_da <= xx_rsc_25_0_da;
  xx_rsc_25_0_comp_db <= xx_rsc_25_0_db;
  xx_rsc_25_0_qa <= xx_rsc_25_0_comp_qa;
  xx_rsc_25_0_qb <= xx_rsc_25_0_comp_qb;

  xx_rsc_26_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_26_0_comp_adra,
      adrb => xx_rsc_26_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_26_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_26_0_clkb_en,
      da => xx_rsc_26_0_comp_da,
      db => xx_rsc_26_0_comp_db,
      qa => xx_rsc_26_0_comp_qa,
      qb => xx_rsc_26_0_comp_qb,
      wea => xx_rsc_26_0_wea,
      web => xx_rsc_26_0_web
    );
  xx_rsc_26_0_comp_adra <= xx_rsc_26_0_adra;
  xx_rsc_26_0_comp_adrb <= xx_rsc_26_0_adrb;
  xx_rsc_26_0_comp_da <= xx_rsc_26_0_da;
  xx_rsc_26_0_comp_db <= xx_rsc_26_0_db;
  xx_rsc_26_0_qa <= xx_rsc_26_0_comp_qa;
  xx_rsc_26_0_qb <= xx_rsc_26_0_comp_qb;

  xx_rsc_27_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_27_0_comp_adra,
      adrb => xx_rsc_27_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_27_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_27_0_clkb_en,
      da => xx_rsc_27_0_comp_da,
      db => xx_rsc_27_0_comp_db,
      qa => xx_rsc_27_0_comp_qa,
      qb => xx_rsc_27_0_comp_qb,
      wea => xx_rsc_27_0_wea,
      web => xx_rsc_27_0_web
    );
  xx_rsc_27_0_comp_adra <= xx_rsc_27_0_adra;
  xx_rsc_27_0_comp_adrb <= xx_rsc_27_0_adrb;
  xx_rsc_27_0_comp_da <= xx_rsc_27_0_da;
  xx_rsc_27_0_comp_db <= xx_rsc_27_0_db;
  xx_rsc_27_0_qa <= xx_rsc_27_0_comp_qa;
  xx_rsc_27_0_qb <= xx_rsc_27_0_comp_qb;

  xx_rsc_28_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_28_0_comp_adra,
      adrb => xx_rsc_28_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_28_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_28_0_clkb_en,
      da => xx_rsc_28_0_comp_da,
      db => xx_rsc_28_0_comp_db,
      qa => xx_rsc_28_0_comp_qa,
      qb => xx_rsc_28_0_comp_qb,
      wea => xx_rsc_28_0_wea,
      web => xx_rsc_28_0_web
    );
  xx_rsc_28_0_comp_adra <= xx_rsc_28_0_adra;
  xx_rsc_28_0_comp_adrb <= xx_rsc_28_0_adrb;
  xx_rsc_28_0_comp_da <= xx_rsc_28_0_da;
  xx_rsc_28_0_comp_db <= xx_rsc_28_0_db;
  xx_rsc_28_0_qa <= xx_rsc_28_0_comp_qa;
  xx_rsc_28_0_qb <= xx_rsc_28_0_comp_qb;

  xx_rsc_29_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_29_0_comp_adra,
      adrb => xx_rsc_29_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_29_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_29_0_clkb_en,
      da => xx_rsc_29_0_comp_da,
      db => xx_rsc_29_0_comp_db,
      qa => xx_rsc_29_0_comp_qa,
      qb => xx_rsc_29_0_comp_qb,
      wea => xx_rsc_29_0_wea,
      web => xx_rsc_29_0_web
    );
  xx_rsc_29_0_comp_adra <= xx_rsc_29_0_adra;
  xx_rsc_29_0_comp_adrb <= xx_rsc_29_0_adrb;
  xx_rsc_29_0_comp_da <= xx_rsc_29_0_da;
  xx_rsc_29_0_comp_db <= xx_rsc_29_0_db;
  xx_rsc_29_0_qa <= xx_rsc_29_0_comp_qa;
  xx_rsc_29_0_qb <= xx_rsc_29_0_comp_qb;

  xx_rsc_30_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_30_0_comp_adra,
      adrb => xx_rsc_30_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_30_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_30_0_clkb_en,
      da => xx_rsc_30_0_comp_da,
      db => xx_rsc_30_0_comp_db,
      qa => xx_rsc_30_0_comp_qa,
      qb => xx_rsc_30_0_comp_qb,
      wea => xx_rsc_30_0_wea,
      web => xx_rsc_30_0_web
    );
  xx_rsc_30_0_comp_adra <= xx_rsc_30_0_adra;
  xx_rsc_30_0_comp_adrb <= xx_rsc_30_0_adrb;
  xx_rsc_30_0_comp_da <= xx_rsc_30_0_da;
  xx_rsc_30_0_comp_db <= xx_rsc_30_0_db;
  xx_rsc_30_0_qa <= xx_rsc_30_0_comp_qa;
  xx_rsc_30_0_qb <= xx_rsc_30_0_comp_qb;

  xx_rsc_31_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => xx_rsc_31_0_comp_adra,
      adrb => xx_rsc_31_0_comp_adrb,
      clka => clk,
      clka_en => xx_rsc_31_0_clkb_en,
      clkb => clk,
      clkb_en => xx_rsc_31_0_clkb_en,
      da => xx_rsc_31_0_comp_da,
      db => xx_rsc_31_0_comp_db,
      qa => xx_rsc_31_0_comp_qa,
      qb => xx_rsc_31_0_comp_qb,
      wea => xx_rsc_31_0_wea,
      web => xx_rsc_31_0_web
    );
  xx_rsc_31_0_comp_adra <= xx_rsc_31_0_adra;
  xx_rsc_31_0_comp_adrb <= xx_rsc_31_0_adrb;
  xx_rsc_31_0_comp_da <= xx_rsc_31_0_da;
  xx_rsc_31_0_comp_db <= xx_rsc_31_0_db;
  xx_rsc_31_0_qa <= xx_rsc_31_0_comp_qa;
  xx_rsc_31_0_qb <= xx_rsc_31_0_comp_qb;

  yy_rsc_0_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_0_0_comp_adra,
      adrb => yy_rsc_0_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_0_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_0_0_clkb_en,
      da => yy_rsc_0_0_comp_da,
      db => yy_rsc_0_0_comp_db,
      qa => yy_rsc_0_0_comp_qa,
      qb => yy_rsc_0_0_comp_qb,
      wea => yy_rsc_0_0_wea,
      web => yy_rsc_0_0_web
    );
  yy_rsc_0_0_comp_adra <= yy_rsc_0_0_adra;
  yy_rsc_0_0_comp_adrb <= yy_rsc_0_0_adrb;
  yy_rsc_0_0_comp_da <= yy_rsc_0_0_da;
  yy_rsc_0_0_comp_db <= yy_rsc_0_0_db;
  yy_rsc_0_0_qa <= yy_rsc_0_0_comp_qa;
  yy_rsc_0_0_qb <= yy_rsc_0_0_comp_qb;

  yy_rsc_1_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_1_0_comp_adra,
      adrb => yy_rsc_1_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_1_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_1_0_clkb_en,
      da => yy_rsc_1_0_comp_da,
      db => yy_rsc_1_0_comp_db,
      qa => yy_rsc_1_0_comp_qa,
      qb => yy_rsc_1_0_comp_qb,
      wea => yy_rsc_1_0_wea,
      web => yy_rsc_1_0_web
    );
  yy_rsc_1_0_comp_adra <= yy_rsc_1_0_adra;
  yy_rsc_1_0_comp_adrb <= yy_rsc_1_0_adrb;
  yy_rsc_1_0_comp_da <= yy_rsc_1_0_da;
  yy_rsc_1_0_comp_db <= yy_rsc_1_0_db;
  yy_rsc_1_0_qa <= yy_rsc_1_0_comp_qa;
  yy_rsc_1_0_qb <= yy_rsc_1_0_comp_qb;

  yy_rsc_2_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_2_0_comp_adra,
      adrb => yy_rsc_2_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_2_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_2_0_clkb_en,
      da => yy_rsc_2_0_comp_da,
      db => yy_rsc_2_0_comp_db,
      qa => yy_rsc_2_0_comp_qa,
      qb => yy_rsc_2_0_comp_qb,
      wea => yy_rsc_2_0_wea,
      web => yy_rsc_2_0_web
    );
  yy_rsc_2_0_comp_adra <= yy_rsc_2_0_adra;
  yy_rsc_2_0_comp_adrb <= yy_rsc_2_0_adrb;
  yy_rsc_2_0_comp_da <= yy_rsc_2_0_da;
  yy_rsc_2_0_comp_db <= yy_rsc_2_0_db;
  yy_rsc_2_0_qa <= yy_rsc_2_0_comp_qa;
  yy_rsc_2_0_qb <= yy_rsc_2_0_comp_qb;

  yy_rsc_3_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_3_0_comp_adra,
      adrb => yy_rsc_3_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_3_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_3_0_clkb_en,
      da => yy_rsc_3_0_comp_da,
      db => yy_rsc_3_0_comp_db,
      qa => yy_rsc_3_0_comp_qa,
      qb => yy_rsc_3_0_comp_qb,
      wea => yy_rsc_3_0_wea,
      web => yy_rsc_3_0_web
    );
  yy_rsc_3_0_comp_adra <= yy_rsc_3_0_adra;
  yy_rsc_3_0_comp_adrb <= yy_rsc_3_0_adrb;
  yy_rsc_3_0_comp_da <= yy_rsc_3_0_da;
  yy_rsc_3_0_comp_db <= yy_rsc_3_0_db;
  yy_rsc_3_0_qa <= yy_rsc_3_0_comp_qa;
  yy_rsc_3_0_qb <= yy_rsc_3_0_comp_qb;

  yy_rsc_4_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_4_0_comp_adra,
      adrb => yy_rsc_4_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_4_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_4_0_clkb_en,
      da => yy_rsc_4_0_comp_da,
      db => yy_rsc_4_0_comp_db,
      qa => yy_rsc_4_0_comp_qa,
      qb => yy_rsc_4_0_comp_qb,
      wea => yy_rsc_4_0_wea,
      web => yy_rsc_4_0_web
    );
  yy_rsc_4_0_comp_adra <= yy_rsc_4_0_adra;
  yy_rsc_4_0_comp_adrb <= yy_rsc_4_0_adrb;
  yy_rsc_4_0_comp_da <= yy_rsc_4_0_da;
  yy_rsc_4_0_comp_db <= yy_rsc_4_0_db;
  yy_rsc_4_0_qa <= yy_rsc_4_0_comp_qa;
  yy_rsc_4_0_qb <= yy_rsc_4_0_comp_qb;

  yy_rsc_5_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_5_0_comp_adra,
      adrb => yy_rsc_5_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_5_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_5_0_clkb_en,
      da => yy_rsc_5_0_comp_da,
      db => yy_rsc_5_0_comp_db,
      qa => yy_rsc_5_0_comp_qa,
      qb => yy_rsc_5_0_comp_qb,
      wea => yy_rsc_5_0_wea,
      web => yy_rsc_5_0_web
    );
  yy_rsc_5_0_comp_adra <= yy_rsc_5_0_adra;
  yy_rsc_5_0_comp_adrb <= yy_rsc_5_0_adrb;
  yy_rsc_5_0_comp_da <= yy_rsc_5_0_da;
  yy_rsc_5_0_comp_db <= yy_rsc_5_0_db;
  yy_rsc_5_0_qa <= yy_rsc_5_0_comp_qa;
  yy_rsc_5_0_qb <= yy_rsc_5_0_comp_qb;

  yy_rsc_6_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_6_0_comp_adra,
      adrb => yy_rsc_6_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_6_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_6_0_clkb_en,
      da => yy_rsc_6_0_comp_da,
      db => yy_rsc_6_0_comp_db,
      qa => yy_rsc_6_0_comp_qa,
      qb => yy_rsc_6_0_comp_qb,
      wea => yy_rsc_6_0_wea,
      web => yy_rsc_6_0_web
    );
  yy_rsc_6_0_comp_adra <= yy_rsc_6_0_adra;
  yy_rsc_6_0_comp_adrb <= yy_rsc_6_0_adrb;
  yy_rsc_6_0_comp_da <= yy_rsc_6_0_da;
  yy_rsc_6_0_comp_db <= yy_rsc_6_0_db;
  yy_rsc_6_0_qa <= yy_rsc_6_0_comp_qa;
  yy_rsc_6_0_qb <= yy_rsc_6_0_comp_qb;

  yy_rsc_7_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_7_0_comp_adra,
      adrb => yy_rsc_7_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_7_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_7_0_clkb_en,
      da => yy_rsc_7_0_comp_da,
      db => yy_rsc_7_0_comp_db,
      qa => yy_rsc_7_0_comp_qa,
      qb => yy_rsc_7_0_comp_qb,
      wea => yy_rsc_7_0_wea,
      web => yy_rsc_7_0_web
    );
  yy_rsc_7_0_comp_adra <= yy_rsc_7_0_adra;
  yy_rsc_7_0_comp_adrb <= yy_rsc_7_0_adrb;
  yy_rsc_7_0_comp_da <= yy_rsc_7_0_da;
  yy_rsc_7_0_comp_db <= yy_rsc_7_0_db;
  yy_rsc_7_0_qa <= yy_rsc_7_0_comp_qa;
  yy_rsc_7_0_qb <= yy_rsc_7_0_comp_qb;

  yy_rsc_8_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_8_0_comp_adra,
      adrb => yy_rsc_8_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_8_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_8_0_clkb_en,
      da => yy_rsc_8_0_comp_da,
      db => yy_rsc_8_0_comp_db,
      qa => yy_rsc_8_0_comp_qa,
      qb => yy_rsc_8_0_comp_qb,
      wea => yy_rsc_8_0_wea,
      web => yy_rsc_8_0_web
    );
  yy_rsc_8_0_comp_adra <= yy_rsc_8_0_adra;
  yy_rsc_8_0_comp_adrb <= yy_rsc_8_0_adrb;
  yy_rsc_8_0_comp_da <= yy_rsc_8_0_da;
  yy_rsc_8_0_comp_db <= yy_rsc_8_0_db;
  yy_rsc_8_0_qa <= yy_rsc_8_0_comp_qa;
  yy_rsc_8_0_qb <= yy_rsc_8_0_comp_qb;

  yy_rsc_9_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_9_0_comp_adra,
      adrb => yy_rsc_9_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_9_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_9_0_clkb_en,
      da => yy_rsc_9_0_comp_da,
      db => yy_rsc_9_0_comp_db,
      qa => yy_rsc_9_0_comp_qa,
      qb => yy_rsc_9_0_comp_qb,
      wea => yy_rsc_9_0_wea,
      web => yy_rsc_9_0_web
    );
  yy_rsc_9_0_comp_adra <= yy_rsc_9_0_adra;
  yy_rsc_9_0_comp_adrb <= yy_rsc_9_0_adrb;
  yy_rsc_9_0_comp_da <= yy_rsc_9_0_da;
  yy_rsc_9_0_comp_db <= yy_rsc_9_0_db;
  yy_rsc_9_0_qa <= yy_rsc_9_0_comp_qa;
  yy_rsc_9_0_qb <= yy_rsc_9_0_comp_qb;

  yy_rsc_10_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_10_0_comp_adra,
      adrb => yy_rsc_10_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_10_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_10_0_clkb_en,
      da => yy_rsc_10_0_comp_da,
      db => yy_rsc_10_0_comp_db,
      qa => yy_rsc_10_0_comp_qa,
      qb => yy_rsc_10_0_comp_qb,
      wea => yy_rsc_10_0_wea,
      web => yy_rsc_10_0_web
    );
  yy_rsc_10_0_comp_adra <= yy_rsc_10_0_adra;
  yy_rsc_10_0_comp_adrb <= yy_rsc_10_0_adrb;
  yy_rsc_10_0_comp_da <= yy_rsc_10_0_da;
  yy_rsc_10_0_comp_db <= yy_rsc_10_0_db;
  yy_rsc_10_0_qa <= yy_rsc_10_0_comp_qa;
  yy_rsc_10_0_qb <= yy_rsc_10_0_comp_qb;

  yy_rsc_11_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_11_0_comp_adra,
      adrb => yy_rsc_11_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_11_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_11_0_clkb_en,
      da => yy_rsc_11_0_comp_da,
      db => yy_rsc_11_0_comp_db,
      qa => yy_rsc_11_0_comp_qa,
      qb => yy_rsc_11_0_comp_qb,
      wea => yy_rsc_11_0_wea,
      web => yy_rsc_11_0_web
    );
  yy_rsc_11_0_comp_adra <= yy_rsc_11_0_adra;
  yy_rsc_11_0_comp_adrb <= yy_rsc_11_0_adrb;
  yy_rsc_11_0_comp_da <= yy_rsc_11_0_da;
  yy_rsc_11_0_comp_db <= yy_rsc_11_0_db;
  yy_rsc_11_0_qa <= yy_rsc_11_0_comp_qa;
  yy_rsc_11_0_qb <= yy_rsc_11_0_comp_qb;

  yy_rsc_12_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_12_0_comp_adra,
      adrb => yy_rsc_12_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_12_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_12_0_clkb_en,
      da => yy_rsc_12_0_comp_da,
      db => yy_rsc_12_0_comp_db,
      qa => yy_rsc_12_0_comp_qa,
      qb => yy_rsc_12_0_comp_qb,
      wea => yy_rsc_12_0_wea,
      web => yy_rsc_12_0_web
    );
  yy_rsc_12_0_comp_adra <= yy_rsc_12_0_adra;
  yy_rsc_12_0_comp_adrb <= yy_rsc_12_0_adrb;
  yy_rsc_12_0_comp_da <= yy_rsc_12_0_da;
  yy_rsc_12_0_comp_db <= yy_rsc_12_0_db;
  yy_rsc_12_0_qa <= yy_rsc_12_0_comp_qa;
  yy_rsc_12_0_qb <= yy_rsc_12_0_comp_qb;

  yy_rsc_13_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_13_0_comp_adra,
      adrb => yy_rsc_13_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_13_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_13_0_clkb_en,
      da => yy_rsc_13_0_comp_da,
      db => yy_rsc_13_0_comp_db,
      qa => yy_rsc_13_0_comp_qa,
      qb => yy_rsc_13_0_comp_qb,
      wea => yy_rsc_13_0_wea,
      web => yy_rsc_13_0_web
    );
  yy_rsc_13_0_comp_adra <= yy_rsc_13_0_adra;
  yy_rsc_13_0_comp_adrb <= yy_rsc_13_0_adrb;
  yy_rsc_13_0_comp_da <= yy_rsc_13_0_da;
  yy_rsc_13_0_comp_db <= yy_rsc_13_0_db;
  yy_rsc_13_0_qa <= yy_rsc_13_0_comp_qa;
  yy_rsc_13_0_qb <= yy_rsc_13_0_comp_qb;

  yy_rsc_14_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_14_0_comp_adra,
      adrb => yy_rsc_14_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_14_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_14_0_clkb_en,
      da => yy_rsc_14_0_comp_da,
      db => yy_rsc_14_0_comp_db,
      qa => yy_rsc_14_0_comp_qa,
      qb => yy_rsc_14_0_comp_qb,
      wea => yy_rsc_14_0_wea,
      web => yy_rsc_14_0_web
    );
  yy_rsc_14_0_comp_adra <= yy_rsc_14_0_adra;
  yy_rsc_14_0_comp_adrb <= yy_rsc_14_0_adrb;
  yy_rsc_14_0_comp_da <= yy_rsc_14_0_da;
  yy_rsc_14_0_comp_db <= yy_rsc_14_0_db;
  yy_rsc_14_0_qa <= yy_rsc_14_0_comp_qa;
  yy_rsc_14_0_qb <= yy_rsc_14_0_comp_qb;

  yy_rsc_15_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_15_0_comp_adra,
      adrb => yy_rsc_15_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_15_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_15_0_clkb_en,
      da => yy_rsc_15_0_comp_da,
      db => yy_rsc_15_0_comp_db,
      qa => yy_rsc_15_0_comp_qa,
      qb => yy_rsc_15_0_comp_qb,
      wea => yy_rsc_15_0_wea,
      web => yy_rsc_15_0_web
    );
  yy_rsc_15_0_comp_adra <= yy_rsc_15_0_adra;
  yy_rsc_15_0_comp_adrb <= yy_rsc_15_0_adrb;
  yy_rsc_15_0_comp_da <= yy_rsc_15_0_da;
  yy_rsc_15_0_comp_db <= yy_rsc_15_0_db;
  yy_rsc_15_0_qa <= yy_rsc_15_0_comp_qa;
  yy_rsc_15_0_qb <= yy_rsc_15_0_comp_qb;

  yy_rsc_16_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_16_0_comp_adra,
      adrb => yy_rsc_16_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_16_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_16_0_clkb_en,
      da => yy_rsc_16_0_comp_da,
      db => yy_rsc_16_0_comp_db,
      qa => yy_rsc_16_0_comp_qa,
      qb => yy_rsc_16_0_comp_qb,
      wea => yy_rsc_16_0_wea,
      web => yy_rsc_16_0_web
    );
  yy_rsc_16_0_comp_adra <= yy_rsc_16_0_adra;
  yy_rsc_16_0_comp_adrb <= yy_rsc_16_0_adrb;
  yy_rsc_16_0_comp_da <= yy_rsc_16_0_da;
  yy_rsc_16_0_comp_db <= yy_rsc_16_0_db;
  yy_rsc_16_0_qa <= yy_rsc_16_0_comp_qa;
  yy_rsc_16_0_qb <= yy_rsc_16_0_comp_qb;

  yy_rsc_17_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_17_0_comp_adra,
      adrb => yy_rsc_17_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_17_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_17_0_clkb_en,
      da => yy_rsc_17_0_comp_da,
      db => yy_rsc_17_0_comp_db,
      qa => yy_rsc_17_0_comp_qa,
      qb => yy_rsc_17_0_comp_qb,
      wea => yy_rsc_17_0_wea,
      web => yy_rsc_17_0_web
    );
  yy_rsc_17_0_comp_adra <= yy_rsc_17_0_adra;
  yy_rsc_17_0_comp_adrb <= yy_rsc_17_0_adrb;
  yy_rsc_17_0_comp_da <= yy_rsc_17_0_da;
  yy_rsc_17_0_comp_db <= yy_rsc_17_0_db;
  yy_rsc_17_0_qa <= yy_rsc_17_0_comp_qa;
  yy_rsc_17_0_qb <= yy_rsc_17_0_comp_qb;

  yy_rsc_18_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_18_0_comp_adra,
      adrb => yy_rsc_18_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_18_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_18_0_clkb_en,
      da => yy_rsc_18_0_comp_da,
      db => yy_rsc_18_0_comp_db,
      qa => yy_rsc_18_0_comp_qa,
      qb => yy_rsc_18_0_comp_qb,
      wea => yy_rsc_18_0_wea,
      web => yy_rsc_18_0_web
    );
  yy_rsc_18_0_comp_adra <= yy_rsc_18_0_adra;
  yy_rsc_18_0_comp_adrb <= yy_rsc_18_0_adrb;
  yy_rsc_18_0_comp_da <= yy_rsc_18_0_da;
  yy_rsc_18_0_comp_db <= yy_rsc_18_0_db;
  yy_rsc_18_0_qa <= yy_rsc_18_0_comp_qa;
  yy_rsc_18_0_qb <= yy_rsc_18_0_comp_qb;

  yy_rsc_19_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_19_0_comp_adra,
      adrb => yy_rsc_19_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_19_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_19_0_clkb_en,
      da => yy_rsc_19_0_comp_da,
      db => yy_rsc_19_0_comp_db,
      qa => yy_rsc_19_0_comp_qa,
      qb => yy_rsc_19_0_comp_qb,
      wea => yy_rsc_19_0_wea,
      web => yy_rsc_19_0_web
    );
  yy_rsc_19_0_comp_adra <= yy_rsc_19_0_adra;
  yy_rsc_19_0_comp_adrb <= yy_rsc_19_0_adrb;
  yy_rsc_19_0_comp_da <= yy_rsc_19_0_da;
  yy_rsc_19_0_comp_db <= yy_rsc_19_0_db;
  yy_rsc_19_0_qa <= yy_rsc_19_0_comp_qa;
  yy_rsc_19_0_qb <= yy_rsc_19_0_comp_qb;

  yy_rsc_20_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_20_0_comp_adra,
      adrb => yy_rsc_20_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_20_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_20_0_clkb_en,
      da => yy_rsc_20_0_comp_da,
      db => yy_rsc_20_0_comp_db,
      qa => yy_rsc_20_0_comp_qa,
      qb => yy_rsc_20_0_comp_qb,
      wea => yy_rsc_20_0_wea,
      web => yy_rsc_20_0_web
    );
  yy_rsc_20_0_comp_adra <= yy_rsc_20_0_adra;
  yy_rsc_20_0_comp_adrb <= yy_rsc_20_0_adrb;
  yy_rsc_20_0_comp_da <= yy_rsc_20_0_da;
  yy_rsc_20_0_comp_db <= yy_rsc_20_0_db;
  yy_rsc_20_0_qa <= yy_rsc_20_0_comp_qa;
  yy_rsc_20_0_qb <= yy_rsc_20_0_comp_qb;

  yy_rsc_21_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_21_0_comp_adra,
      adrb => yy_rsc_21_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_21_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_21_0_clkb_en,
      da => yy_rsc_21_0_comp_da,
      db => yy_rsc_21_0_comp_db,
      qa => yy_rsc_21_0_comp_qa,
      qb => yy_rsc_21_0_comp_qb,
      wea => yy_rsc_21_0_wea,
      web => yy_rsc_21_0_web
    );
  yy_rsc_21_0_comp_adra <= yy_rsc_21_0_adra;
  yy_rsc_21_0_comp_adrb <= yy_rsc_21_0_adrb;
  yy_rsc_21_0_comp_da <= yy_rsc_21_0_da;
  yy_rsc_21_0_comp_db <= yy_rsc_21_0_db;
  yy_rsc_21_0_qa <= yy_rsc_21_0_comp_qa;
  yy_rsc_21_0_qb <= yy_rsc_21_0_comp_qb;

  yy_rsc_22_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_22_0_comp_adra,
      adrb => yy_rsc_22_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_22_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_22_0_clkb_en,
      da => yy_rsc_22_0_comp_da,
      db => yy_rsc_22_0_comp_db,
      qa => yy_rsc_22_0_comp_qa,
      qb => yy_rsc_22_0_comp_qb,
      wea => yy_rsc_22_0_wea,
      web => yy_rsc_22_0_web
    );
  yy_rsc_22_0_comp_adra <= yy_rsc_22_0_adra;
  yy_rsc_22_0_comp_adrb <= yy_rsc_22_0_adrb;
  yy_rsc_22_0_comp_da <= yy_rsc_22_0_da;
  yy_rsc_22_0_comp_db <= yy_rsc_22_0_db;
  yy_rsc_22_0_qa <= yy_rsc_22_0_comp_qa;
  yy_rsc_22_0_qb <= yy_rsc_22_0_comp_qb;

  yy_rsc_23_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_23_0_comp_adra,
      adrb => yy_rsc_23_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_23_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_23_0_clkb_en,
      da => yy_rsc_23_0_comp_da,
      db => yy_rsc_23_0_comp_db,
      qa => yy_rsc_23_0_comp_qa,
      qb => yy_rsc_23_0_comp_qb,
      wea => yy_rsc_23_0_wea,
      web => yy_rsc_23_0_web
    );
  yy_rsc_23_0_comp_adra <= yy_rsc_23_0_adra;
  yy_rsc_23_0_comp_adrb <= yy_rsc_23_0_adrb;
  yy_rsc_23_0_comp_da <= yy_rsc_23_0_da;
  yy_rsc_23_0_comp_db <= yy_rsc_23_0_db;
  yy_rsc_23_0_qa <= yy_rsc_23_0_comp_qa;
  yy_rsc_23_0_qb <= yy_rsc_23_0_comp_qb;

  yy_rsc_24_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_24_0_comp_adra,
      adrb => yy_rsc_24_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_24_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_24_0_clkb_en,
      da => yy_rsc_24_0_comp_da,
      db => yy_rsc_24_0_comp_db,
      qa => yy_rsc_24_0_comp_qa,
      qb => yy_rsc_24_0_comp_qb,
      wea => yy_rsc_24_0_wea,
      web => yy_rsc_24_0_web
    );
  yy_rsc_24_0_comp_adra <= yy_rsc_24_0_adra;
  yy_rsc_24_0_comp_adrb <= yy_rsc_24_0_adrb;
  yy_rsc_24_0_comp_da <= yy_rsc_24_0_da;
  yy_rsc_24_0_comp_db <= yy_rsc_24_0_db;
  yy_rsc_24_0_qa <= yy_rsc_24_0_comp_qa;
  yy_rsc_24_0_qb <= yy_rsc_24_0_comp_qb;

  yy_rsc_25_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_25_0_comp_adra,
      adrb => yy_rsc_25_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_25_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_25_0_clkb_en,
      da => yy_rsc_25_0_comp_da,
      db => yy_rsc_25_0_comp_db,
      qa => yy_rsc_25_0_comp_qa,
      qb => yy_rsc_25_0_comp_qb,
      wea => yy_rsc_25_0_wea,
      web => yy_rsc_25_0_web
    );
  yy_rsc_25_0_comp_adra <= yy_rsc_25_0_adra;
  yy_rsc_25_0_comp_adrb <= yy_rsc_25_0_adrb;
  yy_rsc_25_0_comp_da <= yy_rsc_25_0_da;
  yy_rsc_25_0_comp_db <= yy_rsc_25_0_db;
  yy_rsc_25_0_qa <= yy_rsc_25_0_comp_qa;
  yy_rsc_25_0_qb <= yy_rsc_25_0_comp_qb;

  yy_rsc_26_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_26_0_comp_adra,
      adrb => yy_rsc_26_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_26_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_26_0_clkb_en,
      da => yy_rsc_26_0_comp_da,
      db => yy_rsc_26_0_comp_db,
      qa => yy_rsc_26_0_comp_qa,
      qb => yy_rsc_26_0_comp_qb,
      wea => yy_rsc_26_0_wea,
      web => yy_rsc_26_0_web
    );
  yy_rsc_26_0_comp_adra <= yy_rsc_26_0_adra;
  yy_rsc_26_0_comp_adrb <= yy_rsc_26_0_adrb;
  yy_rsc_26_0_comp_da <= yy_rsc_26_0_da;
  yy_rsc_26_0_comp_db <= yy_rsc_26_0_db;
  yy_rsc_26_0_qa <= yy_rsc_26_0_comp_qa;
  yy_rsc_26_0_qb <= yy_rsc_26_0_comp_qb;

  yy_rsc_27_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_27_0_comp_adra,
      adrb => yy_rsc_27_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_27_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_27_0_clkb_en,
      da => yy_rsc_27_0_comp_da,
      db => yy_rsc_27_0_comp_db,
      qa => yy_rsc_27_0_comp_qa,
      qb => yy_rsc_27_0_comp_qb,
      wea => yy_rsc_27_0_wea,
      web => yy_rsc_27_0_web
    );
  yy_rsc_27_0_comp_adra <= yy_rsc_27_0_adra;
  yy_rsc_27_0_comp_adrb <= yy_rsc_27_0_adrb;
  yy_rsc_27_0_comp_da <= yy_rsc_27_0_da;
  yy_rsc_27_0_comp_db <= yy_rsc_27_0_db;
  yy_rsc_27_0_qa <= yy_rsc_27_0_comp_qa;
  yy_rsc_27_0_qb <= yy_rsc_27_0_comp_qb;

  yy_rsc_28_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_28_0_comp_adra,
      adrb => yy_rsc_28_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_28_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_28_0_clkb_en,
      da => yy_rsc_28_0_comp_da,
      db => yy_rsc_28_0_comp_db,
      qa => yy_rsc_28_0_comp_qa,
      qb => yy_rsc_28_0_comp_qb,
      wea => yy_rsc_28_0_wea,
      web => yy_rsc_28_0_web
    );
  yy_rsc_28_0_comp_adra <= yy_rsc_28_0_adra;
  yy_rsc_28_0_comp_adrb <= yy_rsc_28_0_adrb;
  yy_rsc_28_0_comp_da <= yy_rsc_28_0_da;
  yy_rsc_28_0_comp_db <= yy_rsc_28_0_db;
  yy_rsc_28_0_qa <= yy_rsc_28_0_comp_qa;
  yy_rsc_28_0_qb <= yy_rsc_28_0_comp_qb;

  yy_rsc_29_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_29_0_comp_adra,
      adrb => yy_rsc_29_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_29_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_29_0_clkb_en,
      da => yy_rsc_29_0_comp_da,
      db => yy_rsc_29_0_comp_db,
      qa => yy_rsc_29_0_comp_qa,
      qb => yy_rsc_29_0_comp_qb,
      wea => yy_rsc_29_0_wea,
      web => yy_rsc_29_0_web
    );
  yy_rsc_29_0_comp_adra <= yy_rsc_29_0_adra;
  yy_rsc_29_0_comp_adrb <= yy_rsc_29_0_adrb;
  yy_rsc_29_0_comp_da <= yy_rsc_29_0_da;
  yy_rsc_29_0_comp_db <= yy_rsc_29_0_db;
  yy_rsc_29_0_qa <= yy_rsc_29_0_comp_qa;
  yy_rsc_29_0_qb <= yy_rsc_29_0_comp_qb;

  yy_rsc_30_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_30_0_comp_adra,
      adrb => yy_rsc_30_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_30_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_30_0_clkb_en,
      da => yy_rsc_30_0_comp_da,
      db => yy_rsc_30_0_comp_db,
      qa => yy_rsc_30_0_comp_qa,
      qb => yy_rsc_30_0_comp_qb,
      wea => yy_rsc_30_0_wea,
      web => yy_rsc_30_0_web
    );
  yy_rsc_30_0_comp_adra <= yy_rsc_30_0_adra;
  yy_rsc_30_0_comp_adrb <= yy_rsc_30_0_adrb;
  yy_rsc_30_0_comp_da <= yy_rsc_30_0_da;
  yy_rsc_30_0_comp_db <= yy_rsc_30_0_db;
  yy_rsc_30_0_qa <= yy_rsc_30_0_comp_qa;
  yy_rsc_30_0_qb <= yy_rsc_30_0_comp_qb;

  yy_rsc_31_0_comp : work.block_dpram_rbw_dual_pkg.BLOCK_DPRAM_RBW_DUAL
    GENERIC MAP(
      addr_width => 5,
      data_width => 32,
      depth => 32,
      latency => 1
      )
    PORT MAP(
      adra => yy_rsc_31_0_comp_adra,
      adrb => yy_rsc_31_0_comp_adrb,
      clka => clk,
      clka_en => yy_rsc_31_0_clkb_en,
      clkb => clk,
      clkb_en => yy_rsc_31_0_clkb_en,
      da => yy_rsc_31_0_comp_da,
      db => yy_rsc_31_0_comp_db,
      qa => yy_rsc_31_0_comp_qa,
      qb => yy_rsc_31_0_comp_qb,
      wea => yy_rsc_31_0_wea,
      web => yy_rsc_31_0_web
    );
  yy_rsc_31_0_comp_adra <= yy_rsc_31_0_adra;
  yy_rsc_31_0_comp_adrb <= yy_rsc_31_0_adrb;
  yy_rsc_31_0_comp_da <= yy_rsc_31_0_da;
  yy_rsc_31_0_comp_db <= yy_rsc_31_0_db;
  yy_rsc_31_0_qa <= yy_rsc_31_0_comp_qa;
  yy_rsc_31_0_qb <= yy_rsc_31_0_comp_qb;

  twiddle_rsci : hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_3_5_32_32_32_32_1_gen
    PORT MAP(
      qb => twiddle_rsci_qb,
      adrb => twiddle_rsci_adrb,
      adrb_d => twiddle_rsci_adrb_d_1,
      qb_d => twiddle_rsci_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_rsci_qb <= twiddle_rsc_qb;
  twiddle_rsc_adrb <= twiddle_rsci_adrb;
  twiddle_rsci_adrb_d_1 <= twiddle_rsci_adrb_d;
  twiddle_rsci_qb_d <= twiddle_rsci_qb_d_1;

  twiddle_h_rsci : hybrid_Xilinx_RAMS_BLOCK_2R1W_RBW_rport_4_5_32_32_32_32_1_gen
    PORT MAP(
      qb => twiddle_h_rsci_qb,
      adrb => twiddle_h_rsci_adrb,
      adrb_d => twiddle_h_rsci_adrb_d_1,
      qb_d => twiddle_h_rsci_qb_d_1,
      readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d
    );
  twiddle_h_rsci_qb <= twiddle_h_rsc_qb;
  twiddle_h_rsc_adrb <= twiddle_h_rsci_adrb;
  twiddle_h_rsci_adrb_d_1 <= twiddle_h_rsci_adrb_d;
  twiddle_h_rsci_qb_d <= twiddle_h_rsci_qb_d_1;

  xx_rsc_0_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_0_0_clkb_en,
      clka_en => xx_rsc_0_0_clka_en,
      qb => xx_rsc_0_0_i_qb,
      web => xx_rsc_0_0_web,
      db => xx_rsc_0_0_i_db,
      adrb => xx_rsc_0_0_i_adrb,
      qa => xx_rsc_0_0_i_qa,
      wea => xx_rsc_0_0_wea,
      da => xx_rsc_0_0_i_da,
      adra => xx_rsc_0_0_i_adra,
      adra_d => xx_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_0_0_i_clka_en_d,
      clkb_en_d => xx_rsc_0_0_i_clka_en_d,
      da_d => xx_rsc_0_0_i_da_d,
      qa_d => xx_rsc_0_0_i_qa_d_1,
      wea_d => xx_rsc_0_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_0_0_i_qb <= xx_rsc_0_0_qb;
  xx_rsc_0_0_db <= xx_rsc_0_0_i_db;
  xx_rsc_0_0_adrb <= xx_rsc_0_0_i_adrb;
  xx_rsc_0_0_i_qa <= xx_rsc_0_0_qa;
  xx_rsc_0_0_da <= xx_rsc_0_0_i_da;
  xx_rsc_0_0_adra <= xx_rsc_0_0_i_adra;
  xx_rsc_0_0_i_adra_d_1 <= xx_rsc_0_0_i_adra_d;
  xx_rsc_0_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_0_0_i_qa_d <= xx_rsc_0_0_i_qa_d_1;
  xx_rsc_0_0_i_wea_d_1 <= xx_rsc_0_0_i_wea_d;
  xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_1_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_1_0_clkb_en,
      clka_en => xx_rsc_1_0_clka_en,
      qb => xx_rsc_1_0_i_qb,
      web => xx_rsc_1_0_web,
      db => xx_rsc_1_0_i_db,
      adrb => xx_rsc_1_0_i_adrb,
      qa => xx_rsc_1_0_i_qa,
      wea => xx_rsc_1_0_wea,
      da => xx_rsc_1_0_i_da,
      adra => xx_rsc_1_0_i_adra,
      adra_d => xx_rsc_1_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_1_0_i_clka_en_d,
      clkb_en_d => xx_rsc_1_0_i_clka_en_d,
      da_d => xx_rsc_1_0_i_da_d,
      qa_d => xx_rsc_1_0_i_qa_d_1,
      wea_d => xx_rsc_1_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_1_0_i_qb <= xx_rsc_1_0_qb;
  xx_rsc_1_0_db <= xx_rsc_1_0_i_db;
  xx_rsc_1_0_adrb <= xx_rsc_1_0_i_adrb;
  xx_rsc_1_0_i_qa <= xx_rsc_1_0_qa;
  xx_rsc_1_0_da <= xx_rsc_1_0_i_da;
  xx_rsc_1_0_adra <= xx_rsc_1_0_i_adra;
  xx_rsc_1_0_i_adra_d_1 <= xx_rsc_1_0_i_adra_d;
  xx_rsc_1_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_1_0_i_qa_d <= xx_rsc_1_0_i_qa_d_1;
  xx_rsc_1_0_i_wea_d_1 <= xx_rsc_1_0_i_wea_d;
  xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_2_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_2_0_clkb_en,
      clka_en => xx_rsc_2_0_clka_en,
      qb => xx_rsc_2_0_i_qb,
      web => xx_rsc_2_0_web,
      db => xx_rsc_2_0_i_db,
      adrb => xx_rsc_2_0_i_adrb,
      qa => xx_rsc_2_0_i_qa,
      wea => xx_rsc_2_0_wea,
      da => xx_rsc_2_0_i_da,
      adra => xx_rsc_2_0_i_adra,
      adra_d => xx_rsc_2_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_2_0_i_clka_en_d,
      clkb_en_d => xx_rsc_2_0_i_clka_en_d,
      da_d => xx_rsc_2_0_i_da_d,
      qa_d => xx_rsc_2_0_i_qa_d_1,
      wea_d => xx_rsc_2_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_2_0_i_qb <= xx_rsc_2_0_qb;
  xx_rsc_2_0_db <= xx_rsc_2_0_i_db;
  xx_rsc_2_0_adrb <= xx_rsc_2_0_i_adrb;
  xx_rsc_2_0_i_qa <= xx_rsc_2_0_qa;
  xx_rsc_2_0_da <= xx_rsc_2_0_i_da;
  xx_rsc_2_0_adra <= xx_rsc_2_0_i_adra;
  xx_rsc_2_0_i_adra_d_1 <= xx_rsc_2_0_i_adra_d;
  xx_rsc_2_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_2_0_i_qa_d <= xx_rsc_2_0_i_qa_d_1;
  xx_rsc_2_0_i_wea_d_1 <= xx_rsc_2_0_i_wea_d;
  xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_3_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_3_0_clkb_en,
      clka_en => xx_rsc_3_0_clka_en,
      qb => xx_rsc_3_0_i_qb,
      web => xx_rsc_3_0_web,
      db => xx_rsc_3_0_i_db,
      adrb => xx_rsc_3_0_i_adrb,
      qa => xx_rsc_3_0_i_qa,
      wea => xx_rsc_3_0_wea,
      da => xx_rsc_3_0_i_da,
      adra => xx_rsc_3_0_i_adra,
      adra_d => xx_rsc_3_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_3_0_i_clka_en_d,
      clkb_en_d => xx_rsc_3_0_i_clka_en_d,
      da_d => xx_rsc_3_0_i_da_d,
      qa_d => xx_rsc_3_0_i_qa_d_1,
      wea_d => xx_rsc_3_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_3_0_i_qb <= xx_rsc_3_0_qb;
  xx_rsc_3_0_db <= xx_rsc_3_0_i_db;
  xx_rsc_3_0_adrb <= xx_rsc_3_0_i_adrb;
  xx_rsc_3_0_i_qa <= xx_rsc_3_0_qa;
  xx_rsc_3_0_da <= xx_rsc_3_0_i_da;
  xx_rsc_3_0_adra <= xx_rsc_3_0_i_adra;
  xx_rsc_3_0_i_adra_d_1 <= xx_rsc_3_0_i_adra_d;
  xx_rsc_3_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_3_0_i_qa_d <= xx_rsc_3_0_i_qa_d_1;
  xx_rsc_3_0_i_wea_d_1 <= xx_rsc_3_0_i_wea_d;
  xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_4_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_4_0_clkb_en,
      clka_en => xx_rsc_4_0_clka_en,
      qb => xx_rsc_4_0_i_qb,
      web => xx_rsc_4_0_web,
      db => xx_rsc_4_0_i_db,
      adrb => xx_rsc_4_0_i_adrb,
      qa => xx_rsc_4_0_i_qa,
      wea => xx_rsc_4_0_wea,
      da => xx_rsc_4_0_i_da,
      adra => xx_rsc_4_0_i_adra,
      adra_d => xx_rsc_4_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_4_0_i_clka_en_d,
      clkb_en_d => xx_rsc_4_0_i_clka_en_d,
      da_d => xx_rsc_4_0_i_da_d,
      qa_d => xx_rsc_4_0_i_qa_d_1,
      wea_d => xx_rsc_4_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_4_0_i_qb <= xx_rsc_4_0_qb;
  xx_rsc_4_0_db <= xx_rsc_4_0_i_db;
  xx_rsc_4_0_adrb <= xx_rsc_4_0_i_adrb;
  xx_rsc_4_0_i_qa <= xx_rsc_4_0_qa;
  xx_rsc_4_0_da <= xx_rsc_4_0_i_da;
  xx_rsc_4_0_adra <= xx_rsc_4_0_i_adra;
  xx_rsc_4_0_i_adra_d_1 <= xx_rsc_4_0_i_adra_d;
  xx_rsc_4_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_4_0_i_qa_d <= xx_rsc_4_0_i_qa_d_1;
  xx_rsc_4_0_i_wea_d_1 <= xx_rsc_4_0_i_wea_d;
  xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_5_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_5_0_clkb_en,
      clka_en => xx_rsc_5_0_clka_en,
      qb => xx_rsc_5_0_i_qb,
      web => xx_rsc_5_0_web,
      db => xx_rsc_5_0_i_db,
      adrb => xx_rsc_5_0_i_adrb,
      qa => xx_rsc_5_0_i_qa,
      wea => xx_rsc_5_0_wea,
      da => xx_rsc_5_0_i_da,
      adra => xx_rsc_5_0_i_adra,
      adra_d => xx_rsc_5_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_5_0_i_clka_en_d,
      clkb_en_d => xx_rsc_5_0_i_clka_en_d,
      da_d => xx_rsc_5_0_i_da_d,
      qa_d => xx_rsc_5_0_i_qa_d_1,
      wea_d => xx_rsc_5_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_5_0_i_qb <= xx_rsc_5_0_qb;
  xx_rsc_5_0_db <= xx_rsc_5_0_i_db;
  xx_rsc_5_0_adrb <= xx_rsc_5_0_i_adrb;
  xx_rsc_5_0_i_qa <= xx_rsc_5_0_qa;
  xx_rsc_5_0_da <= xx_rsc_5_0_i_da;
  xx_rsc_5_0_adra <= xx_rsc_5_0_i_adra;
  xx_rsc_5_0_i_adra_d_1 <= xx_rsc_5_0_i_adra_d;
  xx_rsc_5_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_5_0_i_qa_d <= xx_rsc_5_0_i_qa_d_1;
  xx_rsc_5_0_i_wea_d_1 <= xx_rsc_5_0_i_wea_d;
  xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_6_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_6_0_clkb_en,
      clka_en => xx_rsc_6_0_clka_en,
      qb => xx_rsc_6_0_i_qb,
      web => xx_rsc_6_0_web,
      db => xx_rsc_6_0_i_db,
      adrb => xx_rsc_6_0_i_adrb,
      qa => xx_rsc_6_0_i_qa,
      wea => xx_rsc_6_0_wea,
      da => xx_rsc_6_0_i_da,
      adra => xx_rsc_6_0_i_adra,
      adra_d => xx_rsc_6_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_6_0_i_clka_en_d,
      clkb_en_d => xx_rsc_6_0_i_clka_en_d,
      da_d => xx_rsc_6_0_i_da_d,
      qa_d => xx_rsc_6_0_i_qa_d_1,
      wea_d => xx_rsc_6_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_6_0_i_qb <= xx_rsc_6_0_qb;
  xx_rsc_6_0_db <= xx_rsc_6_0_i_db;
  xx_rsc_6_0_adrb <= xx_rsc_6_0_i_adrb;
  xx_rsc_6_0_i_qa <= xx_rsc_6_0_qa;
  xx_rsc_6_0_da <= xx_rsc_6_0_i_da;
  xx_rsc_6_0_adra <= xx_rsc_6_0_i_adra;
  xx_rsc_6_0_i_adra_d_1 <= xx_rsc_6_0_i_adra_d;
  xx_rsc_6_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_6_0_i_qa_d <= xx_rsc_6_0_i_qa_d_1;
  xx_rsc_6_0_i_wea_d_1 <= xx_rsc_6_0_i_wea_d;
  xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_7_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_7_0_clkb_en,
      clka_en => xx_rsc_7_0_clka_en,
      qb => xx_rsc_7_0_i_qb,
      web => xx_rsc_7_0_web,
      db => xx_rsc_7_0_i_db,
      adrb => xx_rsc_7_0_i_adrb,
      qa => xx_rsc_7_0_i_qa,
      wea => xx_rsc_7_0_wea,
      da => xx_rsc_7_0_i_da,
      adra => xx_rsc_7_0_i_adra,
      adra_d => xx_rsc_7_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_7_0_i_clka_en_d,
      clkb_en_d => xx_rsc_7_0_i_clka_en_d,
      da_d => xx_rsc_7_0_i_da_d,
      qa_d => xx_rsc_7_0_i_qa_d_1,
      wea_d => xx_rsc_7_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_7_0_i_qb <= xx_rsc_7_0_qb;
  xx_rsc_7_0_db <= xx_rsc_7_0_i_db;
  xx_rsc_7_0_adrb <= xx_rsc_7_0_i_adrb;
  xx_rsc_7_0_i_qa <= xx_rsc_7_0_qa;
  xx_rsc_7_0_da <= xx_rsc_7_0_i_da;
  xx_rsc_7_0_adra <= xx_rsc_7_0_i_adra;
  xx_rsc_7_0_i_adra_d_1 <= xx_rsc_7_0_i_adra_d;
  xx_rsc_7_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_7_0_i_qa_d <= xx_rsc_7_0_i_qa_d_1;
  xx_rsc_7_0_i_wea_d_1 <= xx_rsc_7_0_i_wea_d;
  xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_8_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_8_0_clkb_en,
      clka_en => xx_rsc_8_0_clka_en,
      qb => xx_rsc_8_0_i_qb,
      web => xx_rsc_8_0_web,
      db => xx_rsc_8_0_i_db,
      adrb => xx_rsc_8_0_i_adrb,
      qa => xx_rsc_8_0_i_qa,
      wea => xx_rsc_8_0_wea,
      da => xx_rsc_8_0_i_da,
      adra => xx_rsc_8_0_i_adra,
      adra_d => xx_rsc_8_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_8_0_i_clka_en_d,
      clkb_en_d => xx_rsc_8_0_i_clka_en_d,
      da_d => xx_rsc_8_0_i_da_d,
      qa_d => xx_rsc_8_0_i_qa_d_1,
      wea_d => xx_rsc_8_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_8_0_i_qb <= xx_rsc_8_0_qb;
  xx_rsc_8_0_db <= xx_rsc_8_0_i_db;
  xx_rsc_8_0_adrb <= xx_rsc_8_0_i_adrb;
  xx_rsc_8_0_i_qa <= xx_rsc_8_0_qa;
  xx_rsc_8_0_da <= xx_rsc_8_0_i_da;
  xx_rsc_8_0_adra <= xx_rsc_8_0_i_adra;
  xx_rsc_8_0_i_adra_d_1 <= xx_rsc_8_0_i_adra_d;
  xx_rsc_8_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_8_0_i_qa_d <= xx_rsc_8_0_i_qa_d_1;
  xx_rsc_8_0_i_wea_d_1 <= xx_rsc_8_0_i_wea_d;
  xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_9_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_9_0_clkb_en,
      clka_en => xx_rsc_9_0_clka_en,
      qb => xx_rsc_9_0_i_qb,
      web => xx_rsc_9_0_web,
      db => xx_rsc_9_0_i_db,
      adrb => xx_rsc_9_0_i_adrb,
      qa => xx_rsc_9_0_i_qa,
      wea => xx_rsc_9_0_wea,
      da => xx_rsc_9_0_i_da,
      adra => xx_rsc_9_0_i_adra,
      adra_d => xx_rsc_9_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_9_0_i_clka_en_d,
      clkb_en_d => xx_rsc_9_0_i_clka_en_d,
      da_d => xx_rsc_9_0_i_da_d,
      qa_d => xx_rsc_9_0_i_qa_d_1,
      wea_d => xx_rsc_9_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_9_0_i_qb <= xx_rsc_9_0_qb;
  xx_rsc_9_0_db <= xx_rsc_9_0_i_db;
  xx_rsc_9_0_adrb <= xx_rsc_9_0_i_adrb;
  xx_rsc_9_0_i_qa <= xx_rsc_9_0_qa;
  xx_rsc_9_0_da <= xx_rsc_9_0_i_da;
  xx_rsc_9_0_adra <= xx_rsc_9_0_i_adra;
  xx_rsc_9_0_i_adra_d_1 <= xx_rsc_9_0_i_adra_d;
  xx_rsc_9_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_9_0_i_qa_d <= xx_rsc_9_0_i_qa_d_1;
  xx_rsc_9_0_i_wea_d_1 <= xx_rsc_9_0_i_wea_d;
  xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_10_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_10_0_clkb_en,
      clka_en => xx_rsc_10_0_clka_en,
      qb => xx_rsc_10_0_i_qb,
      web => xx_rsc_10_0_web,
      db => xx_rsc_10_0_i_db,
      adrb => xx_rsc_10_0_i_adrb,
      qa => xx_rsc_10_0_i_qa,
      wea => xx_rsc_10_0_wea,
      da => xx_rsc_10_0_i_da,
      adra => xx_rsc_10_0_i_adra,
      adra_d => xx_rsc_10_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_10_0_i_clka_en_d,
      clkb_en_d => xx_rsc_10_0_i_clka_en_d,
      da_d => xx_rsc_10_0_i_da_d,
      qa_d => xx_rsc_10_0_i_qa_d_1,
      wea_d => xx_rsc_10_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_10_0_i_qb <= xx_rsc_10_0_qb;
  xx_rsc_10_0_db <= xx_rsc_10_0_i_db;
  xx_rsc_10_0_adrb <= xx_rsc_10_0_i_adrb;
  xx_rsc_10_0_i_qa <= xx_rsc_10_0_qa;
  xx_rsc_10_0_da <= xx_rsc_10_0_i_da;
  xx_rsc_10_0_adra <= xx_rsc_10_0_i_adra;
  xx_rsc_10_0_i_adra_d_1 <= xx_rsc_10_0_i_adra_d;
  xx_rsc_10_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_10_0_i_qa_d <= xx_rsc_10_0_i_qa_d_1;
  xx_rsc_10_0_i_wea_d_1 <= xx_rsc_10_0_i_wea_d;
  xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_11_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_11_0_clkb_en,
      clka_en => xx_rsc_11_0_clka_en,
      qb => xx_rsc_11_0_i_qb,
      web => xx_rsc_11_0_web,
      db => xx_rsc_11_0_i_db,
      adrb => xx_rsc_11_0_i_adrb,
      qa => xx_rsc_11_0_i_qa,
      wea => xx_rsc_11_0_wea,
      da => xx_rsc_11_0_i_da,
      adra => xx_rsc_11_0_i_adra,
      adra_d => xx_rsc_11_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_11_0_i_clka_en_d,
      clkb_en_d => xx_rsc_11_0_i_clka_en_d,
      da_d => xx_rsc_11_0_i_da_d,
      qa_d => xx_rsc_11_0_i_qa_d_1,
      wea_d => xx_rsc_11_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_11_0_i_qb <= xx_rsc_11_0_qb;
  xx_rsc_11_0_db <= xx_rsc_11_0_i_db;
  xx_rsc_11_0_adrb <= xx_rsc_11_0_i_adrb;
  xx_rsc_11_0_i_qa <= xx_rsc_11_0_qa;
  xx_rsc_11_0_da <= xx_rsc_11_0_i_da;
  xx_rsc_11_0_adra <= xx_rsc_11_0_i_adra;
  xx_rsc_11_0_i_adra_d_1 <= xx_rsc_11_0_i_adra_d;
  xx_rsc_11_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_11_0_i_qa_d <= xx_rsc_11_0_i_qa_d_1;
  xx_rsc_11_0_i_wea_d_1 <= xx_rsc_11_0_i_wea_d;
  xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_12_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_12_0_clkb_en,
      clka_en => xx_rsc_12_0_clka_en,
      qb => xx_rsc_12_0_i_qb,
      web => xx_rsc_12_0_web,
      db => xx_rsc_12_0_i_db,
      adrb => xx_rsc_12_0_i_adrb,
      qa => xx_rsc_12_0_i_qa,
      wea => xx_rsc_12_0_wea,
      da => xx_rsc_12_0_i_da,
      adra => xx_rsc_12_0_i_adra,
      adra_d => xx_rsc_12_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_12_0_i_clka_en_d,
      clkb_en_d => xx_rsc_12_0_i_clka_en_d,
      da_d => xx_rsc_12_0_i_da_d,
      qa_d => xx_rsc_12_0_i_qa_d_1,
      wea_d => xx_rsc_12_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_12_0_i_qb <= xx_rsc_12_0_qb;
  xx_rsc_12_0_db <= xx_rsc_12_0_i_db;
  xx_rsc_12_0_adrb <= xx_rsc_12_0_i_adrb;
  xx_rsc_12_0_i_qa <= xx_rsc_12_0_qa;
  xx_rsc_12_0_da <= xx_rsc_12_0_i_da;
  xx_rsc_12_0_adra <= xx_rsc_12_0_i_adra;
  xx_rsc_12_0_i_adra_d_1 <= xx_rsc_12_0_i_adra_d;
  xx_rsc_12_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_12_0_i_qa_d <= xx_rsc_12_0_i_qa_d_1;
  xx_rsc_12_0_i_wea_d_1 <= xx_rsc_12_0_i_wea_d;
  xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_13_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_13_0_clkb_en,
      clka_en => xx_rsc_13_0_clka_en,
      qb => xx_rsc_13_0_i_qb,
      web => xx_rsc_13_0_web,
      db => xx_rsc_13_0_i_db,
      adrb => xx_rsc_13_0_i_adrb,
      qa => xx_rsc_13_0_i_qa,
      wea => xx_rsc_13_0_wea,
      da => xx_rsc_13_0_i_da,
      adra => xx_rsc_13_0_i_adra,
      adra_d => xx_rsc_13_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_13_0_i_clka_en_d,
      clkb_en_d => xx_rsc_13_0_i_clka_en_d,
      da_d => xx_rsc_13_0_i_da_d,
      qa_d => xx_rsc_13_0_i_qa_d_1,
      wea_d => xx_rsc_13_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_13_0_i_qb <= xx_rsc_13_0_qb;
  xx_rsc_13_0_db <= xx_rsc_13_0_i_db;
  xx_rsc_13_0_adrb <= xx_rsc_13_0_i_adrb;
  xx_rsc_13_0_i_qa <= xx_rsc_13_0_qa;
  xx_rsc_13_0_da <= xx_rsc_13_0_i_da;
  xx_rsc_13_0_adra <= xx_rsc_13_0_i_adra;
  xx_rsc_13_0_i_adra_d_1 <= xx_rsc_13_0_i_adra_d;
  xx_rsc_13_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_13_0_i_qa_d <= xx_rsc_13_0_i_qa_d_1;
  xx_rsc_13_0_i_wea_d_1 <= xx_rsc_13_0_i_wea_d;
  xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_14_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_14_0_clkb_en,
      clka_en => xx_rsc_14_0_clka_en,
      qb => xx_rsc_14_0_i_qb,
      web => xx_rsc_14_0_web,
      db => xx_rsc_14_0_i_db,
      adrb => xx_rsc_14_0_i_adrb,
      qa => xx_rsc_14_0_i_qa,
      wea => xx_rsc_14_0_wea,
      da => xx_rsc_14_0_i_da,
      adra => xx_rsc_14_0_i_adra,
      adra_d => xx_rsc_14_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_14_0_i_clka_en_d,
      clkb_en_d => xx_rsc_14_0_i_clka_en_d,
      da_d => xx_rsc_14_0_i_da_d,
      qa_d => xx_rsc_14_0_i_qa_d_1,
      wea_d => xx_rsc_14_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_14_0_i_qb <= xx_rsc_14_0_qb;
  xx_rsc_14_0_db <= xx_rsc_14_0_i_db;
  xx_rsc_14_0_adrb <= xx_rsc_14_0_i_adrb;
  xx_rsc_14_0_i_qa <= xx_rsc_14_0_qa;
  xx_rsc_14_0_da <= xx_rsc_14_0_i_da;
  xx_rsc_14_0_adra <= xx_rsc_14_0_i_adra;
  xx_rsc_14_0_i_adra_d_1 <= xx_rsc_14_0_i_adra_d;
  xx_rsc_14_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_14_0_i_qa_d <= xx_rsc_14_0_i_qa_d_1;
  xx_rsc_14_0_i_wea_d_1 <= xx_rsc_14_0_i_wea_d;
  xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_15_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_15_0_clkb_en,
      clka_en => xx_rsc_15_0_clka_en,
      qb => xx_rsc_15_0_i_qb,
      web => xx_rsc_15_0_web,
      db => xx_rsc_15_0_i_db,
      adrb => xx_rsc_15_0_i_adrb,
      qa => xx_rsc_15_0_i_qa,
      wea => xx_rsc_15_0_wea,
      da => xx_rsc_15_0_i_da,
      adra => xx_rsc_15_0_i_adra,
      adra_d => xx_rsc_15_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_15_0_i_clka_en_d,
      clkb_en_d => xx_rsc_15_0_i_clka_en_d,
      da_d => xx_rsc_15_0_i_da_d,
      qa_d => xx_rsc_15_0_i_qa_d_1,
      wea_d => xx_rsc_15_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_15_0_i_qb <= xx_rsc_15_0_qb;
  xx_rsc_15_0_db <= xx_rsc_15_0_i_db;
  xx_rsc_15_0_adrb <= xx_rsc_15_0_i_adrb;
  xx_rsc_15_0_i_qa <= xx_rsc_15_0_qa;
  xx_rsc_15_0_da <= xx_rsc_15_0_i_da;
  xx_rsc_15_0_adra <= xx_rsc_15_0_i_adra;
  xx_rsc_15_0_i_adra_d_1 <= xx_rsc_15_0_i_adra_d;
  xx_rsc_15_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_15_0_i_qa_d <= xx_rsc_15_0_i_qa_d_1;
  xx_rsc_15_0_i_wea_d_1 <= xx_rsc_15_0_i_wea_d;
  xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_16_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_16_0_clkb_en,
      clka_en => xx_rsc_16_0_clka_en,
      qb => xx_rsc_16_0_i_qb,
      web => xx_rsc_16_0_web,
      db => xx_rsc_16_0_i_db,
      adrb => xx_rsc_16_0_i_adrb,
      qa => xx_rsc_16_0_i_qa,
      wea => xx_rsc_16_0_wea,
      da => xx_rsc_16_0_i_da,
      adra => xx_rsc_16_0_i_adra,
      adra_d => xx_rsc_16_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_16_0_i_clka_en_d,
      clkb_en_d => xx_rsc_16_0_i_clka_en_d,
      da_d => xx_rsc_16_0_i_da_d,
      qa_d => xx_rsc_16_0_i_qa_d_1,
      wea_d => xx_rsc_16_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_16_0_i_qb <= xx_rsc_16_0_qb;
  xx_rsc_16_0_db <= xx_rsc_16_0_i_db;
  xx_rsc_16_0_adrb <= xx_rsc_16_0_i_adrb;
  xx_rsc_16_0_i_qa <= xx_rsc_16_0_qa;
  xx_rsc_16_0_da <= xx_rsc_16_0_i_da;
  xx_rsc_16_0_adra <= xx_rsc_16_0_i_adra;
  xx_rsc_16_0_i_adra_d_1 <= xx_rsc_16_0_i_adra_d;
  xx_rsc_16_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_16_0_i_qa_d <= xx_rsc_16_0_i_qa_d_1;
  xx_rsc_16_0_i_wea_d_1 <= xx_rsc_16_0_i_wea_d;
  xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_17_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_17_0_clkb_en,
      clka_en => xx_rsc_17_0_clka_en,
      qb => xx_rsc_17_0_i_qb,
      web => xx_rsc_17_0_web,
      db => xx_rsc_17_0_i_db,
      adrb => xx_rsc_17_0_i_adrb,
      qa => xx_rsc_17_0_i_qa,
      wea => xx_rsc_17_0_wea,
      da => xx_rsc_17_0_i_da,
      adra => xx_rsc_17_0_i_adra,
      adra_d => xx_rsc_17_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_17_0_i_clka_en_d,
      clkb_en_d => xx_rsc_17_0_i_clka_en_d,
      da_d => xx_rsc_17_0_i_da_d,
      qa_d => xx_rsc_17_0_i_qa_d_1,
      wea_d => xx_rsc_17_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_17_0_i_qb <= xx_rsc_17_0_qb;
  xx_rsc_17_0_db <= xx_rsc_17_0_i_db;
  xx_rsc_17_0_adrb <= xx_rsc_17_0_i_adrb;
  xx_rsc_17_0_i_qa <= xx_rsc_17_0_qa;
  xx_rsc_17_0_da <= xx_rsc_17_0_i_da;
  xx_rsc_17_0_adra <= xx_rsc_17_0_i_adra;
  xx_rsc_17_0_i_adra_d_1 <= xx_rsc_17_0_i_adra_d;
  xx_rsc_17_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_17_0_i_qa_d <= xx_rsc_17_0_i_qa_d_1;
  xx_rsc_17_0_i_wea_d_1 <= xx_rsc_17_0_i_wea_d;
  xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_18_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_18_0_clkb_en,
      clka_en => xx_rsc_18_0_clka_en,
      qb => xx_rsc_18_0_i_qb,
      web => xx_rsc_18_0_web,
      db => xx_rsc_18_0_i_db,
      adrb => xx_rsc_18_0_i_adrb,
      qa => xx_rsc_18_0_i_qa,
      wea => xx_rsc_18_0_wea,
      da => xx_rsc_18_0_i_da,
      adra => xx_rsc_18_0_i_adra,
      adra_d => xx_rsc_18_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_18_0_i_clka_en_d,
      clkb_en_d => xx_rsc_18_0_i_clka_en_d,
      da_d => xx_rsc_18_0_i_da_d,
      qa_d => xx_rsc_18_0_i_qa_d_1,
      wea_d => xx_rsc_18_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_18_0_i_qb <= xx_rsc_18_0_qb;
  xx_rsc_18_0_db <= xx_rsc_18_0_i_db;
  xx_rsc_18_0_adrb <= xx_rsc_18_0_i_adrb;
  xx_rsc_18_0_i_qa <= xx_rsc_18_0_qa;
  xx_rsc_18_0_da <= xx_rsc_18_0_i_da;
  xx_rsc_18_0_adra <= xx_rsc_18_0_i_adra;
  xx_rsc_18_0_i_adra_d_1 <= xx_rsc_18_0_i_adra_d;
  xx_rsc_18_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_18_0_i_qa_d <= xx_rsc_18_0_i_qa_d_1;
  xx_rsc_18_0_i_wea_d_1 <= xx_rsc_18_0_i_wea_d;
  xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_19_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_19_0_clkb_en,
      clka_en => xx_rsc_19_0_clka_en,
      qb => xx_rsc_19_0_i_qb,
      web => xx_rsc_19_0_web,
      db => xx_rsc_19_0_i_db,
      adrb => xx_rsc_19_0_i_adrb,
      qa => xx_rsc_19_0_i_qa,
      wea => xx_rsc_19_0_wea,
      da => xx_rsc_19_0_i_da,
      adra => xx_rsc_19_0_i_adra,
      adra_d => xx_rsc_19_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_19_0_i_clka_en_d,
      clkb_en_d => xx_rsc_19_0_i_clka_en_d,
      da_d => xx_rsc_19_0_i_da_d,
      qa_d => xx_rsc_19_0_i_qa_d_1,
      wea_d => xx_rsc_19_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_19_0_i_qb <= xx_rsc_19_0_qb;
  xx_rsc_19_0_db <= xx_rsc_19_0_i_db;
  xx_rsc_19_0_adrb <= xx_rsc_19_0_i_adrb;
  xx_rsc_19_0_i_qa <= xx_rsc_19_0_qa;
  xx_rsc_19_0_da <= xx_rsc_19_0_i_da;
  xx_rsc_19_0_adra <= xx_rsc_19_0_i_adra;
  xx_rsc_19_0_i_adra_d_1 <= xx_rsc_19_0_i_adra_d;
  xx_rsc_19_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_19_0_i_qa_d <= xx_rsc_19_0_i_qa_d_1;
  xx_rsc_19_0_i_wea_d_1 <= xx_rsc_19_0_i_wea_d;
  xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_20_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_20_0_clkb_en,
      clka_en => xx_rsc_20_0_clka_en,
      qb => xx_rsc_20_0_i_qb,
      web => xx_rsc_20_0_web,
      db => xx_rsc_20_0_i_db,
      adrb => xx_rsc_20_0_i_adrb,
      qa => xx_rsc_20_0_i_qa,
      wea => xx_rsc_20_0_wea,
      da => xx_rsc_20_0_i_da,
      adra => xx_rsc_20_0_i_adra,
      adra_d => xx_rsc_20_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_20_0_i_clka_en_d,
      clkb_en_d => xx_rsc_20_0_i_clka_en_d,
      da_d => xx_rsc_20_0_i_da_d,
      qa_d => xx_rsc_20_0_i_qa_d_1,
      wea_d => xx_rsc_20_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_20_0_i_qb <= xx_rsc_20_0_qb;
  xx_rsc_20_0_db <= xx_rsc_20_0_i_db;
  xx_rsc_20_0_adrb <= xx_rsc_20_0_i_adrb;
  xx_rsc_20_0_i_qa <= xx_rsc_20_0_qa;
  xx_rsc_20_0_da <= xx_rsc_20_0_i_da;
  xx_rsc_20_0_adra <= xx_rsc_20_0_i_adra;
  xx_rsc_20_0_i_adra_d_1 <= xx_rsc_20_0_i_adra_d;
  xx_rsc_20_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_20_0_i_qa_d <= xx_rsc_20_0_i_qa_d_1;
  xx_rsc_20_0_i_wea_d_1 <= xx_rsc_20_0_i_wea_d;
  xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_21_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_21_0_clkb_en,
      clka_en => xx_rsc_21_0_clka_en,
      qb => xx_rsc_21_0_i_qb,
      web => xx_rsc_21_0_web,
      db => xx_rsc_21_0_i_db,
      adrb => xx_rsc_21_0_i_adrb,
      qa => xx_rsc_21_0_i_qa,
      wea => xx_rsc_21_0_wea,
      da => xx_rsc_21_0_i_da,
      adra => xx_rsc_21_0_i_adra,
      adra_d => xx_rsc_21_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_21_0_i_clka_en_d,
      clkb_en_d => xx_rsc_21_0_i_clka_en_d,
      da_d => xx_rsc_21_0_i_da_d,
      qa_d => xx_rsc_21_0_i_qa_d_1,
      wea_d => xx_rsc_21_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_21_0_i_qb <= xx_rsc_21_0_qb;
  xx_rsc_21_0_db <= xx_rsc_21_0_i_db;
  xx_rsc_21_0_adrb <= xx_rsc_21_0_i_adrb;
  xx_rsc_21_0_i_qa <= xx_rsc_21_0_qa;
  xx_rsc_21_0_da <= xx_rsc_21_0_i_da;
  xx_rsc_21_0_adra <= xx_rsc_21_0_i_adra;
  xx_rsc_21_0_i_adra_d_1 <= xx_rsc_21_0_i_adra_d;
  xx_rsc_21_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_21_0_i_qa_d <= xx_rsc_21_0_i_qa_d_1;
  xx_rsc_21_0_i_wea_d_1 <= xx_rsc_21_0_i_wea_d;
  xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_22_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_22_0_clkb_en,
      clka_en => xx_rsc_22_0_clka_en,
      qb => xx_rsc_22_0_i_qb,
      web => xx_rsc_22_0_web,
      db => xx_rsc_22_0_i_db,
      adrb => xx_rsc_22_0_i_adrb,
      qa => xx_rsc_22_0_i_qa,
      wea => xx_rsc_22_0_wea,
      da => xx_rsc_22_0_i_da,
      adra => xx_rsc_22_0_i_adra,
      adra_d => xx_rsc_22_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_22_0_i_clka_en_d,
      clkb_en_d => xx_rsc_22_0_i_clka_en_d,
      da_d => xx_rsc_22_0_i_da_d,
      qa_d => xx_rsc_22_0_i_qa_d_1,
      wea_d => xx_rsc_22_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_22_0_i_qb <= xx_rsc_22_0_qb;
  xx_rsc_22_0_db <= xx_rsc_22_0_i_db;
  xx_rsc_22_0_adrb <= xx_rsc_22_0_i_adrb;
  xx_rsc_22_0_i_qa <= xx_rsc_22_0_qa;
  xx_rsc_22_0_da <= xx_rsc_22_0_i_da;
  xx_rsc_22_0_adra <= xx_rsc_22_0_i_adra;
  xx_rsc_22_0_i_adra_d_1 <= xx_rsc_22_0_i_adra_d;
  xx_rsc_22_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_22_0_i_qa_d <= xx_rsc_22_0_i_qa_d_1;
  xx_rsc_22_0_i_wea_d_1 <= xx_rsc_22_0_i_wea_d;
  xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_23_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_23_0_clkb_en,
      clka_en => xx_rsc_23_0_clka_en,
      qb => xx_rsc_23_0_i_qb,
      web => xx_rsc_23_0_web,
      db => xx_rsc_23_0_i_db,
      adrb => xx_rsc_23_0_i_adrb,
      qa => xx_rsc_23_0_i_qa,
      wea => xx_rsc_23_0_wea,
      da => xx_rsc_23_0_i_da,
      adra => xx_rsc_23_0_i_adra,
      adra_d => xx_rsc_23_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_23_0_i_clka_en_d,
      clkb_en_d => xx_rsc_23_0_i_clka_en_d,
      da_d => xx_rsc_23_0_i_da_d,
      qa_d => xx_rsc_23_0_i_qa_d_1,
      wea_d => xx_rsc_23_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_23_0_i_qb <= xx_rsc_23_0_qb;
  xx_rsc_23_0_db <= xx_rsc_23_0_i_db;
  xx_rsc_23_0_adrb <= xx_rsc_23_0_i_adrb;
  xx_rsc_23_0_i_qa <= xx_rsc_23_0_qa;
  xx_rsc_23_0_da <= xx_rsc_23_0_i_da;
  xx_rsc_23_0_adra <= xx_rsc_23_0_i_adra;
  xx_rsc_23_0_i_adra_d_1 <= xx_rsc_23_0_i_adra_d;
  xx_rsc_23_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_23_0_i_qa_d <= xx_rsc_23_0_i_qa_d_1;
  xx_rsc_23_0_i_wea_d_1 <= xx_rsc_23_0_i_wea_d;
  xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_24_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_24_0_clkb_en,
      clka_en => xx_rsc_24_0_clka_en,
      qb => xx_rsc_24_0_i_qb,
      web => xx_rsc_24_0_web,
      db => xx_rsc_24_0_i_db,
      adrb => xx_rsc_24_0_i_adrb,
      qa => xx_rsc_24_0_i_qa,
      wea => xx_rsc_24_0_wea,
      da => xx_rsc_24_0_i_da,
      adra => xx_rsc_24_0_i_adra,
      adra_d => xx_rsc_24_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_24_0_i_clka_en_d,
      clkb_en_d => xx_rsc_24_0_i_clka_en_d,
      da_d => xx_rsc_24_0_i_da_d,
      qa_d => xx_rsc_24_0_i_qa_d_1,
      wea_d => xx_rsc_24_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_24_0_i_qb <= xx_rsc_24_0_qb;
  xx_rsc_24_0_db <= xx_rsc_24_0_i_db;
  xx_rsc_24_0_adrb <= xx_rsc_24_0_i_adrb;
  xx_rsc_24_0_i_qa <= xx_rsc_24_0_qa;
  xx_rsc_24_0_da <= xx_rsc_24_0_i_da;
  xx_rsc_24_0_adra <= xx_rsc_24_0_i_adra;
  xx_rsc_24_0_i_adra_d_1 <= xx_rsc_24_0_i_adra_d;
  xx_rsc_24_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_24_0_i_qa_d <= xx_rsc_24_0_i_qa_d_1;
  xx_rsc_24_0_i_wea_d_1 <= xx_rsc_24_0_i_wea_d;
  xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_25_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_25_0_clkb_en,
      clka_en => xx_rsc_25_0_clka_en,
      qb => xx_rsc_25_0_i_qb,
      web => xx_rsc_25_0_web,
      db => xx_rsc_25_0_i_db,
      adrb => xx_rsc_25_0_i_adrb,
      qa => xx_rsc_25_0_i_qa,
      wea => xx_rsc_25_0_wea,
      da => xx_rsc_25_0_i_da,
      adra => xx_rsc_25_0_i_adra,
      adra_d => xx_rsc_25_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_25_0_i_clka_en_d,
      clkb_en_d => xx_rsc_25_0_i_clka_en_d,
      da_d => xx_rsc_25_0_i_da_d,
      qa_d => xx_rsc_25_0_i_qa_d_1,
      wea_d => xx_rsc_25_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_25_0_i_qb <= xx_rsc_25_0_qb;
  xx_rsc_25_0_db <= xx_rsc_25_0_i_db;
  xx_rsc_25_0_adrb <= xx_rsc_25_0_i_adrb;
  xx_rsc_25_0_i_qa <= xx_rsc_25_0_qa;
  xx_rsc_25_0_da <= xx_rsc_25_0_i_da;
  xx_rsc_25_0_adra <= xx_rsc_25_0_i_adra;
  xx_rsc_25_0_i_adra_d_1 <= xx_rsc_25_0_i_adra_d;
  xx_rsc_25_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_25_0_i_qa_d <= xx_rsc_25_0_i_qa_d_1;
  xx_rsc_25_0_i_wea_d_1 <= xx_rsc_25_0_i_wea_d;
  xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_26_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_26_0_clkb_en,
      clka_en => xx_rsc_26_0_clka_en,
      qb => xx_rsc_26_0_i_qb,
      web => xx_rsc_26_0_web,
      db => xx_rsc_26_0_i_db,
      adrb => xx_rsc_26_0_i_adrb,
      qa => xx_rsc_26_0_i_qa,
      wea => xx_rsc_26_0_wea,
      da => xx_rsc_26_0_i_da,
      adra => xx_rsc_26_0_i_adra,
      adra_d => xx_rsc_26_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_26_0_i_clka_en_d,
      clkb_en_d => xx_rsc_26_0_i_clka_en_d,
      da_d => xx_rsc_26_0_i_da_d,
      qa_d => xx_rsc_26_0_i_qa_d_1,
      wea_d => xx_rsc_26_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_26_0_i_qb <= xx_rsc_26_0_qb;
  xx_rsc_26_0_db <= xx_rsc_26_0_i_db;
  xx_rsc_26_0_adrb <= xx_rsc_26_0_i_adrb;
  xx_rsc_26_0_i_qa <= xx_rsc_26_0_qa;
  xx_rsc_26_0_da <= xx_rsc_26_0_i_da;
  xx_rsc_26_0_adra <= xx_rsc_26_0_i_adra;
  xx_rsc_26_0_i_adra_d_1 <= xx_rsc_26_0_i_adra_d;
  xx_rsc_26_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_26_0_i_qa_d <= xx_rsc_26_0_i_qa_d_1;
  xx_rsc_26_0_i_wea_d_1 <= xx_rsc_26_0_i_wea_d;
  xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_27_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_27_0_clkb_en,
      clka_en => xx_rsc_27_0_clka_en,
      qb => xx_rsc_27_0_i_qb,
      web => xx_rsc_27_0_web,
      db => xx_rsc_27_0_i_db,
      adrb => xx_rsc_27_0_i_adrb,
      qa => xx_rsc_27_0_i_qa,
      wea => xx_rsc_27_0_wea,
      da => xx_rsc_27_0_i_da,
      adra => xx_rsc_27_0_i_adra,
      adra_d => xx_rsc_27_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_27_0_i_clka_en_d,
      clkb_en_d => xx_rsc_27_0_i_clka_en_d,
      da_d => xx_rsc_27_0_i_da_d,
      qa_d => xx_rsc_27_0_i_qa_d_1,
      wea_d => xx_rsc_27_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_27_0_i_qb <= xx_rsc_27_0_qb;
  xx_rsc_27_0_db <= xx_rsc_27_0_i_db;
  xx_rsc_27_0_adrb <= xx_rsc_27_0_i_adrb;
  xx_rsc_27_0_i_qa <= xx_rsc_27_0_qa;
  xx_rsc_27_0_da <= xx_rsc_27_0_i_da;
  xx_rsc_27_0_adra <= xx_rsc_27_0_i_adra;
  xx_rsc_27_0_i_adra_d_1 <= xx_rsc_27_0_i_adra_d;
  xx_rsc_27_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_27_0_i_qa_d <= xx_rsc_27_0_i_qa_d_1;
  xx_rsc_27_0_i_wea_d_1 <= xx_rsc_27_0_i_wea_d;
  xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_28_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_28_0_clkb_en,
      clka_en => xx_rsc_28_0_clka_en,
      qb => xx_rsc_28_0_i_qb,
      web => xx_rsc_28_0_web,
      db => xx_rsc_28_0_i_db,
      adrb => xx_rsc_28_0_i_adrb,
      qa => xx_rsc_28_0_i_qa,
      wea => xx_rsc_28_0_wea,
      da => xx_rsc_28_0_i_da,
      adra => xx_rsc_28_0_i_adra,
      adra_d => xx_rsc_28_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_28_0_i_clka_en_d,
      clkb_en_d => xx_rsc_28_0_i_clka_en_d,
      da_d => xx_rsc_28_0_i_da_d,
      qa_d => xx_rsc_28_0_i_qa_d_1,
      wea_d => xx_rsc_28_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_28_0_i_qb <= xx_rsc_28_0_qb;
  xx_rsc_28_0_db <= xx_rsc_28_0_i_db;
  xx_rsc_28_0_adrb <= xx_rsc_28_0_i_adrb;
  xx_rsc_28_0_i_qa <= xx_rsc_28_0_qa;
  xx_rsc_28_0_da <= xx_rsc_28_0_i_da;
  xx_rsc_28_0_adra <= xx_rsc_28_0_i_adra;
  xx_rsc_28_0_i_adra_d_1 <= xx_rsc_28_0_i_adra_d;
  xx_rsc_28_0_i_da_d <= xx_rsc_0_0_i_da_d_iff;
  xx_rsc_28_0_i_qa_d <= xx_rsc_28_0_i_qa_d_1;
  xx_rsc_28_0_i_wea_d_1 <= xx_rsc_28_0_i_wea_d;
  xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_29_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_39_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_29_0_clkb_en,
      clka_en => xx_rsc_29_0_clka_en,
      qb => xx_rsc_29_0_i_qb,
      web => xx_rsc_29_0_web,
      db => xx_rsc_29_0_i_db,
      adrb => xx_rsc_29_0_i_adrb,
      qa => xx_rsc_29_0_i_qa,
      wea => xx_rsc_29_0_wea,
      da => xx_rsc_29_0_i_da,
      adra => xx_rsc_29_0_i_adra,
      adra_d => xx_rsc_29_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_29_0_i_clka_en_d,
      clkb_en_d => xx_rsc_29_0_i_clka_en_d,
      da_d => xx_rsc_29_0_i_da_d,
      qa_d => xx_rsc_29_0_i_qa_d_1,
      wea_d => xx_rsc_29_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_29_0_i_qb <= xx_rsc_29_0_qb;
  xx_rsc_29_0_db <= xx_rsc_29_0_i_db;
  xx_rsc_29_0_adrb <= xx_rsc_29_0_i_adrb;
  xx_rsc_29_0_i_qa <= xx_rsc_29_0_qa;
  xx_rsc_29_0_da <= xx_rsc_29_0_i_da;
  xx_rsc_29_0_adra <= xx_rsc_29_0_i_adra;
  xx_rsc_29_0_i_adra_d_1 <= xx_rsc_29_0_i_adra_d;
  xx_rsc_29_0_i_da_d <= xx_rsc_1_0_i_da_d_iff;
  xx_rsc_29_0_i_qa_d <= xx_rsc_29_0_i_qa_d_1;
  xx_rsc_29_0_i_wea_d_1 <= xx_rsc_29_0_i_wea_d;
  xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_30_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_40_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_30_0_clkb_en,
      clka_en => xx_rsc_30_0_clka_en,
      qb => xx_rsc_30_0_i_qb,
      web => xx_rsc_30_0_web,
      db => xx_rsc_30_0_i_db,
      adrb => xx_rsc_30_0_i_adrb,
      qa => xx_rsc_30_0_i_qa,
      wea => xx_rsc_30_0_wea,
      da => xx_rsc_30_0_i_da,
      adra => xx_rsc_30_0_i_adra,
      adra_d => xx_rsc_30_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_30_0_i_clka_en_d,
      clkb_en_d => xx_rsc_30_0_i_clka_en_d,
      da_d => xx_rsc_30_0_i_da_d,
      qa_d => xx_rsc_30_0_i_qa_d_1,
      wea_d => xx_rsc_30_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_30_0_i_qb <= xx_rsc_30_0_qb;
  xx_rsc_30_0_db <= xx_rsc_30_0_i_db;
  xx_rsc_30_0_adrb <= xx_rsc_30_0_i_adrb;
  xx_rsc_30_0_i_qa <= xx_rsc_30_0_qa;
  xx_rsc_30_0_da <= xx_rsc_30_0_i_da;
  xx_rsc_30_0_adra <= xx_rsc_30_0_i_adra;
  xx_rsc_30_0_i_adra_d_1 <= xx_rsc_30_0_i_adra_d;
  xx_rsc_30_0_i_da_d <= xx_rsc_2_0_i_da_d_iff;
  xx_rsc_30_0_i_qa_d <= xx_rsc_30_0_i_qa_d_1;
  xx_rsc_30_0_i_wea_d_1 <= xx_rsc_30_0_i_wea_d;
  xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  xx_rsc_31_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_41_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => xx_rsc_31_0_clkb_en,
      clka_en => xx_rsc_31_0_clka_en,
      qb => xx_rsc_31_0_i_qb,
      web => xx_rsc_31_0_web,
      db => xx_rsc_31_0_i_db,
      adrb => xx_rsc_31_0_i_adrb,
      qa => xx_rsc_31_0_i_qa,
      wea => xx_rsc_31_0_wea,
      da => xx_rsc_31_0_i_da,
      adra => xx_rsc_31_0_i_adra,
      adra_d => xx_rsc_31_0_i_adra_d_1,
      clka => clk,
      clka_en_d => xx_rsc_31_0_i_clka_en_d,
      clkb_en_d => xx_rsc_31_0_i_clka_en_d,
      da_d => xx_rsc_31_0_i_da_d,
      qa_d => xx_rsc_31_0_i_qa_d_1,
      wea_d => xx_rsc_31_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  xx_rsc_31_0_i_qb <= xx_rsc_31_0_qb;
  xx_rsc_31_0_db <= xx_rsc_31_0_i_db;
  xx_rsc_31_0_adrb <= xx_rsc_31_0_i_adrb;
  xx_rsc_31_0_i_qa <= xx_rsc_31_0_qa;
  xx_rsc_31_0_da <= xx_rsc_31_0_i_da;
  xx_rsc_31_0_adra <= xx_rsc_31_0_i_adra;
  xx_rsc_31_0_i_adra_d_1 <= xx_rsc_31_0_i_adra_d;
  xx_rsc_31_0_i_da_d <= xx_rsc_3_0_i_da_d_iff;
  xx_rsc_31_0_i_qa_d <= xx_rsc_31_0_i_qa_d_1;
  xx_rsc_31_0_i_wea_d_1 <= xx_rsc_31_0_i_wea_d;
  xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_0_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_42_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_0_0_clkb_en,
      clka_en => yy_rsc_0_0_clka_en,
      qb => yy_rsc_0_0_i_qb,
      web => yy_rsc_0_0_web,
      db => yy_rsc_0_0_i_db,
      adrb => yy_rsc_0_0_i_adrb,
      qa => yy_rsc_0_0_i_qa,
      wea => yy_rsc_0_0_wea,
      da => yy_rsc_0_0_i_da,
      adra => yy_rsc_0_0_i_adra,
      adra_d => yy_rsc_0_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_0_0_i_clka_en_d,
      clkb_en_d => yy_rsc_0_0_i_clka_en_d,
      da_d => yy_rsc_0_0_i_da_d,
      qa_d => yy_rsc_0_0_i_qa_d_1,
      wea_d => yy_rsc_0_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_0_0_i_qb <= yy_rsc_0_0_qb;
  yy_rsc_0_0_db <= yy_rsc_0_0_i_db;
  yy_rsc_0_0_adrb <= yy_rsc_0_0_i_adrb;
  yy_rsc_0_0_i_qa <= yy_rsc_0_0_qa;
  yy_rsc_0_0_da <= yy_rsc_0_0_i_da;
  yy_rsc_0_0_adra <= yy_rsc_0_0_i_adra;
  yy_rsc_0_0_i_adra_d_1 <= yy_rsc_0_0_i_adra_d;
  yy_rsc_0_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_0_0_i_qa_d <= yy_rsc_0_0_i_qa_d_1;
  yy_rsc_0_0_i_wea_d_1 <= yy_rsc_0_0_i_wea_d;
  yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_1_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_43_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_1_0_clkb_en,
      clka_en => yy_rsc_1_0_clka_en,
      qb => yy_rsc_1_0_i_qb,
      web => yy_rsc_1_0_web,
      db => yy_rsc_1_0_i_db,
      adrb => yy_rsc_1_0_i_adrb,
      qa => yy_rsc_1_0_i_qa,
      wea => yy_rsc_1_0_wea,
      da => yy_rsc_1_0_i_da,
      adra => yy_rsc_1_0_i_adra,
      adra_d => yy_rsc_1_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_1_0_i_clka_en_d,
      clkb_en_d => yy_rsc_1_0_i_clka_en_d,
      da_d => yy_rsc_1_0_i_da_d,
      qa_d => yy_rsc_1_0_i_qa_d_1,
      wea_d => yy_rsc_1_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_1_0_i_qb <= yy_rsc_1_0_qb;
  yy_rsc_1_0_db <= yy_rsc_1_0_i_db;
  yy_rsc_1_0_adrb <= yy_rsc_1_0_i_adrb;
  yy_rsc_1_0_i_qa <= yy_rsc_1_0_qa;
  yy_rsc_1_0_da <= yy_rsc_1_0_i_da;
  yy_rsc_1_0_adra <= yy_rsc_1_0_i_adra;
  yy_rsc_1_0_i_adra_d_1 <= yy_rsc_1_0_i_adra_d;
  yy_rsc_1_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_1_0_i_qa_d <= yy_rsc_1_0_i_qa_d_1;
  yy_rsc_1_0_i_wea_d_1 <= yy_rsc_1_0_i_wea_d;
  yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_2_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_44_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_2_0_clkb_en,
      clka_en => yy_rsc_2_0_clka_en,
      qb => yy_rsc_2_0_i_qb,
      web => yy_rsc_2_0_web,
      db => yy_rsc_2_0_i_db,
      adrb => yy_rsc_2_0_i_adrb,
      qa => yy_rsc_2_0_i_qa,
      wea => yy_rsc_2_0_wea,
      da => yy_rsc_2_0_i_da,
      adra => yy_rsc_2_0_i_adra,
      adra_d => yy_rsc_2_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_2_0_i_clka_en_d,
      clkb_en_d => yy_rsc_2_0_i_clka_en_d,
      da_d => yy_rsc_2_0_i_da_d,
      qa_d => yy_rsc_2_0_i_qa_d_1,
      wea_d => yy_rsc_2_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_2_0_i_qb <= yy_rsc_2_0_qb;
  yy_rsc_2_0_db <= yy_rsc_2_0_i_db;
  yy_rsc_2_0_adrb <= yy_rsc_2_0_i_adrb;
  yy_rsc_2_0_i_qa <= yy_rsc_2_0_qa;
  yy_rsc_2_0_da <= yy_rsc_2_0_i_da;
  yy_rsc_2_0_adra <= yy_rsc_2_0_i_adra;
  yy_rsc_2_0_i_adra_d_1 <= yy_rsc_2_0_i_adra_d;
  yy_rsc_2_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_2_0_i_qa_d <= yy_rsc_2_0_i_qa_d_1;
  yy_rsc_2_0_i_wea_d_1 <= yy_rsc_2_0_i_wea_d;
  yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_3_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_45_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_3_0_clkb_en,
      clka_en => yy_rsc_3_0_clka_en,
      qb => yy_rsc_3_0_i_qb,
      web => yy_rsc_3_0_web,
      db => yy_rsc_3_0_i_db,
      adrb => yy_rsc_3_0_i_adrb,
      qa => yy_rsc_3_0_i_qa,
      wea => yy_rsc_3_0_wea,
      da => yy_rsc_3_0_i_da,
      adra => yy_rsc_3_0_i_adra,
      adra_d => yy_rsc_3_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_3_0_i_clka_en_d,
      clkb_en_d => yy_rsc_3_0_i_clka_en_d,
      da_d => yy_rsc_3_0_i_da_d,
      qa_d => yy_rsc_3_0_i_qa_d_1,
      wea_d => yy_rsc_3_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_3_0_i_qb <= yy_rsc_3_0_qb;
  yy_rsc_3_0_db <= yy_rsc_3_0_i_db;
  yy_rsc_3_0_adrb <= yy_rsc_3_0_i_adrb;
  yy_rsc_3_0_i_qa <= yy_rsc_3_0_qa;
  yy_rsc_3_0_da <= yy_rsc_3_0_i_da;
  yy_rsc_3_0_adra <= yy_rsc_3_0_i_adra;
  yy_rsc_3_0_i_adra_d_1 <= yy_rsc_3_0_i_adra_d;
  yy_rsc_3_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_3_0_i_qa_d <= yy_rsc_3_0_i_qa_d_1;
  yy_rsc_3_0_i_wea_d_1 <= yy_rsc_3_0_i_wea_d;
  yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_4_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_46_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_4_0_clkb_en,
      clka_en => yy_rsc_4_0_clka_en,
      qb => yy_rsc_4_0_i_qb,
      web => yy_rsc_4_0_web,
      db => yy_rsc_4_0_i_db,
      adrb => yy_rsc_4_0_i_adrb,
      qa => yy_rsc_4_0_i_qa,
      wea => yy_rsc_4_0_wea,
      da => yy_rsc_4_0_i_da,
      adra => yy_rsc_4_0_i_adra,
      adra_d => yy_rsc_4_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_4_0_i_clka_en_d,
      clkb_en_d => yy_rsc_4_0_i_clka_en_d,
      da_d => yy_rsc_4_0_i_da_d,
      qa_d => yy_rsc_4_0_i_qa_d_1,
      wea_d => yy_rsc_4_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_4_0_i_qb <= yy_rsc_4_0_qb;
  yy_rsc_4_0_db <= yy_rsc_4_0_i_db;
  yy_rsc_4_0_adrb <= yy_rsc_4_0_i_adrb;
  yy_rsc_4_0_i_qa <= yy_rsc_4_0_qa;
  yy_rsc_4_0_da <= yy_rsc_4_0_i_da;
  yy_rsc_4_0_adra <= yy_rsc_4_0_i_adra;
  yy_rsc_4_0_i_adra_d_1 <= yy_rsc_4_0_i_adra_d;
  yy_rsc_4_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_4_0_i_qa_d <= yy_rsc_4_0_i_qa_d_1;
  yy_rsc_4_0_i_wea_d_1 <= yy_rsc_4_0_i_wea_d;
  yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_5_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_47_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_5_0_clkb_en,
      clka_en => yy_rsc_5_0_clka_en,
      qb => yy_rsc_5_0_i_qb,
      web => yy_rsc_5_0_web,
      db => yy_rsc_5_0_i_db,
      adrb => yy_rsc_5_0_i_adrb,
      qa => yy_rsc_5_0_i_qa,
      wea => yy_rsc_5_0_wea,
      da => yy_rsc_5_0_i_da,
      adra => yy_rsc_5_0_i_adra,
      adra_d => yy_rsc_5_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_5_0_i_clka_en_d,
      clkb_en_d => yy_rsc_5_0_i_clka_en_d,
      da_d => yy_rsc_5_0_i_da_d,
      qa_d => yy_rsc_5_0_i_qa_d_1,
      wea_d => yy_rsc_5_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_5_0_i_qb <= yy_rsc_5_0_qb;
  yy_rsc_5_0_db <= yy_rsc_5_0_i_db;
  yy_rsc_5_0_adrb <= yy_rsc_5_0_i_adrb;
  yy_rsc_5_0_i_qa <= yy_rsc_5_0_qa;
  yy_rsc_5_0_da <= yy_rsc_5_0_i_da;
  yy_rsc_5_0_adra <= yy_rsc_5_0_i_adra;
  yy_rsc_5_0_i_adra_d_1 <= yy_rsc_5_0_i_adra_d;
  yy_rsc_5_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_5_0_i_qa_d <= yy_rsc_5_0_i_qa_d_1;
  yy_rsc_5_0_i_wea_d_1 <= yy_rsc_5_0_i_wea_d;
  yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_6_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_48_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_6_0_clkb_en,
      clka_en => yy_rsc_6_0_clka_en,
      qb => yy_rsc_6_0_i_qb,
      web => yy_rsc_6_0_web,
      db => yy_rsc_6_0_i_db,
      adrb => yy_rsc_6_0_i_adrb,
      qa => yy_rsc_6_0_i_qa,
      wea => yy_rsc_6_0_wea,
      da => yy_rsc_6_0_i_da,
      adra => yy_rsc_6_0_i_adra,
      adra_d => yy_rsc_6_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_6_0_i_clka_en_d,
      clkb_en_d => yy_rsc_6_0_i_clka_en_d,
      da_d => yy_rsc_6_0_i_da_d,
      qa_d => yy_rsc_6_0_i_qa_d_1,
      wea_d => yy_rsc_6_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_6_0_i_qb <= yy_rsc_6_0_qb;
  yy_rsc_6_0_db <= yy_rsc_6_0_i_db;
  yy_rsc_6_0_adrb <= yy_rsc_6_0_i_adrb;
  yy_rsc_6_0_i_qa <= yy_rsc_6_0_qa;
  yy_rsc_6_0_da <= yy_rsc_6_0_i_da;
  yy_rsc_6_0_adra <= yy_rsc_6_0_i_adra;
  yy_rsc_6_0_i_adra_d_1 <= yy_rsc_6_0_i_adra_d;
  yy_rsc_6_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_6_0_i_qa_d <= yy_rsc_6_0_i_qa_d_1;
  yy_rsc_6_0_i_wea_d_1 <= yy_rsc_6_0_i_wea_d;
  yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_7_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_49_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_7_0_clkb_en,
      clka_en => yy_rsc_7_0_clka_en,
      qb => yy_rsc_7_0_i_qb,
      web => yy_rsc_7_0_web,
      db => yy_rsc_7_0_i_db,
      adrb => yy_rsc_7_0_i_adrb,
      qa => yy_rsc_7_0_i_qa,
      wea => yy_rsc_7_0_wea,
      da => yy_rsc_7_0_i_da,
      adra => yy_rsc_7_0_i_adra,
      adra_d => yy_rsc_7_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_7_0_i_clka_en_d,
      clkb_en_d => yy_rsc_7_0_i_clka_en_d,
      da_d => yy_rsc_7_0_i_da_d,
      qa_d => yy_rsc_7_0_i_qa_d_1,
      wea_d => yy_rsc_7_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_7_0_i_qb <= yy_rsc_7_0_qb;
  yy_rsc_7_0_db <= yy_rsc_7_0_i_db;
  yy_rsc_7_0_adrb <= yy_rsc_7_0_i_adrb;
  yy_rsc_7_0_i_qa <= yy_rsc_7_0_qa;
  yy_rsc_7_0_da <= yy_rsc_7_0_i_da;
  yy_rsc_7_0_adra <= yy_rsc_7_0_i_adra;
  yy_rsc_7_0_i_adra_d_1 <= yy_rsc_7_0_i_adra_d;
  yy_rsc_7_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_7_0_i_qa_d <= yy_rsc_7_0_i_qa_d_1;
  yy_rsc_7_0_i_wea_d_1 <= yy_rsc_7_0_i_wea_d;
  yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_8_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_50_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_8_0_clkb_en,
      clka_en => yy_rsc_8_0_clka_en,
      qb => yy_rsc_8_0_i_qb,
      web => yy_rsc_8_0_web,
      db => yy_rsc_8_0_i_db,
      adrb => yy_rsc_8_0_i_adrb,
      qa => yy_rsc_8_0_i_qa,
      wea => yy_rsc_8_0_wea,
      da => yy_rsc_8_0_i_da,
      adra => yy_rsc_8_0_i_adra,
      adra_d => yy_rsc_8_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_8_0_i_clka_en_d,
      clkb_en_d => yy_rsc_8_0_i_clka_en_d,
      da_d => yy_rsc_8_0_i_da_d,
      qa_d => yy_rsc_8_0_i_qa_d_1,
      wea_d => yy_rsc_8_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_8_0_i_qb <= yy_rsc_8_0_qb;
  yy_rsc_8_0_db <= yy_rsc_8_0_i_db;
  yy_rsc_8_0_adrb <= yy_rsc_8_0_i_adrb;
  yy_rsc_8_0_i_qa <= yy_rsc_8_0_qa;
  yy_rsc_8_0_da <= yy_rsc_8_0_i_da;
  yy_rsc_8_0_adra <= yy_rsc_8_0_i_adra;
  yy_rsc_8_0_i_adra_d_1 <= yy_rsc_8_0_i_adra_d;
  yy_rsc_8_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_8_0_i_qa_d <= yy_rsc_8_0_i_qa_d_1;
  yy_rsc_8_0_i_wea_d_1 <= yy_rsc_8_0_i_wea_d;
  yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_9_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_51_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_9_0_clkb_en,
      clka_en => yy_rsc_9_0_clka_en,
      qb => yy_rsc_9_0_i_qb,
      web => yy_rsc_9_0_web,
      db => yy_rsc_9_0_i_db,
      adrb => yy_rsc_9_0_i_adrb,
      qa => yy_rsc_9_0_i_qa,
      wea => yy_rsc_9_0_wea,
      da => yy_rsc_9_0_i_da,
      adra => yy_rsc_9_0_i_adra,
      adra_d => yy_rsc_9_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_9_0_i_clka_en_d,
      clkb_en_d => yy_rsc_9_0_i_clka_en_d,
      da_d => yy_rsc_9_0_i_da_d,
      qa_d => yy_rsc_9_0_i_qa_d_1,
      wea_d => yy_rsc_9_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_9_0_i_qb <= yy_rsc_9_0_qb;
  yy_rsc_9_0_db <= yy_rsc_9_0_i_db;
  yy_rsc_9_0_adrb <= yy_rsc_9_0_i_adrb;
  yy_rsc_9_0_i_qa <= yy_rsc_9_0_qa;
  yy_rsc_9_0_da <= yy_rsc_9_0_i_da;
  yy_rsc_9_0_adra <= yy_rsc_9_0_i_adra;
  yy_rsc_9_0_i_adra_d_1 <= yy_rsc_9_0_i_adra_d;
  yy_rsc_9_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_9_0_i_qa_d <= yy_rsc_9_0_i_qa_d_1;
  yy_rsc_9_0_i_wea_d_1 <= yy_rsc_9_0_i_wea_d;
  yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_10_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_52_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_10_0_clkb_en,
      clka_en => yy_rsc_10_0_clka_en,
      qb => yy_rsc_10_0_i_qb,
      web => yy_rsc_10_0_web,
      db => yy_rsc_10_0_i_db,
      adrb => yy_rsc_10_0_i_adrb,
      qa => yy_rsc_10_0_i_qa,
      wea => yy_rsc_10_0_wea,
      da => yy_rsc_10_0_i_da,
      adra => yy_rsc_10_0_i_adra,
      adra_d => yy_rsc_10_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_10_0_i_clka_en_d,
      clkb_en_d => yy_rsc_10_0_i_clka_en_d,
      da_d => yy_rsc_10_0_i_da_d,
      qa_d => yy_rsc_10_0_i_qa_d_1,
      wea_d => yy_rsc_10_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_10_0_i_qb <= yy_rsc_10_0_qb;
  yy_rsc_10_0_db <= yy_rsc_10_0_i_db;
  yy_rsc_10_0_adrb <= yy_rsc_10_0_i_adrb;
  yy_rsc_10_0_i_qa <= yy_rsc_10_0_qa;
  yy_rsc_10_0_da <= yy_rsc_10_0_i_da;
  yy_rsc_10_0_adra <= yy_rsc_10_0_i_adra;
  yy_rsc_10_0_i_adra_d_1 <= yy_rsc_10_0_i_adra_d;
  yy_rsc_10_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_10_0_i_qa_d <= yy_rsc_10_0_i_qa_d_1;
  yy_rsc_10_0_i_wea_d_1 <= yy_rsc_10_0_i_wea_d;
  yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_11_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_53_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_11_0_clkb_en,
      clka_en => yy_rsc_11_0_clka_en,
      qb => yy_rsc_11_0_i_qb,
      web => yy_rsc_11_0_web,
      db => yy_rsc_11_0_i_db,
      adrb => yy_rsc_11_0_i_adrb,
      qa => yy_rsc_11_0_i_qa,
      wea => yy_rsc_11_0_wea,
      da => yy_rsc_11_0_i_da,
      adra => yy_rsc_11_0_i_adra,
      adra_d => yy_rsc_11_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_11_0_i_clka_en_d,
      clkb_en_d => yy_rsc_11_0_i_clka_en_d,
      da_d => yy_rsc_11_0_i_da_d,
      qa_d => yy_rsc_11_0_i_qa_d_1,
      wea_d => yy_rsc_11_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_11_0_i_qb <= yy_rsc_11_0_qb;
  yy_rsc_11_0_db <= yy_rsc_11_0_i_db;
  yy_rsc_11_0_adrb <= yy_rsc_11_0_i_adrb;
  yy_rsc_11_0_i_qa <= yy_rsc_11_0_qa;
  yy_rsc_11_0_da <= yy_rsc_11_0_i_da;
  yy_rsc_11_0_adra <= yy_rsc_11_0_i_adra;
  yy_rsc_11_0_i_adra_d_1 <= yy_rsc_11_0_i_adra_d;
  yy_rsc_11_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_11_0_i_qa_d <= yy_rsc_11_0_i_qa_d_1;
  yy_rsc_11_0_i_wea_d_1 <= yy_rsc_11_0_i_wea_d;
  yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_12_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_54_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_12_0_clkb_en,
      clka_en => yy_rsc_12_0_clka_en,
      qb => yy_rsc_12_0_i_qb,
      web => yy_rsc_12_0_web,
      db => yy_rsc_12_0_i_db,
      adrb => yy_rsc_12_0_i_adrb,
      qa => yy_rsc_12_0_i_qa,
      wea => yy_rsc_12_0_wea,
      da => yy_rsc_12_0_i_da,
      adra => yy_rsc_12_0_i_adra,
      adra_d => yy_rsc_12_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_12_0_i_clka_en_d,
      clkb_en_d => yy_rsc_12_0_i_clka_en_d,
      da_d => yy_rsc_12_0_i_da_d,
      qa_d => yy_rsc_12_0_i_qa_d_1,
      wea_d => yy_rsc_12_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_12_0_i_qb <= yy_rsc_12_0_qb;
  yy_rsc_12_0_db <= yy_rsc_12_0_i_db;
  yy_rsc_12_0_adrb <= yy_rsc_12_0_i_adrb;
  yy_rsc_12_0_i_qa <= yy_rsc_12_0_qa;
  yy_rsc_12_0_da <= yy_rsc_12_0_i_da;
  yy_rsc_12_0_adra <= yy_rsc_12_0_i_adra;
  yy_rsc_12_0_i_adra_d_1 <= yy_rsc_12_0_i_adra_d;
  yy_rsc_12_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_12_0_i_qa_d <= yy_rsc_12_0_i_qa_d_1;
  yy_rsc_12_0_i_wea_d_1 <= yy_rsc_12_0_i_wea_d;
  yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_13_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_55_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_13_0_clkb_en,
      clka_en => yy_rsc_13_0_clka_en,
      qb => yy_rsc_13_0_i_qb,
      web => yy_rsc_13_0_web,
      db => yy_rsc_13_0_i_db,
      adrb => yy_rsc_13_0_i_adrb,
      qa => yy_rsc_13_0_i_qa,
      wea => yy_rsc_13_0_wea,
      da => yy_rsc_13_0_i_da,
      adra => yy_rsc_13_0_i_adra,
      adra_d => yy_rsc_13_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_13_0_i_clka_en_d,
      clkb_en_d => yy_rsc_13_0_i_clka_en_d,
      da_d => yy_rsc_13_0_i_da_d,
      qa_d => yy_rsc_13_0_i_qa_d_1,
      wea_d => yy_rsc_13_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_13_0_i_qb <= yy_rsc_13_0_qb;
  yy_rsc_13_0_db <= yy_rsc_13_0_i_db;
  yy_rsc_13_0_adrb <= yy_rsc_13_0_i_adrb;
  yy_rsc_13_0_i_qa <= yy_rsc_13_0_qa;
  yy_rsc_13_0_da <= yy_rsc_13_0_i_da;
  yy_rsc_13_0_adra <= yy_rsc_13_0_i_adra;
  yy_rsc_13_0_i_adra_d_1 <= yy_rsc_13_0_i_adra_d;
  yy_rsc_13_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_13_0_i_qa_d <= yy_rsc_13_0_i_qa_d_1;
  yy_rsc_13_0_i_wea_d_1 <= yy_rsc_13_0_i_wea_d;
  yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_14_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_56_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_14_0_clkb_en,
      clka_en => yy_rsc_14_0_clka_en,
      qb => yy_rsc_14_0_i_qb,
      web => yy_rsc_14_0_web,
      db => yy_rsc_14_0_i_db,
      adrb => yy_rsc_14_0_i_adrb,
      qa => yy_rsc_14_0_i_qa,
      wea => yy_rsc_14_0_wea,
      da => yy_rsc_14_0_i_da,
      adra => yy_rsc_14_0_i_adra,
      adra_d => yy_rsc_14_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_14_0_i_clka_en_d,
      clkb_en_d => yy_rsc_14_0_i_clka_en_d,
      da_d => yy_rsc_14_0_i_da_d,
      qa_d => yy_rsc_14_0_i_qa_d_1,
      wea_d => yy_rsc_14_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_14_0_i_qb <= yy_rsc_14_0_qb;
  yy_rsc_14_0_db <= yy_rsc_14_0_i_db;
  yy_rsc_14_0_adrb <= yy_rsc_14_0_i_adrb;
  yy_rsc_14_0_i_qa <= yy_rsc_14_0_qa;
  yy_rsc_14_0_da <= yy_rsc_14_0_i_da;
  yy_rsc_14_0_adra <= yy_rsc_14_0_i_adra;
  yy_rsc_14_0_i_adra_d_1 <= yy_rsc_14_0_i_adra_d;
  yy_rsc_14_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_14_0_i_qa_d <= yy_rsc_14_0_i_qa_d_1;
  yy_rsc_14_0_i_wea_d_1 <= yy_rsc_14_0_i_wea_d;
  yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_15_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_57_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_15_0_clkb_en,
      clka_en => yy_rsc_15_0_clka_en,
      qb => yy_rsc_15_0_i_qb,
      web => yy_rsc_15_0_web,
      db => yy_rsc_15_0_i_db,
      adrb => yy_rsc_15_0_i_adrb,
      qa => yy_rsc_15_0_i_qa,
      wea => yy_rsc_15_0_wea,
      da => yy_rsc_15_0_i_da,
      adra => yy_rsc_15_0_i_adra,
      adra_d => yy_rsc_15_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_15_0_i_clka_en_d,
      clkb_en_d => yy_rsc_15_0_i_clka_en_d,
      da_d => yy_rsc_15_0_i_da_d,
      qa_d => yy_rsc_15_0_i_qa_d_1,
      wea_d => yy_rsc_15_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_15_0_i_qb <= yy_rsc_15_0_qb;
  yy_rsc_15_0_db <= yy_rsc_15_0_i_db;
  yy_rsc_15_0_adrb <= yy_rsc_15_0_i_adrb;
  yy_rsc_15_0_i_qa <= yy_rsc_15_0_qa;
  yy_rsc_15_0_da <= yy_rsc_15_0_i_da;
  yy_rsc_15_0_adra <= yy_rsc_15_0_i_adra;
  yy_rsc_15_0_i_adra_d_1 <= yy_rsc_15_0_i_adra_d;
  yy_rsc_15_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_15_0_i_qa_d <= yy_rsc_15_0_i_qa_d_1;
  yy_rsc_15_0_i_wea_d_1 <= yy_rsc_15_0_i_wea_d;
  yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_16_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_58_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_16_0_clkb_en,
      clka_en => yy_rsc_16_0_clka_en,
      qb => yy_rsc_16_0_i_qb,
      web => yy_rsc_16_0_web,
      db => yy_rsc_16_0_i_db,
      adrb => yy_rsc_16_0_i_adrb,
      qa => yy_rsc_16_0_i_qa,
      wea => yy_rsc_16_0_wea,
      da => yy_rsc_16_0_i_da,
      adra => yy_rsc_16_0_i_adra,
      adra_d => yy_rsc_16_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_16_0_i_clka_en_d,
      clkb_en_d => yy_rsc_16_0_i_clka_en_d,
      da_d => yy_rsc_16_0_i_da_d,
      qa_d => yy_rsc_16_0_i_qa_d_1,
      wea_d => yy_rsc_16_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_16_0_i_qb <= yy_rsc_16_0_qb;
  yy_rsc_16_0_db <= yy_rsc_16_0_i_db;
  yy_rsc_16_0_adrb <= yy_rsc_16_0_i_adrb;
  yy_rsc_16_0_i_qa <= yy_rsc_16_0_qa;
  yy_rsc_16_0_da <= yy_rsc_16_0_i_da;
  yy_rsc_16_0_adra <= yy_rsc_16_0_i_adra;
  yy_rsc_16_0_i_adra_d_1 <= yy_rsc_16_0_i_adra_d;
  yy_rsc_16_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_16_0_i_qa_d <= yy_rsc_16_0_i_qa_d_1;
  yy_rsc_16_0_i_wea_d_1 <= yy_rsc_16_0_i_wea_d;
  yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_17_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_59_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_17_0_clkb_en,
      clka_en => yy_rsc_17_0_clka_en,
      qb => yy_rsc_17_0_i_qb,
      web => yy_rsc_17_0_web,
      db => yy_rsc_17_0_i_db,
      adrb => yy_rsc_17_0_i_adrb,
      qa => yy_rsc_17_0_i_qa,
      wea => yy_rsc_17_0_wea,
      da => yy_rsc_17_0_i_da,
      adra => yy_rsc_17_0_i_adra,
      adra_d => yy_rsc_17_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_17_0_i_clka_en_d,
      clkb_en_d => yy_rsc_17_0_i_clka_en_d,
      da_d => yy_rsc_17_0_i_da_d,
      qa_d => yy_rsc_17_0_i_qa_d_1,
      wea_d => yy_rsc_17_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_17_0_i_qb <= yy_rsc_17_0_qb;
  yy_rsc_17_0_db <= yy_rsc_17_0_i_db;
  yy_rsc_17_0_adrb <= yy_rsc_17_0_i_adrb;
  yy_rsc_17_0_i_qa <= yy_rsc_17_0_qa;
  yy_rsc_17_0_da <= yy_rsc_17_0_i_da;
  yy_rsc_17_0_adra <= yy_rsc_17_0_i_adra;
  yy_rsc_17_0_i_adra_d_1 <= yy_rsc_17_0_i_adra_d;
  yy_rsc_17_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_17_0_i_qa_d <= yy_rsc_17_0_i_qa_d_1;
  yy_rsc_17_0_i_wea_d_1 <= yy_rsc_17_0_i_wea_d;
  yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_18_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_60_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_18_0_clkb_en,
      clka_en => yy_rsc_18_0_clka_en,
      qb => yy_rsc_18_0_i_qb,
      web => yy_rsc_18_0_web,
      db => yy_rsc_18_0_i_db,
      adrb => yy_rsc_18_0_i_adrb,
      qa => yy_rsc_18_0_i_qa,
      wea => yy_rsc_18_0_wea,
      da => yy_rsc_18_0_i_da,
      adra => yy_rsc_18_0_i_adra,
      adra_d => yy_rsc_18_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_18_0_i_clka_en_d,
      clkb_en_d => yy_rsc_18_0_i_clka_en_d,
      da_d => yy_rsc_18_0_i_da_d,
      qa_d => yy_rsc_18_0_i_qa_d_1,
      wea_d => yy_rsc_18_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_18_0_i_qb <= yy_rsc_18_0_qb;
  yy_rsc_18_0_db <= yy_rsc_18_0_i_db;
  yy_rsc_18_0_adrb <= yy_rsc_18_0_i_adrb;
  yy_rsc_18_0_i_qa <= yy_rsc_18_0_qa;
  yy_rsc_18_0_da <= yy_rsc_18_0_i_da;
  yy_rsc_18_0_adra <= yy_rsc_18_0_i_adra;
  yy_rsc_18_0_i_adra_d_1 <= yy_rsc_18_0_i_adra_d;
  yy_rsc_18_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_18_0_i_qa_d <= yy_rsc_18_0_i_qa_d_1;
  yy_rsc_18_0_i_wea_d_1 <= yy_rsc_18_0_i_wea_d;
  yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_19_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_61_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_19_0_clkb_en,
      clka_en => yy_rsc_19_0_clka_en,
      qb => yy_rsc_19_0_i_qb,
      web => yy_rsc_19_0_web,
      db => yy_rsc_19_0_i_db,
      adrb => yy_rsc_19_0_i_adrb,
      qa => yy_rsc_19_0_i_qa,
      wea => yy_rsc_19_0_wea,
      da => yy_rsc_19_0_i_da,
      adra => yy_rsc_19_0_i_adra,
      adra_d => yy_rsc_19_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_19_0_i_clka_en_d,
      clkb_en_d => yy_rsc_19_0_i_clka_en_d,
      da_d => yy_rsc_19_0_i_da_d,
      qa_d => yy_rsc_19_0_i_qa_d_1,
      wea_d => yy_rsc_19_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_19_0_i_qb <= yy_rsc_19_0_qb;
  yy_rsc_19_0_db <= yy_rsc_19_0_i_db;
  yy_rsc_19_0_adrb <= yy_rsc_19_0_i_adrb;
  yy_rsc_19_0_i_qa <= yy_rsc_19_0_qa;
  yy_rsc_19_0_da <= yy_rsc_19_0_i_da;
  yy_rsc_19_0_adra <= yy_rsc_19_0_i_adra;
  yy_rsc_19_0_i_adra_d_1 <= yy_rsc_19_0_i_adra_d;
  yy_rsc_19_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_19_0_i_qa_d <= yy_rsc_19_0_i_qa_d_1;
  yy_rsc_19_0_i_wea_d_1 <= yy_rsc_19_0_i_wea_d;
  yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_20_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_62_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_20_0_clkb_en,
      clka_en => yy_rsc_20_0_clka_en,
      qb => yy_rsc_20_0_i_qb,
      web => yy_rsc_20_0_web,
      db => yy_rsc_20_0_i_db,
      adrb => yy_rsc_20_0_i_adrb,
      qa => yy_rsc_20_0_i_qa,
      wea => yy_rsc_20_0_wea,
      da => yy_rsc_20_0_i_da,
      adra => yy_rsc_20_0_i_adra,
      adra_d => yy_rsc_20_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_20_0_i_clka_en_d,
      clkb_en_d => yy_rsc_20_0_i_clka_en_d,
      da_d => yy_rsc_20_0_i_da_d,
      qa_d => yy_rsc_20_0_i_qa_d_1,
      wea_d => yy_rsc_20_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_20_0_i_qb <= yy_rsc_20_0_qb;
  yy_rsc_20_0_db <= yy_rsc_20_0_i_db;
  yy_rsc_20_0_adrb <= yy_rsc_20_0_i_adrb;
  yy_rsc_20_0_i_qa <= yy_rsc_20_0_qa;
  yy_rsc_20_0_da <= yy_rsc_20_0_i_da;
  yy_rsc_20_0_adra <= yy_rsc_20_0_i_adra;
  yy_rsc_20_0_i_adra_d_1 <= yy_rsc_20_0_i_adra_d;
  yy_rsc_20_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_20_0_i_qa_d <= yy_rsc_20_0_i_qa_d_1;
  yy_rsc_20_0_i_wea_d_1 <= yy_rsc_20_0_i_wea_d;
  yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_21_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_63_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_21_0_clkb_en,
      clka_en => yy_rsc_21_0_clka_en,
      qb => yy_rsc_21_0_i_qb,
      web => yy_rsc_21_0_web,
      db => yy_rsc_21_0_i_db,
      adrb => yy_rsc_21_0_i_adrb,
      qa => yy_rsc_21_0_i_qa,
      wea => yy_rsc_21_0_wea,
      da => yy_rsc_21_0_i_da,
      adra => yy_rsc_21_0_i_adra,
      adra_d => yy_rsc_21_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_21_0_i_clka_en_d,
      clkb_en_d => yy_rsc_21_0_i_clka_en_d,
      da_d => yy_rsc_21_0_i_da_d,
      qa_d => yy_rsc_21_0_i_qa_d_1,
      wea_d => yy_rsc_21_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_21_0_i_qb <= yy_rsc_21_0_qb;
  yy_rsc_21_0_db <= yy_rsc_21_0_i_db;
  yy_rsc_21_0_adrb <= yy_rsc_21_0_i_adrb;
  yy_rsc_21_0_i_qa <= yy_rsc_21_0_qa;
  yy_rsc_21_0_da <= yy_rsc_21_0_i_da;
  yy_rsc_21_0_adra <= yy_rsc_21_0_i_adra;
  yy_rsc_21_0_i_adra_d_1 <= yy_rsc_21_0_i_adra_d;
  yy_rsc_21_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_21_0_i_qa_d <= yy_rsc_21_0_i_qa_d_1;
  yy_rsc_21_0_i_wea_d_1 <= yy_rsc_21_0_i_wea_d;
  yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_22_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_64_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_22_0_clkb_en,
      clka_en => yy_rsc_22_0_clka_en,
      qb => yy_rsc_22_0_i_qb,
      web => yy_rsc_22_0_web,
      db => yy_rsc_22_0_i_db,
      adrb => yy_rsc_22_0_i_adrb,
      qa => yy_rsc_22_0_i_qa,
      wea => yy_rsc_22_0_wea,
      da => yy_rsc_22_0_i_da,
      adra => yy_rsc_22_0_i_adra,
      adra_d => yy_rsc_22_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_22_0_i_clka_en_d,
      clkb_en_d => yy_rsc_22_0_i_clka_en_d,
      da_d => yy_rsc_22_0_i_da_d,
      qa_d => yy_rsc_22_0_i_qa_d_1,
      wea_d => yy_rsc_22_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_22_0_i_qb <= yy_rsc_22_0_qb;
  yy_rsc_22_0_db <= yy_rsc_22_0_i_db;
  yy_rsc_22_0_adrb <= yy_rsc_22_0_i_adrb;
  yy_rsc_22_0_i_qa <= yy_rsc_22_0_qa;
  yy_rsc_22_0_da <= yy_rsc_22_0_i_da;
  yy_rsc_22_0_adra <= yy_rsc_22_0_i_adra;
  yy_rsc_22_0_i_adra_d_1 <= yy_rsc_22_0_i_adra_d;
  yy_rsc_22_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_22_0_i_qa_d <= yy_rsc_22_0_i_qa_d_1;
  yy_rsc_22_0_i_wea_d_1 <= yy_rsc_22_0_i_wea_d;
  yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_23_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_65_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_23_0_clkb_en,
      clka_en => yy_rsc_23_0_clka_en,
      qb => yy_rsc_23_0_i_qb,
      web => yy_rsc_23_0_web,
      db => yy_rsc_23_0_i_db,
      adrb => yy_rsc_23_0_i_adrb,
      qa => yy_rsc_23_0_i_qa,
      wea => yy_rsc_23_0_wea,
      da => yy_rsc_23_0_i_da,
      adra => yy_rsc_23_0_i_adra,
      adra_d => yy_rsc_23_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_23_0_i_clka_en_d,
      clkb_en_d => yy_rsc_23_0_i_clka_en_d,
      da_d => yy_rsc_23_0_i_da_d,
      qa_d => yy_rsc_23_0_i_qa_d_1,
      wea_d => yy_rsc_23_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_23_0_i_qb <= yy_rsc_23_0_qb;
  yy_rsc_23_0_db <= yy_rsc_23_0_i_db;
  yy_rsc_23_0_adrb <= yy_rsc_23_0_i_adrb;
  yy_rsc_23_0_i_qa <= yy_rsc_23_0_qa;
  yy_rsc_23_0_da <= yy_rsc_23_0_i_da;
  yy_rsc_23_0_adra <= yy_rsc_23_0_i_adra;
  yy_rsc_23_0_i_adra_d_1 <= yy_rsc_23_0_i_adra_d;
  yy_rsc_23_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_23_0_i_qa_d <= yy_rsc_23_0_i_qa_d_1;
  yy_rsc_23_0_i_wea_d_1 <= yy_rsc_23_0_i_wea_d;
  yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_24_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_66_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_24_0_clkb_en,
      clka_en => yy_rsc_24_0_clka_en,
      qb => yy_rsc_24_0_i_qb,
      web => yy_rsc_24_0_web,
      db => yy_rsc_24_0_i_db,
      adrb => yy_rsc_24_0_i_adrb,
      qa => yy_rsc_24_0_i_qa,
      wea => yy_rsc_24_0_wea,
      da => yy_rsc_24_0_i_da,
      adra => yy_rsc_24_0_i_adra,
      adra_d => yy_rsc_24_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_24_0_i_clka_en_d,
      clkb_en_d => yy_rsc_24_0_i_clka_en_d,
      da_d => yy_rsc_24_0_i_da_d,
      qa_d => yy_rsc_24_0_i_qa_d_1,
      wea_d => yy_rsc_24_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_24_0_i_qb <= yy_rsc_24_0_qb;
  yy_rsc_24_0_db <= yy_rsc_24_0_i_db;
  yy_rsc_24_0_adrb <= yy_rsc_24_0_i_adrb;
  yy_rsc_24_0_i_qa <= yy_rsc_24_0_qa;
  yy_rsc_24_0_da <= yy_rsc_24_0_i_da;
  yy_rsc_24_0_adra <= yy_rsc_24_0_i_adra;
  yy_rsc_24_0_i_adra_d_1 <= yy_rsc_24_0_i_adra_d;
  yy_rsc_24_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_24_0_i_qa_d <= yy_rsc_24_0_i_qa_d_1;
  yy_rsc_24_0_i_wea_d_1 <= yy_rsc_24_0_i_wea_d;
  yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_25_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_67_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_25_0_clkb_en,
      clka_en => yy_rsc_25_0_clka_en,
      qb => yy_rsc_25_0_i_qb,
      web => yy_rsc_25_0_web,
      db => yy_rsc_25_0_i_db,
      adrb => yy_rsc_25_0_i_adrb,
      qa => yy_rsc_25_0_i_qa,
      wea => yy_rsc_25_0_wea,
      da => yy_rsc_25_0_i_da,
      adra => yy_rsc_25_0_i_adra,
      adra_d => yy_rsc_25_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_25_0_i_clka_en_d,
      clkb_en_d => yy_rsc_25_0_i_clka_en_d,
      da_d => yy_rsc_25_0_i_da_d,
      qa_d => yy_rsc_25_0_i_qa_d_1,
      wea_d => yy_rsc_25_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_25_0_i_qb <= yy_rsc_25_0_qb;
  yy_rsc_25_0_db <= yy_rsc_25_0_i_db;
  yy_rsc_25_0_adrb <= yy_rsc_25_0_i_adrb;
  yy_rsc_25_0_i_qa <= yy_rsc_25_0_qa;
  yy_rsc_25_0_da <= yy_rsc_25_0_i_da;
  yy_rsc_25_0_adra <= yy_rsc_25_0_i_adra;
  yy_rsc_25_0_i_adra_d_1 <= yy_rsc_25_0_i_adra_d;
  yy_rsc_25_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_25_0_i_qa_d <= yy_rsc_25_0_i_qa_d_1;
  yy_rsc_25_0_i_wea_d_1 <= yy_rsc_25_0_i_wea_d;
  yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_26_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_68_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_26_0_clkb_en,
      clka_en => yy_rsc_26_0_clka_en,
      qb => yy_rsc_26_0_i_qb,
      web => yy_rsc_26_0_web,
      db => yy_rsc_26_0_i_db,
      adrb => yy_rsc_26_0_i_adrb,
      qa => yy_rsc_26_0_i_qa,
      wea => yy_rsc_26_0_wea,
      da => yy_rsc_26_0_i_da,
      adra => yy_rsc_26_0_i_adra,
      adra_d => yy_rsc_26_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_26_0_i_clka_en_d,
      clkb_en_d => yy_rsc_26_0_i_clka_en_d,
      da_d => yy_rsc_26_0_i_da_d,
      qa_d => yy_rsc_26_0_i_qa_d_1,
      wea_d => yy_rsc_26_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_26_0_i_qb <= yy_rsc_26_0_qb;
  yy_rsc_26_0_db <= yy_rsc_26_0_i_db;
  yy_rsc_26_0_adrb <= yy_rsc_26_0_i_adrb;
  yy_rsc_26_0_i_qa <= yy_rsc_26_0_qa;
  yy_rsc_26_0_da <= yy_rsc_26_0_i_da;
  yy_rsc_26_0_adra <= yy_rsc_26_0_i_adra;
  yy_rsc_26_0_i_adra_d_1 <= yy_rsc_26_0_i_adra_d;
  yy_rsc_26_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_26_0_i_qa_d <= yy_rsc_26_0_i_qa_d_1;
  yy_rsc_26_0_i_wea_d_1 <= yy_rsc_26_0_i_wea_d;
  yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_27_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_69_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_27_0_clkb_en,
      clka_en => yy_rsc_27_0_clka_en,
      qb => yy_rsc_27_0_i_qb,
      web => yy_rsc_27_0_web,
      db => yy_rsc_27_0_i_db,
      adrb => yy_rsc_27_0_i_adrb,
      qa => yy_rsc_27_0_i_qa,
      wea => yy_rsc_27_0_wea,
      da => yy_rsc_27_0_i_da,
      adra => yy_rsc_27_0_i_adra,
      adra_d => yy_rsc_27_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_27_0_i_clka_en_d,
      clkb_en_d => yy_rsc_27_0_i_clka_en_d,
      da_d => yy_rsc_27_0_i_da_d,
      qa_d => yy_rsc_27_0_i_qa_d_1,
      wea_d => yy_rsc_27_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_27_0_i_qb <= yy_rsc_27_0_qb;
  yy_rsc_27_0_db <= yy_rsc_27_0_i_db;
  yy_rsc_27_0_adrb <= yy_rsc_27_0_i_adrb;
  yy_rsc_27_0_i_qa <= yy_rsc_27_0_qa;
  yy_rsc_27_0_da <= yy_rsc_27_0_i_da;
  yy_rsc_27_0_adra <= yy_rsc_27_0_i_adra;
  yy_rsc_27_0_i_adra_d_1 <= yy_rsc_27_0_i_adra_d;
  yy_rsc_27_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_27_0_i_qa_d <= yy_rsc_27_0_i_qa_d_1;
  yy_rsc_27_0_i_wea_d_1 <= yy_rsc_27_0_i_wea_d;
  yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_28_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_70_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_28_0_clkb_en,
      clka_en => yy_rsc_28_0_clka_en,
      qb => yy_rsc_28_0_i_qb,
      web => yy_rsc_28_0_web,
      db => yy_rsc_28_0_i_db,
      adrb => yy_rsc_28_0_i_adrb,
      qa => yy_rsc_28_0_i_qa,
      wea => yy_rsc_28_0_wea,
      da => yy_rsc_28_0_i_da,
      adra => yy_rsc_28_0_i_adra,
      adra_d => yy_rsc_28_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_28_0_i_clka_en_d,
      clkb_en_d => yy_rsc_28_0_i_clka_en_d,
      da_d => yy_rsc_28_0_i_da_d,
      qa_d => yy_rsc_28_0_i_qa_d_1,
      wea_d => yy_rsc_28_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_28_0_i_qb <= yy_rsc_28_0_qb;
  yy_rsc_28_0_db <= yy_rsc_28_0_i_db;
  yy_rsc_28_0_adrb <= yy_rsc_28_0_i_adrb;
  yy_rsc_28_0_i_qa <= yy_rsc_28_0_qa;
  yy_rsc_28_0_da <= yy_rsc_28_0_i_da;
  yy_rsc_28_0_adra <= yy_rsc_28_0_i_adra;
  yy_rsc_28_0_i_adra_d_1 <= yy_rsc_28_0_i_adra_d;
  yy_rsc_28_0_i_da_d <= yy_rsc_0_0_i_da_d_iff;
  yy_rsc_28_0_i_qa_d <= yy_rsc_28_0_i_qa_d_1;
  yy_rsc_28_0_i_wea_d_1 <= yy_rsc_28_0_i_wea_d;
  yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_29_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_71_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_29_0_clkb_en,
      clka_en => yy_rsc_29_0_clka_en,
      qb => yy_rsc_29_0_i_qb,
      web => yy_rsc_29_0_web,
      db => yy_rsc_29_0_i_db,
      adrb => yy_rsc_29_0_i_adrb,
      qa => yy_rsc_29_0_i_qa,
      wea => yy_rsc_29_0_wea,
      da => yy_rsc_29_0_i_da,
      adra => yy_rsc_29_0_i_adra,
      adra_d => yy_rsc_29_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_29_0_i_clka_en_d,
      clkb_en_d => yy_rsc_29_0_i_clka_en_d,
      da_d => yy_rsc_29_0_i_da_d,
      qa_d => yy_rsc_29_0_i_qa_d_1,
      wea_d => yy_rsc_29_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_29_0_i_qb <= yy_rsc_29_0_qb;
  yy_rsc_29_0_db <= yy_rsc_29_0_i_db;
  yy_rsc_29_0_adrb <= yy_rsc_29_0_i_adrb;
  yy_rsc_29_0_i_qa <= yy_rsc_29_0_qa;
  yy_rsc_29_0_da <= yy_rsc_29_0_i_da;
  yy_rsc_29_0_adra <= yy_rsc_29_0_i_adra;
  yy_rsc_29_0_i_adra_d_1 <= yy_rsc_29_0_i_adra_d;
  yy_rsc_29_0_i_da_d <= yy_rsc_1_0_i_da_d_iff;
  yy_rsc_29_0_i_qa_d <= yy_rsc_29_0_i_qa_d_1;
  yy_rsc_29_0_i_wea_d_1 <= yy_rsc_29_0_i_wea_d;
  yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_30_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_72_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_30_0_clkb_en,
      clka_en => yy_rsc_30_0_clka_en,
      qb => yy_rsc_30_0_i_qb,
      web => yy_rsc_30_0_web,
      db => yy_rsc_30_0_i_db,
      adrb => yy_rsc_30_0_i_adrb,
      qa => yy_rsc_30_0_i_qa,
      wea => yy_rsc_30_0_wea,
      da => yy_rsc_30_0_i_da,
      adra => yy_rsc_30_0_i_adra,
      adra_d => yy_rsc_30_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_30_0_i_clka_en_d,
      clkb_en_d => yy_rsc_30_0_i_clka_en_d,
      da_d => yy_rsc_30_0_i_da_d,
      qa_d => yy_rsc_30_0_i_qa_d_1,
      wea_d => yy_rsc_30_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_30_0_i_qb <= yy_rsc_30_0_qb;
  yy_rsc_30_0_db <= yy_rsc_30_0_i_db;
  yy_rsc_30_0_adrb <= yy_rsc_30_0_i_adrb;
  yy_rsc_30_0_i_qa <= yy_rsc_30_0_qa;
  yy_rsc_30_0_da <= yy_rsc_30_0_i_da;
  yy_rsc_30_0_adra <= yy_rsc_30_0_i_adra;
  yy_rsc_30_0_i_adra_d_1 <= yy_rsc_30_0_i_adra_d;
  yy_rsc_30_0_i_da_d <= yy_rsc_2_0_i_da_d_iff;
  yy_rsc_30_0_i_qa_d <= yy_rsc_30_0_i_qa_d_1;
  yy_rsc_30_0_i_wea_d_1 <= yy_rsc_30_0_i_wea_d;
  yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  yy_rsc_31_0_i : hybrid_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_73_5_32_32_32_32_1_gen
    PORT MAP(
      clkb_en => yy_rsc_31_0_clkb_en,
      clka_en => yy_rsc_31_0_clka_en,
      qb => yy_rsc_31_0_i_qb,
      web => yy_rsc_31_0_web,
      db => yy_rsc_31_0_i_db,
      adrb => yy_rsc_31_0_i_adrb,
      qa => yy_rsc_31_0_i_qa,
      wea => yy_rsc_31_0_wea,
      da => yy_rsc_31_0_i_da,
      adra => yy_rsc_31_0_i_adra,
      adra_d => yy_rsc_31_0_i_adra_d_1,
      clka => clk,
      clka_en_d => yy_rsc_31_0_i_clka_en_d,
      clkb_en_d => yy_rsc_31_0_i_clka_en_d,
      da_d => yy_rsc_31_0_i_da_d,
      qa_d => yy_rsc_31_0_i_qa_d_1,
      wea_d => yy_rsc_31_0_i_wea_d_1,
      rwA_rw_ram_ir_internal_RMASK_B_d => yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1,
      rwA_rw_ram_ir_internal_WMASK_B_d => yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1
    );
  yy_rsc_31_0_i_qb <= yy_rsc_31_0_qb;
  yy_rsc_31_0_db <= yy_rsc_31_0_i_db;
  yy_rsc_31_0_adrb <= yy_rsc_31_0_i_adrb;
  yy_rsc_31_0_i_qa <= yy_rsc_31_0_qa;
  yy_rsc_31_0_da <= yy_rsc_31_0_i_da;
  yy_rsc_31_0_adra <= yy_rsc_31_0_i_adra;
  yy_rsc_31_0_i_adra_d_1 <= yy_rsc_31_0_i_adra_d;
  yy_rsc_31_0_i_da_d <= yy_rsc_3_0_i_da_d_iff;
  yy_rsc_31_0_i_qa_d <= yy_rsc_31_0_i_qa_d_1;
  yy_rsc_31_0_i_wea_d_1 <= yy_rsc_31_0_i_wea_d;
  yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_1 <= yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d_1 <= yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;

  hybrid_core_inst : hybrid_core
    PORT MAP(
      clk => clk,
      rst => rst,
      x_rsc_0_0_s_tdone => x_rsc_0_0_s_tdone,
      x_rsc_0_0_tr_write_done => x_rsc_0_0_tr_write_done,
      x_rsc_0_0_RREADY => x_rsc_0_0_RREADY,
      x_rsc_0_0_RVALID => x_rsc_0_0_RVALID,
      x_rsc_0_0_RUSER => x_rsc_0_0_RUSER,
      x_rsc_0_0_RLAST => x_rsc_0_0_RLAST,
      x_rsc_0_0_RRESP => hybrid_core_inst_x_rsc_0_0_RRESP,
      x_rsc_0_0_RDATA => hybrid_core_inst_x_rsc_0_0_RDATA,
      x_rsc_0_0_RID => x_rsc_0_0_RID,
      x_rsc_0_0_ARREADY => x_rsc_0_0_ARREADY,
      x_rsc_0_0_ARVALID => x_rsc_0_0_ARVALID,
      x_rsc_0_0_ARUSER => x_rsc_0_0_ARUSER,
      x_rsc_0_0_ARREGION => hybrid_core_inst_x_rsc_0_0_ARREGION,
      x_rsc_0_0_ARQOS => hybrid_core_inst_x_rsc_0_0_ARQOS,
      x_rsc_0_0_ARPROT => hybrid_core_inst_x_rsc_0_0_ARPROT,
      x_rsc_0_0_ARCACHE => hybrid_core_inst_x_rsc_0_0_ARCACHE,
      x_rsc_0_0_ARLOCK => x_rsc_0_0_ARLOCK,
      x_rsc_0_0_ARBURST => hybrid_core_inst_x_rsc_0_0_ARBURST,
      x_rsc_0_0_ARSIZE => hybrid_core_inst_x_rsc_0_0_ARSIZE,
      x_rsc_0_0_ARLEN => hybrid_core_inst_x_rsc_0_0_ARLEN,
      x_rsc_0_0_ARADDR => hybrid_core_inst_x_rsc_0_0_ARADDR,
      x_rsc_0_0_ARID => x_rsc_0_0_ARID,
      x_rsc_0_0_BREADY => x_rsc_0_0_BREADY,
      x_rsc_0_0_BVALID => x_rsc_0_0_BVALID,
      x_rsc_0_0_BUSER => x_rsc_0_0_BUSER,
      x_rsc_0_0_BRESP => hybrid_core_inst_x_rsc_0_0_BRESP,
      x_rsc_0_0_BID => x_rsc_0_0_BID,
      x_rsc_0_0_WREADY => x_rsc_0_0_WREADY,
      x_rsc_0_0_WVALID => x_rsc_0_0_WVALID,
      x_rsc_0_0_WUSER => x_rsc_0_0_WUSER,
      x_rsc_0_0_WLAST => x_rsc_0_0_WLAST,
      x_rsc_0_0_WSTRB => hybrid_core_inst_x_rsc_0_0_WSTRB,
      x_rsc_0_0_WDATA => hybrid_core_inst_x_rsc_0_0_WDATA,
      x_rsc_0_0_AWREADY => x_rsc_0_0_AWREADY,
      x_rsc_0_0_AWVALID => x_rsc_0_0_AWVALID,
      x_rsc_0_0_AWUSER => x_rsc_0_0_AWUSER,
      x_rsc_0_0_AWREGION => hybrid_core_inst_x_rsc_0_0_AWREGION,
      x_rsc_0_0_AWQOS => hybrid_core_inst_x_rsc_0_0_AWQOS,
      x_rsc_0_0_AWPROT => hybrid_core_inst_x_rsc_0_0_AWPROT,
      x_rsc_0_0_AWCACHE => hybrid_core_inst_x_rsc_0_0_AWCACHE,
      x_rsc_0_0_AWLOCK => x_rsc_0_0_AWLOCK,
      x_rsc_0_0_AWBURST => hybrid_core_inst_x_rsc_0_0_AWBURST,
      x_rsc_0_0_AWSIZE => hybrid_core_inst_x_rsc_0_0_AWSIZE,
      x_rsc_0_0_AWLEN => hybrid_core_inst_x_rsc_0_0_AWLEN,
      x_rsc_0_0_AWADDR => hybrid_core_inst_x_rsc_0_0_AWADDR,
      x_rsc_0_0_AWID => x_rsc_0_0_AWID,
      x_rsc_triosy_0_0_lz => x_rsc_triosy_0_0_lz,
      x_rsc_1_0_s_tdone => x_rsc_1_0_s_tdone,
      x_rsc_1_0_tr_write_done => x_rsc_1_0_tr_write_done,
      x_rsc_1_0_RREADY => x_rsc_1_0_RREADY,
      x_rsc_1_0_RVALID => x_rsc_1_0_RVALID,
      x_rsc_1_0_RUSER => x_rsc_1_0_RUSER,
      x_rsc_1_0_RLAST => x_rsc_1_0_RLAST,
      x_rsc_1_0_RRESP => hybrid_core_inst_x_rsc_1_0_RRESP,
      x_rsc_1_0_RDATA => hybrid_core_inst_x_rsc_1_0_RDATA,
      x_rsc_1_0_RID => x_rsc_1_0_RID,
      x_rsc_1_0_ARREADY => x_rsc_1_0_ARREADY,
      x_rsc_1_0_ARVALID => x_rsc_1_0_ARVALID,
      x_rsc_1_0_ARUSER => x_rsc_1_0_ARUSER,
      x_rsc_1_0_ARREGION => hybrid_core_inst_x_rsc_1_0_ARREGION,
      x_rsc_1_0_ARQOS => hybrid_core_inst_x_rsc_1_0_ARQOS,
      x_rsc_1_0_ARPROT => hybrid_core_inst_x_rsc_1_0_ARPROT,
      x_rsc_1_0_ARCACHE => hybrid_core_inst_x_rsc_1_0_ARCACHE,
      x_rsc_1_0_ARLOCK => x_rsc_1_0_ARLOCK,
      x_rsc_1_0_ARBURST => hybrid_core_inst_x_rsc_1_0_ARBURST,
      x_rsc_1_0_ARSIZE => hybrid_core_inst_x_rsc_1_0_ARSIZE,
      x_rsc_1_0_ARLEN => hybrid_core_inst_x_rsc_1_0_ARLEN,
      x_rsc_1_0_ARADDR => hybrid_core_inst_x_rsc_1_0_ARADDR,
      x_rsc_1_0_ARID => x_rsc_1_0_ARID,
      x_rsc_1_0_BREADY => x_rsc_1_0_BREADY,
      x_rsc_1_0_BVALID => x_rsc_1_0_BVALID,
      x_rsc_1_0_BUSER => x_rsc_1_0_BUSER,
      x_rsc_1_0_BRESP => hybrid_core_inst_x_rsc_1_0_BRESP,
      x_rsc_1_0_BID => x_rsc_1_0_BID,
      x_rsc_1_0_WREADY => x_rsc_1_0_WREADY,
      x_rsc_1_0_WVALID => x_rsc_1_0_WVALID,
      x_rsc_1_0_WUSER => x_rsc_1_0_WUSER,
      x_rsc_1_0_WLAST => x_rsc_1_0_WLAST,
      x_rsc_1_0_WSTRB => hybrid_core_inst_x_rsc_1_0_WSTRB,
      x_rsc_1_0_WDATA => hybrid_core_inst_x_rsc_1_0_WDATA,
      x_rsc_1_0_AWREADY => x_rsc_1_0_AWREADY,
      x_rsc_1_0_AWVALID => x_rsc_1_0_AWVALID,
      x_rsc_1_0_AWUSER => x_rsc_1_0_AWUSER,
      x_rsc_1_0_AWREGION => hybrid_core_inst_x_rsc_1_0_AWREGION,
      x_rsc_1_0_AWQOS => hybrid_core_inst_x_rsc_1_0_AWQOS,
      x_rsc_1_0_AWPROT => hybrid_core_inst_x_rsc_1_0_AWPROT,
      x_rsc_1_0_AWCACHE => hybrid_core_inst_x_rsc_1_0_AWCACHE,
      x_rsc_1_0_AWLOCK => x_rsc_1_0_AWLOCK,
      x_rsc_1_0_AWBURST => hybrid_core_inst_x_rsc_1_0_AWBURST,
      x_rsc_1_0_AWSIZE => hybrid_core_inst_x_rsc_1_0_AWSIZE,
      x_rsc_1_0_AWLEN => hybrid_core_inst_x_rsc_1_0_AWLEN,
      x_rsc_1_0_AWADDR => hybrid_core_inst_x_rsc_1_0_AWADDR,
      x_rsc_1_0_AWID => x_rsc_1_0_AWID,
      x_rsc_triosy_1_0_lz => x_rsc_triosy_1_0_lz,
      x_rsc_2_0_s_tdone => x_rsc_2_0_s_tdone,
      x_rsc_2_0_tr_write_done => x_rsc_2_0_tr_write_done,
      x_rsc_2_0_RREADY => x_rsc_2_0_RREADY,
      x_rsc_2_0_RVALID => x_rsc_2_0_RVALID,
      x_rsc_2_0_RUSER => x_rsc_2_0_RUSER,
      x_rsc_2_0_RLAST => x_rsc_2_0_RLAST,
      x_rsc_2_0_RRESP => hybrid_core_inst_x_rsc_2_0_RRESP,
      x_rsc_2_0_RDATA => hybrid_core_inst_x_rsc_2_0_RDATA,
      x_rsc_2_0_RID => x_rsc_2_0_RID,
      x_rsc_2_0_ARREADY => x_rsc_2_0_ARREADY,
      x_rsc_2_0_ARVALID => x_rsc_2_0_ARVALID,
      x_rsc_2_0_ARUSER => x_rsc_2_0_ARUSER,
      x_rsc_2_0_ARREGION => hybrid_core_inst_x_rsc_2_0_ARREGION,
      x_rsc_2_0_ARQOS => hybrid_core_inst_x_rsc_2_0_ARQOS,
      x_rsc_2_0_ARPROT => hybrid_core_inst_x_rsc_2_0_ARPROT,
      x_rsc_2_0_ARCACHE => hybrid_core_inst_x_rsc_2_0_ARCACHE,
      x_rsc_2_0_ARLOCK => x_rsc_2_0_ARLOCK,
      x_rsc_2_0_ARBURST => hybrid_core_inst_x_rsc_2_0_ARBURST,
      x_rsc_2_0_ARSIZE => hybrid_core_inst_x_rsc_2_0_ARSIZE,
      x_rsc_2_0_ARLEN => hybrid_core_inst_x_rsc_2_0_ARLEN,
      x_rsc_2_0_ARADDR => hybrid_core_inst_x_rsc_2_0_ARADDR,
      x_rsc_2_0_ARID => x_rsc_2_0_ARID,
      x_rsc_2_0_BREADY => x_rsc_2_0_BREADY,
      x_rsc_2_0_BVALID => x_rsc_2_0_BVALID,
      x_rsc_2_0_BUSER => x_rsc_2_0_BUSER,
      x_rsc_2_0_BRESP => hybrid_core_inst_x_rsc_2_0_BRESP,
      x_rsc_2_0_BID => x_rsc_2_0_BID,
      x_rsc_2_0_WREADY => x_rsc_2_0_WREADY,
      x_rsc_2_0_WVALID => x_rsc_2_0_WVALID,
      x_rsc_2_0_WUSER => x_rsc_2_0_WUSER,
      x_rsc_2_0_WLAST => x_rsc_2_0_WLAST,
      x_rsc_2_0_WSTRB => hybrid_core_inst_x_rsc_2_0_WSTRB,
      x_rsc_2_0_WDATA => hybrid_core_inst_x_rsc_2_0_WDATA,
      x_rsc_2_0_AWREADY => x_rsc_2_0_AWREADY,
      x_rsc_2_0_AWVALID => x_rsc_2_0_AWVALID,
      x_rsc_2_0_AWUSER => x_rsc_2_0_AWUSER,
      x_rsc_2_0_AWREGION => hybrid_core_inst_x_rsc_2_0_AWREGION,
      x_rsc_2_0_AWQOS => hybrid_core_inst_x_rsc_2_0_AWQOS,
      x_rsc_2_0_AWPROT => hybrid_core_inst_x_rsc_2_0_AWPROT,
      x_rsc_2_0_AWCACHE => hybrid_core_inst_x_rsc_2_0_AWCACHE,
      x_rsc_2_0_AWLOCK => x_rsc_2_0_AWLOCK,
      x_rsc_2_0_AWBURST => hybrid_core_inst_x_rsc_2_0_AWBURST,
      x_rsc_2_0_AWSIZE => hybrid_core_inst_x_rsc_2_0_AWSIZE,
      x_rsc_2_0_AWLEN => hybrid_core_inst_x_rsc_2_0_AWLEN,
      x_rsc_2_0_AWADDR => hybrid_core_inst_x_rsc_2_0_AWADDR,
      x_rsc_2_0_AWID => x_rsc_2_0_AWID,
      x_rsc_triosy_2_0_lz => x_rsc_triosy_2_0_lz,
      x_rsc_3_0_s_tdone => x_rsc_3_0_s_tdone,
      x_rsc_3_0_tr_write_done => x_rsc_3_0_tr_write_done,
      x_rsc_3_0_RREADY => x_rsc_3_0_RREADY,
      x_rsc_3_0_RVALID => x_rsc_3_0_RVALID,
      x_rsc_3_0_RUSER => x_rsc_3_0_RUSER,
      x_rsc_3_0_RLAST => x_rsc_3_0_RLAST,
      x_rsc_3_0_RRESP => hybrid_core_inst_x_rsc_3_0_RRESP,
      x_rsc_3_0_RDATA => hybrid_core_inst_x_rsc_3_0_RDATA,
      x_rsc_3_0_RID => x_rsc_3_0_RID,
      x_rsc_3_0_ARREADY => x_rsc_3_0_ARREADY,
      x_rsc_3_0_ARVALID => x_rsc_3_0_ARVALID,
      x_rsc_3_0_ARUSER => x_rsc_3_0_ARUSER,
      x_rsc_3_0_ARREGION => hybrid_core_inst_x_rsc_3_0_ARREGION,
      x_rsc_3_0_ARQOS => hybrid_core_inst_x_rsc_3_0_ARQOS,
      x_rsc_3_0_ARPROT => hybrid_core_inst_x_rsc_3_0_ARPROT,
      x_rsc_3_0_ARCACHE => hybrid_core_inst_x_rsc_3_0_ARCACHE,
      x_rsc_3_0_ARLOCK => x_rsc_3_0_ARLOCK,
      x_rsc_3_0_ARBURST => hybrid_core_inst_x_rsc_3_0_ARBURST,
      x_rsc_3_0_ARSIZE => hybrid_core_inst_x_rsc_3_0_ARSIZE,
      x_rsc_3_0_ARLEN => hybrid_core_inst_x_rsc_3_0_ARLEN,
      x_rsc_3_0_ARADDR => hybrid_core_inst_x_rsc_3_0_ARADDR,
      x_rsc_3_0_ARID => x_rsc_3_0_ARID,
      x_rsc_3_0_BREADY => x_rsc_3_0_BREADY,
      x_rsc_3_0_BVALID => x_rsc_3_0_BVALID,
      x_rsc_3_0_BUSER => x_rsc_3_0_BUSER,
      x_rsc_3_0_BRESP => hybrid_core_inst_x_rsc_3_0_BRESP,
      x_rsc_3_0_BID => x_rsc_3_0_BID,
      x_rsc_3_0_WREADY => x_rsc_3_0_WREADY,
      x_rsc_3_0_WVALID => x_rsc_3_0_WVALID,
      x_rsc_3_0_WUSER => x_rsc_3_0_WUSER,
      x_rsc_3_0_WLAST => x_rsc_3_0_WLAST,
      x_rsc_3_0_WSTRB => hybrid_core_inst_x_rsc_3_0_WSTRB,
      x_rsc_3_0_WDATA => hybrid_core_inst_x_rsc_3_0_WDATA,
      x_rsc_3_0_AWREADY => x_rsc_3_0_AWREADY,
      x_rsc_3_0_AWVALID => x_rsc_3_0_AWVALID,
      x_rsc_3_0_AWUSER => x_rsc_3_0_AWUSER,
      x_rsc_3_0_AWREGION => hybrid_core_inst_x_rsc_3_0_AWREGION,
      x_rsc_3_0_AWQOS => hybrid_core_inst_x_rsc_3_0_AWQOS,
      x_rsc_3_0_AWPROT => hybrid_core_inst_x_rsc_3_0_AWPROT,
      x_rsc_3_0_AWCACHE => hybrid_core_inst_x_rsc_3_0_AWCACHE,
      x_rsc_3_0_AWLOCK => x_rsc_3_0_AWLOCK,
      x_rsc_3_0_AWBURST => hybrid_core_inst_x_rsc_3_0_AWBURST,
      x_rsc_3_0_AWSIZE => hybrid_core_inst_x_rsc_3_0_AWSIZE,
      x_rsc_3_0_AWLEN => hybrid_core_inst_x_rsc_3_0_AWLEN,
      x_rsc_3_0_AWADDR => hybrid_core_inst_x_rsc_3_0_AWADDR,
      x_rsc_3_0_AWID => x_rsc_3_0_AWID,
      x_rsc_triosy_3_0_lz => x_rsc_triosy_3_0_lz,
      x_rsc_4_0_s_tdone => x_rsc_4_0_s_tdone,
      x_rsc_4_0_tr_write_done => x_rsc_4_0_tr_write_done,
      x_rsc_4_0_RREADY => x_rsc_4_0_RREADY,
      x_rsc_4_0_RVALID => x_rsc_4_0_RVALID,
      x_rsc_4_0_RUSER => x_rsc_4_0_RUSER,
      x_rsc_4_0_RLAST => x_rsc_4_0_RLAST,
      x_rsc_4_0_RRESP => hybrid_core_inst_x_rsc_4_0_RRESP,
      x_rsc_4_0_RDATA => hybrid_core_inst_x_rsc_4_0_RDATA,
      x_rsc_4_0_RID => x_rsc_4_0_RID,
      x_rsc_4_0_ARREADY => x_rsc_4_0_ARREADY,
      x_rsc_4_0_ARVALID => x_rsc_4_0_ARVALID,
      x_rsc_4_0_ARUSER => x_rsc_4_0_ARUSER,
      x_rsc_4_0_ARREGION => hybrid_core_inst_x_rsc_4_0_ARREGION,
      x_rsc_4_0_ARQOS => hybrid_core_inst_x_rsc_4_0_ARQOS,
      x_rsc_4_0_ARPROT => hybrid_core_inst_x_rsc_4_0_ARPROT,
      x_rsc_4_0_ARCACHE => hybrid_core_inst_x_rsc_4_0_ARCACHE,
      x_rsc_4_0_ARLOCK => x_rsc_4_0_ARLOCK,
      x_rsc_4_0_ARBURST => hybrid_core_inst_x_rsc_4_0_ARBURST,
      x_rsc_4_0_ARSIZE => hybrid_core_inst_x_rsc_4_0_ARSIZE,
      x_rsc_4_0_ARLEN => hybrid_core_inst_x_rsc_4_0_ARLEN,
      x_rsc_4_0_ARADDR => hybrid_core_inst_x_rsc_4_0_ARADDR,
      x_rsc_4_0_ARID => x_rsc_4_0_ARID,
      x_rsc_4_0_BREADY => x_rsc_4_0_BREADY,
      x_rsc_4_0_BVALID => x_rsc_4_0_BVALID,
      x_rsc_4_0_BUSER => x_rsc_4_0_BUSER,
      x_rsc_4_0_BRESP => hybrid_core_inst_x_rsc_4_0_BRESP,
      x_rsc_4_0_BID => x_rsc_4_0_BID,
      x_rsc_4_0_WREADY => x_rsc_4_0_WREADY,
      x_rsc_4_0_WVALID => x_rsc_4_0_WVALID,
      x_rsc_4_0_WUSER => x_rsc_4_0_WUSER,
      x_rsc_4_0_WLAST => x_rsc_4_0_WLAST,
      x_rsc_4_0_WSTRB => hybrid_core_inst_x_rsc_4_0_WSTRB,
      x_rsc_4_0_WDATA => hybrid_core_inst_x_rsc_4_0_WDATA,
      x_rsc_4_0_AWREADY => x_rsc_4_0_AWREADY,
      x_rsc_4_0_AWVALID => x_rsc_4_0_AWVALID,
      x_rsc_4_0_AWUSER => x_rsc_4_0_AWUSER,
      x_rsc_4_0_AWREGION => hybrid_core_inst_x_rsc_4_0_AWREGION,
      x_rsc_4_0_AWQOS => hybrid_core_inst_x_rsc_4_0_AWQOS,
      x_rsc_4_0_AWPROT => hybrid_core_inst_x_rsc_4_0_AWPROT,
      x_rsc_4_0_AWCACHE => hybrid_core_inst_x_rsc_4_0_AWCACHE,
      x_rsc_4_0_AWLOCK => x_rsc_4_0_AWLOCK,
      x_rsc_4_0_AWBURST => hybrid_core_inst_x_rsc_4_0_AWBURST,
      x_rsc_4_0_AWSIZE => hybrid_core_inst_x_rsc_4_0_AWSIZE,
      x_rsc_4_0_AWLEN => hybrid_core_inst_x_rsc_4_0_AWLEN,
      x_rsc_4_0_AWADDR => hybrid_core_inst_x_rsc_4_0_AWADDR,
      x_rsc_4_0_AWID => x_rsc_4_0_AWID,
      x_rsc_triosy_4_0_lz => x_rsc_triosy_4_0_lz,
      x_rsc_5_0_s_tdone => x_rsc_5_0_s_tdone,
      x_rsc_5_0_tr_write_done => x_rsc_5_0_tr_write_done,
      x_rsc_5_0_RREADY => x_rsc_5_0_RREADY,
      x_rsc_5_0_RVALID => x_rsc_5_0_RVALID,
      x_rsc_5_0_RUSER => x_rsc_5_0_RUSER,
      x_rsc_5_0_RLAST => x_rsc_5_0_RLAST,
      x_rsc_5_0_RRESP => hybrid_core_inst_x_rsc_5_0_RRESP,
      x_rsc_5_0_RDATA => hybrid_core_inst_x_rsc_5_0_RDATA,
      x_rsc_5_0_RID => x_rsc_5_0_RID,
      x_rsc_5_0_ARREADY => x_rsc_5_0_ARREADY,
      x_rsc_5_0_ARVALID => x_rsc_5_0_ARVALID,
      x_rsc_5_0_ARUSER => x_rsc_5_0_ARUSER,
      x_rsc_5_0_ARREGION => hybrid_core_inst_x_rsc_5_0_ARREGION,
      x_rsc_5_0_ARQOS => hybrid_core_inst_x_rsc_5_0_ARQOS,
      x_rsc_5_0_ARPROT => hybrid_core_inst_x_rsc_5_0_ARPROT,
      x_rsc_5_0_ARCACHE => hybrid_core_inst_x_rsc_5_0_ARCACHE,
      x_rsc_5_0_ARLOCK => x_rsc_5_0_ARLOCK,
      x_rsc_5_0_ARBURST => hybrid_core_inst_x_rsc_5_0_ARBURST,
      x_rsc_5_0_ARSIZE => hybrid_core_inst_x_rsc_5_0_ARSIZE,
      x_rsc_5_0_ARLEN => hybrid_core_inst_x_rsc_5_0_ARLEN,
      x_rsc_5_0_ARADDR => hybrid_core_inst_x_rsc_5_0_ARADDR,
      x_rsc_5_0_ARID => x_rsc_5_0_ARID,
      x_rsc_5_0_BREADY => x_rsc_5_0_BREADY,
      x_rsc_5_0_BVALID => x_rsc_5_0_BVALID,
      x_rsc_5_0_BUSER => x_rsc_5_0_BUSER,
      x_rsc_5_0_BRESP => hybrid_core_inst_x_rsc_5_0_BRESP,
      x_rsc_5_0_BID => x_rsc_5_0_BID,
      x_rsc_5_0_WREADY => x_rsc_5_0_WREADY,
      x_rsc_5_0_WVALID => x_rsc_5_0_WVALID,
      x_rsc_5_0_WUSER => x_rsc_5_0_WUSER,
      x_rsc_5_0_WLAST => x_rsc_5_0_WLAST,
      x_rsc_5_0_WSTRB => hybrid_core_inst_x_rsc_5_0_WSTRB,
      x_rsc_5_0_WDATA => hybrid_core_inst_x_rsc_5_0_WDATA,
      x_rsc_5_0_AWREADY => x_rsc_5_0_AWREADY,
      x_rsc_5_0_AWVALID => x_rsc_5_0_AWVALID,
      x_rsc_5_0_AWUSER => x_rsc_5_0_AWUSER,
      x_rsc_5_0_AWREGION => hybrid_core_inst_x_rsc_5_0_AWREGION,
      x_rsc_5_0_AWQOS => hybrid_core_inst_x_rsc_5_0_AWQOS,
      x_rsc_5_0_AWPROT => hybrid_core_inst_x_rsc_5_0_AWPROT,
      x_rsc_5_0_AWCACHE => hybrid_core_inst_x_rsc_5_0_AWCACHE,
      x_rsc_5_0_AWLOCK => x_rsc_5_0_AWLOCK,
      x_rsc_5_0_AWBURST => hybrid_core_inst_x_rsc_5_0_AWBURST,
      x_rsc_5_0_AWSIZE => hybrid_core_inst_x_rsc_5_0_AWSIZE,
      x_rsc_5_0_AWLEN => hybrid_core_inst_x_rsc_5_0_AWLEN,
      x_rsc_5_0_AWADDR => hybrid_core_inst_x_rsc_5_0_AWADDR,
      x_rsc_5_0_AWID => x_rsc_5_0_AWID,
      x_rsc_triosy_5_0_lz => x_rsc_triosy_5_0_lz,
      x_rsc_6_0_s_tdone => x_rsc_6_0_s_tdone,
      x_rsc_6_0_tr_write_done => x_rsc_6_0_tr_write_done,
      x_rsc_6_0_RREADY => x_rsc_6_0_RREADY,
      x_rsc_6_0_RVALID => x_rsc_6_0_RVALID,
      x_rsc_6_0_RUSER => x_rsc_6_0_RUSER,
      x_rsc_6_0_RLAST => x_rsc_6_0_RLAST,
      x_rsc_6_0_RRESP => hybrid_core_inst_x_rsc_6_0_RRESP,
      x_rsc_6_0_RDATA => hybrid_core_inst_x_rsc_6_0_RDATA,
      x_rsc_6_0_RID => x_rsc_6_0_RID,
      x_rsc_6_0_ARREADY => x_rsc_6_0_ARREADY,
      x_rsc_6_0_ARVALID => x_rsc_6_0_ARVALID,
      x_rsc_6_0_ARUSER => x_rsc_6_0_ARUSER,
      x_rsc_6_0_ARREGION => hybrid_core_inst_x_rsc_6_0_ARREGION,
      x_rsc_6_0_ARQOS => hybrid_core_inst_x_rsc_6_0_ARQOS,
      x_rsc_6_0_ARPROT => hybrid_core_inst_x_rsc_6_0_ARPROT,
      x_rsc_6_0_ARCACHE => hybrid_core_inst_x_rsc_6_0_ARCACHE,
      x_rsc_6_0_ARLOCK => x_rsc_6_0_ARLOCK,
      x_rsc_6_0_ARBURST => hybrid_core_inst_x_rsc_6_0_ARBURST,
      x_rsc_6_0_ARSIZE => hybrid_core_inst_x_rsc_6_0_ARSIZE,
      x_rsc_6_0_ARLEN => hybrid_core_inst_x_rsc_6_0_ARLEN,
      x_rsc_6_0_ARADDR => hybrid_core_inst_x_rsc_6_0_ARADDR,
      x_rsc_6_0_ARID => x_rsc_6_0_ARID,
      x_rsc_6_0_BREADY => x_rsc_6_0_BREADY,
      x_rsc_6_0_BVALID => x_rsc_6_0_BVALID,
      x_rsc_6_0_BUSER => x_rsc_6_0_BUSER,
      x_rsc_6_0_BRESP => hybrid_core_inst_x_rsc_6_0_BRESP,
      x_rsc_6_0_BID => x_rsc_6_0_BID,
      x_rsc_6_0_WREADY => x_rsc_6_0_WREADY,
      x_rsc_6_0_WVALID => x_rsc_6_0_WVALID,
      x_rsc_6_0_WUSER => x_rsc_6_0_WUSER,
      x_rsc_6_0_WLAST => x_rsc_6_0_WLAST,
      x_rsc_6_0_WSTRB => hybrid_core_inst_x_rsc_6_0_WSTRB,
      x_rsc_6_0_WDATA => hybrid_core_inst_x_rsc_6_0_WDATA,
      x_rsc_6_0_AWREADY => x_rsc_6_0_AWREADY,
      x_rsc_6_0_AWVALID => x_rsc_6_0_AWVALID,
      x_rsc_6_0_AWUSER => x_rsc_6_0_AWUSER,
      x_rsc_6_0_AWREGION => hybrid_core_inst_x_rsc_6_0_AWREGION,
      x_rsc_6_0_AWQOS => hybrid_core_inst_x_rsc_6_0_AWQOS,
      x_rsc_6_0_AWPROT => hybrid_core_inst_x_rsc_6_0_AWPROT,
      x_rsc_6_0_AWCACHE => hybrid_core_inst_x_rsc_6_0_AWCACHE,
      x_rsc_6_0_AWLOCK => x_rsc_6_0_AWLOCK,
      x_rsc_6_0_AWBURST => hybrid_core_inst_x_rsc_6_0_AWBURST,
      x_rsc_6_0_AWSIZE => hybrid_core_inst_x_rsc_6_0_AWSIZE,
      x_rsc_6_0_AWLEN => hybrid_core_inst_x_rsc_6_0_AWLEN,
      x_rsc_6_0_AWADDR => hybrid_core_inst_x_rsc_6_0_AWADDR,
      x_rsc_6_0_AWID => x_rsc_6_0_AWID,
      x_rsc_triosy_6_0_lz => x_rsc_triosy_6_0_lz,
      x_rsc_7_0_s_tdone => x_rsc_7_0_s_tdone,
      x_rsc_7_0_tr_write_done => x_rsc_7_0_tr_write_done,
      x_rsc_7_0_RREADY => x_rsc_7_0_RREADY,
      x_rsc_7_0_RVALID => x_rsc_7_0_RVALID,
      x_rsc_7_0_RUSER => x_rsc_7_0_RUSER,
      x_rsc_7_0_RLAST => x_rsc_7_0_RLAST,
      x_rsc_7_0_RRESP => hybrid_core_inst_x_rsc_7_0_RRESP,
      x_rsc_7_0_RDATA => hybrid_core_inst_x_rsc_7_0_RDATA,
      x_rsc_7_0_RID => x_rsc_7_0_RID,
      x_rsc_7_0_ARREADY => x_rsc_7_0_ARREADY,
      x_rsc_7_0_ARVALID => x_rsc_7_0_ARVALID,
      x_rsc_7_0_ARUSER => x_rsc_7_0_ARUSER,
      x_rsc_7_0_ARREGION => hybrid_core_inst_x_rsc_7_0_ARREGION,
      x_rsc_7_0_ARQOS => hybrid_core_inst_x_rsc_7_0_ARQOS,
      x_rsc_7_0_ARPROT => hybrid_core_inst_x_rsc_7_0_ARPROT,
      x_rsc_7_0_ARCACHE => hybrid_core_inst_x_rsc_7_0_ARCACHE,
      x_rsc_7_0_ARLOCK => x_rsc_7_0_ARLOCK,
      x_rsc_7_0_ARBURST => hybrid_core_inst_x_rsc_7_0_ARBURST,
      x_rsc_7_0_ARSIZE => hybrid_core_inst_x_rsc_7_0_ARSIZE,
      x_rsc_7_0_ARLEN => hybrid_core_inst_x_rsc_7_0_ARLEN,
      x_rsc_7_0_ARADDR => hybrid_core_inst_x_rsc_7_0_ARADDR,
      x_rsc_7_0_ARID => x_rsc_7_0_ARID,
      x_rsc_7_0_BREADY => x_rsc_7_0_BREADY,
      x_rsc_7_0_BVALID => x_rsc_7_0_BVALID,
      x_rsc_7_0_BUSER => x_rsc_7_0_BUSER,
      x_rsc_7_0_BRESP => hybrid_core_inst_x_rsc_7_0_BRESP,
      x_rsc_7_0_BID => x_rsc_7_0_BID,
      x_rsc_7_0_WREADY => x_rsc_7_0_WREADY,
      x_rsc_7_0_WVALID => x_rsc_7_0_WVALID,
      x_rsc_7_0_WUSER => x_rsc_7_0_WUSER,
      x_rsc_7_0_WLAST => x_rsc_7_0_WLAST,
      x_rsc_7_0_WSTRB => hybrid_core_inst_x_rsc_7_0_WSTRB,
      x_rsc_7_0_WDATA => hybrid_core_inst_x_rsc_7_0_WDATA,
      x_rsc_7_0_AWREADY => x_rsc_7_0_AWREADY,
      x_rsc_7_0_AWVALID => x_rsc_7_0_AWVALID,
      x_rsc_7_0_AWUSER => x_rsc_7_0_AWUSER,
      x_rsc_7_0_AWREGION => hybrid_core_inst_x_rsc_7_0_AWREGION,
      x_rsc_7_0_AWQOS => hybrid_core_inst_x_rsc_7_0_AWQOS,
      x_rsc_7_0_AWPROT => hybrid_core_inst_x_rsc_7_0_AWPROT,
      x_rsc_7_0_AWCACHE => hybrid_core_inst_x_rsc_7_0_AWCACHE,
      x_rsc_7_0_AWLOCK => x_rsc_7_0_AWLOCK,
      x_rsc_7_0_AWBURST => hybrid_core_inst_x_rsc_7_0_AWBURST,
      x_rsc_7_0_AWSIZE => hybrid_core_inst_x_rsc_7_0_AWSIZE,
      x_rsc_7_0_AWLEN => hybrid_core_inst_x_rsc_7_0_AWLEN,
      x_rsc_7_0_AWADDR => hybrid_core_inst_x_rsc_7_0_AWADDR,
      x_rsc_7_0_AWID => x_rsc_7_0_AWID,
      x_rsc_triosy_7_0_lz => x_rsc_triosy_7_0_lz,
      x_rsc_8_0_s_tdone => x_rsc_8_0_s_tdone,
      x_rsc_8_0_tr_write_done => x_rsc_8_0_tr_write_done,
      x_rsc_8_0_RREADY => x_rsc_8_0_RREADY,
      x_rsc_8_0_RVALID => x_rsc_8_0_RVALID,
      x_rsc_8_0_RUSER => x_rsc_8_0_RUSER,
      x_rsc_8_0_RLAST => x_rsc_8_0_RLAST,
      x_rsc_8_0_RRESP => hybrid_core_inst_x_rsc_8_0_RRESP,
      x_rsc_8_0_RDATA => hybrid_core_inst_x_rsc_8_0_RDATA,
      x_rsc_8_0_RID => x_rsc_8_0_RID,
      x_rsc_8_0_ARREADY => x_rsc_8_0_ARREADY,
      x_rsc_8_0_ARVALID => x_rsc_8_0_ARVALID,
      x_rsc_8_0_ARUSER => x_rsc_8_0_ARUSER,
      x_rsc_8_0_ARREGION => hybrid_core_inst_x_rsc_8_0_ARREGION,
      x_rsc_8_0_ARQOS => hybrid_core_inst_x_rsc_8_0_ARQOS,
      x_rsc_8_0_ARPROT => hybrid_core_inst_x_rsc_8_0_ARPROT,
      x_rsc_8_0_ARCACHE => hybrid_core_inst_x_rsc_8_0_ARCACHE,
      x_rsc_8_0_ARLOCK => x_rsc_8_0_ARLOCK,
      x_rsc_8_0_ARBURST => hybrid_core_inst_x_rsc_8_0_ARBURST,
      x_rsc_8_0_ARSIZE => hybrid_core_inst_x_rsc_8_0_ARSIZE,
      x_rsc_8_0_ARLEN => hybrid_core_inst_x_rsc_8_0_ARLEN,
      x_rsc_8_0_ARADDR => hybrid_core_inst_x_rsc_8_0_ARADDR,
      x_rsc_8_0_ARID => x_rsc_8_0_ARID,
      x_rsc_8_0_BREADY => x_rsc_8_0_BREADY,
      x_rsc_8_0_BVALID => x_rsc_8_0_BVALID,
      x_rsc_8_0_BUSER => x_rsc_8_0_BUSER,
      x_rsc_8_0_BRESP => hybrid_core_inst_x_rsc_8_0_BRESP,
      x_rsc_8_0_BID => x_rsc_8_0_BID,
      x_rsc_8_0_WREADY => x_rsc_8_0_WREADY,
      x_rsc_8_0_WVALID => x_rsc_8_0_WVALID,
      x_rsc_8_0_WUSER => x_rsc_8_0_WUSER,
      x_rsc_8_0_WLAST => x_rsc_8_0_WLAST,
      x_rsc_8_0_WSTRB => hybrid_core_inst_x_rsc_8_0_WSTRB,
      x_rsc_8_0_WDATA => hybrid_core_inst_x_rsc_8_0_WDATA,
      x_rsc_8_0_AWREADY => x_rsc_8_0_AWREADY,
      x_rsc_8_0_AWVALID => x_rsc_8_0_AWVALID,
      x_rsc_8_0_AWUSER => x_rsc_8_0_AWUSER,
      x_rsc_8_0_AWREGION => hybrid_core_inst_x_rsc_8_0_AWREGION,
      x_rsc_8_0_AWQOS => hybrid_core_inst_x_rsc_8_0_AWQOS,
      x_rsc_8_0_AWPROT => hybrid_core_inst_x_rsc_8_0_AWPROT,
      x_rsc_8_0_AWCACHE => hybrid_core_inst_x_rsc_8_0_AWCACHE,
      x_rsc_8_0_AWLOCK => x_rsc_8_0_AWLOCK,
      x_rsc_8_0_AWBURST => hybrid_core_inst_x_rsc_8_0_AWBURST,
      x_rsc_8_0_AWSIZE => hybrid_core_inst_x_rsc_8_0_AWSIZE,
      x_rsc_8_0_AWLEN => hybrid_core_inst_x_rsc_8_0_AWLEN,
      x_rsc_8_0_AWADDR => hybrid_core_inst_x_rsc_8_0_AWADDR,
      x_rsc_8_0_AWID => x_rsc_8_0_AWID,
      x_rsc_triosy_8_0_lz => x_rsc_triosy_8_0_lz,
      x_rsc_9_0_s_tdone => x_rsc_9_0_s_tdone,
      x_rsc_9_0_tr_write_done => x_rsc_9_0_tr_write_done,
      x_rsc_9_0_RREADY => x_rsc_9_0_RREADY,
      x_rsc_9_0_RVALID => x_rsc_9_0_RVALID,
      x_rsc_9_0_RUSER => x_rsc_9_0_RUSER,
      x_rsc_9_0_RLAST => x_rsc_9_0_RLAST,
      x_rsc_9_0_RRESP => hybrid_core_inst_x_rsc_9_0_RRESP,
      x_rsc_9_0_RDATA => hybrid_core_inst_x_rsc_9_0_RDATA,
      x_rsc_9_0_RID => x_rsc_9_0_RID,
      x_rsc_9_0_ARREADY => x_rsc_9_0_ARREADY,
      x_rsc_9_0_ARVALID => x_rsc_9_0_ARVALID,
      x_rsc_9_0_ARUSER => x_rsc_9_0_ARUSER,
      x_rsc_9_0_ARREGION => hybrid_core_inst_x_rsc_9_0_ARREGION,
      x_rsc_9_0_ARQOS => hybrid_core_inst_x_rsc_9_0_ARQOS,
      x_rsc_9_0_ARPROT => hybrid_core_inst_x_rsc_9_0_ARPROT,
      x_rsc_9_0_ARCACHE => hybrid_core_inst_x_rsc_9_0_ARCACHE,
      x_rsc_9_0_ARLOCK => x_rsc_9_0_ARLOCK,
      x_rsc_9_0_ARBURST => hybrid_core_inst_x_rsc_9_0_ARBURST,
      x_rsc_9_0_ARSIZE => hybrid_core_inst_x_rsc_9_0_ARSIZE,
      x_rsc_9_0_ARLEN => hybrid_core_inst_x_rsc_9_0_ARLEN,
      x_rsc_9_0_ARADDR => hybrid_core_inst_x_rsc_9_0_ARADDR,
      x_rsc_9_0_ARID => x_rsc_9_0_ARID,
      x_rsc_9_0_BREADY => x_rsc_9_0_BREADY,
      x_rsc_9_0_BVALID => x_rsc_9_0_BVALID,
      x_rsc_9_0_BUSER => x_rsc_9_0_BUSER,
      x_rsc_9_0_BRESP => hybrid_core_inst_x_rsc_9_0_BRESP,
      x_rsc_9_0_BID => x_rsc_9_0_BID,
      x_rsc_9_0_WREADY => x_rsc_9_0_WREADY,
      x_rsc_9_0_WVALID => x_rsc_9_0_WVALID,
      x_rsc_9_0_WUSER => x_rsc_9_0_WUSER,
      x_rsc_9_0_WLAST => x_rsc_9_0_WLAST,
      x_rsc_9_0_WSTRB => hybrid_core_inst_x_rsc_9_0_WSTRB,
      x_rsc_9_0_WDATA => hybrid_core_inst_x_rsc_9_0_WDATA,
      x_rsc_9_0_AWREADY => x_rsc_9_0_AWREADY,
      x_rsc_9_0_AWVALID => x_rsc_9_0_AWVALID,
      x_rsc_9_0_AWUSER => x_rsc_9_0_AWUSER,
      x_rsc_9_0_AWREGION => hybrid_core_inst_x_rsc_9_0_AWREGION,
      x_rsc_9_0_AWQOS => hybrid_core_inst_x_rsc_9_0_AWQOS,
      x_rsc_9_0_AWPROT => hybrid_core_inst_x_rsc_9_0_AWPROT,
      x_rsc_9_0_AWCACHE => hybrid_core_inst_x_rsc_9_0_AWCACHE,
      x_rsc_9_0_AWLOCK => x_rsc_9_0_AWLOCK,
      x_rsc_9_0_AWBURST => hybrid_core_inst_x_rsc_9_0_AWBURST,
      x_rsc_9_0_AWSIZE => hybrid_core_inst_x_rsc_9_0_AWSIZE,
      x_rsc_9_0_AWLEN => hybrid_core_inst_x_rsc_9_0_AWLEN,
      x_rsc_9_0_AWADDR => hybrid_core_inst_x_rsc_9_0_AWADDR,
      x_rsc_9_0_AWID => x_rsc_9_0_AWID,
      x_rsc_triosy_9_0_lz => x_rsc_triosy_9_0_lz,
      x_rsc_10_0_s_tdone => x_rsc_10_0_s_tdone,
      x_rsc_10_0_tr_write_done => x_rsc_10_0_tr_write_done,
      x_rsc_10_0_RREADY => x_rsc_10_0_RREADY,
      x_rsc_10_0_RVALID => x_rsc_10_0_RVALID,
      x_rsc_10_0_RUSER => x_rsc_10_0_RUSER,
      x_rsc_10_0_RLAST => x_rsc_10_0_RLAST,
      x_rsc_10_0_RRESP => hybrid_core_inst_x_rsc_10_0_RRESP,
      x_rsc_10_0_RDATA => hybrid_core_inst_x_rsc_10_0_RDATA,
      x_rsc_10_0_RID => x_rsc_10_0_RID,
      x_rsc_10_0_ARREADY => x_rsc_10_0_ARREADY,
      x_rsc_10_0_ARVALID => x_rsc_10_0_ARVALID,
      x_rsc_10_0_ARUSER => x_rsc_10_0_ARUSER,
      x_rsc_10_0_ARREGION => hybrid_core_inst_x_rsc_10_0_ARREGION,
      x_rsc_10_0_ARQOS => hybrid_core_inst_x_rsc_10_0_ARQOS,
      x_rsc_10_0_ARPROT => hybrid_core_inst_x_rsc_10_0_ARPROT,
      x_rsc_10_0_ARCACHE => hybrid_core_inst_x_rsc_10_0_ARCACHE,
      x_rsc_10_0_ARLOCK => x_rsc_10_0_ARLOCK,
      x_rsc_10_0_ARBURST => hybrid_core_inst_x_rsc_10_0_ARBURST,
      x_rsc_10_0_ARSIZE => hybrid_core_inst_x_rsc_10_0_ARSIZE,
      x_rsc_10_0_ARLEN => hybrid_core_inst_x_rsc_10_0_ARLEN,
      x_rsc_10_0_ARADDR => hybrid_core_inst_x_rsc_10_0_ARADDR,
      x_rsc_10_0_ARID => x_rsc_10_0_ARID,
      x_rsc_10_0_BREADY => x_rsc_10_0_BREADY,
      x_rsc_10_0_BVALID => x_rsc_10_0_BVALID,
      x_rsc_10_0_BUSER => x_rsc_10_0_BUSER,
      x_rsc_10_0_BRESP => hybrid_core_inst_x_rsc_10_0_BRESP,
      x_rsc_10_0_BID => x_rsc_10_0_BID,
      x_rsc_10_0_WREADY => x_rsc_10_0_WREADY,
      x_rsc_10_0_WVALID => x_rsc_10_0_WVALID,
      x_rsc_10_0_WUSER => x_rsc_10_0_WUSER,
      x_rsc_10_0_WLAST => x_rsc_10_0_WLAST,
      x_rsc_10_0_WSTRB => hybrid_core_inst_x_rsc_10_0_WSTRB,
      x_rsc_10_0_WDATA => hybrid_core_inst_x_rsc_10_0_WDATA,
      x_rsc_10_0_AWREADY => x_rsc_10_0_AWREADY,
      x_rsc_10_0_AWVALID => x_rsc_10_0_AWVALID,
      x_rsc_10_0_AWUSER => x_rsc_10_0_AWUSER,
      x_rsc_10_0_AWREGION => hybrid_core_inst_x_rsc_10_0_AWREGION,
      x_rsc_10_0_AWQOS => hybrid_core_inst_x_rsc_10_0_AWQOS,
      x_rsc_10_0_AWPROT => hybrid_core_inst_x_rsc_10_0_AWPROT,
      x_rsc_10_0_AWCACHE => hybrid_core_inst_x_rsc_10_0_AWCACHE,
      x_rsc_10_0_AWLOCK => x_rsc_10_0_AWLOCK,
      x_rsc_10_0_AWBURST => hybrid_core_inst_x_rsc_10_0_AWBURST,
      x_rsc_10_0_AWSIZE => hybrid_core_inst_x_rsc_10_0_AWSIZE,
      x_rsc_10_0_AWLEN => hybrid_core_inst_x_rsc_10_0_AWLEN,
      x_rsc_10_0_AWADDR => hybrid_core_inst_x_rsc_10_0_AWADDR,
      x_rsc_10_0_AWID => x_rsc_10_0_AWID,
      x_rsc_triosy_10_0_lz => x_rsc_triosy_10_0_lz,
      x_rsc_11_0_s_tdone => x_rsc_11_0_s_tdone,
      x_rsc_11_0_tr_write_done => x_rsc_11_0_tr_write_done,
      x_rsc_11_0_RREADY => x_rsc_11_0_RREADY,
      x_rsc_11_0_RVALID => x_rsc_11_0_RVALID,
      x_rsc_11_0_RUSER => x_rsc_11_0_RUSER,
      x_rsc_11_0_RLAST => x_rsc_11_0_RLAST,
      x_rsc_11_0_RRESP => hybrid_core_inst_x_rsc_11_0_RRESP,
      x_rsc_11_0_RDATA => hybrid_core_inst_x_rsc_11_0_RDATA,
      x_rsc_11_0_RID => x_rsc_11_0_RID,
      x_rsc_11_0_ARREADY => x_rsc_11_0_ARREADY,
      x_rsc_11_0_ARVALID => x_rsc_11_0_ARVALID,
      x_rsc_11_0_ARUSER => x_rsc_11_0_ARUSER,
      x_rsc_11_0_ARREGION => hybrid_core_inst_x_rsc_11_0_ARREGION,
      x_rsc_11_0_ARQOS => hybrid_core_inst_x_rsc_11_0_ARQOS,
      x_rsc_11_0_ARPROT => hybrid_core_inst_x_rsc_11_0_ARPROT,
      x_rsc_11_0_ARCACHE => hybrid_core_inst_x_rsc_11_0_ARCACHE,
      x_rsc_11_0_ARLOCK => x_rsc_11_0_ARLOCK,
      x_rsc_11_0_ARBURST => hybrid_core_inst_x_rsc_11_0_ARBURST,
      x_rsc_11_0_ARSIZE => hybrid_core_inst_x_rsc_11_0_ARSIZE,
      x_rsc_11_0_ARLEN => hybrid_core_inst_x_rsc_11_0_ARLEN,
      x_rsc_11_0_ARADDR => hybrid_core_inst_x_rsc_11_0_ARADDR,
      x_rsc_11_0_ARID => x_rsc_11_0_ARID,
      x_rsc_11_0_BREADY => x_rsc_11_0_BREADY,
      x_rsc_11_0_BVALID => x_rsc_11_0_BVALID,
      x_rsc_11_0_BUSER => x_rsc_11_0_BUSER,
      x_rsc_11_0_BRESP => hybrid_core_inst_x_rsc_11_0_BRESP,
      x_rsc_11_0_BID => x_rsc_11_0_BID,
      x_rsc_11_0_WREADY => x_rsc_11_0_WREADY,
      x_rsc_11_0_WVALID => x_rsc_11_0_WVALID,
      x_rsc_11_0_WUSER => x_rsc_11_0_WUSER,
      x_rsc_11_0_WLAST => x_rsc_11_0_WLAST,
      x_rsc_11_0_WSTRB => hybrid_core_inst_x_rsc_11_0_WSTRB,
      x_rsc_11_0_WDATA => hybrid_core_inst_x_rsc_11_0_WDATA,
      x_rsc_11_0_AWREADY => x_rsc_11_0_AWREADY,
      x_rsc_11_0_AWVALID => x_rsc_11_0_AWVALID,
      x_rsc_11_0_AWUSER => x_rsc_11_0_AWUSER,
      x_rsc_11_0_AWREGION => hybrid_core_inst_x_rsc_11_0_AWREGION,
      x_rsc_11_0_AWQOS => hybrid_core_inst_x_rsc_11_0_AWQOS,
      x_rsc_11_0_AWPROT => hybrid_core_inst_x_rsc_11_0_AWPROT,
      x_rsc_11_0_AWCACHE => hybrid_core_inst_x_rsc_11_0_AWCACHE,
      x_rsc_11_0_AWLOCK => x_rsc_11_0_AWLOCK,
      x_rsc_11_0_AWBURST => hybrid_core_inst_x_rsc_11_0_AWBURST,
      x_rsc_11_0_AWSIZE => hybrid_core_inst_x_rsc_11_0_AWSIZE,
      x_rsc_11_0_AWLEN => hybrid_core_inst_x_rsc_11_0_AWLEN,
      x_rsc_11_0_AWADDR => hybrid_core_inst_x_rsc_11_0_AWADDR,
      x_rsc_11_0_AWID => x_rsc_11_0_AWID,
      x_rsc_triosy_11_0_lz => x_rsc_triosy_11_0_lz,
      x_rsc_12_0_s_tdone => x_rsc_12_0_s_tdone,
      x_rsc_12_0_tr_write_done => x_rsc_12_0_tr_write_done,
      x_rsc_12_0_RREADY => x_rsc_12_0_RREADY,
      x_rsc_12_0_RVALID => x_rsc_12_0_RVALID,
      x_rsc_12_0_RUSER => x_rsc_12_0_RUSER,
      x_rsc_12_0_RLAST => x_rsc_12_0_RLAST,
      x_rsc_12_0_RRESP => hybrid_core_inst_x_rsc_12_0_RRESP,
      x_rsc_12_0_RDATA => hybrid_core_inst_x_rsc_12_0_RDATA,
      x_rsc_12_0_RID => x_rsc_12_0_RID,
      x_rsc_12_0_ARREADY => x_rsc_12_0_ARREADY,
      x_rsc_12_0_ARVALID => x_rsc_12_0_ARVALID,
      x_rsc_12_0_ARUSER => x_rsc_12_0_ARUSER,
      x_rsc_12_0_ARREGION => hybrid_core_inst_x_rsc_12_0_ARREGION,
      x_rsc_12_0_ARQOS => hybrid_core_inst_x_rsc_12_0_ARQOS,
      x_rsc_12_0_ARPROT => hybrid_core_inst_x_rsc_12_0_ARPROT,
      x_rsc_12_0_ARCACHE => hybrid_core_inst_x_rsc_12_0_ARCACHE,
      x_rsc_12_0_ARLOCK => x_rsc_12_0_ARLOCK,
      x_rsc_12_0_ARBURST => hybrid_core_inst_x_rsc_12_0_ARBURST,
      x_rsc_12_0_ARSIZE => hybrid_core_inst_x_rsc_12_0_ARSIZE,
      x_rsc_12_0_ARLEN => hybrid_core_inst_x_rsc_12_0_ARLEN,
      x_rsc_12_0_ARADDR => hybrid_core_inst_x_rsc_12_0_ARADDR,
      x_rsc_12_0_ARID => x_rsc_12_0_ARID,
      x_rsc_12_0_BREADY => x_rsc_12_0_BREADY,
      x_rsc_12_0_BVALID => x_rsc_12_0_BVALID,
      x_rsc_12_0_BUSER => x_rsc_12_0_BUSER,
      x_rsc_12_0_BRESP => hybrid_core_inst_x_rsc_12_0_BRESP,
      x_rsc_12_0_BID => x_rsc_12_0_BID,
      x_rsc_12_0_WREADY => x_rsc_12_0_WREADY,
      x_rsc_12_0_WVALID => x_rsc_12_0_WVALID,
      x_rsc_12_0_WUSER => x_rsc_12_0_WUSER,
      x_rsc_12_0_WLAST => x_rsc_12_0_WLAST,
      x_rsc_12_0_WSTRB => hybrid_core_inst_x_rsc_12_0_WSTRB,
      x_rsc_12_0_WDATA => hybrid_core_inst_x_rsc_12_0_WDATA,
      x_rsc_12_0_AWREADY => x_rsc_12_0_AWREADY,
      x_rsc_12_0_AWVALID => x_rsc_12_0_AWVALID,
      x_rsc_12_0_AWUSER => x_rsc_12_0_AWUSER,
      x_rsc_12_0_AWREGION => hybrid_core_inst_x_rsc_12_0_AWREGION,
      x_rsc_12_0_AWQOS => hybrid_core_inst_x_rsc_12_0_AWQOS,
      x_rsc_12_0_AWPROT => hybrid_core_inst_x_rsc_12_0_AWPROT,
      x_rsc_12_0_AWCACHE => hybrid_core_inst_x_rsc_12_0_AWCACHE,
      x_rsc_12_0_AWLOCK => x_rsc_12_0_AWLOCK,
      x_rsc_12_0_AWBURST => hybrid_core_inst_x_rsc_12_0_AWBURST,
      x_rsc_12_0_AWSIZE => hybrid_core_inst_x_rsc_12_0_AWSIZE,
      x_rsc_12_0_AWLEN => hybrid_core_inst_x_rsc_12_0_AWLEN,
      x_rsc_12_0_AWADDR => hybrid_core_inst_x_rsc_12_0_AWADDR,
      x_rsc_12_0_AWID => x_rsc_12_0_AWID,
      x_rsc_triosy_12_0_lz => x_rsc_triosy_12_0_lz,
      x_rsc_13_0_s_tdone => x_rsc_13_0_s_tdone,
      x_rsc_13_0_tr_write_done => x_rsc_13_0_tr_write_done,
      x_rsc_13_0_RREADY => x_rsc_13_0_RREADY,
      x_rsc_13_0_RVALID => x_rsc_13_0_RVALID,
      x_rsc_13_0_RUSER => x_rsc_13_0_RUSER,
      x_rsc_13_0_RLAST => x_rsc_13_0_RLAST,
      x_rsc_13_0_RRESP => hybrid_core_inst_x_rsc_13_0_RRESP,
      x_rsc_13_0_RDATA => hybrid_core_inst_x_rsc_13_0_RDATA,
      x_rsc_13_0_RID => x_rsc_13_0_RID,
      x_rsc_13_0_ARREADY => x_rsc_13_0_ARREADY,
      x_rsc_13_0_ARVALID => x_rsc_13_0_ARVALID,
      x_rsc_13_0_ARUSER => x_rsc_13_0_ARUSER,
      x_rsc_13_0_ARREGION => hybrid_core_inst_x_rsc_13_0_ARREGION,
      x_rsc_13_0_ARQOS => hybrid_core_inst_x_rsc_13_0_ARQOS,
      x_rsc_13_0_ARPROT => hybrid_core_inst_x_rsc_13_0_ARPROT,
      x_rsc_13_0_ARCACHE => hybrid_core_inst_x_rsc_13_0_ARCACHE,
      x_rsc_13_0_ARLOCK => x_rsc_13_0_ARLOCK,
      x_rsc_13_0_ARBURST => hybrid_core_inst_x_rsc_13_0_ARBURST,
      x_rsc_13_0_ARSIZE => hybrid_core_inst_x_rsc_13_0_ARSIZE,
      x_rsc_13_0_ARLEN => hybrid_core_inst_x_rsc_13_0_ARLEN,
      x_rsc_13_0_ARADDR => hybrid_core_inst_x_rsc_13_0_ARADDR,
      x_rsc_13_0_ARID => x_rsc_13_0_ARID,
      x_rsc_13_0_BREADY => x_rsc_13_0_BREADY,
      x_rsc_13_0_BVALID => x_rsc_13_0_BVALID,
      x_rsc_13_0_BUSER => x_rsc_13_0_BUSER,
      x_rsc_13_0_BRESP => hybrid_core_inst_x_rsc_13_0_BRESP,
      x_rsc_13_0_BID => x_rsc_13_0_BID,
      x_rsc_13_0_WREADY => x_rsc_13_0_WREADY,
      x_rsc_13_0_WVALID => x_rsc_13_0_WVALID,
      x_rsc_13_0_WUSER => x_rsc_13_0_WUSER,
      x_rsc_13_0_WLAST => x_rsc_13_0_WLAST,
      x_rsc_13_0_WSTRB => hybrid_core_inst_x_rsc_13_0_WSTRB,
      x_rsc_13_0_WDATA => hybrid_core_inst_x_rsc_13_0_WDATA,
      x_rsc_13_0_AWREADY => x_rsc_13_0_AWREADY,
      x_rsc_13_0_AWVALID => x_rsc_13_0_AWVALID,
      x_rsc_13_0_AWUSER => x_rsc_13_0_AWUSER,
      x_rsc_13_0_AWREGION => hybrid_core_inst_x_rsc_13_0_AWREGION,
      x_rsc_13_0_AWQOS => hybrid_core_inst_x_rsc_13_0_AWQOS,
      x_rsc_13_0_AWPROT => hybrid_core_inst_x_rsc_13_0_AWPROT,
      x_rsc_13_0_AWCACHE => hybrid_core_inst_x_rsc_13_0_AWCACHE,
      x_rsc_13_0_AWLOCK => x_rsc_13_0_AWLOCK,
      x_rsc_13_0_AWBURST => hybrid_core_inst_x_rsc_13_0_AWBURST,
      x_rsc_13_0_AWSIZE => hybrid_core_inst_x_rsc_13_0_AWSIZE,
      x_rsc_13_0_AWLEN => hybrid_core_inst_x_rsc_13_0_AWLEN,
      x_rsc_13_0_AWADDR => hybrid_core_inst_x_rsc_13_0_AWADDR,
      x_rsc_13_0_AWID => x_rsc_13_0_AWID,
      x_rsc_triosy_13_0_lz => x_rsc_triosy_13_0_lz,
      x_rsc_14_0_s_tdone => x_rsc_14_0_s_tdone,
      x_rsc_14_0_tr_write_done => x_rsc_14_0_tr_write_done,
      x_rsc_14_0_RREADY => x_rsc_14_0_RREADY,
      x_rsc_14_0_RVALID => x_rsc_14_0_RVALID,
      x_rsc_14_0_RUSER => x_rsc_14_0_RUSER,
      x_rsc_14_0_RLAST => x_rsc_14_0_RLAST,
      x_rsc_14_0_RRESP => hybrid_core_inst_x_rsc_14_0_RRESP,
      x_rsc_14_0_RDATA => hybrid_core_inst_x_rsc_14_0_RDATA,
      x_rsc_14_0_RID => x_rsc_14_0_RID,
      x_rsc_14_0_ARREADY => x_rsc_14_0_ARREADY,
      x_rsc_14_0_ARVALID => x_rsc_14_0_ARVALID,
      x_rsc_14_0_ARUSER => x_rsc_14_0_ARUSER,
      x_rsc_14_0_ARREGION => hybrid_core_inst_x_rsc_14_0_ARREGION,
      x_rsc_14_0_ARQOS => hybrid_core_inst_x_rsc_14_0_ARQOS,
      x_rsc_14_0_ARPROT => hybrid_core_inst_x_rsc_14_0_ARPROT,
      x_rsc_14_0_ARCACHE => hybrid_core_inst_x_rsc_14_0_ARCACHE,
      x_rsc_14_0_ARLOCK => x_rsc_14_0_ARLOCK,
      x_rsc_14_0_ARBURST => hybrid_core_inst_x_rsc_14_0_ARBURST,
      x_rsc_14_0_ARSIZE => hybrid_core_inst_x_rsc_14_0_ARSIZE,
      x_rsc_14_0_ARLEN => hybrid_core_inst_x_rsc_14_0_ARLEN,
      x_rsc_14_0_ARADDR => hybrid_core_inst_x_rsc_14_0_ARADDR,
      x_rsc_14_0_ARID => x_rsc_14_0_ARID,
      x_rsc_14_0_BREADY => x_rsc_14_0_BREADY,
      x_rsc_14_0_BVALID => x_rsc_14_0_BVALID,
      x_rsc_14_0_BUSER => x_rsc_14_0_BUSER,
      x_rsc_14_0_BRESP => hybrid_core_inst_x_rsc_14_0_BRESP,
      x_rsc_14_0_BID => x_rsc_14_0_BID,
      x_rsc_14_0_WREADY => x_rsc_14_0_WREADY,
      x_rsc_14_0_WVALID => x_rsc_14_0_WVALID,
      x_rsc_14_0_WUSER => x_rsc_14_0_WUSER,
      x_rsc_14_0_WLAST => x_rsc_14_0_WLAST,
      x_rsc_14_0_WSTRB => hybrid_core_inst_x_rsc_14_0_WSTRB,
      x_rsc_14_0_WDATA => hybrid_core_inst_x_rsc_14_0_WDATA,
      x_rsc_14_0_AWREADY => x_rsc_14_0_AWREADY,
      x_rsc_14_0_AWVALID => x_rsc_14_0_AWVALID,
      x_rsc_14_0_AWUSER => x_rsc_14_0_AWUSER,
      x_rsc_14_0_AWREGION => hybrid_core_inst_x_rsc_14_0_AWREGION,
      x_rsc_14_0_AWQOS => hybrid_core_inst_x_rsc_14_0_AWQOS,
      x_rsc_14_0_AWPROT => hybrid_core_inst_x_rsc_14_0_AWPROT,
      x_rsc_14_0_AWCACHE => hybrid_core_inst_x_rsc_14_0_AWCACHE,
      x_rsc_14_0_AWLOCK => x_rsc_14_0_AWLOCK,
      x_rsc_14_0_AWBURST => hybrid_core_inst_x_rsc_14_0_AWBURST,
      x_rsc_14_0_AWSIZE => hybrid_core_inst_x_rsc_14_0_AWSIZE,
      x_rsc_14_0_AWLEN => hybrid_core_inst_x_rsc_14_0_AWLEN,
      x_rsc_14_0_AWADDR => hybrid_core_inst_x_rsc_14_0_AWADDR,
      x_rsc_14_0_AWID => x_rsc_14_0_AWID,
      x_rsc_triosy_14_0_lz => x_rsc_triosy_14_0_lz,
      x_rsc_15_0_s_tdone => x_rsc_15_0_s_tdone,
      x_rsc_15_0_tr_write_done => x_rsc_15_0_tr_write_done,
      x_rsc_15_0_RREADY => x_rsc_15_0_RREADY,
      x_rsc_15_0_RVALID => x_rsc_15_0_RVALID,
      x_rsc_15_0_RUSER => x_rsc_15_0_RUSER,
      x_rsc_15_0_RLAST => x_rsc_15_0_RLAST,
      x_rsc_15_0_RRESP => hybrid_core_inst_x_rsc_15_0_RRESP,
      x_rsc_15_0_RDATA => hybrid_core_inst_x_rsc_15_0_RDATA,
      x_rsc_15_0_RID => x_rsc_15_0_RID,
      x_rsc_15_0_ARREADY => x_rsc_15_0_ARREADY,
      x_rsc_15_0_ARVALID => x_rsc_15_0_ARVALID,
      x_rsc_15_0_ARUSER => x_rsc_15_0_ARUSER,
      x_rsc_15_0_ARREGION => hybrid_core_inst_x_rsc_15_0_ARREGION,
      x_rsc_15_0_ARQOS => hybrid_core_inst_x_rsc_15_0_ARQOS,
      x_rsc_15_0_ARPROT => hybrid_core_inst_x_rsc_15_0_ARPROT,
      x_rsc_15_0_ARCACHE => hybrid_core_inst_x_rsc_15_0_ARCACHE,
      x_rsc_15_0_ARLOCK => x_rsc_15_0_ARLOCK,
      x_rsc_15_0_ARBURST => hybrid_core_inst_x_rsc_15_0_ARBURST,
      x_rsc_15_0_ARSIZE => hybrid_core_inst_x_rsc_15_0_ARSIZE,
      x_rsc_15_0_ARLEN => hybrid_core_inst_x_rsc_15_0_ARLEN,
      x_rsc_15_0_ARADDR => hybrid_core_inst_x_rsc_15_0_ARADDR,
      x_rsc_15_0_ARID => x_rsc_15_0_ARID,
      x_rsc_15_0_BREADY => x_rsc_15_0_BREADY,
      x_rsc_15_0_BVALID => x_rsc_15_0_BVALID,
      x_rsc_15_0_BUSER => x_rsc_15_0_BUSER,
      x_rsc_15_0_BRESP => hybrid_core_inst_x_rsc_15_0_BRESP,
      x_rsc_15_0_BID => x_rsc_15_0_BID,
      x_rsc_15_0_WREADY => x_rsc_15_0_WREADY,
      x_rsc_15_0_WVALID => x_rsc_15_0_WVALID,
      x_rsc_15_0_WUSER => x_rsc_15_0_WUSER,
      x_rsc_15_0_WLAST => x_rsc_15_0_WLAST,
      x_rsc_15_0_WSTRB => hybrid_core_inst_x_rsc_15_0_WSTRB,
      x_rsc_15_0_WDATA => hybrid_core_inst_x_rsc_15_0_WDATA,
      x_rsc_15_0_AWREADY => x_rsc_15_0_AWREADY,
      x_rsc_15_0_AWVALID => x_rsc_15_0_AWVALID,
      x_rsc_15_0_AWUSER => x_rsc_15_0_AWUSER,
      x_rsc_15_0_AWREGION => hybrid_core_inst_x_rsc_15_0_AWREGION,
      x_rsc_15_0_AWQOS => hybrid_core_inst_x_rsc_15_0_AWQOS,
      x_rsc_15_0_AWPROT => hybrid_core_inst_x_rsc_15_0_AWPROT,
      x_rsc_15_0_AWCACHE => hybrid_core_inst_x_rsc_15_0_AWCACHE,
      x_rsc_15_0_AWLOCK => x_rsc_15_0_AWLOCK,
      x_rsc_15_0_AWBURST => hybrid_core_inst_x_rsc_15_0_AWBURST,
      x_rsc_15_0_AWSIZE => hybrid_core_inst_x_rsc_15_0_AWSIZE,
      x_rsc_15_0_AWLEN => hybrid_core_inst_x_rsc_15_0_AWLEN,
      x_rsc_15_0_AWADDR => hybrid_core_inst_x_rsc_15_0_AWADDR,
      x_rsc_15_0_AWID => x_rsc_15_0_AWID,
      x_rsc_triosy_15_0_lz => x_rsc_triosy_15_0_lz,
      x_rsc_16_0_s_tdone => x_rsc_16_0_s_tdone,
      x_rsc_16_0_tr_write_done => x_rsc_16_0_tr_write_done,
      x_rsc_16_0_RREADY => x_rsc_16_0_RREADY,
      x_rsc_16_0_RVALID => x_rsc_16_0_RVALID,
      x_rsc_16_0_RUSER => x_rsc_16_0_RUSER,
      x_rsc_16_0_RLAST => x_rsc_16_0_RLAST,
      x_rsc_16_0_RRESP => hybrid_core_inst_x_rsc_16_0_RRESP,
      x_rsc_16_0_RDATA => hybrid_core_inst_x_rsc_16_0_RDATA,
      x_rsc_16_0_RID => x_rsc_16_0_RID,
      x_rsc_16_0_ARREADY => x_rsc_16_0_ARREADY,
      x_rsc_16_0_ARVALID => x_rsc_16_0_ARVALID,
      x_rsc_16_0_ARUSER => x_rsc_16_0_ARUSER,
      x_rsc_16_0_ARREGION => hybrid_core_inst_x_rsc_16_0_ARREGION,
      x_rsc_16_0_ARQOS => hybrid_core_inst_x_rsc_16_0_ARQOS,
      x_rsc_16_0_ARPROT => hybrid_core_inst_x_rsc_16_0_ARPROT,
      x_rsc_16_0_ARCACHE => hybrid_core_inst_x_rsc_16_0_ARCACHE,
      x_rsc_16_0_ARLOCK => x_rsc_16_0_ARLOCK,
      x_rsc_16_0_ARBURST => hybrid_core_inst_x_rsc_16_0_ARBURST,
      x_rsc_16_0_ARSIZE => hybrid_core_inst_x_rsc_16_0_ARSIZE,
      x_rsc_16_0_ARLEN => hybrid_core_inst_x_rsc_16_0_ARLEN,
      x_rsc_16_0_ARADDR => hybrid_core_inst_x_rsc_16_0_ARADDR,
      x_rsc_16_0_ARID => x_rsc_16_0_ARID,
      x_rsc_16_0_BREADY => x_rsc_16_0_BREADY,
      x_rsc_16_0_BVALID => x_rsc_16_0_BVALID,
      x_rsc_16_0_BUSER => x_rsc_16_0_BUSER,
      x_rsc_16_0_BRESP => hybrid_core_inst_x_rsc_16_0_BRESP,
      x_rsc_16_0_BID => x_rsc_16_0_BID,
      x_rsc_16_0_WREADY => x_rsc_16_0_WREADY,
      x_rsc_16_0_WVALID => x_rsc_16_0_WVALID,
      x_rsc_16_0_WUSER => x_rsc_16_0_WUSER,
      x_rsc_16_0_WLAST => x_rsc_16_0_WLAST,
      x_rsc_16_0_WSTRB => hybrid_core_inst_x_rsc_16_0_WSTRB,
      x_rsc_16_0_WDATA => hybrid_core_inst_x_rsc_16_0_WDATA,
      x_rsc_16_0_AWREADY => x_rsc_16_0_AWREADY,
      x_rsc_16_0_AWVALID => x_rsc_16_0_AWVALID,
      x_rsc_16_0_AWUSER => x_rsc_16_0_AWUSER,
      x_rsc_16_0_AWREGION => hybrid_core_inst_x_rsc_16_0_AWREGION,
      x_rsc_16_0_AWQOS => hybrid_core_inst_x_rsc_16_0_AWQOS,
      x_rsc_16_0_AWPROT => hybrid_core_inst_x_rsc_16_0_AWPROT,
      x_rsc_16_0_AWCACHE => hybrid_core_inst_x_rsc_16_0_AWCACHE,
      x_rsc_16_0_AWLOCK => x_rsc_16_0_AWLOCK,
      x_rsc_16_0_AWBURST => hybrid_core_inst_x_rsc_16_0_AWBURST,
      x_rsc_16_0_AWSIZE => hybrid_core_inst_x_rsc_16_0_AWSIZE,
      x_rsc_16_0_AWLEN => hybrid_core_inst_x_rsc_16_0_AWLEN,
      x_rsc_16_0_AWADDR => hybrid_core_inst_x_rsc_16_0_AWADDR,
      x_rsc_16_0_AWID => x_rsc_16_0_AWID,
      x_rsc_triosy_16_0_lz => x_rsc_triosy_16_0_lz,
      x_rsc_17_0_s_tdone => x_rsc_17_0_s_tdone,
      x_rsc_17_0_tr_write_done => x_rsc_17_0_tr_write_done,
      x_rsc_17_0_RREADY => x_rsc_17_0_RREADY,
      x_rsc_17_0_RVALID => x_rsc_17_0_RVALID,
      x_rsc_17_0_RUSER => x_rsc_17_0_RUSER,
      x_rsc_17_0_RLAST => x_rsc_17_0_RLAST,
      x_rsc_17_0_RRESP => hybrid_core_inst_x_rsc_17_0_RRESP,
      x_rsc_17_0_RDATA => hybrid_core_inst_x_rsc_17_0_RDATA,
      x_rsc_17_0_RID => x_rsc_17_0_RID,
      x_rsc_17_0_ARREADY => x_rsc_17_0_ARREADY,
      x_rsc_17_0_ARVALID => x_rsc_17_0_ARVALID,
      x_rsc_17_0_ARUSER => x_rsc_17_0_ARUSER,
      x_rsc_17_0_ARREGION => hybrid_core_inst_x_rsc_17_0_ARREGION,
      x_rsc_17_0_ARQOS => hybrid_core_inst_x_rsc_17_0_ARQOS,
      x_rsc_17_0_ARPROT => hybrid_core_inst_x_rsc_17_0_ARPROT,
      x_rsc_17_0_ARCACHE => hybrid_core_inst_x_rsc_17_0_ARCACHE,
      x_rsc_17_0_ARLOCK => x_rsc_17_0_ARLOCK,
      x_rsc_17_0_ARBURST => hybrid_core_inst_x_rsc_17_0_ARBURST,
      x_rsc_17_0_ARSIZE => hybrid_core_inst_x_rsc_17_0_ARSIZE,
      x_rsc_17_0_ARLEN => hybrid_core_inst_x_rsc_17_0_ARLEN,
      x_rsc_17_0_ARADDR => hybrid_core_inst_x_rsc_17_0_ARADDR,
      x_rsc_17_0_ARID => x_rsc_17_0_ARID,
      x_rsc_17_0_BREADY => x_rsc_17_0_BREADY,
      x_rsc_17_0_BVALID => x_rsc_17_0_BVALID,
      x_rsc_17_0_BUSER => x_rsc_17_0_BUSER,
      x_rsc_17_0_BRESP => hybrid_core_inst_x_rsc_17_0_BRESP,
      x_rsc_17_0_BID => x_rsc_17_0_BID,
      x_rsc_17_0_WREADY => x_rsc_17_0_WREADY,
      x_rsc_17_0_WVALID => x_rsc_17_0_WVALID,
      x_rsc_17_0_WUSER => x_rsc_17_0_WUSER,
      x_rsc_17_0_WLAST => x_rsc_17_0_WLAST,
      x_rsc_17_0_WSTRB => hybrid_core_inst_x_rsc_17_0_WSTRB,
      x_rsc_17_0_WDATA => hybrid_core_inst_x_rsc_17_0_WDATA,
      x_rsc_17_0_AWREADY => x_rsc_17_0_AWREADY,
      x_rsc_17_0_AWVALID => x_rsc_17_0_AWVALID,
      x_rsc_17_0_AWUSER => x_rsc_17_0_AWUSER,
      x_rsc_17_0_AWREGION => hybrid_core_inst_x_rsc_17_0_AWREGION,
      x_rsc_17_0_AWQOS => hybrid_core_inst_x_rsc_17_0_AWQOS,
      x_rsc_17_0_AWPROT => hybrid_core_inst_x_rsc_17_0_AWPROT,
      x_rsc_17_0_AWCACHE => hybrid_core_inst_x_rsc_17_0_AWCACHE,
      x_rsc_17_0_AWLOCK => x_rsc_17_0_AWLOCK,
      x_rsc_17_0_AWBURST => hybrid_core_inst_x_rsc_17_0_AWBURST,
      x_rsc_17_0_AWSIZE => hybrid_core_inst_x_rsc_17_0_AWSIZE,
      x_rsc_17_0_AWLEN => hybrid_core_inst_x_rsc_17_0_AWLEN,
      x_rsc_17_0_AWADDR => hybrid_core_inst_x_rsc_17_0_AWADDR,
      x_rsc_17_0_AWID => x_rsc_17_0_AWID,
      x_rsc_triosy_17_0_lz => x_rsc_triosy_17_0_lz,
      x_rsc_18_0_s_tdone => x_rsc_18_0_s_tdone,
      x_rsc_18_0_tr_write_done => x_rsc_18_0_tr_write_done,
      x_rsc_18_0_RREADY => x_rsc_18_0_RREADY,
      x_rsc_18_0_RVALID => x_rsc_18_0_RVALID,
      x_rsc_18_0_RUSER => x_rsc_18_0_RUSER,
      x_rsc_18_0_RLAST => x_rsc_18_0_RLAST,
      x_rsc_18_0_RRESP => hybrid_core_inst_x_rsc_18_0_RRESP,
      x_rsc_18_0_RDATA => hybrid_core_inst_x_rsc_18_0_RDATA,
      x_rsc_18_0_RID => x_rsc_18_0_RID,
      x_rsc_18_0_ARREADY => x_rsc_18_0_ARREADY,
      x_rsc_18_0_ARVALID => x_rsc_18_0_ARVALID,
      x_rsc_18_0_ARUSER => x_rsc_18_0_ARUSER,
      x_rsc_18_0_ARREGION => hybrid_core_inst_x_rsc_18_0_ARREGION,
      x_rsc_18_0_ARQOS => hybrid_core_inst_x_rsc_18_0_ARQOS,
      x_rsc_18_0_ARPROT => hybrid_core_inst_x_rsc_18_0_ARPROT,
      x_rsc_18_0_ARCACHE => hybrid_core_inst_x_rsc_18_0_ARCACHE,
      x_rsc_18_0_ARLOCK => x_rsc_18_0_ARLOCK,
      x_rsc_18_0_ARBURST => hybrid_core_inst_x_rsc_18_0_ARBURST,
      x_rsc_18_0_ARSIZE => hybrid_core_inst_x_rsc_18_0_ARSIZE,
      x_rsc_18_0_ARLEN => hybrid_core_inst_x_rsc_18_0_ARLEN,
      x_rsc_18_0_ARADDR => hybrid_core_inst_x_rsc_18_0_ARADDR,
      x_rsc_18_0_ARID => x_rsc_18_0_ARID,
      x_rsc_18_0_BREADY => x_rsc_18_0_BREADY,
      x_rsc_18_0_BVALID => x_rsc_18_0_BVALID,
      x_rsc_18_0_BUSER => x_rsc_18_0_BUSER,
      x_rsc_18_0_BRESP => hybrid_core_inst_x_rsc_18_0_BRESP,
      x_rsc_18_0_BID => x_rsc_18_0_BID,
      x_rsc_18_0_WREADY => x_rsc_18_0_WREADY,
      x_rsc_18_0_WVALID => x_rsc_18_0_WVALID,
      x_rsc_18_0_WUSER => x_rsc_18_0_WUSER,
      x_rsc_18_0_WLAST => x_rsc_18_0_WLAST,
      x_rsc_18_0_WSTRB => hybrid_core_inst_x_rsc_18_0_WSTRB,
      x_rsc_18_0_WDATA => hybrid_core_inst_x_rsc_18_0_WDATA,
      x_rsc_18_0_AWREADY => x_rsc_18_0_AWREADY,
      x_rsc_18_0_AWVALID => x_rsc_18_0_AWVALID,
      x_rsc_18_0_AWUSER => x_rsc_18_0_AWUSER,
      x_rsc_18_0_AWREGION => hybrid_core_inst_x_rsc_18_0_AWREGION,
      x_rsc_18_0_AWQOS => hybrid_core_inst_x_rsc_18_0_AWQOS,
      x_rsc_18_0_AWPROT => hybrid_core_inst_x_rsc_18_0_AWPROT,
      x_rsc_18_0_AWCACHE => hybrid_core_inst_x_rsc_18_0_AWCACHE,
      x_rsc_18_0_AWLOCK => x_rsc_18_0_AWLOCK,
      x_rsc_18_0_AWBURST => hybrid_core_inst_x_rsc_18_0_AWBURST,
      x_rsc_18_0_AWSIZE => hybrid_core_inst_x_rsc_18_0_AWSIZE,
      x_rsc_18_0_AWLEN => hybrid_core_inst_x_rsc_18_0_AWLEN,
      x_rsc_18_0_AWADDR => hybrid_core_inst_x_rsc_18_0_AWADDR,
      x_rsc_18_0_AWID => x_rsc_18_0_AWID,
      x_rsc_triosy_18_0_lz => x_rsc_triosy_18_0_lz,
      x_rsc_19_0_s_tdone => x_rsc_19_0_s_tdone,
      x_rsc_19_0_tr_write_done => x_rsc_19_0_tr_write_done,
      x_rsc_19_0_RREADY => x_rsc_19_0_RREADY,
      x_rsc_19_0_RVALID => x_rsc_19_0_RVALID,
      x_rsc_19_0_RUSER => x_rsc_19_0_RUSER,
      x_rsc_19_0_RLAST => x_rsc_19_0_RLAST,
      x_rsc_19_0_RRESP => hybrid_core_inst_x_rsc_19_0_RRESP,
      x_rsc_19_0_RDATA => hybrid_core_inst_x_rsc_19_0_RDATA,
      x_rsc_19_0_RID => x_rsc_19_0_RID,
      x_rsc_19_0_ARREADY => x_rsc_19_0_ARREADY,
      x_rsc_19_0_ARVALID => x_rsc_19_0_ARVALID,
      x_rsc_19_0_ARUSER => x_rsc_19_0_ARUSER,
      x_rsc_19_0_ARREGION => hybrid_core_inst_x_rsc_19_0_ARREGION,
      x_rsc_19_0_ARQOS => hybrid_core_inst_x_rsc_19_0_ARQOS,
      x_rsc_19_0_ARPROT => hybrid_core_inst_x_rsc_19_0_ARPROT,
      x_rsc_19_0_ARCACHE => hybrid_core_inst_x_rsc_19_0_ARCACHE,
      x_rsc_19_0_ARLOCK => x_rsc_19_0_ARLOCK,
      x_rsc_19_0_ARBURST => hybrid_core_inst_x_rsc_19_0_ARBURST,
      x_rsc_19_0_ARSIZE => hybrid_core_inst_x_rsc_19_0_ARSIZE,
      x_rsc_19_0_ARLEN => hybrid_core_inst_x_rsc_19_0_ARLEN,
      x_rsc_19_0_ARADDR => hybrid_core_inst_x_rsc_19_0_ARADDR,
      x_rsc_19_0_ARID => x_rsc_19_0_ARID,
      x_rsc_19_0_BREADY => x_rsc_19_0_BREADY,
      x_rsc_19_0_BVALID => x_rsc_19_0_BVALID,
      x_rsc_19_0_BUSER => x_rsc_19_0_BUSER,
      x_rsc_19_0_BRESP => hybrid_core_inst_x_rsc_19_0_BRESP,
      x_rsc_19_0_BID => x_rsc_19_0_BID,
      x_rsc_19_0_WREADY => x_rsc_19_0_WREADY,
      x_rsc_19_0_WVALID => x_rsc_19_0_WVALID,
      x_rsc_19_0_WUSER => x_rsc_19_0_WUSER,
      x_rsc_19_0_WLAST => x_rsc_19_0_WLAST,
      x_rsc_19_0_WSTRB => hybrid_core_inst_x_rsc_19_0_WSTRB,
      x_rsc_19_0_WDATA => hybrid_core_inst_x_rsc_19_0_WDATA,
      x_rsc_19_0_AWREADY => x_rsc_19_0_AWREADY,
      x_rsc_19_0_AWVALID => x_rsc_19_0_AWVALID,
      x_rsc_19_0_AWUSER => x_rsc_19_0_AWUSER,
      x_rsc_19_0_AWREGION => hybrid_core_inst_x_rsc_19_0_AWREGION,
      x_rsc_19_0_AWQOS => hybrid_core_inst_x_rsc_19_0_AWQOS,
      x_rsc_19_0_AWPROT => hybrid_core_inst_x_rsc_19_0_AWPROT,
      x_rsc_19_0_AWCACHE => hybrid_core_inst_x_rsc_19_0_AWCACHE,
      x_rsc_19_0_AWLOCK => x_rsc_19_0_AWLOCK,
      x_rsc_19_0_AWBURST => hybrid_core_inst_x_rsc_19_0_AWBURST,
      x_rsc_19_0_AWSIZE => hybrid_core_inst_x_rsc_19_0_AWSIZE,
      x_rsc_19_0_AWLEN => hybrid_core_inst_x_rsc_19_0_AWLEN,
      x_rsc_19_0_AWADDR => hybrid_core_inst_x_rsc_19_0_AWADDR,
      x_rsc_19_0_AWID => x_rsc_19_0_AWID,
      x_rsc_triosy_19_0_lz => x_rsc_triosy_19_0_lz,
      x_rsc_20_0_s_tdone => x_rsc_20_0_s_tdone,
      x_rsc_20_0_tr_write_done => x_rsc_20_0_tr_write_done,
      x_rsc_20_0_RREADY => x_rsc_20_0_RREADY,
      x_rsc_20_0_RVALID => x_rsc_20_0_RVALID,
      x_rsc_20_0_RUSER => x_rsc_20_0_RUSER,
      x_rsc_20_0_RLAST => x_rsc_20_0_RLAST,
      x_rsc_20_0_RRESP => hybrid_core_inst_x_rsc_20_0_RRESP,
      x_rsc_20_0_RDATA => hybrid_core_inst_x_rsc_20_0_RDATA,
      x_rsc_20_0_RID => x_rsc_20_0_RID,
      x_rsc_20_0_ARREADY => x_rsc_20_0_ARREADY,
      x_rsc_20_0_ARVALID => x_rsc_20_0_ARVALID,
      x_rsc_20_0_ARUSER => x_rsc_20_0_ARUSER,
      x_rsc_20_0_ARREGION => hybrid_core_inst_x_rsc_20_0_ARREGION,
      x_rsc_20_0_ARQOS => hybrid_core_inst_x_rsc_20_0_ARQOS,
      x_rsc_20_0_ARPROT => hybrid_core_inst_x_rsc_20_0_ARPROT,
      x_rsc_20_0_ARCACHE => hybrid_core_inst_x_rsc_20_0_ARCACHE,
      x_rsc_20_0_ARLOCK => x_rsc_20_0_ARLOCK,
      x_rsc_20_0_ARBURST => hybrid_core_inst_x_rsc_20_0_ARBURST,
      x_rsc_20_0_ARSIZE => hybrid_core_inst_x_rsc_20_0_ARSIZE,
      x_rsc_20_0_ARLEN => hybrid_core_inst_x_rsc_20_0_ARLEN,
      x_rsc_20_0_ARADDR => hybrid_core_inst_x_rsc_20_0_ARADDR,
      x_rsc_20_0_ARID => x_rsc_20_0_ARID,
      x_rsc_20_0_BREADY => x_rsc_20_0_BREADY,
      x_rsc_20_0_BVALID => x_rsc_20_0_BVALID,
      x_rsc_20_0_BUSER => x_rsc_20_0_BUSER,
      x_rsc_20_0_BRESP => hybrid_core_inst_x_rsc_20_0_BRESP,
      x_rsc_20_0_BID => x_rsc_20_0_BID,
      x_rsc_20_0_WREADY => x_rsc_20_0_WREADY,
      x_rsc_20_0_WVALID => x_rsc_20_0_WVALID,
      x_rsc_20_0_WUSER => x_rsc_20_0_WUSER,
      x_rsc_20_0_WLAST => x_rsc_20_0_WLAST,
      x_rsc_20_0_WSTRB => hybrid_core_inst_x_rsc_20_0_WSTRB,
      x_rsc_20_0_WDATA => hybrid_core_inst_x_rsc_20_0_WDATA,
      x_rsc_20_0_AWREADY => x_rsc_20_0_AWREADY,
      x_rsc_20_0_AWVALID => x_rsc_20_0_AWVALID,
      x_rsc_20_0_AWUSER => x_rsc_20_0_AWUSER,
      x_rsc_20_0_AWREGION => hybrid_core_inst_x_rsc_20_0_AWREGION,
      x_rsc_20_0_AWQOS => hybrid_core_inst_x_rsc_20_0_AWQOS,
      x_rsc_20_0_AWPROT => hybrid_core_inst_x_rsc_20_0_AWPROT,
      x_rsc_20_0_AWCACHE => hybrid_core_inst_x_rsc_20_0_AWCACHE,
      x_rsc_20_0_AWLOCK => x_rsc_20_0_AWLOCK,
      x_rsc_20_0_AWBURST => hybrid_core_inst_x_rsc_20_0_AWBURST,
      x_rsc_20_0_AWSIZE => hybrid_core_inst_x_rsc_20_0_AWSIZE,
      x_rsc_20_0_AWLEN => hybrid_core_inst_x_rsc_20_0_AWLEN,
      x_rsc_20_0_AWADDR => hybrid_core_inst_x_rsc_20_0_AWADDR,
      x_rsc_20_0_AWID => x_rsc_20_0_AWID,
      x_rsc_triosy_20_0_lz => x_rsc_triosy_20_0_lz,
      x_rsc_21_0_s_tdone => x_rsc_21_0_s_tdone,
      x_rsc_21_0_tr_write_done => x_rsc_21_0_tr_write_done,
      x_rsc_21_0_RREADY => x_rsc_21_0_RREADY,
      x_rsc_21_0_RVALID => x_rsc_21_0_RVALID,
      x_rsc_21_0_RUSER => x_rsc_21_0_RUSER,
      x_rsc_21_0_RLAST => x_rsc_21_0_RLAST,
      x_rsc_21_0_RRESP => hybrid_core_inst_x_rsc_21_0_RRESP,
      x_rsc_21_0_RDATA => hybrid_core_inst_x_rsc_21_0_RDATA,
      x_rsc_21_0_RID => x_rsc_21_0_RID,
      x_rsc_21_0_ARREADY => x_rsc_21_0_ARREADY,
      x_rsc_21_0_ARVALID => x_rsc_21_0_ARVALID,
      x_rsc_21_0_ARUSER => x_rsc_21_0_ARUSER,
      x_rsc_21_0_ARREGION => hybrid_core_inst_x_rsc_21_0_ARREGION,
      x_rsc_21_0_ARQOS => hybrid_core_inst_x_rsc_21_0_ARQOS,
      x_rsc_21_0_ARPROT => hybrid_core_inst_x_rsc_21_0_ARPROT,
      x_rsc_21_0_ARCACHE => hybrid_core_inst_x_rsc_21_0_ARCACHE,
      x_rsc_21_0_ARLOCK => x_rsc_21_0_ARLOCK,
      x_rsc_21_0_ARBURST => hybrid_core_inst_x_rsc_21_0_ARBURST,
      x_rsc_21_0_ARSIZE => hybrid_core_inst_x_rsc_21_0_ARSIZE,
      x_rsc_21_0_ARLEN => hybrid_core_inst_x_rsc_21_0_ARLEN,
      x_rsc_21_0_ARADDR => hybrid_core_inst_x_rsc_21_0_ARADDR,
      x_rsc_21_0_ARID => x_rsc_21_0_ARID,
      x_rsc_21_0_BREADY => x_rsc_21_0_BREADY,
      x_rsc_21_0_BVALID => x_rsc_21_0_BVALID,
      x_rsc_21_0_BUSER => x_rsc_21_0_BUSER,
      x_rsc_21_0_BRESP => hybrid_core_inst_x_rsc_21_0_BRESP,
      x_rsc_21_0_BID => x_rsc_21_0_BID,
      x_rsc_21_0_WREADY => x_rsc_21_0_WREADY,
      x_rsc_21_0_WVALID => x_rsc_21_0_WVALID,
      x_rsc_21_0_WUSER => x_rsc_21_0_WUSER,
      x_rsc_21_0_WLAST => x_rsc_21_0_WLAST,
      x_rsc_21_0_WSTRB => hybrid_core_inst_x_rsc_21_0_WSTRB,
      x_rsc_21_0_WDATA => hybrid_core_inst_x_rsc_21_0_WDATA,
      x_rsc_21_0_AWREADY => x_rsc_21_0_AWREADY,
      x_rsc_21_0_AWVALID => x_rsc_21_0_AWVALID,
      x_rsc_21_0_AWUSER => x_rsc_21_0_AWUSER,
      x_rsc_21_0_AWREGION => hybrid_core_inst_x_rsc_21_0_AWREGION,
      x_rsc_21_0_AWQOS => hybrid_core_inst_x_rsc_21_0_AWQOS,
      x_rsc_21_0_AWPROT => hybrid_core_inst_x_rsc_21_0_AWPROT,
      x_rsc_21_0_AWCACHE => hybrid_core_inst_x_rsc_21_0_AWCACHE,
      x_rsc_21_0_AWLOCK => x_rsc_21_0_AWLOCK,
      x_rsc_21_0_AWBURST => hybrid_core_inst_x_rsc_21_0_AWBURST,
      x_rsc_21_0_AWSIZE => hybrid_core_inst_x_rsc_21_0_AWSIZE,
      x_rsc_21_0_AWLEN => hybrid_core_inst_x_rsc_21_0_AWLEN,
      x_rsc_21_0_AWADDR => hybrid_core_inst_x_rsc_21_0_AWADDR,
      x_rsc_21_0_AWID => x_rsc_21_0_AWID,
      x_rsc_triosy_21_0_lz => x_rsc_triosy_21_0_lz,
      x_rsc_22_0_s_tdone => x_rsc_22_0_s_tdone,
      x_rsc_22_0_tr_write_done => x_rsc_22_0_tr_write_done,
      x_rsc_22_0_RREADY => x_rsc_22_0_RREADY,
      x_rsc_22_0_RVALID => x_rsc_22_0_RVALID,
      x_rsc_22_0_RUSER => x_rsc_22_0_RUSER,
      x_rsc_22_0_RLAST => x_rsc_22_0_RLAST,
      x_rsc_22_0_RRESP => hybrid_core_inst_x_rsc_22_0_RRESP,
      x_rsc_22_0_RDATA => hybrid_core_inst_x_rsc_22_0_RDATA,
      x_rsc_22_0_RID => x_rsc_22_0_RID,
      x_rsc_22_0_ARREADY => x_rsc_22_0_ARREADY,
      x_rsc_22_0_ARVALID => x_rsc_22_0_ARVALID,
      x_rsc_22_0_ARUSER => x_rsc_22_0_ARUSER,
      x_rsc_22_0_ARREGION => hybrid_core_inst_x_rsc_22_0_ARREGION,
      x_rsc_22_0_ARQOS => hybrid_core_inst_x_rsc_22_0_ARQOS,
      x_rsc_22_0_ARPROT => hybrid_core_inst_x_rsc_22_0_ARPROT,
      x_rsc_22_0_ARCACHE => hybrid_core_inst_x_rsc_22_0_ARCACHE,
      x_rsc_22_0_ARLOCK => x_rsc_22_0_ARLOCK,
      x_rsc_22_0_ARBURST => hybrid_core_inst_x_rsc_22_0_ARBURST,
      x_rsc_22_0_ARSIZE => hybrid_core_inst_x_rsc_22_0_ARSIZE,
      x_rsc_22_0_ARLEN => hybrid_core_inst_x_rsc_22_0_ARLEN,
      x_rsc_22_0_ARADDR => hybrid_core_inst_x_rsc_22_0_ARADDR,
      x_rsc_22_0_ARID => x_rsc_22_0_ARID,
      x_rsc_22_0_BREADY => x_rsc_22_0_BREADY,
      x_rsc_22_0_BVALID => x_rsc_22_0_BVALID,
      x_rsc_22_0_BUSER => x_rsc_22_0_BUSER,
      x_rsc_22_0_BRESP => hybrid_core_inst_x_rsc_22_0_BRESP,
      x_rsc_22_0_BID => x_rsc_22_0_BID,
      x_rsc_22_0_WREADY => x_rsc_22_0_WREADY,
      x_rsc_22_0_WVALID => x_rsc_22_0_WVALID,
      x_rsc_22_0_WUSER => x_rsc_22_0_WUSER,
      x_rsc_22_0_WLAST => x_rsc_22_0_WLAST,
      x_rsc_22_0_WSTRB => hybrid_core_inst_x_rsc_22_0_WSTRB,
      x_rsc_22_0_WDATA => hybrid_core_inst_x_rsc_22_0_WDATA,
      x_rsc_22_0_AWREADY => x_rsc_22_0_AWREADY,
      x_rsc_22_0_AWVALID => x_rsc_22_0_AWVALID,
      x_rsc_22_0_AWUSER => x_rsc_22_0_AWUSER,
      x_rsc_22_0_AWREGION => hybrid_core_inst_x_rsc_22_0_AWREGION,
      x_rsc_22_0_AWQOS => hybrid_core_inst_x_rsc_22_0_AWQOS,
      x_rsc_22_0_AWPROT => hybrid_core_inst_x_rsc_22_0_AWPROT,
      x_rsc_22_0_AWCACHE => hybrid_core_inst_x_rsc_22_0_AWCACHE,
      x_rsc_22_0_AWLOCK => x_rsc_22_0_AWLOCK,
      x_rsc_22_0_AWBURST => hybrid_core_inst_x_rsc_22_0_AWBURST,
      x_rsc_22_0_AWSIZE => hybrid_core_inst_x_rsc_22_0_AWSIZE,
      x_rsc_22_0_AWLEN => hybrid_core_inst_x_rsc_22_0_AWLEN,
      x_rsc_22_0_AWADDR => hybrid_core_inst_x_rsc_22_0_AWADDR,
      x_rsc_22_0_AWID => x_rsc_22_0_AWID,
      x_rsc_triosy_22_0_lz => x_rsc_triosy_22_0_lz,
      x_rsc_23_0_s_tdone => x_rsc_23_0_s_tdone,
      x_rsc_23_0_tr_write_done => x_rsc_23_0_tr_write_done,
      x_rsc_23_0_RREADY => x_rsc_23_0_RREADY,
      x_rsc_23_0_RVALID => x_rsc_23_0_RVALID,
      x_rsc_23_0_RUSER => x_rsc_23_0_RUSER,
      x_rsc_23_0_RLAST => x_rsc_23_0_RLAST,
      x_rsc_23_0_RRESP => hybrid_core_inst_x_rsc_23_0_RRESP,
      x_rsc_23_0_RDATA => hybrid_core_inst_x_rsc_23_0_RDATA,
      x_rsc_23_0_RID => x_rsc_23_0_RID,
      x_rsc_23_0_ARREADY => x_rsc_23_0_ARREADY,
      x_rsc_23_0_ARVALID => x_rsc_23_0_ARVALID,
      x_rsc_23_0_ARUSER => x_rsc_23_0_ARUSER,
      x_rsc_23_0_ARREGION => hybrid_core_inst_x_rsc_23_0_ARREGION,
      x_rsc_23_0_ARQOS => hybrid_core_inst_x_rsc_23_0_ARQOS,
      x_rsc_23_0_ARPROT => hybrid_core_inst_x_rsc_23_0_ARPROT,
      x_rsc_23_0_ARCACHE => hybrid_core_inst_x_rsc_23_0_ARCACHE,
      x_rsc_23_0_ARLOCK => x_rsc_23_0_ARLOCK,
      x_rsc_23_0_ARBURST => hybrid_core_inst_x_rsc_23_0_ARBURST,
      x_rsc_23_0_ARSIZE => hybrid_core_inst_x_rsc_23_0_ARSIZE,
      x_rsc_23_0_ARLEN => hybrid_core_inst_x_rsc_23_0_ARLEN,
      x_rsc_23_0_ARADDR => hybrid_core_inst_x_rsc_23_0_ARADDR,
      x_rsc_23_0_ARID => x_rsc_23_0_ARID,
      x_rsc_23_0_BREADY => x_rsc_23_0_BREADY,
      x_rsc_23_0_BVALID => x_rsc_23_0_BVALID,
      x_rsc_23_0_BUSER => x_rsc_23_0_BUSER,
      x_rsc_23_0_BRESP => hybrid_core_inst_x_rsc_23_0_BRESP,
      x_rsc_23_0_BID => x_rsc_23_0_BID,
      x_rsc_23_0_WREADY => x_rsc_23_0_WREADY,
      x_rsc_23_0_WVALID => x_rsc_23_0_WVALID,
      x_rsc_23_0_WUSER => x_rsc_23_0_WUSER,
      x_rsc_23_0_WLAST => x_rsc_23_0_WLAST,
      x_rsc_23_0_WSTRB => hybrid_core_inst_x_rsc_23_0_WSTRB,
      x_rsc_23_0_WDATA => hybrid_core_inst_x_rsc_23_0_WDATA,
      x_rsc_23_0_AWREADY => x_rsc_23_0_AWREADY,
      x_rsc_23_0_AWVALID => x_rsc_23_0_AWVALID,
      x_rsc_23_0_AWUSER => x_rsc_23_0_AWUSER,
      x_rsc_23_0_AWREGION => hybrid_core_inst_x_rsc_23_0_AWREGION,
      x_rsc_23_0_AWQOS => hybrid_core_inst_x_rsc_23_0_AWQOS,
      x_rsc_23_0_AWPROT => hybrid_core_inst_x_rsc_23_0_AWPROT,
      x_rsc_23_0_AWCACHE => hybrid_core_inst_x_rsc_23_0_AWCACHE,
      x_rsc_23_0_AWLOCK => x_rsc_23_0_AWLOCK,
      x_rsc_23_0_AWBURST => hybrid_core_inst_x_rsc_23_0_AWBURST,
      x_rsc_23_0_AWSIZE => hybrid_core_inst_x_rsc_23_0_AWSIZE,
      x_rsc_23_0_AWLEN => hybrid_core_inst_x_rsc_23_0_AWLEN,
      x_rsc_23_0_AWADDR => hybrid_core_inst_x_rsc_23_0_AWADDR,
      x_rsc_23_0_AWID => x_rsc_23_0_AWID,
      x_rsc_triosy_23_0_lz => x_rsc_triosy_23_0_lz,
      x_rsc_24_0_s_tdone => x_rsc_24_0_s_tdone,
      x_rsc_24_0_tr_write_done => x_rsc_24_0_tr_write_done,
      x_rsc_24_0_RREADY => x_rsc_24_0_RREADY,
      x_rsc_24_0_RVALID => x_rsc_24_0_RVALID,
      x_rsc_24_0_RUSER => x_rsc_24_0_RUSER,
      x_rsc_24_0_RLAST => x_rsc_24_0_RLAST,
      x_rsc_24_0_RRESP => hybrid_core_inst_x_rsc_24_0_RRESP,
      x_rsc_24_0_RDATA => hybrid_core_inst_x_rsc_24_0_RDATA,
      x_rsc_24_0_RID => x_rsc_24_0_RID,
      x_rsc_24_0_ARREADY => x_rsc_24_0_ARREADY,
      x_rsc_24_0_ARVALID => x_rsc_24_0_ARVALID,
      x_rsc_24_0_ARUSER => x_rsc_24_0_ARUSER,
      x_rsc_24_0_ARREGION => hybrid_core_inst_x_rsc_24_0_ARREGION,
      x_rsc_24_0_ARQOS => hybrid_core_inst_x_rsc_24_0_ARQOS,
      x_rsc_24_0_ARPROT => hybrid_core_inst_x_rsc_24_0_ARPROT,
      x_rsc_24_0_ARCACHE => hybrid_core_inst_x_rsc_24_0_ARCACHE,
      x_rsc_24_0_ARLOCK => x_rsc_24_0_ARLOCK,
      x_rsc_24_0_ARBURST => hybrid_core_inst_x_rsc_24_0_ARBURST,
      x_rsc_24_0_ARSIZE => hybrid_core_inst_x_rsc_24_0_ARSIZE,
      x_rsc_24_0_ARLEN => hybrid_core_inst_x_rsc_24_0_ARLEN,
      x_rsc_24_0_ARADDR => hybrid_core_inst_x_rsc_24_0_ARADDR,
      x_rsc_24_0_ARID => x_rsc_24_0_ARID,
      x_rsc_24_0_BREADY => x_rsc_24_0_BREADY,
      x_rsc_24_0_BVALID => x_rsc_24_0_BVALID,
      x_rsc_24_0_BUSER => x_rsc_24_0_BUSER,
      x_rsc_24_0_BRESP => hybrid_core_inst_x_rsc_24_0_BRESP,
      x_rsc_24_0_BID => x_rsc_24_0_BID,
      x_rsc_24_0_WREADY => x_rsc_24_0_WREADY,
      x_rsc_24_0_WVALID => x_rsc_24_0_WVALID,
      x_rsc_24_0_WUSER => x_rsc_24_0_WUSER,
      x_rsc_24_0_WLAST => x_rsc_24_0_WLAST,
      x_rsc_24_0_WSTRB => hybrid_core_inst_x_rsc_24_0_WSTRB,
      x_rsc_24_0_WDATA => hybrid_core_inst_x_rsc_24_0_WDATA,
      x_rsc_24_0_AWREADY => x_rsc_24_0_AWREADY,
      x_rsc_24_0_AWVALID => x_rsc_24_0_AWVALID,
      x_rsc_24_0_AWUSER => x_rsc_24_0_AWUSER,
      x_rsc_24_0_AWREGION => hybrid_core_inst_x_rsc_24_0_AWREGION,
      x_rsc_24_0_AWQOS => hybrid_core_inst_x_rsc_24_0_AWQOS,
      x_rsc_24_0_AWPROT => hybrid_core_inst_x_rsc_24_0_AWPROT,
      x_rsc_24_0_AWCACHE => hybrid_core_inst_x_rsc_24_0_AWCACHE,
      x_rsc_24_0_AWLOCK => x_rsc_24_0_AWLOCK,
      x_rsc_24_0_AWBURST => hybrid_core_inst_x_rsc_24_0_AWBURST,
      x_rsc_24_0_AWSIZE => hybrid_core_inst_x_rsc_24_0_AWSIZE,
      x_rsc_24_0_AWLEN => hybrid_core_inst_x_rsc_24_0_AWLEN,
      x_rsc_24_0_AWADDR => hybrid_core_inst_x_rsc_24_0_AWADDR,
      x_rsc_24_0_AWID => x_rsc_24_0_AWID,
      x_rsc_triosy_24_0_lz => x_rsc_triosy_24_0_lz,
      x_rsc_25_0_s_tdone => x_rsc_25_0_s_tdone,
      x_rsc_25_0_tr_write_done => x_rsc_25_0_tr_write_done,
      x_rsc_25_0_RREADY => x_rsc_25_0_RREADY,
      x_rsc_25_0_RVALID => x_rsc_25_0_RVALID,
      x_rsc_25_0_RUSER => x_rsc_25_0_RUSER,
      x_rsc_25_0_RLAST => x_rsc_25_0_RLAST,
      x_rsc_25_0_RRESP => hybrid_core_inst_x_rsc_25_0_RRESP,
      x_rsc_25_0_RDATA => hybrid_core_inst_x_rsc_25_0_RDATA,
      x_rsc_25_0_RID => x_rsc_25_0_RID,
      x_rsc_25_0_ARREADY => x_rsc_25_0_ARREADY,
      x_rsc_25_0_ARVALID => x_rsc_25_0_ARVALID,
      x_rsc_25_0_ARUSER => x_rsc_25_0_ARUSER,
      x_rsc_25_0_ARREGION => hybrid_core_inst_x_rsc_25_0_ARREGION,
      x_rsc_25_0_ARQOS => hybrid_core_inst_x_rsc_25_0_ARQOS,
      x_rsc_25_0_ARPROT => hybrid_core_inst_x_rsc_25_0_ARPROT,
      x_rsc_25_0_ARCACHE => hybrid_core_inst_x_rsc_25_0_ARCACHE,
      x_rsc_25_0_ARLOCK => x_rsc_25_0_ARLOCK,
      x_rsc_25_0_ARBURST => hybrid_core_inst_x_rsc_25_0_ARBURST,
      x_rsc_25_0_ARSIZE => hybrid_core_inst_x_rsc_25_0_ARSIZE,
      x_rsc_25_0_ARLEN => hybrid_core_inst_x_rsc_25_0_ARLEN,
      x_rsc_25_0_ARADDR => hybrid_core_inst_x_rsc_25_0_ARADDR,
      x_rsc_25_0_ARID => x_rsc_25_0_ARID,
      x_rsc_25_0_BREADY => x_rsc_25_0_BREADY,
      x_rsc_25_0_BVALID => x_rsc_25_0_BVALID,
      x_rsc_25_0_BUSER => x_rsc_25_0_BUSER,
      x_rsc_25_0_BRESP => hybrid_core_inst_x_rsc_25_0_BRESP,
      x_rsc_25_0_BID => x_rsc_25_0_BID,
      x_rsc_25_0_WREADY => x_rsc_25_0_WREADY,
      x_rsc_25_0_WVALID => x_rsc_25_0_WVALID,
      x_rsc_25_0_WUSER => x_rsc_25_0_WUSER,
      x_rsc_25_0_WLAST => x_rsc_25_0_WLAST,
      x_rsc_25_0_WSTRB => hybrid_core_inst_x_rsc_25_0_WSTRB,
      x_rsc_25_0_WDATA => hybrid_core_inst_x_rsc_25_0_WDATA,
      x_rsc_25_0_AWREADY => x_rsc_25_0_AWREADY,
      x_rsc_25_0_AWVALID => x_rsc_25_0_AWVALID,
      x_rsc_25_0_AWUSER => x_rsc_25_0_AWUSER,
      x_rsc_25_0_AWREGION => hybrid_core_inst_x_rsc_25_0_AWREGION,
      x_rsc_25_0_AWQOS => hybrid_core_inst_x_rsc_25_0_AWQOS,
      x_rsc_25_0_AWPROT => hybrid_core_inst_x_rsc_25_0_AWPROT,
      x_rsc_25_0_AWCACHE => hybrid_core_inst_x_rsc_25_0_AWCACHE,
      x_rsc_25_0_AWLOCK => x_rsc_25_0_AWLOCK,
      x_rsc_25_0_AWBURST => hybrid_core_inst_x_rsc_25_0_AWBURST,
      x_rsc_25_0_AWSIZE => hybrid_core_inst_x_rsc_25_0_AWSIZE,
      x_rsc_25_0_AWLEN => hybrid_core_inst_x_rsc_25_0_AWLEN,
      x_rsc_25_0_AWADDR => hybrid_core_inst_x_rsc_25_0_AWADDR,
      x_rsc_25_0_AWID => x_rsc_25_0_AWID,
      x_rsc_triosy_25_0_lz => x_rsc_triosy_25_0_lz,
      x_rsc_26_0_s_tdone => x_rsc_26_0_s_tdone,
      x_rsc_26_0_tr_write_done => x_rsc_26_0_tr_write_done,
      x_rsc_26_0_RREADY => x_rsc_26_0_RREADY,
      x_rsc_26_0_RVALID => x_rsc_26_0_RVALID,
      x_rsc_26_0_RUSER => x_rsc_26_0_RUSER,
      x_rsc_26_0_RLAST => x_rsc_26_0_RLAST,
      x_rsc_26_0_RRESP => hybrid_core_inst_x_rsc_26_0_RRESP,
      x_rsc_26_0_RDATA => hybrid_core_inst_x_rsc_26_0_RDATA,
      x_rsc_26_0_RID => x_rsc_26_0_RID,
      x_rsc_26_0_ARREADY => x_rsc_26_0_ARREADY,
      x_rsc_26_0_ARVALID => x_rsc_26_0_ARVALID,
      x_rsc_26_0_ARUSER => x_rsc_26_0_ARUSER,
      x_rsc_26_0_ARREGION => hybrid_core_inst_x_rsc_26_0_ARREGION,
      x_rsc_26_0_ARQOS => hybrid_core_inst_x_rsc_26_0_ARQOS,
      x_rsc_26_0_ARPROT => hybrid_core_inst_x_rsc_26_0_ARPROT,
      x_rsc_26_0_ARCACHE => hybrid_core_inst_x_rsc_26_0_ARCACHE,
      x_rsc_26_0_ARLOCK => x_rsc_26_0_ARLOCK,
      x_rsc_26_0_ARBURST => hybrid_core_inst_x_rsc_26_0_ARBURST,
      x_rsc_26_0_ARSIZE => hybrid_core_inst_x_rsc_26_0_ARSIZE,
      x_rsc_26_0_ARLEN => hybrid_core_inst_x_rsc_26_0_ARLEN,
      x_rsc_26_0_ARADDR => hybrid_core_inst_x_rsc_26_0_ARADDR,
      x_rsc_26_0_ARID => x_rsc_26_0_ARID,
      x_rsc_26_0_BREADY => x_rsc_26_0_BREADY,
      x_rsc_26_0_BVALID => x_rsc_26_0_BVALID,
      x_rsc_26_0_BUSER => x_rsc_26_0_BUSER,
      x_rsc_26_0_BRESP => hybrid_core_inst_x_rsc_26_0_BRESP,
      x_rsc_26_0_BID => x_rsc_26_0_BID,
      x_rsc_26_0_WREADY => x_rsc_26_0_WREADY,
      x_rsc_26_0_WVALID => x_rsc_26_0_WVALID,
      x_rsc_26_0_WUSER => x_rsc_26_0_WUSER,
      x_rsc_26_0_WLAST => x_rsc_26_0_WLAST,
      x_rsc_26_0_WSTRB => hybrid_core_inst_x_rsc_26_0_WSTRB,
      x_rsc_26_0_WDATA => hybrid_core_inst_x_rsc_26_0_WDATA,
      x_rsc_26_0_AWREADY => x_rsc_26_0_AWREADY,
      x_rsc_26_0_AWVALID => x_rsc_26_0_AWVALID,
      x_rsc_26_0_AWUSER => x_rsc_26_0_AWUSER,
      x_rsc_26_0_AWREGION => hybrid_core_inst_x_rsc_26_0_AWREGION,
      x_rsc_26_0_AWQOS => hybrid_core_inst_x_rsc_26_0_AWQOS,
      x_rsc_26_0_AWPROT => hybrid_core_inst_x_rsc_26_0_AWPROT,
      x_rsc_26_0_AWCACHE => hybrid_core_inst_x_rsc_26_0_AWCACHE,
      x_rsc_26_0_AWLOCK => x_rsc_26_0_AWLOCK,
      x_rsc_26_0_AWBURST => hybrid_core_inst_x_rsc_26_0_AWBURST,
      x_rsc_26_0_AWSIZE => hybrid_core_inst_x_rsc_26_0_AWSIZE,
      x_rsc_26_0_AWLEN => hybrid_core_inst_x_rsc_26_0_AWLEN,
      x_rsc_26_0_AWADDR => hybrid_core_inst_x_rsc_26_0_AWADDR,
      x_rsc_26_0_AWID => x_rsc_26_0_AWID,
      x_rsc_triosy_26_0_lz => x_rsc_triosy_26_0_lz,
      x_rsc_27_0_s_tdone => x_rsc_27_0_s_tdone,
      x_rsc_27_0_tr_write_done => x_rsc_27_0_tr_write_done,
      x_rsc_27_0_RREADY => x_rsc_27_0_RREADY,
      x_rsc_27_0_RVALID => x_rsc_27_0_RVALID,
      x_rsc_27_0_RUSER => x_rsc_27_0_RUSER,
      x_rsc_27_0_RLAST => x_rsc_27_0_RLAST,
      x_rsc_27_0_RRESP => hybrid_core_inst_x_rsc_27_0_RRESP,
      x_rsc_27_0_RDATA => hybrid_core_inst_x_rsc_27_0_RDATA,
      x_rsc_27_0_RID => x_rsc_27_0_RID,
      x_rsc_27_0_ARREADY => x_rsc_27_0_ARREADY,
      x_rsc_27_0_ARVALID => x_rsc_27_0_ARVALID,
      x_rsc_27_0_ARUSER => x_rsc_27_0_ARUSER,
      x_rsc_27_0_ARREGION => hybrid_core_inst_x_rsc_27_0_ARREGION,
      x_rsc_27_0_ARQOS => hybrid_core_inst_x_rsc_27_0_ARQOS,
      x_rsc_27_0_ARPROT => hybrid_core_inst_x_rsc_27_0_ARPROT,
      x_rsc_27_0_ARCACHE => hybrid_core_inst_x_rsc_27_0_ARCACHE,
      x_rsc_27_0_ARLOCK => x_rsc_27_0_ARLOCK,
      x_rsc_27_0_ARBURST => hybrid_core_inst_x_rsc_27_0_ARBURST,
      x_rsc_27_0_ARSIZE => hybrid_core_inst_x_rsc_27_0_ARSIZE,
      x_rsc_27_0_ARLEN => hybrid_core_inst_x_rsc_27_0_ARLEN,
      x_rsc_27_0_ARADDR => hybrid_core_inst_x_rsc_27_0_ARADDR,
      x_rsc_27_0_ARID => x_rsc_27_0_ARID,
      x_rsc_27_0_BREADY => x_rsc_27_0_BREADY,
      x_rsc_27_0_BVALID => x_rsc_27_0_BVALID,
      x_rsc_27_0_BUSER => x_rsc_27_0_BUSER,
      x_rsc_27_0_BRESP => hybrid_core_inst_x_rsc_27_0_BRESP,
      x_rsc_27_0_BID => x_rsc_27_0_BID,
      x_rsc_27_0_WREADY => x_rsc_27_0_WREADY,
      x_rsc_27_0_WVALID => x_rsc_27_0_WVALID,
      x_rsc_27_0_WUSER => x_rsc_27_0_WUSER,
      x_rsc_27_0_WLAST => x_rsc_27_0_WLAST,
      x_rsc_27_0_WSTRB => hybrid_core_inst_x_rsc_27_0_WSTRB,
      x_rsc_27_0_WDATA => hybrid_core_inst_x_rsc_27_0_WDATA,
      x_rsc_27_0_AWREADY => x_rsc_27_0_AWREADY,
      x_rsc_27_0_AWVALID => x_rsc_27_0_AWVALID,
      x_rsc_27_0_AWUSER => x_rsc_27_0_AWUSER,
      x_rsc_27_0_AWREGION => hybrid_core_inst_x_rsc_27_0_AWREGION,
      x_rsc_27_0_AWQOS => hybrid_core_inst_x_rsc_27_0_AWQOS,
      x_rsc_27_0_AWPROT => hybrid_core_inst_x_rsc_27_0_AWPROT,
      x_rsc_27_0_AWCACHE => hybrid_core_inst_x_rsc_27_0_AWCACHE,
      x_rsc_27_0_AWLOCK => x_rsc_27_0_AWLOCK,
      x_rsc_27_0_AWBURST => hybrid_core_inst_x_rsc_27_0_AWBURST,
      x_rsc_27_0_AWSIZE => hybrid_core_inst_x_rsc_27_0_AWSIZE,
      x_rsc_27_0_AWLEN => hybrid_core_inst_x_rsc_27_0_AWLEN,
      x_rsc_27_0_AWADDR => hybrid_core_inst_x_rsc_27_0_AWADDR,
      x_rsc_27_0_AWID => x_rsc_27_0_AWID,
      x_rsc_triosy_27_0_lz => x_rsc_triosy_27_0_lz,
      x_rsc_28_0_s_tdone => x_rsc_28_0_s_tdone,
      x_rsc_28_0_tr_write_done => x_rsc_28_0_tr_write_done,
      x_rsc_28_0_RREADY => x_rsc_28_0_RREADY,
      x_rsc_28_0_RVALID => x_rsc_28_0_RVALID,
      x_rsc_28_0_RUSER => x_rsc_28_0_RUSER,
      x_rsc_28_0_RLAST => x_rsc_28_0_RLAST,
      x_rsc_28_0_RRESP => hybrid_core_inst_x_rsc_28_0_RRESP,
      x_rsc_28_0_RDATA => hybrid_core_inst_x_rsc_28_0_RDATA,
      x_rsc_28_0_RID => x_rsc_28_0_RID,
      x_rsc_28_0_ARREADY => x_rsc_28_0_ARREADY,
      x_rsc_28_0_ARVALID => x_rsc_28_0_ARVALID,
      x_rsc_28_0_ARUSER => x_rsc_28_0_ARUSER,
      x_rsc_28_0_ARREGION => hybrid_core_inst_x_rsc_28_0_ARREGION,
      x_rsc_28_0_ARQOS => hybrid_core_inst_x_rsc_28_0_ARQOS,
      x_rsc_28_0_ARPROT => hybrid_core_inst_x_rsc_28_0_ARPROT,
      x_rsc_28_0_ARCACHE => hybrid_core_inst_x_rsc_28_0_ARCACHE,
      x_rsc_28_0_ARLOCK => x_rsc_28_0_ARLOCK,
      x_rsc_28_0_ARBURST => hybrid_core_inst_x_rsc_28_0_ARBURST,
      x_rsc_28_0_ARSIZE => hybrid_core_inst_x_rsc_28_0_ARSIZE,
      x_rsc_28_0_ARLEN => hybrid_core_inst_x_rsc_28_0_ARLEN,
      x_rsc_28_0_ARADDR => hybrid_core_inst_x_rsc_28_0_ARADDR,
      x_rsc_28_0_ARID => x_rsc_28_0_ARID,
      x_rsc_28_0_BREADY => x_rsc_28_0_BREADY,
      x_rsc_28_0_BVALID => x_rsc_28_0_BVALID,
      x_rsc_28_0_BUSER => x_rsc_28_0_BUSER,
      x_rsc_28_0_BRESP => hybrid_core_inst_x_rsc_28_0_BRESP,
      x_rsc_28_0_BID => x_rsc_28_0_BID,
      x_rsc_28_0_WREADY => x_rsc_28_0_WREADY,
      x_rsc_28_0_WVALID => x_rsc_28_0_WVALID,
      x_rsc_28_0_WUSER => x_rsc_28_0_WUSER,
      x_rsc_28_0_WLAST => x_rsc_28_0_WLAST,
      x_rsc_28_0_WSTRB => hybrid_core_inst_x_rsc_28_0_WSTRB,
      x_rsc_28_0_WDATA => hybrid_core_inst_x_rsc_28_0_WDATA,
      x_rsc_28_0_AWREADY => x_rsc_28_0_AWREADY,
      x_rsc_28_0_AWVALID => x_rsc_28_0_AWVALID,
      x_rsc_28_0_AWUSER => x_rsc_28_0_AWUSER,
      x_rsc_28_0_AWREGION => hybrid_core_inst_x_rsc_28_0_AWREGION,
      x_rsc_28_0_AWQOS => hybrid_core_inst_x_rsc_28_0_AWQOS,
      x_rsc_28_0_AWPROT => hybrid_core_inst_x_rsc_28_0_AWPROT,
      x_rsc_28_0_AWCACHE => hybrid_core_inst_x_rsc_28_0_AWCACHE,
      x_rsc_28_0_AWLOCK => x_rsc_28_0_AWLOCK,
      x_rsc_28_0_AWBURST => hybrid_core_inst_x_rsc_28_0_AWBURST,
      x_rsc_28_0_AWSIZE => hybrid_core_inst_x_rsc_28_0_AWSIZE,
      x_rsc_28_0_AWLEN => hybrid_core_inst_x_rsc_28_0_AWLEN,
      x_rsc_28_0_AWADDR => hybrid_core_inst_x_rsc_28_0_AWADDR,
      x_rsc_28_0_AWID => x_rsc_28_0_AWID,
      x_rsc_triosy_28_0_lz => x_rsc_triosy_28_0_lz,
      x_rsc_29_0_s_tdone => x_rsc_29_0_s_tdone,
      x_rsc_29_0_tr_write_done => x_rsc_29_0_tr_write_done,
      x_rsc_29_0_RREADY => x_rsc_29_0_RREADY,
      x_rsc_29_0_RVALID => x_rsc_29_0_RVALID,
      x_rsc_29_0_RUSER => x_rsc_29_0_RUSER,
      x_rsc_29_0_RLAST => x_rsc_29_0_RLAST,
      x_rsc_29_0_RRESP => hybrid_core_inst_x_rsc_29_0_RRESP,
      x_rsc_29_0_RDATA => hybrid_core_inst_x_rsc_29_0_RDATA,
      x_rsc_29_0_RID => x_rsc_29_0_RID,
      x_rsc_29_0_ARREADY => x_rsc_29_0_ARREADY,
      x_rsc_29_0_ARVALID => x_rsc_29_0_ARVALID,
      x_rsc_29_0_ARUSER => x_rsc_29_0_ARUSER,
      x_rsc_29_0_ARREGION => hybrid_core_inst_x_rsc_29_0_ARREGION,
      x_rsc_29_0_ARQOS => hybrid_core_inst_x_rsc_29_0_ARQOS,
      x_rsc_29_0_ARPROT => hybrid_core_inst_x_rsc_29_0_ARPROT,
      x_rsc_29_0_ARCACHE => hybrid_core_inst_x_rsc_29_0_ARCACHE,
      x_rsc_29_0_ARLOCK => x_rsc_29_0_ARLOCK,
      x_rsc_29_0_ARBURST => hybrid_core_inst_x_rsc_29_0_ARBURST,
      x_rsc_29_0_ARSIZE => hybrid_core_inst_x_rsc_29_0_ARSIZE,
      x_rsc_29_0_ARLEN => hybrid_core_inst_x_rsc_29_0_ARLEN,
      x_rsc_29_0_ARADDR => hybrid_core_inst_x_rsc_29_0_ARADDR,
      x_rsc_29_0_ARID => x_rsc_29_0_ARID,
      x_rsc_29_0_BREADY => x_rsc_29_0_BREADY,
      x_rsc_29_0_BVALID => x_rsc_29_0_BVALID,
      x_rsc_29_0_BUSER => x_rsc_29_0_BUSER,
      x_rsc_29_0_BRESP => hybrid_core_inst_x_rsc_29_0_BRESP,
      x_rsc_29_0_BID => x_rsc_29_0_BID,
      x_rsc_29_0_WREADY => x_rsc_29_0_WREADY,
      x_rsc_29_0_WVALID => x_rsc_29_0_WVALID,
      x_rsc_29_0_WUSER => x_rsc_29_0_WUSER,
      x_rsc_29_0_WLAST => x_rsc_29_0_WLAST,
      x_rsc_29_0_WSTRB => hybrid_core_inst_x_rsc_29_0_WSTRB,
      x_rsc_29_0_WDATA => hybrid_core_inst_x_rsc_29_0_WDATA,
      x_rsc_29_0_AWREADY => x_rsc_29_0_AWREADY,
      x_rsc_29_0_AWVALID => x_rsc_29_0_AWVALID,
      x_rsc_29_0_AWUSER => x_rsc_29_0_AWUSER,
      x_rsc_29_0_AWREGION => hybrid_core_inst_x_rsc_29_0_AWREGION,
      x_rsc_29_0_AWQOS => hybrid_core_inst_x_rsc_29_0_AWQOS,
      x_rsc_29_0_AWPROT => hybrid_core_inst_x_rsc_29_0_AWPROT,
      x_rsc_29_0_AWCACHE => hybrid_core_inst_x_rsc_29_0_AWCACHE,
      x_rsc_29_0_AWLOCK => x_rsc_29_0_AWLOCK,
      x_rsc_29_0_AWBURST => hybrid_core_inst_x_rsc_29_0_AWBURST,
      x_rsc_29_0_AWSIZE => hybrid_core_inst_x_rsc_29_0_AWSIZE,
      x_rsc_29_0_AWLEN => hybrid_core_inst_x_rsc_29_0_AWLEN,
      x_rsc_29_0_AWADDR => hybrid_core_inst_x_rsc_29_0_AWADDR,
      x_rsc_29_0_AWID => x_rsc_29_0_AWID,
      x_rsc_triosy_29_0_lz => x_rsc_triosy_29_0_lz,
      x_rsc_30_0_s_tdone => x_rsc_30_0_s_tdone,
      x_rsc_30_0_tr_write_done => x_rsc_30_0_tr_write_done,
      x_rsc_30_0_RREADY => x_rsc_30_0_RREADY,
      x_rsc_30_0_RVALID => x_rsc_30_0_RVALID,
      x_rsc_30_0_RUSER => x_rsc_30_0_RUSER,
      x_rsc_30_0_RLAST => x_rsc_30_0_RLAST,
      x_rsc_30_0_RRESP => hybrid_core_inst_x_rsc_30_0_RRESP,
      x_rsc_30_0_RDATA => hybrid_core_inst_x_rsc_30_0_RDATA,
      x_rsc_30_0_RID => x_rsc_30_0_RID,
      x_rsc_30_0_ARREADY => x_rsc_30_0_ARREADY,
      x_rsc_30_0_ARVALID => x_rsc_30_0_ARVALID,
      x_rsc_30_0_ARUSER => x_rsc_30_0_ARUSER,
      x_rsc_30_0_ARREGION => hybrid_core_inst_x_rsc_30_0_ARREGION,
      x_rsc_30_0_ARQOS => hybrid_core_inst_x_rsc_30_0_ARQOS,
      x_rsc_30_0_ARPROT => hybrid_core_inst_x_rsc_30_0_ARPROT,
      x_rsc_30_0_ARCACHE => hybrid_core_inst_x_rsc_30_0_ARCACHE,
      x_rsc_30_0_ARLOCK => x_rsc_30_0_ARLOCK,
      x_rsc_30_0_ARBURST => hybrid_core_inst_x_rsc_30_0_ARBURST,
      x_rsc_30_0_ARSIZE => hybrid_core_inst_x_rsc_30_0_ARSIZE,
      x_rsc_30_0_ARLEN => hybrid_core_inst_x_rsc_30_0_ARLEN,
      x_rsc_30_0_ARADDR => hybrid_core_inst_x_rsc_30_0_ARADDR,
      x_rsc_30_0_ARID => x_rsc_30_0_ARID,
      x_rsc_30_0_BREADY => x_rsc_30_0_BREADY,
      x_rsc_30_0_BVALID => x_rsc_30_0_BVALID,
      x_rsc_30_0_BUSER => x_rsc_30_0_BUSER,
      x_rsc_30_0_BRESP => hybrid_core_inst_x_rsc_30_0_BRESP,
      x_rsc_30_0_BID => x_rsc_30_0_BID,
      x_rsc_30_0_WREADY => x_rsc_30_0_WREADY,
      x_rsc_30_0_WVALID => x_rsc_30_0_WVALID,
      x_rsc_30_0_WUSER => x_rsc_30_0_WUSER,
      x_rsc_30_0_WLAST => x_rsc_30_0_WLAST,
      x_rsc_30_0_WSTRB => hybrid_core_inst_x_rsc_30_0_WSTRB,
      x_rsc_30_0_WDATA => hybrid_core_inst_x_rsc_30_0_WDATA,
      x_rsc_30_0_AWREADY => x_rsc_30_0_AWREADY,
      x_rsc_30_0_AWVALID => x_rsc_30_0_AWVALID,
      x_rsc_30_0_AWUSER => x_rsc_30_0_AWUSER,
      x_rsc_30_0_AWREGION => hybrid_core_inst_x_rsc_30_0_AWREGION,
      x_rsc_30_0_AWQOS => hybrid_core_inst_x_rsc_30_0_AWQOS,
      x_rsc_30_0_AWPROT => hybrid_core_inst_x_rsc_30_0_AWPROT,
      x_rsc_30_0_AWCACHE => hybrid_core_inst_x_rsc_30_0_AWCACHE,
      x_rsc_30_0_AWLOCK => x_rsc_30_0_AWLOCK,
      x_rsc_30_0_AWBURST => hybrid_core_inst_x_rsc_30_0_AWBURST,
      x_rsc_30_0_AWSIZE => hybrid_core_inst_x_rsc_30_0_AWSIZE,
      x_rsc_30_0_AWLEN => hybrid_core_inst_x_rsc_30_0_AWLEN,
      x_rsc_30_0_AWADDR => hybrid_core_inst_x_rsc_30_0_AWADDR,
      x_rsc_30_0_AWID => x_rsc_30_0_AWID,
      x_rsc_triosy_30_0_lz => x_rsc_triosy_30_0_lz,
      x_rsc_31_0_s_tdone => x_rsc_31_0_s_tdone,
      x_rsc_31_0_tr_write_done => x_rsc_31_0_tr_write_done,
      x_rsc_31_0_RREADY => x_rsc_31_0_RREADY,
      x_rsc_31_0_RVALID => x_rsc_31_0_RVALID,
      x_rsc_31_0_RUSER => x_rsc_31_0_RUSER,
      x_rsc_31_0_RLAST => x_rsc_31_0_RLAST,
      x_rsc_31_0_RRESP => hybrid_core_inst_x_rsc_31_0_RRESP,
      x_rsc_31_0_RDATA => hybrid_core_inst_x_rsc_31_0_RDATA,
      x_rsc_31_0_RID => x_rsc_31_0_RID,
      x_rsc_31_0_ARREADY => x_rsc_31_0_ARREADY,
      x_rsc_31_0_ARVALID => x_rsc_31_0_ARVALID,
      x_rsc_31_0_ARUSER => x_rsc_31_0_ARUSER,
      x_rsc_31_0_ARREGION => hybrid_core_inst_x_rsc_31_0_ARREGION,
      x_rsc_31_0_ARQOS => hybrid_core_inst_x_rsc_31_0_ARQOS,
      x_rsc_31_0_ARPROT => hybrid_core_inst_x_rsc_31_0_ARPROT,
      x_rsc_31_0_ARCACHE => hybrid_core_inst_x_rsc_31_0_ARCACHE,
      x_rsc_31_0_ARLOCK => x_rsc_31_0_ARLOCK,
      x_rsc_31_0_ARBURST => hybrid_core_inst_x_rsc_31_0_ARBURST,
      x_rsc_31_0_ARSIZE => hybrid_core_inst_x_rsc_31_0_ARSIZE,
      x_rsc_31_0_ARLEN => hybrid_core_inst_x_rsc_31_0_ARLEN,
      x_rsc_31_0_ARADDR => hybrid_core_inst_x_rsc_31_0_ARADDR,
      x_rsc_31_0_ARID => x_rsc_31_0_ARID,
      x_rsc_31_0_BREADY => x_rsc_31_0_BREADY,
      x_rsc_31_0_BVALID => x_rsc_31_0_BVALID,
      x_rsc_31_0_BUSER => x_rsc_31_0_BUSER,
      x_rsc_31_0_BRESP => hybrid_core_inst_x_rsc_31_0_BRESP,
      x_rsc_31_0_BID => x_rsc_31_0_BID,
      x_rsc_31_0_WREADY => x_rsc_31_0_WREADY,
      x_rsc_31_0_WVALID => x_rsc_31_0_WVALID,
      x_rsc_31_0_WUSER => x_rsc_31_0_WUSER,
      x_rsc_31_0_WLAST => x_rsc_31_0_WLAST,
      x_rsc_31_0_WSTRB => hybrid_core_inst_x_rsc_31_0_WSTRB,
      x_rsc_31_0_WDATA => hybrid_core_inst_x_rsc_31_0_WDATA,
      x_rsc_31_0_AWREADY => x_rsc_31_0_AWREADY,
      x_rsc_31_0_AWVALID => x_rsc_31_0_AWVALID,
      x_rsc_31_0_AWUSER => x_rsc_31_0_AWUSER,
      x_rsc_31_0_AWREGION => hybrid_core_inst_x_rsc_31_0_AWREGION,
      x_rsc_31_0_AWQOS => hybrid_core_inst_x_rsc_31_0_AWQOS,
      x_rsc_31_0_AWPROT => hybrid_core_inst_x_rsc_31_0_AWPROT,
      x_rsc_31_0_AWCACHE => hybrid_core_inst_x_rsc_31_0_AWCACHE,
      x_rsc_31_0_AWLOCK => x_rsc_31_0_AWLOCK,
      x_rsc_31_0_AWBURST => hybrid_core_inst_x_rsc_31_0_AWBURST,
      x_rsc_31_0_AWSIZE => hybrid_core_inst_x_rsc_31_0_AWSIZE,
      x_rsc_31_0_AWLEN => hybrid_core_inst_x_rsc_31_0_AWLEN,
      x_rsc_31_0_AWADDR => hybrid_core_inst_x_rsc_31_0_AWADDR,
      x_rsc_31_0_AWID => x_rsc_31_0_AWID,
      x_rsc_triosy_31_0_lz => x_rsc_triosy_31_0_lz,
      m_rsc_dat => hybrid_core_inst_m_rsc_dat,
      m_rsc_triosy_lz => m_rsc_triosy_lz,
      twiddle_rsc_triosy_lz => twiddle_rsc_triosy_lz,
      twiddle_h_rsc_triosy_lz => twiddle_h_rsc_triosy_lz,
      revArr_rsc_s_tdone => revArr_rsc_s_tdone,
      revArr_rsc_tr_write_done => revArr_rsc_tr_write_done,
      revArr_rsc_RREADY => revArr_rsc_RREADY,
      revArr_rsc_RVALID => revArr_rsc_RVALID,
      revArr_rsc_RUSER => revArr_rsc_RUSER,
      revArr_rsc_RLAST => revArr_rsc_RLAST,
      revArr_rsc_RRESP => hybrid_core_inst_revArr_rsc_RRESP,
      revArr_rsc_RDATA => hybrid_core_inst_revArr_rsc_RDATA,
      revArr_rsc_RID => revArr_rsc_RID,
      revArr_rsc_ARREADY => revArr_rsc_ARREADY,
      revArr_rsc_ARVALID => revArr_rsc_ARVALID,
      revArr_rsc_ARUSER => revArr_rsc_ARUSER,
      revArr_rsc_ARREGION => hybrid_core_inst_revArr_rsc_ARREGION,
      revArr_rsc_ARQOS => hybrid_core_inst_revArr_rsc_ARQOS,
      revArr_rsc_ARPROT => hybrid_core_inst_revArr_rsc_ARPROT,
      revArr_rsc_ARCACHE => hybrid_core_inst_revArr_rsc_ARCACHE,
      revArr_rsc_ARLOCK => revArr_rsc_ARLOCK,
      revArr_rsc_ARBURST => hybrid_core_inst_revArr_rsc_ARBURST,
      revArr_rsc_ARSIZE => hybrid_core_inst_revArr_rsc_ARSIZE,
      revArr_rsc_ARLEN => hybrid_core_inst_revArr_rsc_ARLEN,
      revArr_rsc_ARADDR => hybrid_core_inst_revArr_rsc_ARADDR,
      revArr_rsc_ARID => revArr_rsc_ARID,
      revArr_rsc_BREADY => revArr_rsc_BREADY,
      revArr_rsc_BVALID => revArr_rsc_BVALID,
      revArr_rsc_BUSER => revArr_rsc_BUSER,
      revArr_rsc_BRESP => hybrid_core_inst_revArr_rsc_BRESP,
      revArr_rsc_BID => revArr_rsc_BID,
      revArr_rsc_WREADY => revArr_rsc_WREADY,
      revArr_rsc_WVALID => revArr_rsc_WVALID,
      revArr_rsc_WUSER => revArr_rsc_WUSER,
      revArr_rsc_WLAST => revArr_rsc_WLAST,
      revArr_rsc_WSTRB => hybrid_core_inst_revArr_rsc_WSTRB,
      revArr_rsc_WDATA => hybrid_core_inst_revArr_rsc_WDATA,
      revArr_rsc_AWREADY => revArr_rsc_AWREADY,
      revArr_rsc_AWVALID => revArr_rsc_AWVALID,
      revArr_rsc_AWUSER => revArr_rsc_AWUSER,
      revArr_rsc_AWREGION => hybrid_core_inst_revArr_rsc_AWREGION,
      revArr_rsc_AWQOS => hybrid_core_inst_revArr_rsc_AWQOS,
      revArr_rsc_AWPROT => hybrid_core_inst_revArr_rsc_AWPROT,
      revArr_rsc_AWCACHE => hybrid_core_inst_revArr_rsc_AWCACHE,
      revArr_rsc_AWLOCK => revArr_rsc_AWLOCK,
      revArr_rsc_AWBURST => hybrid_core_inst_revArr_rsc_AWBURST,
      revArr_rsc_AWSIZE => hybrid_core_inst_revArr_rsc_AWSIZE,
      revArr_rsc_AWLEN => hybrid_core_inst_revArr_rsc_AWLEN,
      revArr_rsc_AWADDR => hybrid_core_inst_revArr_rsc_AWADDR,
      revArr_rsc_AWID => revArr_rsc_AWID,
      revArr_rsc_triosy_lz => revArr_rsc_triosy_lz,
      tw_rsc_s_tdone => tw_rsc_s_tdone,
      tw_rsc_tr_write_done => tw_rsc_tr_write_done,
      tw_rsc_RREADY => tw_rsc_RREADY,
      tw_rsc_RVALID => tw_rsc_RVALID,
      tw_rsc_RUSER => tw_rsc_RUSER,
      tw_rsc_RLAST => tw_rsc_RLAST,
      tw_rsc_RRESP => hybrid_core_inst_tw_rsc_RRESP,
      tw_rsc_RDATA => hybrid_core_inst_tw_rsc_RDATA,
      tw_rsc_RID => tw_rsc_RID,
      tw_rsc_ARREADY => tw_rsc_ARREADY,
      tw_rsc_ARVALID => tw_rsc_ARVALID,
      tw_rsc_ARUSER => tw_rsc_ARUSER,
      tw_rsc_ARREGION => hybrid_core_inst_tw_rsc_ARREGION,
      tw_rsc_ARQOS => hybrid_core_inst_tw_rsc_ARQOS,
      tw_rsc_ARPROT => hybrid_core_inst_tw_rsc_ARPROT,
      tw_rsc_ARCACHE => hybrid_core_inst_tw_rsc_ARCACHE,
      tw_rsc_ARLOCK => tw_rsc_ARLOCK,
      tw_rsc_ARBURST => hybrid_core_inst_tw_rsc_ARBURST,
      tw_rsc_ARSIZE => hybrid_core_inst_tw_rsc_ARSIZE,
      tw_rsc_ARLEN => hybrid_core_inst_tw_rsc_ARLEN,
      tw_rsc_ARADDR => hybrid_core_inst_tw_rsc_ARADDR,
      tw_rsc_ARID => tw_rsc_ARID,
      tw_rsc_BREADY => tw_rsc_BREADY,
      tw_rsc_BVALID => tw_rsc_BVALID,
      tw_rsc_BUSER => tw_rsc_BUSER,
      tw_rsc_BRESP => hybrid_core_inst_tw_rsc_BRESP,
      tw_rsc_BID => tw_rsc_BID,
      tw_rsc_WREADY => tw_rsc_WREADY,
      tw_rsc_WVALID => tw_rsc_WVALID,
      tw_rsc_WUSER => tw_rsc_WUSER,
      tw_rsc_WLAST => tw_rsc_WLAST,
      tw_rsc_WSTRB => hybrid_core_inst_tw_rsc_WSTRB,
      tw_rsc_WDATA => hybrid_core_inst_tw_rsc_WDATA,
      tw_rsc_AWREADY => tw_rsc_AWREADY,
      tw_rsc_AWVALID => tw_rsc_AWVALID,
      tw_rsc_AWUSER => tw_rsc_AWUSER,
      tw_rsc_AWREGION => hybrid_core_inst_tw_rsc_AWREGION,
      tw_rsc_AWQOS => hybrid_core_inst_tw_rsc_AWQOS,
      tw_rsc_AWPROT => hybrid_core_inst_tw_rsc_AWPROT,
      tw_rsc_AWCACHE => hybrid_core_inst_tw_rsc_AWCACHE,
      tw_rsc_AWLOCK => tw_rsc_AWLOCK,
      tw_rsc_AWBURST => hybrid_core_inst_tw_rsc_AWBURST,
      tw_rsc_AWSIZE => hybrid_core_inst_tw_rsc_AWSIZE,
      tw_rsc_AWLEN => hybrid_core_inst_tw_rsc_AWLEN,
      tw_rsc_AWADDR => hybrid_core_inst_tw_rsc_AWADDR,
      tw_rsc_AWID => tw_rsc_AWID,
      tw_rsc_triosy_lz => tw_rsc_triosy_lz,
      tw_h_rsc_s_tdone => tw_h_rsc_s_tdone,
      tw_h_rsc_tr_write_done => tw_h_rsc_tr_write_done,
      tw_h_rsc_RREADY => tw_h_rsc_RREADY,
      tw_h_rsc_RVALID => tw_h_rsc_RVALID,
      tw_h_rsc_RUSER => tw_h_rsc_RUSER,
      tw_h_rsc_RLAST => tw_h_rsc_RLAST,
      tw_h_rsc_RRESP => hybrid_core_inst_tw_h_rsc_RRESP,
      tw_h_rsc_RDATA => hybrid_core_inst_tw_h_rsc_RDATA,
      tw_h_rsc_RID => tw_h_rsc_RID,
      tw_h_rsc_ARREADY => tw_h_rsc_ARREADY,
      tw_h_rsc_ARVALID => tw_h_rsc_ARVALID,
      tw_h_rsc_ARUSER => tw_h_rsc_ARUSER,
      tw_h_rsc_ARREGION => hybrid_core_inst_tw_h_rsc_ARREGION,
      tw_h_rsc_ARQOS => hybrid_core_inst_tw_h_rsc_ARQOS,
      tw_h_rsc_ARPROT => hybrid_core_inst_tw_h_rsc_ARPROT,
      tw_h_rsc_ARCACHE => hybrid_core_inst_tw_h_rsc_ARCACHE,
      tw_h_rsc_ARLOCK => tw_h_rsc_ARLOCK,
      tw_h_rsc_ARBURST => hybrid_core_inst_tw_h_rsc_ARBURST,
      tw_h_rsc_ARSIZE => hybrid_core_inst_tw_h_rsc_ARSIZE,
      tw_h_rsc_ARLEN => hybrid_core_inst_tw_h_rsc_ARLEN,
      tw_h_rsc_ARADDR => hybrid_core_inst_tw_h_rsc_ARADDR,
      tw_h_rsc_ARID => tw_h_rsc_ARID,
      tw_h_rsc_BREADY => tw_h_rsc_BREADY,
      tw_h_rsc_BVALID => tw_h_rsc_BVALID,
      tw_h_rsc_BUSER => tw_h_rsc_BUSER,
      tw_h_rsc_BRESP => hybrid_core_inst_tw_h_rsc_BRESP,
      tw_h_rsc_BID => tw_h_rsc_BID,
      tw_h_rsc_WREADY => tw_h_rsc_WREADY,
      tw_h_rsc_WVALID => tw_h_rsc_WVALID,
      tw_h_rsc_WUSER => tw_h_rsc_WUSER,
      tw_h_rsc_WLAST => tw_h_rsc_WLAST,
      tw_h_rsc_WSTRB => hybrid_core_inst_tw_h_rsc_WSTRB,
      tw_h_rsc_WDATA => hybrid_core_inst_tw_h_rsc_WDATA,
      tw_h_rsc_AWREADY => tw_h_rsc_AWREADY,
      tw_h_rsc_AWVALID => tw_h_rsc_AWVALID,
      tw_h_rsc_AWUSER => tw_h_rsc_AWUSER,
      tw_h_rsc_AWREGION => hybrid_core_inst_tw_h_rsc_AWREGION,
      tw_h_rsc_AWQOS => hybrid_core_inst_tw_h_rsc_AWQOS,
      tw_h_rsc_AWPROT => hybrid_core_inst_tw_h_rsc_AWPROT,
      tw_h_rsc_AWCACHE => hybrid_core_inst_tw_h_rsc_AWCACHE,
      tw_h_rsc_AWLOCK => tw_h_rsc_AWLOCK,
      tw_h_rsc_AWBURST => hybrid_core_inst_tw_h_rsc_AWBURST,
      tw_h_rsc_AWSIZE => hybrid_core_inst_tw_h_rsc_AWSIZE,
      tw_h_rsc_AWLEN => hybrid_core_inst_tw_h_rsc_AWLEN,
      tw_h_rsc_AWADDR => hybrid_core_inst_tw_h_rsc_AWADDR,
      tw_h_rsc_AWID => tw_h_rsc_AWID,
      tw_h_rsc_triosy_lz => tw_h_rsc_triosy_lz,
      twiddle_rsci_adrb_d => hybrid_core_inst_twiddle_rsci_adrb_d,
      twiddle_rsci_qb_d => hybrid_core_inst_twiddle_rsci_qb_d,
      twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d => twiddle_rsci_readB_r_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsci_adrb_d => hybrid_core_inst_twiddle_h_rsci_adrb_d,
      twiddle_h_rsci_qb_d => hybrid_core_inst_twiddle_h_rsci_qb_d,
      twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d => twiddle_h_rsci_readB_r_ram_ir_internal_RMASK_B_d,
      xx_rsc_0_0_i_adra_d => hybrid_core_inst_xx_rsc_0_0_i_adra_d,
      xx_rsc_0_0_i_clka_en_d => xx_rsc_0_0_i_clka_en_d,
      xx_rsc_0_0_i_qa_d => hybrid_core_inst_xx_rsc_0_0_i_qa_d,
      xx_rsc_0_0_i_wea_d => hybrid_core_inst_xx_rsc_0_0_i_wea_d,
      xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_1_0_i_adra_d => hybrid_core_inst_xx_rsc_1_0_i_adra_d,
      xx_rsc_1_0_i_clka_en_d => xx_rsc_1_0_i_clka_en_d,
      xx_rsc_1_0_i_qa_d => hybrid_core_inst_xx_rsc_1_0_i_qa_d,
      xx_rsc_1_0_i_wea_d => hybrid_core_inst_xx_rsc_1_0_i_wea_d,
      xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_2_0_i_adra_d => hybrid_core_inst_xx_rsc_2_0_i_adra_d,
      xx_rsc_2_0_i_clka_en_d => xx_rsc_2_0_i_clka_en_d,
      xx_rsc_2_0_i_qa_d => hybrid_core_inst_xx_rsc_2_0_i_qa_d,
      xx_rsc_2_0_i_wea_d => hybrid_core_inst_xx_rsc_2_0_i_wea_d,
      xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_3_0_i_adra_d => hybrid_core_inst_xx_rsc_3_0_i_adra_d,
      xx_rsc_3_0_i_clka_en_d => xx_rsc_3_0_i_clka_en_d,
      xx_rsc_3_0_i_qa_d => hybrid_core_inst_xx_rsc_3_0_i_qa_d,
      xx_rsc_3_0_i_wea_d => hybrid_core_inst_xx_rsc_3_0_i_wea_d,
      xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_4_0_i_adra_d => hybrid_core_inst_xx_rsc_4_0_i_adra_d,
      xx_rsc_4_0_i_clka_en_d => xx_rsc_4_0_i_clka_en_d,
      xx_rsc_4_0_i_qa_d => hybrid_core_inst_xx_rsc_4_0_i_qa_d,
      xx_rsc_4_0_i_wea_d => hybrid_core_inst_xx_rsc_4_0_i_wea_d,
      xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_5_0_i_adra_d => hybrid_core_inst_xx_rsc_5_0_i_adra_d,
      xx_rsc_5_0_i_clka_en_d => xx_rsc_5_0_i_clka_en_d,
      xx_rsc_5_0_i_qa_d => hybrid_core_inst_xx_rsc_5_0_i_qa_d,
      xx_rsc_5_0_i_wea_d => hybrid_core_inst_xx_rsc_5_0_i_wea_d,
      xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_6_0_i_adra_d => hybrid_core_inst_xx_rsc_6_0_i_adra_d,
      xx_rsc_6_0_i_clka_en_d => xx_rsc_6_0_i_clka_en_d,
      xx_rsc_6_0_i_qa_d => hybrid_core_inst_xx_rsc_6_0_i_qa_d,
      xx_rsc_6_0_i_wea_d => hybrid_core_inst_xx_rsc_6_0_i_wea_d,
      xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_7_0_i_adra_d => hybrid_core_inst_xx_rsc_7_0_i_adra_d,
      xx_rsc_7_0_i_clka_en_d => xx_rsc_7_0_i_clka_en_d,
      xx_rsc_7_0_i_qa_d => hybrid_core_inst_xx_rsc_7_0_i_qa_d,
      xx_rsc_7_0_i_wea_d => hybrid_core_inst_xx_rsc_7_0_i_wea_d,
      xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_8_0_i_adra_d => hybrid_core_inst_xx_rsc_8_0_i_adra_d,
      xx_rsc_8_0_i_clka_en_d => xx_rsc_8_0_i_clka_en_d,
      xx_rsc_8_0_i_qa_d => hybrid_core_inst_xx_rsc_8_0_i_qa_d,
      xx_rsc_8_0_i_wea_d => hybrid_core_inst_xx_rsc_8_0_i_wea_d,
      xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_9_0_i_adra_d => hybrid_core_inst_xx_rsc_9_0_i_adra_d,
      xx_rsc_9_0_i_clka_en_d => xx_rsc_9_0_i_clka_en_d,
      xx_rsc_9_0_i_qa_d => hybrid_core_inst_xx_rsc_9_0_i_qa_d,
      xx_rsc_9_0_i_wea_d => hybrid_core_inst_xx_rsc_9_0_i_wea_d,
      xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_10_0_i_adra_d => hybrid_core_inst_xx_rsc_10_0_i_adra_d,
      xx_rsc_10_0_i_clka_en_d => xx_rsc_10_0_i_clka_en_d,
      xx_rsc_10_0_i_qa_d => hybrid_core_inst_xx_rsc_10_0_i_qa_d,
      xx_rsc_10_0_i_wea_d => hybrid_core_inst_xx_rsc_10_0_i_wea_d,
      xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_11_0_i_adra_d => hybrid_core_inst_xx_rsc_11_0_i_adra_d,
      xx_rsc_11_0_i_clka_en_d => xx_rsc_11_0_i_clka_en_d,
      xx_rsc_11_0_i_qa_d => hybrid_core_inst_xx_rsc_11_0_i_qa_d,
      xx_rsc_11_0_i_wea_d => hybrid_core_inst_xx_rsc_11_0_i_wea_d,
      xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_12_0_i_adra_d => hybrid_core_inst_xx_rsc_12_0_i_adra_d,
      xx_rsc_12_0_i_clka_en_d => xx_rsc_12_0_i_clka_en_d,
      xx_rsc_12_0_i_qa_d => hybrid_core_inst_xx_rsc_12_0_i_qa_d,
      xx_rsc_12_0_i_wea_d => hybrid_core_inst_xx_rsc_12_0_i_wea_d,
      xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_13_0_i_adra_d => hybrid_core_inst_xx_rsc_13_0_i_adra_d,
      xx_rsc_13_0_i_clka_en_d => xx_rsc_13_0_i_clka_en_d,
      xx_rsc_13_0_i_qa_d => hybrid_core_inst_xx_rsc_13_0_i_qa_d,
      xx_rsc_13_0_i_wea_d => hybrid_core_inst_xx_rsc_13_0_i_wea_d,
      xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_14_0_i_adra_d => hybrid_core_inst_xx_rsc_14_0_i_adra_d,
      xx_rsc_14_0_i_clka_en_d => xx_rsc_14_0_i_clka_en_d,
      xx_rsc_14_0_i_qa_d => hybrid_core_inst_xx_rsc_14_0_i_qa_d,
      xx_rsc_14_0_i_wea_d => hybrid_core_inst_xx_rsc_14_0_i_wea_d,
      xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_15_0_i_adra_d => hybrid_core_inst_xx_rsc_15_0_i_adra_d,
      xx_rsc_15_0_i_clka_en_d => xx_rsc_15_0_i_clka_en_d,
      xx_rsc_15_0_i_qa_d => hybrid_core_inst_xx_rsc_15_0_i_qa_d,
      xx_rsc_15_0_i_wea_d => hybrid_core_inst_xx_rsc_15_0_i_wea_d,
      xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_16_0_i_adra_d => hybrid_core_inst_xx_rsc_16_0_i_adra_d,
      xx_rsc_16_0_i_clka_en_d => xx_rsc_16_0_i_clka_en_d,
      xx_rsc_16_0_i_qa_d => hybrid_core_inst_xx_rsc_16_0_i_qa_d,
      xx_rsc_16_0_i_wea_d => hybrid_core_inst_xx_rsc_16_0_i_wea_d,
      xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_17_0_i_adra_d => hybrid_core_inst_xx_rsc_17_0_i_adra_d,
      xx_rsc_17_0_i_clka_en_d => xx_rsc_17_0_i_clka_en_d,
      xx_rsc_17_0_i_qa_d => hybrid_core_inst_xx_rsc_17_0_i_qa_d,
      xx_rsc_17_0_i_wea_d => hybrid_core_inst_xx_rsc_17_0_i_wea_d,
      xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_18_0_i_adra_d => hybrid_core_inst_xx_rsc_18_0_i_adra_d,
      xx_rsc_18_0_i_clka_en_d => xx_rsc_18_0_i_clka_en_d,
      xx_rsc_18_0_i_qa_d => hybrid_core_inst_xx_rsc_18_0_i_qa_d,
      xx_rsc_18_0_i_wea_d => hybrid_core_inst_xx_rsc_18_0_i_wea_d,
      xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_19_0_i_adra_d => hybrid_core_inst_xx_rsc_19_0_i_adra_d,
      xx_rsc_19_0_i_clka_en_d => xx_rsc_19_0_i_clka_en_d,
      xx_rsc_19_0_i_qa_d => hybrid_core_inst_xx_rsc_19_0_i_qa_d,
      xx_rsc_19_0_i_wea_d => hybrid_core_inst_xx_rsc_19_0_i_wea_d,
      xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_20_0_i_adra_d => hybrid_core_inst_xx_rsc_20_0_i_adra_d,
      xx_rsc_20_0_i_clka_en_d => xx_rsc_20_0_i_clka_en_d,
      xx_rsc_20_0_i_qa_d => hybrid_core_inst_xx_rsc_20_0_i_qa_d,
      xx_rsc_20_0_i_wea_d => hybrid_core_inst_xx_rsc_20_0_i_wea_d,
      xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_21_0_i_adra_d => hybrid_core_inst_xx_rsc_21_0_i_adra_d,
      xx_rsc_21_0_i_clka_en_d => xx_rsc_21_0_i_clka_en_d,
      xx_rsc_21_0_i_qa_d => hybrid_core_inst_xx_rsc_21_0_i_qa_d,
      xx_rsc_21_0_i_wea_d => hybrid_core_inst_xx_rsc_21_0_i_wea_d,
      xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_22_0_i_adra_d => hybrid_core_inst_xx_rsc_22_0_i_adra_d,
      xx_rsc_22_0_i_clka_en_d => xx_rsc_22_0_i_clka_en_d,
      xx_rsc_22_0_i_qa_d => hybrid_core_inst_xx_rsc_22_0_i_qa_d,
      xx_rsc_22_0_i_wea_d => hybrid_core_inst_xx_rsc_22_0_i_wea_d,
      xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_23_0_i_adra_d => hybrid_core_inst_xx_rsc_23_0_i_adra_d,
      xx_rsc_23_0_i_clka_en_d => xx_rsc_23_0_i_clka_en_d,
      xx_rsc_23_0_i_qa_d => hybrid_core_inst_xx_rsc_23_0_i_qa_d,
      xx_rsc_23_0_i_wea_d => hybrid_core_inst_xx_rsc_23_0_i_wea_d,
      xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_24_0_i_adra_d => hybrid_core_inst_xx_rsc_24_0_i_adra_d,
      xx_rsc_24_0_i_clka_en_d => xx_rsc_24_0_i_clka_en_d,
      xx_rsc_24_0_i_qa_d => hybrid_core_inst_xx_rsc_24_0_i_qa_d,
      xx_rsc_24_0_i_wea_d => hybrid_core_inst_xx_rsc_24_0_i_wea_d,
      xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_25_0_i_adra_d => hybrid_core_inst_xx_rsc_25_0_i_adra_d,
      xx_rsc_25_0_i_clka_en_d => xx_rsc_25_0_i_clka_en_d,
      xx_rsc_25_0_i_qa_d => hybrid_core_inst_xx_rsc_25_0_i_qa_d,
      xx_rsc_25_0_i_wea_d => hybrid_core_inst_xx_rsc_25_0_i_wea_d,
      xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_26_0_i_adra_d => hybrid_core_inst_xx_rsc_26_0_i_adra_d,
      xx_rsc_26_0_i_clka_en_d => xx_rsc_26_0_i_clka_en_d,
      xx_rsc_26_0_i_qa_d => hybrid_core_inst_xx_rsc_26_0_i_qa_d,
      xx_rsc_26_0_i_wea_d => hybrid_core_inst_xx_rsc_26_0_i_wea_d,
      xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_27_0_i_adra_d => hybrid_core_inst_xx_rsc_27_0_i_adra_d,
      xx_rsc_27_0_i_clka_en_d => xx_rsc_27_0_i_clka_en_d,
      xx_rsc_27_0_i_qa_d => hybrid_core_inst_xx_rsc_27_0_i_qa_d,
      xx_rsc_27_0_i_wea_d => hybrid_core_inst_xx_rsc_27_0_i_wea_d,
      xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_28_0_i_adra_d => hybrid_core_inst_xx_rsc_28_0_i_adra_d,
      xx_rsc_28_0_i_clka_en_d => xx_rsc_28_0_i_clka_en_d,
      xx_rsc_28_0_i_qa_d => hybrid_core_inst_xx_rsc_28_0_i_qa_d,
      xx_rsc_28_0_i_wea_d => hybrid_core_inst_xx_rsc_28_0_i_wea_d,
      xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_29_0_i_adra_d => hybrid_core_inst_xx_rsc_29_0_i_adra_d,
      xx_rsc_29_0_i_clka_en_d => xx_rsc_29_0_i_clka_en_d,
      xx_rsc_29_0_i_qa_d => hybrid_core_inst_xx_rsc_29_0_i_qa_d,
      xx_rsc_29_0_i_wea_d => hybrid_core_inst_xx_rsc_29_0_i_wea_d,
      xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_30_0_i_adra_d => hybrid_core_inst_xx_rsc_30_0_i_adra_d,
      xx_rsc_30_0_i_clka_en_d => xx_rsc_30_0_i_clka_en_d,
      xx_rsc_30_0_i_qa_d => hybrid_core_inst_xx_rsc_30_0_i_qa_d,
      xx_rsc_30_0_i_wea_d => hybrid_core_inst_xx_rsc_30_0_i_wea_d,
      xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      xx_rsc_31_0_i_adra_d => hybrid_core_inst_xx_rsc_31_0_i_adra_d,
      xx_rsc_31_0_i_clka_en_d => xx_rsc_31_0_i_clka_en_d,
      xx_rsc_31_0_i_qa_d => hybrid_core_inst_xx_rsc_31_0_i_qa_d,
      xx_rsc_31_0_i_wea_d => hybrid_core_inst_xx_rsc_31_0_i_wea_d,
      xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_0_0_i_adra_d => hybrid_core_inst_yy_rsc_0_0_i_adra_d,
      yy_rsc_0_0_i_clka_en_d => yy_rsc_0_0_i_clka_en_d,
      yy_rsc_0_0_i_qa_d => hybrid_core_inst_yy_rsc_0_0_i_qa_d,
      yy_rsc_0_0_i_wea_d => hybrid_core_inst_yy_rsc_0_0_i_wea_d,
      yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_1_0_i_adra_d => hybrid_core_inst_yy_rsc_1_0_i_adra_d,
      yy_rsc_1_0_i_clka_en_d => yy_rsc_1_0_i_clka_en_d,
      yy_rsc_1_0_i_qa_d => hybrid_core_inst_yy_rsc_1_0_i_qa_d,
      yy_rsc_1_0_i_wea_d => hybrid_core_inst_yy_rsc_1_0_i_wea_d,
      yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_2_0_i_adra_d => hybrid_core_inst_yy_rsc_2_0_i_adra_d,
      yy_rsc_2_0_i_clka_en_d => yy_rsc_2_0_i_clka_en_d,
      yy_rsc_2_0_i_qa_d => hybrid_core_inst_yy_rsc_2_0_i_qa_d,
      yy_rsc_2_0_i_wea_d => hybrid_core_inst_yy_rsc_2_0_i_wea_d,
      yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_3_0_i_adra_d => hybrid_core_inst_yy_rsc_3_0_i_adra_d,
      yy_rsc_3_0_i_clka_en_d => yy_rsc_3_0_i_clka_en_d,
      yy_rsc_3_0_i_qa_d => hybrid_core_inst_yy_rsc_3_0_i_qa_d,
      yy_rsc_3_0_i_wea_d => hybrid_core_inst_yy_rsc_3_0_i_wea_d,
      yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_4_0_i_adra_d => hybrid_core_inst_yy_rsc_4_0_i_adra_d,
      yy_rsc_4_0_i_clka_en_d => yy_rsc_4_0_i_clka_en_d,
      yy_rsc_4_0_i_qa_d => hybrid_core_inst_yy_rsc_4_0_i_qa_d,
      yy_rsc_4_0_i_wea_d => hybrid_core_inst_yy_rsc_4_0_i_wea_d,
      yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_5_0_i_adra_d => hybrid_core_inst_yy_rsc_5_0_i_adra_d,
      yy_rsc_5_0_i_clka_en_d => yy_rsc_5_0_i_clka_en_d,
      yy_rsc_5_0_i_qa_d => hybrid_core_inst_yy_rsc_5_0_i_qa_d,
      yy_rsc_5_0_i_wea_d => hybrid_core_inst_yy_rsc_5_0_i_wea_d,
      yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_6_0_i_adra_d => hybrid_core_inst_yy_rsc_6_0_i_adra_d,
      yy_rsc_6_0_i_clka_en_d => yy_rsc_6_0_i_clka_en_d,
      yy_rsc_6_0_i_qa_d => hybrid_core_inst_yy_rsc_6_0_i_qa_d,
      yy_rsc_6_0_i_wea_d => hybrid_core_inst_yy_rsc_6_0_i_wea_d,
      yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_7_0_i_adra_d => hybrid_core_inst_yy_rsc_7_0_i_adra_d,
      yy_rsc_7_0_i_clka_en_d => yy_rsc_7_0_i_clka_en_d,
      yy_rsc_7_0_i_qa_d => hybrid_core_inst_yy_rsc_7_0_i_qa_d,
      yy_rsc_7_0_i_wea_d => hybrid_core_inst_yy_rsc_7_0_i_wea_d,
      yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_8_0_i_adra_d => hybrid_core_inst_yy_rsc_8_0_i_adra_d,
      yy_rsc_8_0_i_clka_en_d => yy_rsc_8_0_i_clka_en_d,
      yy_rsc_8_0_i_qa_d => hybrid_core_inst_yy_rsc_8_0_i_qa_d,
      yy_rsc_8_0_i_wea_d => hybrid_core_inst_yy_rsc_8_0_i_wea_d,
      yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_9_0_i_adra_d => hybrid_core_inst_yy_rsc_9_0_i_adra_d,
      yy_rsc_9_0_i_clka_en_d => yy_rsc_9_0_i_clka_en_d,
      yy_rsc_9_0_i_qa_d => hybrid_core_inst_yy_rsc_9_0_i_qa_d,
      yy_rsc_9_0_i_wea_d => hybrid_core_inst_yy_rsc_9_0_i_wea_d,
      yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_10_0_i_adra_d => hybrid_core_inst_yy_rsc_10_0_i_adra_d,
      yy_rsc_10_0_i_clka_en_d => yy_rsc_10_0_i_clka_en_d,
      yy_rsc_10_0_i_qa_d => hybrid_core_inst_yy_rsc_10_0_i_qa_d,
      yy_rsc_10_0_i_wea_d => hybrid_core_inst_yy_rsc_10_0_i_wea_d,
      yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_11_0_i_adra_d => hybrid_core_inst_yy_rsc_11_0_i_adra_d,
      yy_rsc_11_0_i_clka_en_d => yy_rsc_11_0_i_clka_en_d,
      yy_rsc_11_0_i_qa_d => hybrid_core_inst_yy_rsc_11_0_i_qa_d,
      yy_rsc_11_0_i_wea_d => hybrid_core_inst_yy_rsc_11_0_i_wea_d,
      yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_12_0_i_adra_d => hybrid_core_inst_yy_rsc_12_0_i_adra_d,
      yy_rsc_12_0_i_clka_en_d => yy_rsc_12_0_i_clka_en_d,
      yy_rsc_12_0_i_qa_d => hybrid_core_inst_yy_rsc_12_0_i_qa_d,
      yy_rsc_12_0_i_wea_d => hybrid_core_inst_yy_rsc_12_0_i_wea_d,
      yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_13_0_i_adra_d => hybrid_core_inst_yy_rsc_13_0_i_adra_d,
      yy_rsc_13_0_i_clka_en_d => yy_rsc_13_0_i_clka_en_d,
      yy_rsc_13_0_i_qa_d => hybrid_core_inst_yy_rsc_13_0_i_qa_d,
      yy_rsc_13_0_i_wea_d => hybrid_core_inst_yy_rsc_13_0_i_wea_d,
      yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_14_0_i_adra_d => hybrid_core_inst_yy_rsc_14_0_i_adra_d,
      yy_rsc_14_0_i_clka_en_d => yy_rsc_14_0_i_clka_en_d,
      yy_rsc_14_0_i_qa_d => hybrid_core_inst_yy_rsc_14_0_i_qa_d,
      yy_rsc_14_0_i_wea_d => hybrid_core_inst_yy_rsc_14_0_i_wea_d,
      yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_15_0_i_adra_d => hybrid_core_inst_yy_rsc_15_0_i_adra_d,
      yy_rsc_15_0_i_clka_en_d => yy_rsc_15_0_i_clka_en_d,
      yy_rsc_15_0_i_qa_d => hybrid_core_inst_yy_rsc_15_0_i_qa_d,
      yy_rsc_15_0_i_wea_d => hybrid_core_inst_yy_rsc_15_0_i_wea_d,
      yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_16_0_i_adra_d => hybrid_core_inst_yy_rsc_16_0_i_adra_d,
      yy_rsc_16_0_i_clka_en_d => yy_rsc_16_0_i_clka_en_d,
      yy_rsc_16_0_i_qa_d => hybrid_core_inst_yy_rsc_16_0_i_qa_d,
      yy_rsc_16_0_i_wea_d => hybrid_core_inst_yy_rsc_16_0_i_wea_d,
      yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_17_0_i_adra_d => hybrid_core_inst_yy_rsc_17_0_i_adra_d,
      yy_rsc_17_0_i_clka_en_d => yy_rsc_17_0_i_clka_en_d,
      yy_rsc_17_0_i_qa_d => hybrid_core_inst_yy_rsc_17_0_i_qa_d,
      yy_rsc_17_0_i_wea_d => hybrid_core_inst_yy_rsc_17_0_i_wea_d,
      yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_18_0_i_adra_d => hybrid_core_inst_yy_rsc_18_0_i_adra_d,
      yy_rsc_18_0_i_clka_en_d => yy_rsc_18_0_i_clka_en_d,
      yy_rsc_18_0_i_qa_d => hybrid_core_inst_yy_rsc_18_0_i_qa_d,
      yy_rsc_18_0_i_wea_d => hybrid_core_inst_yy_rsc_18_0_i_wea_d,
      yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_19_0_i_adra_d => hybrid_core_inst_yy_rsc_19_0_i_adra_d,
      yy_rsc_19_0_i_clka_en_d => yy_rsc_19_0_i_clka_en_d,
      yy_rsc_19_0_i_qa_d => hybrid_core_inst_yy_rsc_19_0_i_qa_d,
      yy_rsc_19_0_i_wea_d => hybrid_core_inst_yy_rsc_19_0_i_wea_d,
      yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_20_0_i_adra_d => hybrid_core_inst_yy_rsc_20_0_i_adra_d,
      yy_rsc_20_0_i_clka_en_d => yy_rsc_20_0_i_clka_en_d,
      yy_rsc_20_0_i_qa_d => hybrid_core_inst_yy_rsc_20_0_i_qa_d,
      yy_rsc_20_0_i_wea_d => hybrid_core_inst_yy_rsc_20_0_i_wea_d,
      yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_21_0_i_adra_d => hybrid_core_inst_yy_rsc_21_0_i_adra_d,
      yy_rsc_21_0_i_clka_en_d => yy_rsc_21_0_i_clka_en_d,
      yy_rsc_21_0_i_qa_d => hybrid_core_inst_yy_rsc_21_0_i_qa_d,
      yy_rsc_21_0_i_wea_d => hybrid_core_inst_yy_rsc_21_0_i_wea_d,
      yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_22_0_i_adra_d => hybrid_core_inst_yy_rsc_22_0_i_adra_d,
      yy_rsc_22_0_i_clka_en_d => yy_rsc_22_0_i_clka_en_d,
      yy_rsc_22_0_i_qa_d => hybrid_core_inst_yy_rsc_22_0_i_qa_d,
      yy_rsc_22_0_i_wea_d => hybrid_core_inst_yy_rsc_22_0_i_wea_d,
      yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_23_0_i_adra_d => hybrid_core_inst_yy_rsc_23_0_i_adra_d,
      yy_rsc_23_0_i_clka_en_d => yy_rsc_23_0_i_clka_en_d,
      yy_rsc_23_0_i_qa_d => hybrid_core_inst_yy_rsc_23_0_i_qa_d,
      yy_rsc_23_0_i_wea_d => hybrid_core_inst_yy_rsc_23_0_i_wea_d,
      yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_24_0_i_adra_d => hybrid_core_inst_yy_rsc_24_0_i_adra_d,
      yy_rsc_24_0_i_clka_en_d => yy_rsc_24_0_i_clka_en_d,
      yy_rsc_24_0_i_qa_d => hybrid_core_inst_yy_rsc_24_0_i_qa_d,
      yy_rsc_24_0_i_wea_d => hybrid_core_inst_yy_rsc_24_0_i_wea_d,
      yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_25_0_i_adra_d => hybrid_core_inst_yy_rsc_25_0_i_adra_d,
      yy_rsc_25_0_i_clka_en_d => yy_rsc_25_0_i_clka_en_d,
      yy_rsc_25_0_i_qa_d => hybrid_core_inst_yy_rsc_25_0_i_qa_d,
      yy_rsc_25_0_i_wea_d => hybrid_core_inst_yy_rsc_25_0_i_wea_d,
      yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_26_0_i_adra_d => hybrid_core_inst_yy_rsc_26_0_i_adra_d,
      yy_rsc_26_0_i_clka_en_d => yy_rsc_26_0_i_clka_en_d,
      yy_rsc_26_0_i_qa_d => hybrid_core_inst_yy_rsc_26_0_i_qa_d,
      yy_rsc_26_0_i_wea_d => hybrid_core_inst_yy_rsc_26_0_i_wea_d,
      yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_27_0_i_adra_d => hybrid_core_inst_yy_rsc_27_0_i_adra_d,
      yy_rsc_27_0_i_clka_en_d => yy_rsc_27_0_i_clka_en_d,
      yy_rsc_27_0_i_qa_d => hybrid_core_inst_yy_rsc_27_0_i_qa_d,
      yy_rsc_27_0_i_wea_d => hybrid_core_inst_yy_rsc_27_0_i_wea_d,
      yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_28_0_i_adra_d => hybrid_core_inst_yy_rsc_28_0_i_adra_d,
      yy_rsc_28_0_i_clka_en_d => yy_rsc_28_0_i_clka_en_d,
      yy_rsc_28_0_i_qa_d => hybrid_core_inst_yy_rsc_28_0_i_qa_d,
      yy_rsc_28_0_i_wea_d => hybrid_core_inst_yy_rsc_28_0_i_wea_d,
      yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_29_0_i_adra_d => hybrid_core_inst_yy_rsc_29_0_i_adra_d,
      yy_rsc_29_0_i_clka_en_d => yy_rsc_29_0_i_clka_en_d,
      yy_rsc_29_0_i_qa_d => hybrid_core_inst_yy_rsc_29_0_i_qa_d,
      yy_rsc_29_0_i_wea_d => hybrid_core_inst_yy_rsc_29_0_i_wea_d,
      yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_30_0_i_adra_d => hybrid_core_inst_yy_rsc_30_0_i_adra_d,
      yy_rsc_30_0_i_clka_en_d => yy_rsc_30_0_i_clka_en_d,
      yy_rsc_30_0_i_qa_d => hybrid_core_inst_yy_rsc_30_0_i_qa_d,
      yy_rsc_30_0_i_wea_d => hybrid_core_inst_yy_rsc_30_0_i_wea_d,
      yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      yy_rsc_31_0_i_adra_d => hybrid_core_inst_yy_rsc_31_0_i_adra_d,
      yy_rsc_31_0_i_clka_en_d => yy_rsc_31_0_i_clka_en_d,
      yy_rsc_31_0_i_qa_d => hybrid_core_inst_yy_rsc_31_0_i_qa_d,
      yy_rsc_31_0_i_wea_d => hybrid_core_inst_yy_rsc_31_0_i_wea_d,
      yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => hybrid_core_inst_yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d => hybrid_core_inst_yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d,
      S34_OUTER_LOOP_for_tf_mul_cmp_a => hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_a,
      S34_OUTER_LOOP_for_tf_mul_cmp_b => hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_b,
      S34_OUTER_LOOP_for_tf_mul_cmp_z => hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z,
      xx_rsc_0_0_i_da_d_pff => hybrid_core_inst_xx_rsc_0_0_i_da_d_pff,
      xx_rsc_1_0_i_da_d_pff => hybrid_core_inst_xx_rsc_1_0_i_da_d_pff,
      xx_rsc_2_0_i_da_d_pff => hybrid_core_inst_xx_rsc_2_0_i_da_d_pff,
      xx_rsc_3_0_i_da_d_pff => hybrid_core_inst_xx_rsc_3_0_i_da_d_pff,
      yy_rsc_0_0_i_da_d_pff => hybrid_core_inst_yy_rsc_0_0_i_da_d_pff,
      yy_rsc_1_0_i_da_d_pff => hybrid_core_inst_yy_rsc_1_0_i_da_d_pff,
      yy_rsc_2_0_i_da_d_pff => hybrid_core_inst_yy_rsc_2_0_i_da_d_pff,
      yy_rsc_3_0_i_da_d_pff => hybrid_core_inst_yy_rsc_3_0_i_da_d_pff
    );
  x_rsc_0_0_RRESP <= hybrid_core_inst_x_rsc_0_0_RRESP;
  x_rsc_0_0_RDATA <= hybrid_core_inst_x_rsc_0_0_RDATA;
  hybrid_core_inst_x_rsc_0_0_ARREGION <= x_rsc_0_0_ARREGION;
  hybrid_core_inst_x_rsc_0_0_ARQOS <= x_rsc_0_0_ARQOS;
  hybrid_core_inst_x_rsc_0_0_ARPROT <= x_rsc_0_0_ARPROT;
  hybrid_core_inst_x_rsc_0_0_ARCACHE <= x_rsc_0_0_ARCACHE;
  hybrid_core_inst_x_rsc_0_0_ARBURST <= x_rsc_0_0_ARBURST;
  hybrid_core_inst_x_rsc_0_0_ARSIZE <= x_rsc_0_0_ARSIZE;
  hybrid_core_inst_x_rsc_0_0_ARLEN <= x_rsc_0_0_ARLEN;
  hybrid_core_inst_x_rsc_0_0_ARADDR <= x_rsc_0_0_ARADDR;
  x_rsc_0_0_BRESP <= hybrid_core_inst_x_rsc_0_0_BRESP;
  hybrid_core_inst_x_rsc_0_0_WSTRB <= x_rsc_0_0_WSTRB;
  hybrid_core_inst_x_rsc_0_0_WDATA <= x_rsc_0_0_WDATA;
  hybrid_core_inst_x_rsc_0_0_AWREGION <= x_rsc_0_0_AWREGION;
  hybrid_core_inst_x_rsc_0_0_AWQOS <= x_rsc_0_0_AWQOS;
  hybrid_core_inst_x_rsc_0_0_AWPROT <= x_rsc_0_0_AWPROT;
  hybrid_core_inst_x_rsc_0_0_AWCACHE <= x_rsc_0_0_AWCACHE;
  hybrid_core_inst_x_rsc_0_0_AWBURST <= x_rsc_0_0_AWBURST;
  hybrid_core_inst_x_rsc_0_0_AWSIZE <= x_rsc_0_0_AWSIZE;
  hybrid_core_inst_x_rsc_0_0_AWLEN <= x_rsc_0_0_AWLEN;
  hybrid_core_inst_x_rsc_0_0_AWADDR <= x_rsc_0_0_AWADDR;
  x_rsc_1_0_RRESP <= hybrid_core_inst_x_rsc_1_0_RRESP;
  x_rsc_1_0_RDATA <= hybrid_core_inst_x_rsc_1_0_RDATA;
  hybrid_core_inst_x_rsc_1_0_ARREGION <= x_rsc_1_0_ARREGION;
  hybrid_core_inst_x_rsc_1_0_ARQOS <= x_rsc_1_0_ARQOS;
  hybrid_core_inst_x_rsc_1_0_ARPROT <= x_rsc_1_0_ARPROT;
  hybrid_core_inst_x_rsc_1_0_ARCACHE <= x_rsc_1_0_ARCACHE;
  hybrid_core_inst_x_rsc_1_0_ARBURST <= x_rsc_1_0_ARBURST;
  hybrid_core_inst_x_rsc_1_0_ARSIZE <= x_rsc_1_0_ARSIZE;
  hybrid_core_inst_x_rsc_1_0_ARLEN <= x_rsc_1_0_ARLEN;
  hybrid_core_inst_x_rsc_1_0_ARADDR <= x_rsc_1_0_ARADDR;
  x_rsc_1_0_BRESP <= hybrid_core_inst_x_rsc_1_0_BRESP;
  hybrid_core_inst_x_rsc_1_0_WSTRB <= x_rsc_1_0_WSTRB;
  hybrid_core_inst_x_rsc_1_0_WDATA <= x_rsc_1_0_WDATA;
  hybrid_core_inst_x_rsc_1_0_AWREGION <= x_rsc_1_0_AWREGION;
  hybrid_core_inst_x_rsc_1_0_AWQOS <= x_rsc_1_0_AWQOS;
  hybrid_core_inst_x_rsc_1_0_AWPROT <= x_rsc_1_0_AWPROT;
  hybrid_core_inst_x_rsc_1_0_AWCACHE <= x_rsc_1_0_AWCACHE;
  hybrid_core_inst_x_rsc_1_0_AWBURST <= x_rsc_1_0_AWBURST;
  hybrid_core_inst_x_rsc_1_0_AWSIZE <= x_rsc_1_0_AWSIZE;
  hybrid_core_inst_x_rsc_1_0_AWLEN <= x_rsc_1_0_AWLEN;
  hybrid_core_inst_x_rsc_1_0_AWADDR <= x_rsc_1_0_AWADDR;
  x_rsc_2_0_RRESP <= hybrid_core_inst_x_rsc_2_0_RRESP;
  x_rsc_2_0_RDATA <= hybrid_core_inst_x_rsc_2_0_RDATA;
  hybrid_core_inst_x_rsc_2_0_ARREGION <= x_rsc_2_0_ARREGION;
  hybrid_core_inst_x_rsc_2_0_ARQOS <= x_rsc_2_0_ARQOS;
  hybrid_core_inst_x_rsc_2_0_ARPROT <= x_rsc_2_0_ARPROT;
  hybrid_core_inst_x_rsc_2_0_ARCACHE <= x_rsc_2_0_ARCACHE;
  hybrid_core_inst_x_rsc_2_0_ARBURST <= x_rsc_2_0_ARBURST;
  hybrid_core_inst_x_rsc_2_0_ARSIZE <= x_rsc_2_0_ARSIZE;
  hybrid_core_inst_x_rsc_2_0_ARLEN <= x_rsc_2_0_ARLEN;
  hybrid_core_inst_x_rsc_2_0_ARADDR <= x_rsc_2_0_ARADDR;
  x_rsc_2_0_BRESP <= hybrid_core_inst_x_rsc_2_0_BRESP;
  hybrid_core_inst_x_rsc_2_0_WSTRB <= x_rsc_2_0_WSTRB;
  hybrid_core_inst_x_rsc_2_0_WDATA <= x_rsc_2_0_WDATA;
  hybrid_core_inst_x_rsc_2_0_AWREGION <= x_rsc_2_0_AWREGION;
  hybrid_core_inst_x_rsc_2_0_AWQOS <= x_rsc_2_0_AWQOS;
  hybrid_core_inst_x_rsc_2_0_AWPROT <= x_rsc_2_0_AWPROT;
  hybrid_core_inst_x_rsc_2_0_AWCACHE <= x_rsc_2_0_AWCACHE;
  hybrid_core_inst_x_rsc_2_0_AWBURST <= x_rsc_2_0_AWBURST;
  hybrid_core_inst_x_rsc_2_0_AWSIZE <= x_rsc_2_0_AWSIZE;
  hybrid_core_inst_x_rsc_2_0_AWLEN <= x_rsc_2_0_AWLEN;
  hybrid_core_inst_x_rsc_2_0_AWADDR <= x_rsc_2_0_AWADDR;
  x_rsc_3_0_RRESP <= hybrid_core_inst_x_rsc_3_0_RRESP;
  x_rsc_3_0_RDATA <= hybrid_core_inst_x_rsc_3_0_RDATA;
  hybrid_core_inst_x_rsc_3_0_ARREGION <= x_rsc_3_0_ARREGION;
  hybrid_core_inst_x_rsc_3_0_ARQOS <= x_rsc_3_0_ARQOS;
  hybrid_core_inst_x_rsc_3_0_ARPROT <= x_rsc_3_0_ARPROT;
  hybrid_core_inst_x_rsc_3_0_ARCACHE <= x_rsc_3_0_ARCACHE;
  hybrid_core_inst_x_rsc_3_0_ARBURST <= x_rsc_3_0_ARBURST;
  hybrid_core_inst_x_rsc_3_0_ARSIZE <= x_rsc_3_0_ARSIZE;
  hybrid_core_inst_x_rsc_3_0_ARLEN <= x_rsc_3_0_ARLEN;
  hybrid_core_inst_x_rsc_3_0_ARADDR <= x_rsc_3_0_ARADDR;
  x_rsc_3_0_BRESP <= hybrid_core_inst_x_rsc_3_0_BRESP;
  hybrid_core_inst_x_rsc_3_0_WSTRB <= x_rsc_3_0_WSTRB;
  hybrid_core_inst_x_rsc_3_0_WDATA <= x_rsc_3_0_WDATA;
  hybrid_core_inst_x_rsc_3_0_AWREGION <= x_rsc_3_0_AWREGION;
  hybrid_core_inst_x_rsc_3_0_AWQOS <= x_rsc_3_0_AWQOS;
  hybrid_core_inst_x_rsc_3_0_AWPROT <= x_rsc_3_0_AWPROT;
  hybrid_core_inst_x_rsc_3_0_AWCACHE <= x_rsc_3_0_AWCACHE;
  hybrid_core_inst_x_rsc_3_0_AWBURST <= x_rsc_3_0_AWBURST;
  hybrid_core_inst_x_rsc_3_0_AWSIZE <= x_rsc_3_0_AWSIZE;
  hybrid_core_inst_x_rsc_3_0_AWLEN <= x_rsc_3_0_AWLEN;
  hybrid_core_inst_x_rsc_3_0_AWADDR <= x_rsc_3_0_AWADDR;
  x_rsc_4_0_RRESP <= hybrid_core_inst_x_rsc_4_0_RRESP;
  x_rsc_4_0_RDATA <= hybrid_core_inst_x_rsc_4_0_RDATA;
  hybrid_core_inst_x_rsc_4_0_ARREGION <= x_rsc_4_0_ARREGION;
  hybrid_core_inst_x_rsc_4_0_ARQOS <= x_rsc_4_0_ARQOS;
  hybrid_core_inst_x_rsc_4_0_ARPROT <= x_rsc_4_0_ARPROT;
  hybrid_core_inst_x_rsc_4_0_ARCACHE <= x_rsc_4_0_ARCACHE;
  hybrid_core_inst_x_rsc_4_0_ARBURST <= x_rsc_4_0_ARBURST;
  hybrid_core_inst_x_rsc_4_0_ARSIZE <= x_rsc_4_0_ARSIZE;
  hybrid_core_inst_x_rsc_4_0_ARLEN <= x_rsc_4_0_ARLEN;
  hybrid_core_inst_x_rsc_4_0_ARADDR <= x_rsc_4_0_ARADDR;
  x_rsc_4_0_BRESP <= hybrid_core_inst_x_rsc_4_0_BRESP;
  hybrid_core_inst_x_rsc_4_0_WSTRB <= x_rsc_4_0_WSTRB;
  hybrid_core_inst_x_rsc_4_0_WDATA <= x_rsc_4_0_WDATA;
  hybrid_core_inst_x_rsc_4_0_AWREGION <= x_rsc_4_0_AWREGION;
  hybrid_core_inst_x_rsc_4_0_AWQOS <= x_rsc_4_0_AWQOS;
  hybrid_core_inst_x_rsc_4_0_AWPROT <= x_rsc_4_0_AWPROT;
  hybrid_core_inst_x_rsc_4_0_AWCACHE <= x_rsc_4_0_AWCACHE;
  hybrid_core_inst_x_rsc_4_0_AWBURST <= x_rsc_4_0_AWBURST;
  hybrid_core_inst_x_rsc_4_0_AWSIZE <= x_rsc_4_0_AWSIZE;
  hybrid_core_inst_x_rsc_4_0_AWLEN <= x_rsc_4_0_AWLEN;
  hybrid_core_inst_x_rsc_4_0_AWADDR <= x_rsc_4_0_AWADDR;
  x_rsc_5_0_RRESP <= hybrid_core_inst_x_rsc_5_0_RRESP;
  x_rsc_5_0_RDATA <= hybrid_core_inst_x_rsc_5_0_RDATA;
  hybrid_core_inst_x_rsc_5_0_ARREGION <= x_rsc_5_0_ARREGION;
  hybrid_core_inst_x_rsc_5_0_ARQOS <= x_rsc_5_0_ARQOS;
  hybrid_core_inst_x_rsc_5_0_ARPROT <= x_rsc_5_0_ARPROT;
  hybrid_core_inst_x_rsc_5_0_ARCACHE <= x_rsc_5_0_ARCACHE;
  hybrid_core_inst_x_rsc_5_0_ARBURST <= x_rsc_5_0_ARBURST;
  hybrid_core_inst_x_rsc_5_0_ARSIZE <= x_rsc_5_0_ARSIZE;
  hybrid_core_inst_x_rsc_5_0_ARLEN <= x_rsc_5_0_ARLEN;
  hybrid_core_inst_x_rsc_5_0_ARADDR <= x_rsc_5_0_ARADDR;
  x_rsc_5_0_BRESP <= hybrid_core_inst_x_rsc_5_0_BRESP;
  hybrid_core_inst_x_rsc_5_0_WSTRB <= x_rsc_5_0_WSTRB;
  hybrid_core_inst_x_rsc_5_0_WDATA <= x_rsc_5_0_WDATA;
  hybrid_core_inst_x_rsc_5_0_AWREGION <= x_rsc_5_0_AWREGION;
  hybrid_core_inst_x_rsc_5_0_AWQOS <= x_rsc_5_0_AWQOS;
  hybrid_core_inst_x_rsc_5_0_AWPROT <= x_rsc_5_0_AWPROT;
  hybrid_core_inst_x_rsc_5_0_AWCACHE <= x_rsc_5_0_AWCACHE;
  hybrid_core_inst_x_rsc_5_0_AWBURST <= x_rsc_5_0_AWBURST;
  hybrid_core_inst_x_rsc_5_0_AWSIZE <= x_rsc_5_0_AWSIZE;
  hybrid_core_inst_x_rsc_5_0_AWLEN <= x_rsc_5_0_AWLEN;
  hybrid_core_inst_x_rsc_5_0_AWADDR <= x_rsc_5_0_AWADDR;
  x_rsc_6_0_RRESP <= hybrid_core_inst_x_rsc_6_0_RRESP;
  x_rsc_6_0_RDATA <= hybrid_core_inst_x_rsc_6_0_RDATA;
  hybrid_core_inst_x_rsc_6_0_ARREGION <= x_rsc_6_0_ARREGION;
  hybrid_core_inst_x_rsc_6_0_ARQOS <= x_rsc_6_0_ARQOS;
  hybrid_core_inst_x_rsc_6_0_ARPROT <= x_rsc_6_0_ARPROT;
  hybrid_core_inst_x_rsc_6_0_ARCACHE <= x_rsc_6_0_ARCACHE;
  hybrid_core_inst_x_rsc_6_0_ARBURST <= x_rsc_6_0_ARBURST;
  hybrid_core_inst_x_rsc_6_0_ARSIZE <= x_rsc_6_0_ARSIZE;
  hybrid_core_inst_x_rsc_6_0_ARLEN <= x_rsc_6_0_ARLEN;
  hybrid_core_inst_x_rsc_6_0_ARADDR <= x_rsc_6_0_ARADDR;
  x_rsc_6_0_BRESP <= hybrid_core_inst_x_rsc_6_0_BRESP;
  hybrid_core_inst_x_rsc_6_0_WSTRB <= x_rsc_6_0_WSTRB;
  hybrid_core_inst_x_rsc_6_0_WDATA <= x_rsc_6_0_WDATA;
  hybrid_core_inst_x_rsc_6_0_AWREGION <= x_rsc_6_0_AWREGION;
  hybrid_core_inst_x_rsc_6_0_AWQOS <= x_rsc_6_0_AWQOS;
  hybrid_core_inst_x_rsc_6_0_AWPROT <= x_rsc_6_0_AWPROT;
  hybrid_core_inst_x_rsc_6_0_AWCACHE <= x_rsc_6_0_AWCACHE;
  hybrid_core_inst_x_rsc_6_0_AWBURST <= x_rsc_6_0_AWBURST;
  hybrid_core_inst_x_rsc_6_0_AWSIZE <= x_rsc_6_0_AWSIZE;
  hybrid_core_inst_x_rsc_6_0_AWLEN <= x_rsc_6_0_AWLEN;
  hybrid_core_inst_x_rsc_6_0_AWADDR <= x_rsc_6_0_AWADDR;
  x_rsc_7_0_RRESP <= hybrid_core_inst_x_rsc_7_0_RRESP;
  x_rsc_7_0_RDATA <= hybrid_core_inst_x_rsc_7_0_RDATA;
  hybrid_core_inst_x_rsc_7_0_ARREGION <= x_rsc_7_0_ARREGION;
  hybrid_core_inst_x_rsc_7_0_ARQOS <= x_rsc_7_0_ARQOS;
  hybrid_core_inst_x_rsc_7_0_ARPROT <= x_rsc_7_0_ARPROT;
  hybrid_core_inst_x_rsc_7_0_ARCACHE <= x_rsc_7_0_ARCACHE;
  hybrid_core_inst_x_rsc_7_0_ARBURST <= x_rsc_7_0_ARBURST;
  hybrid_core_inst_x_rsc_7_0_ARSIZE <= x_rsc_7_0_ARSIZE;
  hybrid_core_inst_x_rsc_7_0_ARLEN <= x_rsc_7_0_ARLEN;
  hybrid_core_inst_x_rsc_7_0_ARADDR <= x_rsc_7_0_ARADDR;
  x_rsc_7_0_BRESP <= hybrid_core_inst_x_rsc_7_0_BRESP;
  hybrid_core_inst_x_rsc_7_0_WSTRB <= x_rsc_7_0_WSTRB;
  hybrid_core_inst_x_rsc_7_0_WDATA <= x_rsc_7_0_WDATA;
  hybrid_core_inst_x_rsc_7_0_AWREGION <= x_rsc_7_0_AWREGION;
  hybrid_core_inst_x_rsc_7_0_AWQOS <= x_rsc_7_0_AWQOS;
  hybrid_core_inst_x_rsc_7_0_AWPROT <= x_rsc_7_0_AWPROT;
  hybrid_core_inst_x_rsc_7_0_AWCACHE <= x_rsc_7_0_AWCACHE;
  hybrid_core_inst_x_rsc_7_0_AWBURST <= x_rsc_7_0_AWBURST;
  hybrid_core_inst_x_rsc_7_0_AWSIZE <= x_rsc_7_0_AWSIZE;
  hybrid_core_inst_x_rsc_7_0_AWLEN <= x_rsc_7_0_AWLEN;
  hybrid_core_inst_x_rsc_7_0_AWADDR <= x_rsc_7_0_AWADDR;
  x_rsc_8_0_RRESP <= hybrid_core_inst_x_rsc_8_0_RRESP;
  x_rsc_8_0_RDATA <= hybrid_core_inst_x_rsc_8_0_RDATA;
  hybrid_core_inst_x_rsc_8_0_ARREGION <= x_rsc_8_0_ARREGION;
  hybrid_core_inst_x_rsc_8_0_ARQOS <= x_rsc_8_0_ARQOS;
  hybrid_core_inst_x_rsc_8_0_ARPROT <= x_rsc_8_0_ARPROT;
  hybrid_core_inst_x_rsc_8_0_ARCACHE <= x_rsc_8_0_ARCACHE;
  hybrid_core_inst_x_rsc_8_0_ARBURST <= x_rsc_8_0_ARBURST;
  hybrid_core_inst_x_rsc_8_0_ARSIZE <= x_rsc_8_0_ARSIZE;
  hybrid_core_inst_x_rsc_8_0_ARLEN <= x_rsc_8_0_ARLEN;
  hybrid_core_inst_x_rsc_8_0_ARADDR <= x_rsc_8_0_ARADDR;
  x_rsc_8_0_BRESP <= hybrid_core_inst_x_rsc_8_0_BRESP;
  hybrid_core_inst_x_rsc_8_0_WSTRB <= x_rsc_8_0_WSTRB;
  hybrid_core_inst_x_rsc_8_0_WDATA <= x_rsc_8_0_WDATA;
  hybrid_core_inst_x_rsc_8_0_AWREGION <= x_rsc_8_0_AWREGION;
  hybrid_core_inst_x_rsc_8_0_AWQOS <= x_rsc_8_0_AWQOS;
  hybrid_core_inst_x_rsc_8_0_AWPROT <= x_rsc_8_0_AWPROT;
  hybrid_core_inst_x_rsc_8_0_AWCACHE <= x_rsc_8_0_AWCACHE;
  hybrid_core_inst_x_rsc_8_0_AWBURST <= x_rsc_8_0_AWBURST;
  hybrid_core_inst_x_rsc_8_0_AWSIZE <= x_rsc_8_0_AWSIZE;
  hybrid_core_inst_x_rsc_8_0_AWLEN <= x_rsc_8_0_AWLEN;
  hybrid_core_inst_x_rsc_8_0_AWADDR <= x_rsc_8_0_AWADDR;
  x_rsc_9_0_RRESP <= hybrid_core_inst_x_rsc_9_0_RRESP;
  x_rsc_9_0_RDATA <= hybrid_core_inst_x_rsc_9_0_RDATA;
  hybrid_core_inst_x_rsc_9_0_ARREGION <= x_rsc_9_0_ARREGION;
  hybrid_core_inst_x_rsc_9_0_ARQOS <= x_rsc_9_0_ARQOS;
  hybrid_core_inst_x_rsc_9_0_ARPROT <= x_rsc_9_0_ARPROT;
  hybrid_core_inst_x_rsc_9_0_ARCACHE <= x_rsc_9_0_ARCACHE;
  hybrid_core_inst_x_rsc_9_0_ARBURST <= x_rsc_9_0_ARBURST;
  hybrid_core_inst_x_rsc_9_0_ARSIZE <= x_rsc_9_0_ARSIZE;
  hybrid_core_inst_x_rsc_9_0_ARLEN <= x_rsc_9_0_ARLEN;
  hybrid_core_inst_x_rsc_9_0_ARADDR <= x_rsc_9_0_ARADDR;
  x_rsc_9_0_BRESP <= hybrid_core_inst_x_rsc_9_0_BRESP;
  hybrid_core_inst_x_rsc_9_0_WSTRB <= x_rsc_9_0_WSTRB;
  hybrid_core_inst_x_rsc_9_0_WDATA <= x_rsc_9_0_WDATA;
  hybrid_core_inst_x_rsc_9_0_AWREGION <= x_rsc_9_0_AWREGION;
  hybrid_core_inst_x_rsc_9_0_AWQOS <= x_rsc_9_0_AWQOS;
  hybrid_core_inst_x_rsc_9_0_AWPROT <= x_rsc_9_0_AWPROT;
  hybrid_core_inst_x_rsc_9_0_AWCACHE <= x_rsc_9_0_AWCACHE;
  hybrid_core_inst_x_rsc_9_0_AWBURST <= x_rsc_9_0_AWBURST;
  hybrid_core_inst_x_rsc_9_0_AWSIZE <= x_rsc_9_0_AWSIZE;
  hybrid_core_inst_x_rsc_9_0_AWLEN <= x_rsc_9_0_AWLEN;
  hybrid_core_inst_x_rsc_9_0_AWADDR <= x_rsc_9_0_AWADDR;
  x_rsc_10_0_RRESP <= hybrid_core_inst_x_rsc_10_0_RRESP;
  x_rsc_10_0_RDATA <= hybrid_core_inst_x_rsc_10_0_RDATA;
  hybrid_core_inst_x_rsc_10_0_ARREGION <= x_rsc_10_0_ARREGION;
  hybrid_core_inst_x_rsc_10_0_ARQOS <= x_rsc_10_0_ARQOS;
  hybrid_core_inst_x_rsc_10_0_ARPROT <= x_rsc_10_0_ARPROT;
  hybrid_core_inst_x_rsc_10_0_ARCACHE <= x_rsc_10_0_ARCACHE;
  hybrid_core_inst_x_rsc_10_0_ARBURST <= x_rsc_10_0_ARBURST;
  hybrid_core_inst_x_rsc_10_0_ARSIZE <= x_rsc_10_0_ARSIZE;
  hybrid_core_inst_x_rsc_10_0_ARLEN <= x_rsc_10_0_ARLEN;
  hybrid_core_inst_x_rsc_10_0_ARADDR <= x_rsc_10_0_ARADDR;
  x_rsc_10_0_BRESP <= hybrid_core_inst_x_rsc_10_0_BRESP;
  hybrid_core_inst_x_rsc_10_0_WSTRB <= x_rsc_10_0_WSTRB;
  hybrid_core_inst_x_rsc_10_0_WDATA <= x_rsc_10_0_WDATA;
  hybrid_core_inst_x_rsc_10_0_AWREGION <= x_rsc_10_0_AWREGION;
  hybrid_core_inst_x_rsc_10_0_AWQOS <= x_rsc_10_0_AWQOS;
  hybrid_core_inst_x_rsc_10_0_AWPROT <= x_rsc_10_0_AWPROT;
  hybrid_core_inst_x_rsc_10_0_AWCACHE <= x_rsc_10_0_AWCACHE;
  hybrid_core_inst_x_rsc_10_0_AWBURST <= x_rsc_10_0_AWBURST;
  hybrid_core_inst_x_rsc_10_0_AWSIZE <= x_rsc_10_0_AWSIZE;
  hybrid_core_inst_x_rsc_10_0_AWLEN <= x_rsc_10_0_AWLEN;
  hybrid_core_inst_x_rsc_10_0_AWADDR <= x_rsc_10_0_AWADDR;
  x_rsc_11_0_RRESP <= hybrid_core_inst_x_rsc_11_0_RRESP;
  x_rsc_11_0_RDATA <= hybrid_core_inst_x_rsc_11_0_RDATA;
  hybrid_core_inst_x_rsc_11_0_ARREGION <= x_rsc_11_0_ARREGION;
  hybrid_core_inst_x_rsc_11_0_ARQOS <= x_rsc_11_0_ARQOS;
  hybrid_core_inst_x_rsc_11_0_ARPROT <= x_rsc_11_0_ARPROT;
  hybrid_core_inst_x_rsc_11_0_ARCACHE <= x_rsc_11_0_ARCACHE;
  hybrid_core_inst_x_rsc_11_0_ARBURST <= x_rsc_11_0_ARBURST;
  hybrid_core_inst_x_rsc_11_0_ARSIZE <= x_rsc_11_0_ARSIZE;
  hybrid_core_inst_x_rsc_11_0_ARLEN <= x_rsc_11_0_ARLEN;
  hybrid_core_inst_x_rsc_11_0_ARADDR <= x_rsc_11_0_ARADDR;
  x_rsc_11_0_BRESP <= hybrid_core_inst_x_rsc_11_0_BRESP;
  hybrid_core_inst_x_rsc_11_0_WSTRB <= x_rsc_11_0_WSTRB;
  hybrid_core_inst_x_rsc_11_0_WDATA <= x_rsc_11_0_WDATA;
  hybrid_core_inst_x_rsc_11_0_AWREGION <= x_rsc_11_0_AWREGION;
  hybrid_core_inst_x_rsc_11_0_AWQOS <= x_rsc_11_0_AWQOS;
  hybrid_core_inst_x_rsc_11_0_AWPROT <= x_rsc_11_0_AWPROT;
  hybrid_core_inst_x_rsc_11_0_AWCACHE <= x_rsc_11_0_AWCACHE;
  hybrid_core_inst_x_rsc_11_0_AWBURST <= x_rsc_11_0_AWBURST;
  hybrid_core_inst_x_rsc_11_0_AWSIZE <= x_rsc_11_0_AWSIZE;
  hybrid_core_inst_x_rsc_11_0_AWLEN <= x_rsc_11_0_AWLEN;
  hybrid_core_inst_x_rsc_11_0_AWADDR <= x_rsc_11_0_AWADDR;
  x_rsc_12_0_RRESP <= hybrid_core_inst_x_rsc_12_0_RRESP;
  x_rsc_12_0_RDATA <= hybrid_core_inst_x_rsc_12_0_RDATA;
  hybrid_core_inst_x_rsc_12_0_ARREGION <= x_rsc_12_0_ARREGION;
  hybrid_core_inst_x_rsc_12_0_ARQOS <= x_rsc_12_0_ARQOS;
  hybrid_core_inst_x_rsc_12_0_ARPROT <= x_rsc_12_0_ARPROT;
  hybrid_core_inst_x_rsc_12_0_ARCACHE <= x_rsc_12_0_ARCACHE;
  hybrid_core_inst_x_rsc_12_0_ARBURST <= x_rsc_12_0_ARBURST;
  hybrid_core_inst_x_rsc_12_0_ARSIZE <= x_rsc_12_0_ARSIZE;
  hybrid_core_inst_x_rsc_12_0_ARLEN <= x_rsc_12_0_ARLEN;
  hybrid_core_inst_x_rsc_12_0_ARADDR <= x_rsc_12_0_ARADDR;
  x_rsc_12_0_BRESP <= hybrid_core_inst_x_rsc_12_0_BRESP;
  hybrid_core_inst_x_rsc_12_0_WSTRB <= x_rsc_12_0_WSTRB;
  hybrid_core_inst_x_rsc_12_0_WDATA <= x_rsc_12_0_WDATA;
  hybrid_core_inst_x_rsc_12_0_AWREGION <= x_rsc_12_0_AWREGION;
  hybrid_core_inst_x_rsc_12_0_AWQOS <= x_rsc_12_0_AWQOS;
  hybrid_core_inst_x_rsc_12_0_AWPROT <= x_rsc_12_0_AWPROT;
  hybrid_core_inst_x_rsc_12_0_AWCACHE <= x_rsc_12_0_AWCACHE;
  hybrid_core_inst_x_rsc_12_0_AWBURST <= x_rsc_12_0_AWBURST;
  hybrid_core_inst_x_rsc_12_0_AWSIZE <= x_rsc_12_0_AWSIZE;
  hybrid_core_inst_x_rsc_12_0_AWLEN <= x_rsc_12_0_AWLEN;
  hybrid_core_inst_x_rsc_12_0_AWADDR <= x_rsc_12_0_AWADDR;
  x_rsc_13_0_RRESP <= hybrid_core_inst_x_rsc_13_0_RRESP;
  x_rsc_13_0_RDATA <= hybrid_core_inst_x_rsc_13_0_RDATA;
  hybrid_core_inst_x_rsc_13_0_ARREGION <= x_rsc_13_0_ARREGION;
  hybrid_core_inst_x_rsc_13_0_ARQOS <= x_rsc_13_0_ARQOS;
  hybrid_core_inst_x_rsc_13_0_ARPROT <= x_rsc_13_0_ARPROT;
  hybrid_core_inst_x_rsc_13_0_ARCACHE <= x_rsc_13_0_ARCACHE;
  hybrid_core_inst_x_rsc_13_0_ARBURST <= x_rsc_13_0_ARBURST;
  hybrid_core_inst_x_rsc_13_0_ARSIZE <= x_rsc_13_0_ARSIZE;
  hybrid_core_inst_x_rsc_13_0_ARLEN <= x_rsc_13_0_ARLEN;
  hybrid_core_inst_x_rsc_13_0_ARADDR <= x_rsc_13_0_ARADDR;
  x_rsc_13_0_BRESP <= hybrid_core_inst_x_rsc_13_0_BRESP;
  hybrid_core_inst_x_rsc_13_0_WSTRB <= x_rsc_13_0_WSTRB;
  hybrid_core_inst_x_rsc_13_0_WDATA <= x_rsc_13_0_WDATA;
  hybrid_core_inst_x_rsc_13_0_AWREGION <= x_rsc_13_0_AWREGION;
  hybrid_core_inst_x_rsc_13_0_AWQOS <= x_rsc_13_0_AWQOS;
  hybrid_core_inst_x_rsc_13_0_AWPROT <= x_rsc_13_0_AWPROT;
  hybrid_core_inst_x_rsc_13_0_AWCACHE <= x_rsc_13_0_AWCACHE;
  hybrid_core_inst_x_rsc_13_0_AWBURST <= x_rsc_13_0_AWBURST;
  hybrid_core_inst_x_rsc_13_0_AWSIZE <= x_rsc_13_0_AWSIZE;
  hybrid_core_inst_x_rsc_13_0_AWLEN <= x_rsc_13_0_AWLEN;
  hybrid_core_inst_x_rsc_13_0_AWADDR <= x_rsc_13_0_AWADDR;
  x_rsc_14_0_RRESP <= hybrid_core_inst_x_rsc_14_0_RRESP;
  x_rsc_14_0_RDATA <= hybrid_core_inst_x_rsc_14_0_RDATA;
  hybrid_core_inst_x_rsc_14_0_ARREGION <= x_rsc_14_0_ARREGION;
  hybrid_core_inst_x_rsc_14_0_ARQOS <= x_rsc_14_0_ARQOS;
  hybrid_core_inst_x_rsc_14_0_ARPROT <= x_rsc_14_0_ARPROT;
  hybrid_core_inst_x_rsc_14_0_ARCACHE <= x_rsc_14_0_ARCACHE;
  hybrid_core_inst_x_rsc_14_0_ARBURST <= x_rsc_14_0_ARBURST;
  hybrid_core_inst_x_rsc_14_0_ARSIZE <= x_rsc_14_0_ARSIZE;
  hybrid_core_inst_x_rsc_14_0_ARLEN <= x_rsc_14_0_ARLEN;
  hybrid_core_inst_x_rsc_14_0_ARADDR <= x_rsc_14_0_ARADDR;
  x_rsc_14_0_BRESP <= hybrid_core_inst_x_rsc_14_0_BRESP;
  hybrid_core_inst_x_rsc_14_0_WSTRB <= x_rsc_14_0_WSTRB;
  hybrid_core_inst_x_rsc_14_0_WDATA <= x_rsc_14_0_WDATA;
  hybrid_core_inst_x_rsc_14_0_AWREGION <= x_rsc_14_0_AWREGION;
  hybrid_core_inst_x_rsc_14_0_AWQOS <= x_rsc_14_0_AWQOS;
  hybrid_core_inst_x_rsc_14_0_AWPROT <= x_rsc_14_0_AWPROT;
  hybrid_core_inst_x_rsc_14_0_AWCACHE <= x_rsc_14_0_AWCACHE;
  hybrid_core_inst_x_rsc_14_0_AWBURST <= x_rsc_14_0_AWBURST;
  hybrid_core_inst_x_rsc_14_0_AWSIZE <= x_rsc_14_0_AWSIZE;
  hybrid_core_inst_x_rsc_14_0_AWLEN <= x_rsc_14_0_AWLEN;
  hybrid_core_inst_x_rsc_14_0_AWADDR <= x_rsc_14_0_AWADDR;
  x_rsc_15_0_RRESP <= hybrid_core_inst_x_rsc_15_0_RRESP;
  x_rsc_15_0_RDATA <= hybrid_core_inst_x_rsc_15_0_RDATA;
  hybrid_core_inst_x_rsc_15_0_ARREGION <= x_rsc_15_0_ARREGION;
  hybrid_core_inst_x_rsc_15_0_ARQOS <= x_rsc_15_0_ARQOS;
  hybrid_core_inst_x_rsc_15_0_ARPROT <= x_rsc_15_0_ARPROT;
  hybrid_core_inst_x_rsc_15_0_ARCACHE <= x_rsc_15_0_ARCACHE;
  hybrid_core_inst_x_rsc_15_0_ARBURST <= x_rsc_15_0_ARBURST;
  hybrid_core_inst_x_rsc_15_0_ARSIZE <= x_rsc_15_0_ARSIZE;
  hybrid_core_inst_x_rsc_15_0_ARLEN <= x_rsc_15_0_ARLEN;
  hybrid_core_inst_x_rsc_15_0_ARADDR <= x_rsc_15_0_ARADDR;
  x_rsc_15_0_BRESP <= hybrid_core_inst_x_rsc_15_0_BRESP;
  hybrid_core_inst_x_rsc_15_0_WSTRB <= x_rsc_15_0_WSTRB;
  hybrid_core_inst_x_rsc_15_0_WDATA <= x_rsc_15_0_WDATA;
  hybrid_core_inst_x_rsc_15_0_AWREGION <= x_rsc_15_0_AWREGION;
  hybrid_core_inst_x_rsc_15_0_AWQOS <= x_rsc_15_0_AWQOS;
  hybrid_core_inst_x_rsc_15_0_AWPROT <= x_rsc_15_0_AWPROT;
  hybrid_core_inst_x_rsc_15_0_AWCACHE <= x_rsc_15_0_AWCACHE;
  hybrid_core_inst_x_rsc_15_0_AWBURST <= x_rsc_15_0_AWBURST;
  hybrid_core_inst_x_rsc_15_0_AWSIZE <= x_rsc_15_0_AWSIZE;
  hybrid_core_inst_x_rsc_15_0_AWLEN <= x_rsc_15_0_AWLEN;
  hybrid_core_inst_x_rsc_15_0_AWADDR <= x_rsc_15_0_AWADDR;
  x_rsc_16_0_RRESP <= hybrid_core_inst_x_rsc_16_0_RRESP;
  x_rsc_16_0_RDATA <= hybrid_core_inst_x_rsc_16_0_RDATA;
  hybrid_core_inst_x_rsc_16_0_ARREGION <= x_rsc_16_0_ARREGION;
  hybrid_core_inst_x_rsc_16_0_ARQOS <= x_rsc_16_0_ARQOS;
  hybrid_core_inst_x_rsc_16_0_ARPROT <= x_rsc_16_0_ARPROT;
  hybrid_core_inst_x_rsc_16_0_ARCACHE <= x_rsc_16_0_ARCACHE;
  hybrid_core_inst_x_rsc_16_0_ARBURST <= x_rsc_16_0_ARBURST;
  hybrid_core_inst_x_rsc_16_0_ARSIZE <= x_rsc_16_0_ARSIZE;
  hybrid_core_inst_x_rsc_16_0_ARLEN <= x_rsc_16_0_ARLEN;
  hybrid_core_inst_x_rsc_16_0_ARADDR <= x_rsc_16_0_ARADDR;
  x_rsc_16_0_BRESP <= hybrid_core_inst_x_rsc_16_0_BRESP;
  hybrid_core_inst_x_rsc_16_0_WSTRB <= x_rsc_16_0_WSTRB;
  hybrid_core_inst_x_rsc_16_0_WDATA <= x_rsc_16_0_WDATA;
  hybrid_core_inst_x_rsc_16_0_AWREGION <= x_rsc_16_0_AWREGION;
  hybrid_core_inst_x_rsc_16_0_AWQOS <= x_rsc_16_0_AWQOS;
  hybrid_core_inst_x_rsc_16_0_AWPROT <= x_rsc_16_0_AWPROT;
  hybrid_core_inst_x_rsc_16_0_AWCACHE <= x_rsc_16_0_AWCACHE;
  hybrid_core_inst_x_rsc_16_0_AWBURST <= x_rsc_16_0_AWBURST;
  hybrid_core_inst_x_rsc_16_0_AWSIZE <= x_rsc_16_0_AWSIZE;
  hybrid_core_inst_x_rsc_16_0_AWLEN <= x_rsc_16_0_AWLEN;
  hybrid_core_inst_x_rsc_16_0_AWADDR <= x_rsc_16_0_AWADDR;
  x_rsc_17_0_RRESP <= hybrid_core_inst_x_rsc_17_0_RRESP;
  x_rsc_17_0_RDATA <= hybrid_core_inst_x_rsc_17_0_RDATA;
  hybrid_core_inst_x_rsc_17_0_ARREGION <= x_rsc_17_0_ARREGION;
  hybrid_core_inst_x_rsc_17_0_ARQOS <= x_rsc_17_0_ARQOS;
  hybrid_core_inst_x_rsc_17_0_ARPROT <= x_rsc_17_0_ARPROT;
  hybrid_core_inst_x_rsc_17_0_ARCACHE <= x_rsc_17_0_ARCACHE;
  hybrid_core_inst_x_rsc_17_0_ARBURST <= x_rsc_17_0_ARBURST;
  hybrid_core_inst_x_rsc_17_0_ARSIZE <= x_rsc_17_0_ARSIZE;
  hybrid_core_inst_x_rsc_17_0_ARLEN <= x_rsc_17_0_ARLEN;
  hybrid_core_inst_x_rsc_17_0_ARADDR <= x_rsc_17_0_ARADDR;
  x_rsc_17_0_BRESP <= hybrid_core_inst_x_rsc_17_0_BRESP;
  hybrid_core_inst_x_rsc_17_0_WSTRB <= x_rsc_17_0_WSTRB;
  hybrid_core_inst_x_rsc_17_0_WDATA <= x_rsc_17_0_WDATA;
  hybrid_core_inst_x_rsc_17_0_AWREGION <= x_rsc_17_0_AWREGION;
  hybrid_core_inst_x_rsc_17_0_AWQOS <= x_rsc_17_0_AWQOS;
  hybrid_core_inst_x_rsc_17_0_AWPROT <= x_rsc_17_0_AWPROT;
  hybrid_core_inst_x_rsc_17_0_AWCACHE <= x_rsc_17_0_AWCACHE;
  hybrid_core_inst_x_rsc_17_0_AWBURST <= x_rsc_17_0_AWBURST;
  hybrid_core_inst_x_rsc_17_0_AWSIZE <= x_rsc_17_0_AWSIZE;
  hybrid_core_inst_x_rsc_17_0_AWLEN <= x_rsc_17_0_AWLEN;
  hybrid_core_inst_x_rsc_17_0_AWADDR <= x_rsc_17_0_AWADDR;
  x_rsc_18_0_RRESP <= hybrid_core_inst_x_rsc_18_0_RRESP;
  x_rsc_18_0_RDATA <= hybrid_core_inst_x_rsc_18_0_RDATA;
  hybrid_core_inst_x_rsc_18_0_ARREGION <= x_rsc_18_0_ARREGION;
  hybrid_core_inst_x_rsc_18_0_ARQOS <= x_rsc_18_0_ARQOS;
  hybrid_core_inst_x_rsc_18_0_ARPROT <= x_rsc_18_0_ARPROT;
  hybrid_core_inst_x_rsc_18_0_ARCACHE <= x_rsc_18_0_ARCACHE;
  hybrid_core_inst_x_rsc_18_0_ARBURST <= x_rsc_18_0_ARBURST;
  hybrid_core_inst_x_rsc_18_0_ARSIZE <= x_rsc_18_0_ARSIZE;
  hybrid_core_inst_x_rsc_18_0_ARLEN <= x_rsc_18_0_ARLEN;
  hybrid_core_inst_x_rsc_18_0_ARADDR <= x_rsc_18_0_ARADDR;
  x_rsc_18_0_BRESP <= hybrid_core_inst_x_rsc_18_0_BRESP;
  hybrid_core_inst_x_rsc_18_0_WSTRB <= x_rsc_18_0_WSTRB;
  hybrid_core_inst_x_rsc_18_0_WDATA <= x_rsc_18_0_WDATA;
  hybrid_core_inst_x_rsc_18_0_AWREGION <= x_rsc_18_0_AWREGION;
  hybrid_core_inst_x_rsc_18_0_AWQOS <= x_rsc_18_0_AWQOS;
  hybrid_core_inst_x_rsc_18_0_AWPROT <= x_rsc_18_0_AWPROT;
  hybrid_core_inst_x_rsc_18_0_AWCACHE <= x_rsc_18_0_AWCACHE;
  hybrid_core_inst_x_rsc_18_0_AWBURST <= x_rsc_18_0_AWBURST;
  hybrid_core_inst_x_rsc_18_0_AWSIZE <= x_rsc_18_0_AWSIZE;
  hybrid_core_inst_x_rsc_18_0_AWLEN <= x_rsc_18_0_AWLEN;
  hybrid_core_inst_x_rsc_18_0_AWADDR <= x_rsc_18_0_AWADDR;
  x_rsc_19_0_RRESP <= hybrid_core_inst_x_rsc_19_0_RRESP;
  x_rsc_19_0_RDATA <= hybrid_core_inst_x_rsc_19_0_RDATA;
  hybrid_core_inst_x_rsc_19_0_ARREGION <= x_rsc_19_0_ARREGION;
  hybrid_core_inst_x_rsc_19_0_ARQOS <= x_rsc_19_0_ARQOS;
  hybrid_core_inst_x_rsc_19_0_ARPROT <= x_rsc_19_0_ARPROT;
  hybrid_core_inst_x_rsc_19_0_ARCACHE <= x_rsc_19_0_ARCACHE;
  hybrid_core_inst_x_rsc_19_0_ARBURST <= x_rsc_19_0_ARBURST;
  hybrid_core_inst_x_rsc_19_0_ARSIZE <= x_rsc_19_0_ARSIZE;
  hybrid_core_inst_x_rsc_19_0_ARLEN <= x_rsc_19_0_ARLEN;
  hybrid_core_inst_x_rsc_19_0_ARADDR <= x_rsc_19_0_ARADDR;
  x_rsc_19_0_BRESP <= hybrid_core_inst_x_rsc_19_0_BRESP;
  hybrid_core_inst_x_rsc_19_0_WSTRB <= x_rsc_19_0_WSTRB;
  hybrid_core_inst_x_rsc_19_0_WDATA <= x_rsc_19_0_WDATA;
  hybrid_core_inst_x_rsc_19_0_AWREGION <= x_rsc_19_0_AWREGION;
  hybrid_core_inst_x_rsc_19_0_AWQOS <= x_rsc_19_0_AWQOS;
  hybrid_core_inst_x_rsc_19_0_AWPROT <= x_rsc_19_0_AWPROT;
  hybrid_core_inst_x_rsc_19_0_AWCACHE <= x_rsc_19_0_AWCACHE;
  hybrid_core_inst_x_rsc_19_0_AWBURST <= x_rsc_19_0_AWBURST;
  hybrid_core_inst_x_rsc_19_0_AWSIZE <= x_rsc_19_0_AWSIZE;
  hybrid_core_inst_x_rsc_19_0_AWLEN <= x_rsc_19_0_AWLEN;
  hybrid_core_inst_x_rsc_19_0_AWADDR <= x_rsc_19_0_AWADDR;
  x_rsc_20_0_RRESP <= hybrid_core_inst_x_rsc_20_0_RRESP;
  x_rsc_20_0_RDATA <= hybrid_core_inst_x_rsc_20_0_RDATA;
  hybrid_core_inst_x_rsc_20_0_ARREGION <= x_rsc_20_0_ARREGION;
  hybrid_core_inst_x_rsc_20_0_ARQOS <= x_rsc_20_0_ARQOS;
  hybrid_core_inst_x_rsc_20_0_ARPROT <= x_rsc_20_0_ARPROT;
  hybrid_core_inst_x_rsc_20_0_ARCACHE <= x_rsc_20_0_ARCACHE;
  hybrid_core_inst_x_rsc_20_0_ARBURST <= x_rsc_20_0_ARBURST;
  hybrid_core_inst_x_rsc_20_0_ARSIZE <= x_rsc_20_0_ARSIZE;
  hybrid_core_inst_x_rsc_20_0_ARLEN <= x_rsc_20_0_ARLEN;
  hybrid_core_inst_x_rsc_20_0_ARADDR <= x_rsc_20_0_ARADDR;
  x_rsc_20_0_BRESP <= hybrid_core_inst_x_rsc_20_0_BRESP;
  hybrid_core_inst_x_rsc_20_0_WSTRB <= x_rsc_20_0_WSTRB;
  hybrid_core_inst_x_rsc_20_0_WDATA <= x_rsc_20_0_WDATA;
  hybrid_core_inst_x_rsc_20_0_AWREGION <= x_rsc_20_0_AWREGION;
  hybrid_core_inst_x_rsc_20_0_AWQOS <= x_rsc_20_0_AWQOS;
  hybrid_core_inst_x_rsc_20_0_AWPROT <= x_rsc_20_0_AWPROT;
  hybrid_core_inst_x_rsc_20_0_AWCACHE <= x_rsc_20_0_AWCACHE;
  hybrid_core_inst_x_rsc_20_0_AWBURST <= x_rsc_20_0_AWBURST;
  hybrid_core_inst_x_rsc_20_0_AWSIZE <= x_rsc_20_0_AWSIZE;
  hybrid_core_inst_x_rsc_20_0_AWLEN <= x_rsc_20_0_AWLEN;
  hybrid_core_inst_x_rsc_20_0_AWADDR <= x_rsc_20_0_AWADDR;
  x_rsc_21_0_RRESP <= hybrid_core_inst_x_rsc_21_0_RRESP;
  x_rsc_21_0_RDATA <= hybrid_core_inst_x_rsc_21_0_RDATA;
  hybrid_core_inst_x_rsc_21_0_ARREGION <= x_rsc_21_0_ARREGION;
  hybrid_core_inst_x_rsc_21_0_ARQOS <= x_rsc_21_0_ARQOS;
  hybrid_core_inst_x_rsc_21_0_ARPROT <= x_rsc_21_0_ARPROT;
  hybrid_core_inst_x_rsc_21_0_ARCACHE <= x_rsc_21_0_ARCACHE;
  hybrid_core_inst_x_rsc_21_0_ARBURST <= x_rsc_21_0_ARBURST;
  hybrid_core_inst_x_rsc_21_0_ARSIZE <= x_rsc_21_0_ARSIZE;
  hybrid_core_inst_x_rsc_21_0_ARLEN <= x_rsc_21_0_ARLEN;
  hybrid_core_inst_x_rsc_21_0_ARADDR <= x_rsc_21_0_ARADDR;
  x_rsc_21_0_BRESP <= hybrid_core_inst_x_rsc_21_0_BRESP;
  hybrid_core_inst_x_rsc_21_0_WSTRB <= x_rsc_21_0_WSTRB;
  hybrid_core_inst_x_rsc_21_0_WDATA <= x_rsc_21_0_WDATA;
  hybrid_core_inst_x_rsc_21_0_AWREGION <= x_rsc_21_0_AWREGION;
  hybrid_core_inst_x_rsc_21_0_AWQOS <= x_rsc_21_0_AWQOS;
  hybrid_core_inst_x_rsc_21_0_AWPROT <= x_rsc_21_0_AWPROT;
  hybrid_core_inst_x_rsc_21_0_AWCACHE <= x_rsc_21_0_AWCACHE;
  hybrid_core_inst_x_rsc_21_0_AWBURST <= x_rsc_21_0_AWBURST;
  hybrid_core_inst_x_rsc_21_0_AWSIZE <= x_rsc_21_0_AWSIZE;
  hybrid_core_inst_x_rsc_21_0_AWLEN <= x_rsc_21_0_AWLEN;
  hybrid_core_inst_x_rsc_21_0_AWADDR <= x_rsc_21_0_AWADDR;
  x_rsc_22_0_RRESP <= hybrid_core_inst_x_rsc_22_0_RRESP;
  x_rsc_22_0_RDATA <= hybrid_core_inst_x_rsc_22_0_RDATA;
  hybrid_core_inst_x_rsc_22_0_ARREGION <= x_rsc_22_0_ARREGION;
  hybrid_core_inst_x_rsc_22_0_ARQOS <= x_rsc_22_0_ARQOS;
  hybrid_core_inst_x_rsc_22_0_ARPROT <= x_rsc_22_0_ARPROT;
  hybrid_core_inst_x_rsc_22_0_ARCACHE <= x_rsc_22_0_ARCACHE;
  hybrid_core_inst_x_rsc_22_0_ARBURST <= x_rsc_22_0_ARBURST;
  hybrid_core_inst_x_rsc_22_0_ARSIZE <= x_rsc_22_0_ARSIZE;
  hybrid_core_inst_x_rsc_22_0_ARLEN <= x_rsc_22_0_ARLEN;
  hybrid_core_inst_x_rsc_22_0_ARADDR <= x_rsc_22_0_ARADDR;
  x_rsc_22_0_BRESP <= hybrid_core_inst_x_rsc_22_0_BRESP;
  hybrid_core_inst_x_rsc_22_0_WSTRB <= x_rsc_22_0_WSTRB;
  hybrid_core_inst_x_rsc_22_0_WDATA <= x_rsc_22_0_WDATA;
  hybrid_core_inst_x_rsc_22_0_AWREGION <= x_rsc_22_0_AWREGION;
  hybrid_core_inst_x_rsc_22_0_AWQOS <= x_rsc_22_0_AWQOS;
  hybrid_core_inst_x_rsc_22_0_AWPROT <= x_rsc_22_0_AWPROT;
  hybrid_core_inst_x_rsc_22_0_AWCACHE <= x_rsc_22_0_AWCACHE;
  hybrid_core_inst_x_rsc_22_0_AWBURST <= x_rsc_22_0_AWBURST;
  hybrid_core_inst_x_rsc_22_0_AWSIZE <= x_rsc_22_0_AWSIZE;
  hybrid_core_inst_x_rsc_22_0_AWLEN <= x_rsc_22_0_AWLEN;
  hybrid_core_inst_x_rsc_22_0_AWADDR <= x_rsc_22_0_AWADDR;
  x_rsc_23_0_RRESP <= hybrid_core_inst_x_rsc_23_0_RRESP;
  x_rsc_23_0_RDATA <= hybrid_core_inst_x_rsc_23_0_RDATA;
  hybrid_core_inst_x_rsc_23_0_ARREGION <= x_rsc_23_0_ARREGION;
  hybrid_core_inst_x_rsc_23_0_ARQOS <= x_rsc_23_0_ARQOS;
  hybrid_core_inst_x_rsc_23_0_ARPROT <= x_rsc_23_0_ARPROT;
  hybrid_core_inst_x_rsc_23_0_ARCACHE <= x_rsc_23_0_ARCACHE;
  hybrid_core_inst_x_rsc_23_0_ARBURST <= x_rsc_23_0_ARBURST;
  hybrid_core_inst_x_rsc_23_0_ARSIZE <= x_rsc_23_0_ARSIZE;
  hybrid_core_inst_x_rsc_23_0_ARLEN <= x_rsc_23_0_ARLEN;
  hybrid_core_inst_x_rsc_23_0_ARADDR <= x_rsc_23_0_ARADDR;
  x_rsc_23_0_BRESP <= hybrid_core_inst_x_rsc_23_0_BRESP;
  hybrid_core_inst_x_rsc_23_0_WSTRB <= x_rsc_23_0_WSTRB;
  hybrid_core_inst_x_rsc_23_0_WDATA <= x_rsc_23_0_WDATA;
  hybrid_core_inst_x_rsc_23_0_AWREGION <= x_rsc_23_0_AWREGION;
  hybrid_core_inst_x_rsc_23_0_AWQOS <= x_rsc_23_0_AWQOS;
  hybrid_core_inst_x_rsc_23_0_AWPROT <= x_rsc_23_0_AWPROT;
  hybrid_core_inst_x_rsc_23_0_AWCACHE <= x_rsc_23_0_AWCACHE;
  hybrid_core_inst_x_rsc_23_0_AWBURST <= x_rsc_23_0_AWBURST;
  hybrid_core_inst_x_rsc_23_0_AWSIZE <= x_rsc_23_0_AWSIZE;
  hybrid_core_inst_x_rsc_23_0_AWLEN <= x_rsc_23_0_AWLEN;
  hybrid_core_inst_x_rsc_23_0_AWADDR <= x_rsc_23_0_AWADDR;
  x_rsc_24_0_RRESP <= hybrid_core_inst_x_rsc_24_0_RRESP;
  x_rsc_24_0_RDATA <= hybrid_core_inst_x_rsc_24_0_RDATA;
  hybrid_core_inst_x_rsc_24_0_ARREGION <= x_rsc_24_0_ARREGION;
  hybrid_core_inst_x_rsc_24_0_ARQOS <= x_rsc_24_0_ARQOS;
  hybrid_core_inst_x_rsc_24_0_ARPROT <= x_rsc_24_0_ARPROT;
  hybrid_core_inst_x_rsc_24_0_ARCACHE <= x_rsc_24_0_ARCACHE;
  hybrid_core_inst_x_rsc_24_0_ARBURST <= x_rsc_24_0_ARBURST;
  hybrid_core_inst_x_rsc_24_0_ARSIZE <= x_rsc_24_0_ARSIZE;
  hybrid_core_inst_x_rsc_24_0_ARLEN <= x_rsc_24_0_ARLEN;
  hybrid_core_inst_x_rsc_24_0_ARADDR <= x_rsc_24_0_ARADDR;
  x_rsc_24_0_BRESP <= hybrid_core_inst_x_rsc_24_0_BRESP;
  hybrid_core_inst_x_rsc_24_0_WSTRB <= x_rsc_24_0_WSTRB;
  hybrid_core_inst_x_rsc_24_0_WDATA <= x_rsc_24_0_WDATA;
  hybrid_core_inst_x_rsc_24_0_AWREGION <= x_rsc_24_0_AWREGION;
  hybrid_core_inst_x_rsc_24_0_AWQOS <= x_rsc_24_0_AWQOS;
  hybrid_core_inst_x_rsc_24_0_AWPROT <= x_rsc_24_0_AWPROT;
  hybrid_core_inst_x_rsc_24_0_AWCACHE <= x_rsc_24_0_AWCACHE;
  hybrid_core_inst_x_rsc_24_0_AWBURST <= x_rsc_24_0_AWBURST;
  hybrid_core_inst_x_rsc_24_0_AWSIZE <= x_rsc_24_0_AWSIZE;
  hybrid_core_inst_x_rsc_24_0_AWLEN <= x_rsc_24_0_AWLEN;
  hybrid_core_inst_x_rsc_24_0_AWADDR <= x_rsc_24_0_AWADDR;
  x_rsc_25_0_RRESP <= hybrid_core_inst_x_rsc_25_0_RRESP;
  x_rsc_25_0_RDATA <= hybrid_core_inst_x_rsc_25_0_RDATA;
  hybrid_core_inst_x_rsc_25_0_ARREGION <= x_rsc_25_0_ARREGION;
  hybrid_core_inst_x_rsc_25_0_ARQOS <= x_rsc_25_0_ARQOS;
  hybrid_core_inst_x_rsc_25_0_ARPROT <= x_rsc_25_0_ARPROT;
  hybrid_core_inst_x_rsc_25_0_ARCACHE <= x_rsc_25_0_ARCACHE;
  hybrid_core_inst_x_rsc_25_0_ARBURST <= x_rsc_25_0_ARBURST;
  hybrid_core_inst_x_rsc_25_0_ARSIZE <= x_rsc_25_0_ARSIZE;
  hybrid_core_inst_x_rsc_25_0_ARLEN <= x_rsc_25_0_ARLEN;
  hybrid_core_inst_x_rsc_25_0_ARADDR <= x_rsc_25_0_ARADDR;
  x_rsc_25_0_BRESP <= hybrid_core_inst_x_rsc_25_0_BRESP;
  hybrid_core_inst_x_rsc_25_0_WSTRB <= x_rsc_25_0_WSTRB;
  hybrid_core_inst_x_rsc_25_0_WDATA <= x_rsc_25_0_WDATA;
  hybrid_core_inst_x_rsc_25_0_AWREGION <= x_rsc_25_0_AWREGION;
  hybrid_core_inst_x_rsc_25_0_AWQOS <= x_rsc_25_0_AWQOS;
  hybrid_core_inst_x_rsc_25_0_AWPROT <= x_rsc_25_0_AWPROT;
  hybrid_core_inst_x_rsc_25_0_AWCACHE <= x_rsc_25_0_AWCACHE;
  hybrid_core_inst_x_rsc_25_0_AWBURST <= x_rsc_25_0_AWBURST;
  hybrid_core_inst_x_rsc_25_0_AWSIZE <= x_rsc_25_0_AWSIZE;
  hybrid_core_inst_x_rsc_25_0_AWLEN <= x_rsc_25_0_AWLEN;
  hybrid_core_inst_x_rsc_25_0_AWADDR <= x_rsc_25_0_AWADDR;
  x_rsc_26_0_RRESP <= hybrid_core_inst_x_rsc_26_0_RRESP;
  x_rsc_26_0_RDATA <= hybrid_core_inst_x_rsc_26_0_RDATA;
  hybrid_core_inst_x_rsc_26_0_ARREGION <= x_rsc_26_0_ARREGION;
  hybrid_core_inst_x_rsc_26_0_ARQOS <= x_rsc_26_0_ARQOS;
  hybrid_core_inst_x_rsc_26_0_ARPROT <= x_rsc_26_0_ARPROT;
  hybrid_core_inst_x_rsc_26_0_ARCACHE <= x_rsc_26_0_ARCACHE;
  hybrid_core_inst_x_rsc_26_0_ARBURST <= x_rsc_26_0_ARBURST;
  hybrid_core_inst_x_rsc_26_0_ARSIZE <= x_rsc_26_0_ARSIZE;
  hybrid_core_inst_x_rsc_26_0_ARLEN <= x_rsc_26_0_ARLEN;
  hybrid_core_inst_x_rsc_26_0_ARADDR <= x_rsc_26_0_ARADDR;
  x_rsc_26_0_BRESP <= hybrid_core_inst_x_rsc_26_0_BRESP;
  hybrid_core_inst_x_rsc_26_0_WSTRB <= x_rsc_26_0_WSTRB;
  hybrid_core_inst_x_rsc_26_0_WDATA <= x_rsc_26_0_WDATA;
  hybrid_core_inst_x_rsc_26_0_AWREGION <= x_rsc_26_0_AWREGION;
  hybrid_core_inst_x_rsc_26_0_AWQOS <= x_rsc_26_0_AWQOS;
  hybrid_core_inst_x_rsc_26_0_AWPROT <= x_rsc_26_0_AWPROT;
  hybrid_core_inst_x_rsc_26_0_AWCACHE <= x_rsc_26_0_AWCACHE;
  hybrid_core_inst_x_rsc_26_0_AWBURST <= x_rsc_26_0_AWBURST;
  hybrid_core_inst_x_rsc_26_0_AWSIZE <= x_rsc_26_0_AWSIZE;
  hybrid_core_inst_x_rsc_26_0_AWLEN <= x_rsc_26_0_AWLEN;
  hybrid_core_inst_x_rsc_26_0_AWADDR <= x_rsc_26_0_AWADDR;
  x_rsc_27_0_RRESP <= hybrid_core_inst_x_rsc_27_0_RRESP;
  x_rsc_27_0_RDATA <= hybrid_core_inst_x_rsc_27_0_RDATA;
  hybrid_core_inst_x_rsc_27_0_ARREGION <= x_rsc_27_0_ARREGION;
  hybrid_core_inst_x_rsc_27_0_ARQOS <= x_rsc_27_0_ARQOS;
  hybrid_core_inst_x_rsc_27_0_ARPROT <= x_rsc_27_0_ARPROT;
  hybrid_core_inst_x_rsc_27_0_ARCACHE <= x_rsc_27_0_ARCACHE;
  hybrid_core_inst_x_rsc_27_0_ARBURST <= x_rsc_27_0_ARBURST;
  hybrid_core_inst_x_rsc_27_0_ARSIZE <= x_rsc_27_0_ARSIZE;
  hybrid_core_inst_x_rsc_27_0_ARLEN <= x_rsc_27_0_ARLEN;
  hybrid_core_inst_x_rsc_27_0_ARADDR <= x_rsc_27_0_ARADDR;
  x_rsc_27_0_BRESP <= hybrid_core_inst_x_rsc_27_0_BRESP;
  hybrid_core_inst_x_rsc_27_0_WSTRB <= x_rsc_27_0_WSTRB;
  hybrid_core_inst_x_rsc_27_0_WDATA <= x_rsc_27_0_WDATA;
  hybrid_core_inst_x_rsc_27_0_AWREGION <= x_rsc_27_0_AWREGION;
  hybrid_core_inst_x_rsc_27_0_AWQOS <= x_rsc_27_0_AWQOS;
  hybrid_core_inst_x_rsc_27_0_AWPROT <= x_rsc_27_0_AWPROT;
  hybrid_core_inst_x_rsc_27_0_AWCACHE <= x_rsc_27_0_AWCACHE;
  hybrid_core_inst_x_rsc_27_0_AWBURST <= x_rsc_27_0_AWBURST;
  hybrid_core_inst_x_rsc_27_0_AWSIZE <= x_rsc_27_0_AWSIZE;
  hybrid_core_inst_x_rsc_27_0_AWLEN <= x_rsc_27_0_AWLEN;
  hybrid_core_inst_x_rsc_27_0_AWADDR <= x_rsc_27_0_AWADDR;
  x_rsc_28_0_RRESP <= hybrid_core_inst_x_rsc_28_0_RRESP;
  x_rsc_28_0_RDATA <= hybrid_core_inst_x_rsc_28_0_RDATA;
  hybrid_core_inst_x_rsc_28_0_ARREGION <= x_rsc_28_0_ARREGION;
  hybrid_core_inst_x_rsc_28_0_ARQOS <= x_rsc_28_0_ARQOS;
  hybrid_core_inst_x_rsc_28_0_ARPROT <= x_rsc_28_0_ARPROT;
  hybrid_core_inst_x_rsc_28_0_ARCACHE <= x_rsc_28_0_ARCACHE;
  hybrid_core_inst_x_rsc_28_0_ARBURST <= x_rsc_28_0_ARBURST;
  hybrid_core_inst_x_rsc_28_0_ARSIZE <= x_rsc_28_0_ARSIZE;
  hybrid_core_inst_x_rsc_28_0_ARLEN <= x_rsc_28_0_ARLEN;
  hybrid_core_inst_x_rsc_28_0_ARADDR <= x_rsc_28_0_ARADDR;
  x_rsc_28_0_BRESP <= hybrid_core_inst_x_rsc_28_0_BRESP;
  hybrid_core_inst_x_rsc_28_0_WSTRB <= x_rsc_28_0_WSTRB;
  hybrid_core_inst_x_rsc_28_0_WDATA <= x_rsc_28_0_WDATA;
  hybrid_core_inst_x_rsc_28_0_AWREGION <= x_rsc_28_0_AWREGION;
  hybrid_core_inst_x_rsc_28_0_AWQOS <= x_rsc_28_0_AWQOS;
  hybrid_core_inst_x_rsc_28_0_AWPROT <= x_rsc_28_0_AWPROT;
  hybrid_core_inst_x_rsc_28_0_AWCACHE <= x_rsc_28_0_AWCACHE;
  hybrid_core_inst_x_rsc_28_0_AWBURST <= x_rsc_28_0_AWBURST;
  hybrid_core_inst_x_rsc_28_0_AWSIZE <= x_rsc_28_0_AWSIZE;
  hybrid_core_inst_x_rsc_28_0_AWLEN <= x_rsc_28_0_AWLEN;
  hybrid_core_inst_x_rsc_28_0_AWADDR <= x_rsc_28_0_AWADDR;
  x_rsc_29_0_RRESP <= hybrid_core_inst_x_rsc_29_0_RRESP;
  x_rsc_29_0_RDATA <= hybrid_core_inst_x_rsc_29_0_RDATA;
  hybrid_core_inst_x_rsc_29_0_ARREGION <= x_rsc_29_0_ARREGION;
  hybrid_core_inst_x_rsc_29_0_ARQOS <= x_rsc_29_0_ARQOS;
  hybrid_core_inst_x_rsc_29_0_ARPROT <= x_rsc_29_0_ARPROT;
  hybrid_core_inst_x_rsc_29_0_ARCACHE <= x_rsc_29_0_ARCACHE;
  hybrid_core_inst_x_rsc_29_0_ARBURST <= x_rsc_29_0_ARBURST;
  hybrid_core_inst_x_rsc_29_0_ARSIZE <= x_rsc_29_0_ARSIZE;
  hybrid_core_inst_x_rsc_29_0_ARLEN <= x_rsc_29_0_ARLEN;
  hybrid_core_inst_x_rsc_29_0_ARADDR <= x_rsc_29_0_ARADDR;
  x_rsc_29_0_BRESP <= hybrid_core_inst_x_rsc_29_0_BRESP;
  hybrid_core_inst_x_rsc_29_0_WSTRB <= x_rsc_29_0_WSTRB;
  hybrid_core_inst_x_rsc_29_0_WDATA <= x_rsc_29_0_WDATA;
  hybrid_core_inst_x_rsc_29_0_AWREGION <= x_rsc_29_0_AWREGION;
  hybrid_core_inst_x_rsc_29_0_AWQOS <= x_rsc_29_0_AWQOS;
  hybrid_core_inst_x_rsc_29_0_AWPROT <= x_rsc_29_0_AWPROT;
  hybrid_core_inst_x_rsc_29_0_AWCACHE <= x_rsc_29_0_AWCACHE;
  hybrid_core_inst_x_rsc_29_0_AWBURST <= x_rsc_29_0_AWBURST;
  hybrid_core_inst_x_rsc_29_0_AWSIZE <= x_rsc_29_0_AWSIZE;
  hybrid_core_inst_x_rsc_29_0_AWLEN <= x_rsc_29_0_AWLEN;
  hybrid_core_inst_x_rsc_29_0_AWADDR <= x_rsc_29_0_AWADDR;
  x_rsc_30_0_RRESP <= hybrid_core_inst_x_rsc_30_0_RRESP;
  x_rsc_30_0_RDATA <= hybrid_core_inst_x_rsc_30_0_RDATA;
  hybrid_core_inst_x_rsc_30_0_ARREGION <= x_rsc_30_0_ARREGION;
  hybrid_core_inst_x_rsc_30_0_ARQOS <= x_rsc_30_0_ARQOS;
  hybrid_core_inst_x_rsc_30_0_ARPROT <= x_rsc_30_0_ARPROT;
  hybrid_core_inst_x_rsc_30_0_ARCACHE <= x_rsc_30_0_ARCACHE;
  hybrid_core_inst_x_rsc_30_0_ARBURST <= x_rsc_30_0_ARBURST;
  hybrid_core_inst_x_rsc_30_0_ARSIZE <= x_rsc_30_0_ARSIZE;
  hybrid_core_inst_x_rsc_30_0_ARLEN <= x_rsc_30_0_ARLEN;
  hybrid_core_inst_x_rsc_30_0_ARADDR <= x_rsc_30_0_ARADDR;
  x_rsc_30_0_BRESP <= hybrid_core_inst_x_rsc_30_0_BRESP;
  hybrid_core_inst_x_rsc_30_0_WSTRB <= x_rsc_30_0_WSTRB;
  hybrid_core_inst_x_rsc_30_0_WDATA <= x_rsc_30_0_WDATA;
  hybrid_core_inst_x_rsc_30_0_AWREGION <= x_rsc_30_0_AWREGION;
  hybrid_core_inst_x_rsc_30_0_AWQOS <= x_rsc_30_0_AWQOS;
  hybrid_core_inst_x_rsc_30_0_AWPROT <= x_rsc_30_0_AWPROT;
  hybrid_core_inst_x_rsc_30_0_AWCACHE <= x_rsc_30_0_AWCACHE;
  hybrid_core_inst_x_rsc_30_0_AWBURST <= x_rsc_30_0_AWBURST;
  hybrid_core_inst_x_rsc_30_0_AWSIZE <= x_rsc_30_0_AWSIZE;
  hybrid_core_inst_x_rsc_30_0_AWLEN <= x_rsc_30_0_AWLEN;
  hybrid_core_inst_x_rsc_30_0_AWADDR <= x_rsc_30_0_AWADDR;
  x_rsc_31_0_RRESP <= hybrid_core_inst_x_rsc_31_0_RRESP;
  x_rsc_31_0_RDATA <= hybrid_core_inst_x_rsc_31_0_RDATA;
  hybrid_core_inst_x_rsc_31_0_ARREGION <= x_rsc_31_0_ARREGION;
  hybrid_core_inst_x_rsc_31_0_ARQOS <= x_rsc_31_0_ARQOS;
  hybrid_core_inst_x_rsc_31_0_ARPROT <= x_rsc_31_0_ARPROT;
  hybrid_core_inst_x_rsc_31_0_ARCACHE <= x_rsc_31_0_ARCACHE;
  hybrid_core_inst_x_rsc_31_0_ARBURST <= x_rsc_31_0_ARBURST;
  hybrid_core_inst_x_rsc_31_0_ARSIZE <= x_rsc_31_0_ARSIZE;
  hybrid_core_inst_x_rsc_31_0_ARLEN <= x_rsc_31_0_ARLEN;
  hybrid_core_inst_x_rsc_31_0_ARADDR <= x_rsc_31_0_ARADDR;
  x_rsc_31_0_BRESP <= hybrid_core_inst_x_rsc_31_0_BRESP;
  hybrid_core_inst_x_rsc_31_0_WSTRB <= x_rsc_31_0_WSTRB;
  hybrid_core_inst_x_rsc_31_0_WDATA <= x_rsc_31_0_WDATA;
  hybrid_core_inst_x_rsc_31_0_AWREGION <= x_rsc_31_0_AWREGION;
  hybrid_core_inst_x_rsc_31_0_AWQOS <= x_rsc_31_0_AWQOS;
  hybrid_core_inst_x_rsc_31_0_AWPROT <= x_rsc_31_0_AWPROT;
  hybrid_core_inst_x_rsc_31_0_AWCACHE <= x_rsc_31_0_AWCACHE;
  hybrid_core_inst_x_rsc_31_0_AWBURST <= x_rsc_31_0_AWBURST;
  hybrid_core_inst_x_rsc_31_0_AWSIZE <= x_rsc_31_0_AWSIZE;
  hybrid_core_inst_x_rsc_31_0_AWLEN <= x_rsc_31_0_AWLEN;
  hybrid_core_inst_x_rsc_31_0_AWADDR <= x_rsc_31_0_AWADDR;
  hybrid_core_inst_m_rsc_dat <= m_rsc_dat;
  revArr_rsc_RRESP <= hybrid_core_inst_revArr_rsc_RRESP;
  revArr_rsc_RDATA <= hybrid_core_inst_revArr_rsc_RDATA;
  hybrid_core_inst_revArr_rsc_ARREGION <= revArr_rsc_ARREGION;
  hybrid_core_inst_revArr_rsc_ARQOS <= revArr_rsc_ARQOS;
  hybrid_core_inst_revArr_rsc_ARPROT <= revArr_rsc_ARPROT;
  hybrid_core_inst_revArr_rsc_ARCACHE <= revArr_rsc_ARCACHE;
  hybrid_core_inst_revArr_rsc_ARBURST <= revArr_rsc_ARBURST;
  hybrid_core_inst_revArr_rsc_ARSIZE <= revArr_rsc_ARSIZE;
  hybrid_core_inst_revArr_rsc_ARLEN <= revArr_rsc_ARLEN;
  hybrid_core_inst_revArr_rsc_ARADDR <= revArr_rsc_ARADDR;
  revArr_rsc_BRESP <= hybrid_core_inst_revArr_rsc_BRESP;
  hybrid_core_inst_revArr_rsc_WSTRB <= revArr_rsc_WSTRB;
  hybrid_core_inst_revArr_rsc_WDATA <= revArr_rsc_WDATA;
  hybrid_core_inst_revArr_rsc_AWREGION <= revArr_rsc_AWREGION;
  hybrid_core_inst_revArr_rsc_AWQOS <= revArr_rsc_AWQOS;
  hybrid_core_inst_revArr_rsc_AWPROT <= revArr_rsc_AWPROT;
  hybrid_core_inst_revArr_rsc_AWCACHE <= revArr_rsc_AWCACHE;
  hybrid_core_inst_revArr_rsc_AWBURST <= revArr_rsc_AWBURST;
  hybrid_core_inst_revArr_rsc_AWSIZE <= revArr_rsc_AWSIZE;
  hybrid_core_inst_revArr_rsc_AWLEN <= revArr_rsc_AWLEN;
  hybrid_core_inst_revArr_rsc_AWADDR <= revArr_rsc_AWADDR;
  tw_rsc_RRESP <= hybrid_core_inst_tw_rsc_RRESP;
  tw_rsc_RDATA <= hybrid_core_inst_tw_rsc_RDATA;
  hybrid_core_inst_tw_rsc_ARREGION <= tw_rsc_ARREGION;
  hybrid_core_inst_tw_rsc_ARQOS <= tw_rsc_ARQOS;
  hybrid_core_inst_tw_rsc_ARPROT <= tw_rsc_ARPROT;
  hybrid_core_inst_tw_rsc_ARCACHE <= tw_rsc_ARCACHE;
  hybrid_core_inst_tw_rsc_ARBURST <= tw_rsc_ARBURST;
  hybrid_core_inst_tw_rsc_ARSIZE <= tw_rsc_ARSIZE;
  hybrid_core_inst_tw_rsc_ARLEN <= tw_rsc_ARLEN;
  hybrid_core_inst_tw_rsc_ARADDR <= tw_rsc_ARADDR;
  tw_rsc_BRESP <= hybrid_core_inst_tw_rsc_BRESP;
  hybrid_core_inst_tw_rsc_WSTRB <= tw_rsc_WSTRB;
  hybrid_core_inst_tw_rsc_WDATA <= tw_rsc_WDATA;
  hybrid_core_inst_tw_rsc_AWREGION <= tw_rsc_AWREGION;
  hybrid_core_inst_tw_rsc_AWQOS <= tw_rsc_AWQOS;
  hybrid_core_inst_tw_rsc_AWPROT <= tw_rsc_AWPROT;
  hybrid_core_inst_tw_rsc_AWCACHE <= tw_rsc_AWCACHE;
  hybrid_core_inst_tw_rsc_AWBURST <= tw_rsc_AWBURST;
  hybrid_core_inst_tw_rsc_AWSIZE <= tw_rsc_AWSIZE;
  hybrid_core_inst_tw_rsc_AWLEN <= tw_rsc_AWLEN;
  hybrid_core_inst_tw_rsc_AWADDR <= tw_rsc_AWADDR;
  tw_h_rsc_RRESP <= hybrid_core_inst_tw_h_rsc_RRESP;
  tw_h_rsc_RDATA <= hybrid_core_inst_tw_h_rsc_RDATA;
  hybrid_core_inst_tw_h_rsc_ARREGION <= tw_h_rsc_ARREGION;
  hybrid_core_inst_tw_h_rsc_ARQOS <= tw_h_rsc_ARQOS;
  hybrid_core_inst_tw_h_rsc_ARPROT <= tw_h_rsc_ARPROT;
  hybrid_core_inst_tw_h_rsc_ARCACHE <= tw_h_rsc_ARCACHE;
  hybrid_core_inst_tw_h_rsc_ARBURST <= tw_h_rsc_ARBURST;
  hybrid_core_inst_tw_h_rsc_ARSIZE <= tw_h_rsc_ARSIZE;
  hybrid_core_inst_tw_h_rsc_ARLEN <= tw_h_rsc_ARLEN;
  hybrid_core_inst_tw_h_rsc_ARADDR <= tw_h_rsc_ARADDR;
  tw_h_rsc_BRESP <= hybrid_core_inst_tw_h_rsc_BRESP;
  hybrid_core_inst_tw_h_rsc_WSTRB <= tw_h_rsc_WSTRB;
  hybrid_core_inst_tw_h_rsc_WDATA <= tw_h_rsc_WDATA;
  hybrid_core_inst_tw_h_rsc_AWREGION <= tw_h_rsc_AWREGION;
  hybrid_core_inst_tw_h_rsc_AWQOS <= tw_h_rsc_AWQOS;
  hybrid_core_inst_tw_h_rsc_AWPROT <= tw_h_rsc_AWPROT;
  hybrid_core_inst_tw_h_rsc_AWCACHE <= tw_h_rsc_AWCACHE;
  hybrid_core_inst_tw_h_rsc_AWBURST <= tw_h_rsc_AWBURST;
  hybrid_core_inst_tw_h_rsc_AWSIZE <= tw_h_rsc_AWSIZE;
  hybrid_core_inst_tw_h_rsc_AWLEN <= tw_h_rsc_AWLEN;
  hybrid_core_inst_tw_h_rsc_AWADDR <= tw_h_rsc_AWADDR;
  twiddle_rsci_adrb_d <= hybrid_core_inst_twiddle_rsci_adrb_d;
  hybrid_core_inst_twiddle_rsci_qb_d <= twiddle_rsci_qb_d;
  twiddle_h_rsci_adrb_d <= hybrid_core_inst_twiddle_h_rsci_adrb_d;
  hybrid_core_inst_twiddle_h_rsci_qb_d <= twiddle_h_rsci_qb_d;
  xx_rsc_0_0_i_adra_d <= hybrid_core_inst_xx_rsc_0_0_i_adra_d;
  hybrid_core_inst_xx_rsc_0_0_i_qa_d <= xx_rsc_0_0_i_qa_d;
  xx_rsc_0_0_i_wea_d <= hybrid_core_inst_xx_rsc_0_0_i_wea_d;
  xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_1_0_i_adra_d <= hybrid_core_inst_xx_rsc_1_0_i_adra_d;
  hybrid_core_inst_xx_rsc_1_0_i_qa_d <= xx_rsc_1_0_i_qa_d;
  xx_rsc_1_0_i_wea_d <= hybrid_core_inst_xx_rsc_1_0_i_wea_d;
  xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_2_0_i_adra_d <= hybrid_core_inst_xx_rsc_2_0_i_adra_d;
  hybrid_core_inst_xx_rsc_2_0_i_qa_d <= xx_rsc_2_0_i_qa_d;
  xx_rsc_2_0_i_wea_d <= hybrid_core_inst_xx_rsc_2_0_i_wea_d;
  xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_3_0_i_adra_d <= hybrid_core_inst_xx_rsc_3_0_i_adra_d;
  hybrid_core_inst_xx_rsc_3_0_i_qa_d <= xx_rsc_3_0_i_qa_d;
  xx_rsc_3_0_i_wea_d <= hybrid_core_inst_xx_rsc_3_0_i_wea_d;
  xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_4_0_i_adra_d <= hybrid_core_inst_xx_rsc_4_0_i_adra_d;
  hybrid_core_inst_xx_rsc_4_0_i_qa_d <= xx_rsc_4_0_i_qa_d;
  xx_rsc_4_0_i_wea_d <= hybrid_core_inst_xx_rsc_4_0_i_wea_d;
  xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_5_0_i_adra_d <= hybrid_core_inst_xx_rsc_5_0_i_adra_d;
  hybrid_core_inst_xx_rsc_5_0_i_qa_d <= xx_rsc_5_0_i_qa_d;
  xx_rsc_5_0_i_wea_d <= hybrid_core_inst_xx_rsc_5_0_i_wea_d;
  xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_6_0_i_adra_d <= hybrid_core_inst_xx_rsc_6_0_i_adra_d;
  hybrid_core_inst_xx_rsc_6_0_i_qa_d <= xx_rsc_6_0_i_qa_d;
  xx_rsc_6_0_i_wea_d <= hybrid_core_inst_xx_rsc_6_0_i_wea_d;
  xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_7_0_i_adra_d <= hybrid_core_inst_xx_rsc_7_0_i_adra_d;
  hybrid_core_inst_xx_rsc_7_0_i_qa_d <= xx_rsc_7_0_i_qa_d;
  xx_rsc_7_0_i_wea_d <= hybrid_core_inst_xx_rsc_7_0_i_wea_d;
  xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_8_0_i_adra_d <= hybrid_core_inst_xx_rsc_8_0_i_adra_d;
  hybrid_core_inst_xx_rsc_8_0_i_qa_d <= xx_rsc_8_0_i_qa_d;
  xx_rsc_8_0_i_wea_d <= hybrid_core_inst_xx_rsc_8_0_i_wea_d;
  xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_9_0_i_adra_d <= hybrid_core_inst_xx_rsc_9_0_i_adra_d;
  hybrid_core_inst_xx_rsc_9_0_i_qa_d <= xx_rsc_9_0_i_qa_d;
  xx_rsc_9_0_i_wea_d <= hybrid_core_inst_xx_rsc_9_0_i_wea_d;
  xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_10_0_i_adra_d <= hybrid_core_inst_xx_rsc_10_0_i_adra_d;
  hybrid_core_inst_xx_rsc_10_0_i_qa_d <= xx_rsc_10_0_i_qa_d;
  xx_rsc_10_0_i_wea_d <= hybrid_core_inst_xx_rsc_10_0_i_wea_d;
  xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_11_0_i_adra_d <= hybrid_core_inst_xx_rsc_11_0_i_adra_d;
  hybrid_core_inst_xx_rsc_11_0_i_qa_d <= xx_rsc_11_0_i_qa_d;
  xx_rsc_11_0_i_wea_d <= hybrid_core_inst_xx_rsc_11_0_i_wea_d;
  xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_12_0_i_adra_d <= hybrid_core_inst_xx_rsc_12_0_i_adra_d;
  hybrid_core_inst_xx_rsc_12_0_i_qa_d <= xx_rsc_12_0_i_qa_d;
  xx_rsc_12_0_i_wea_d <= hybrid_core_inst_xx_rsc_12_0_i_wea_d;
  xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_13_0_i_adra_d <= hybrid_core_inst_xx_rsc_13_0_i_adra_d;
  hybrid_core_inst_xx_rsc_13_0_i_qa_d <= xx_rsc_13_0_i_qa_d;
  xx_rsc_13_0_i_wea_d <= hybrid_core_inst_xx_rsc_13_0_i_wea_d;
  xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_14_0_i_adra_d <= hybrid_core_inst_xx_rsc_14_0_i_adra_d;
  hybrid_core_inst_xx_rsc_14_0_i_qa_d <= xx_rsc_14_0_i_qa_d;
  xx_rsc_14_0_i_wea_d <= hybrid_core_inst_xx_rsc_14_0_i_wea_d;
  xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_15_0_i_adra_d <= hybrid_core_inst_xx_rsc_15_0_i_adra_d;
  hybrid_core_inst_xx_rsc_15_0_i_qa_d <= xx_rsc_15_0_i_qa_d;
  xx_rsc_15_0_i_wea_d <= hybrid_core_inst_xx_rsc_15_0_i_wea_d;
  xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_16_0_i_adra_d <= hybrid_core_inst_xx_rsc_16_0_i_adra_d;
  hybrid_core_inst_xx_rsc_16_0_i_qa_d <= xx_rsc_16_0_i_qa_d;
  xx_rsc_16_0_i_wea_d <= hybrid_core_inst_xx_rsc_16_0_i_wea_d;
  xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_17_0_i_adra_d <= hybrid_core_inst_xx_rsc_17_0_i_adra_d;
  hybrid_core_inst_xx_rsc_17_0_i_qa_d <= xx_rsc_17_0_i_qa_d;
  xx_rsc_17_0_i_wea_d <= hybrid_core_inst_xx_rsc_17_0_i_wea_d;
  xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_18_0_i_adra_d <= hybrid_core_inst_xx_rsc_18_0_i_adra_d;
  hybrid_core_inst_xx_rsc_18_0_i_qa_d <= xx_rsc_18_0_i_qa_d;
  xx_rsc_18_0_i_wea_d <= hybrid_core_inst_xx_rsc_18_0_i_wea_d;
  xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_19_0_i_adra_d <= hybrid_core_inst_xx_rsc_19_0_i_adra_d;
  hybrid_core_inst_xx_rsc_19_0_i_qa_d <= xx_rsc_19_0_i_qa_d;
  xx_rsc_19_0_i_wea_d <= hybrid_core_inst_xx_rsc_19_0_i_wea_d;
  xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_20_0_i_adra_d <= hybrid_core_inst_xx_rsc_20_0_i_adra_d;
  hybrid_core_inst_xx_rsc_20_0_i_qa_d <= xx_rsc_20_0_i_qa_d;
  xx_rsc_20_0_i_wea_d <= hybrid_core_inst_xx_rsc_20_0_i_wea_d;
  xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_21_0_i_adra_d <= hybrid_core_inst_xx_rsc_21_0_i_adra_d;
  hybrid_core_inst_xx_rsc_21_0_i_qa_d <= xx_rsc_21_0_i_qa_d;
  xx_rsc_21_0_i_wea_d <= hybrid_core_inst_xx_rsc_21_0_i_wea_d;
  xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_22_0_i_adra_d <= hybrid_core_inst_xx_rsc_22_0_i_adra_d;
  hybrid_core_inst_xx_rsc_22_0_i_qa_d <= xx_rsc_22_0_i_qa_d;
  xx_rsc_22_0_i_wea_d <= hybrid_core_inst_xx_rsc_22_0_i_wea_d;
  xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_23_0_i_adra_d <= hybrid_core_inst_xx_rsc_23_0_i_adra_d;
  hybrid_core_inst_xx_rsc_23_0_i_qa_d <= xx_rsc_23_0_i_qa_d;
  xx_rsc_23_0_i_wea_d <= hybrid_core_inst_xx_rsc_23_0_i_wea_d;
  xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_24_0_i_adra_d <= hybrid_core_inst_xx_rsc_24_0_i_adra_d;
  hybrid_core_inst_xx_rsc_24_0_i_qa_d <= xx_rsc_24_0_i_qa_d;
  xx_rsc_24_0_i_wea_d <= hybrid_core_inst_xx_rsc_24_0_i_wea_d;
  xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_25_0_i_adra_d <= hybrid_core_inst_xx_rsc_25_0_i_adra_d;
  hybrid_core_inst_xx_rsc_25_0_i_qa_d <= xx_rsc_25_0_i_qa_d;
  xx_rsc_25_0_i_wea_d <= hybrid_core_inst_xx_rsc_25_0_i_wea_d;
  xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_26_0_i_adra_d <= hybrid_core_inst_xx_rsc_26_0_i_adra_d;
  hybrid_core_inst_xx_rsc_26_0_i_qa_d <= xx_rsc_26_0_i_qa_d;
  xx_rsc_26_0_i_wea_d <= hybrid_core_inst_xx_rsc_26_0_i_wea_d;
  xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_27_0_i_adra_d <= hybrid_core_inst_xx_rsc_27_0_i_adra_d;
  hybrid_core_inst_xx_rsc_27_0_i_qa_d <= xx_rsc_27_0_i_qa_d;
  xx_rsc_27_0_i_wea_d <= hybrid_core_inst_xx_rsc_27_0_i_wea_d;
  xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_28_0_i_adra_d <= hybrid_core_inst_xx_rsc_28_0_i_adra_d;
  hybrid_core_inst_xx_rsc_28_0_i_qa_d <= xx_rsc_28_0_i_qa_d;
  xx_rsc_28_0_i_wea_d <= hybrid_core_inst_xx_rsc_28_0_i_wea_d;
  xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_29_0_i_adra_d <= hybrid_core_inst_xx_rsc_29_0_i_adra_d;
  hybrid_core_inst_xx_rsc_29_0_i_qa_d <= xx_rsc_29_0_i_qa_d;
  xx_rsc_29_0_i_wea_d <= hybrid_core_inst_xx_rsc_29_0_i_wea_d;
  xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_30_0_i_adra_d <= hybrid_core_inst_xx_rsc_30_0_i_adra_d;
  hybrid_core_inst_xx_rsc_30_0_i_qa_d <= xx_rsc_30_0_i_qa_d;
  xx_rsc_30_0_i_wea_d <= hybrid_core_inst_xx_rsc_30_0_i_wea_d;
  xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  xx_rsc_31_0_i_adra_d <= hybrid_core_inst_xx_rsc_31_0_i_adra_d;
  hybrid_core_inst_xx_rsc_31_0_i_qa_d <= xx_rsc_31_0_i_qa_d;
  xx_rsc_31_0_i_wea_d <= hybrid_core_inst_xx_rsc_31_0_i_wea_d;
  xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_xx_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_xx_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_0_0_i_adra_d <= hybrid_core_inst_yy_rsc_0_0_i_adra_d;
  hybrid_core_inst_yy_rsc_0_0_i_qa_d <= yy_rsc_0_0_i_qa_d;
  yy_rsc_0_0_i_wea_d <= hybrid_core_inst_yy_rsc_0_0_i_wea_d;
  yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_0_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_1_0_i_adra_d <= hybrid_core_inst_yy_rsc_1_0_i_adra_d;
  hybrid_core_inst_yy_rsc_1_0_i_qa_d <= yy_rsc_1_0_i_qa_d;
  yy_rsc_1_0_i_wea_d <= hybrid_core_inst_yy_rsc_1_0_i_wea_d;
  yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_1_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_2_0_i_adra_d <= hybrid_core_inst_yy_rsc_2_0_i_adra_d;
  hybrid_core_inst_yy_rsc_2_0_i_qa_d <= yy_rsc_2_0_i_qa_d;
  yy_rsc_2_0_i_wea_d <= hybrid_core_inst_yy_rsc_2_0_i_wea_d;
  yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_2_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_2_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_3_0_i_adra_d <= hybrid_core_inst_yy_rsc_3_0_i_adra_d;
  hybrid_core_inst_yy_rsc_3_0_i_qa_d <= yy_rsc_3_0_i_qa_d;
  yy_rsc_3_0_i_wea_d <= hybrid_core_inst_yy_rsc_3_0_i_wea_d;
  yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_3_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_3_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_4_0_i_adra_d <= hybrid_core_inst_yy_rsc_4_0_i_adra_d;
  hybrid_core_inst_yy_rsc_4_0_i_qa_d <= yy_rsc_4_0_i_qa_d;
  yy_rsc_4_0_i_wea_d <= hybrid_core_inst_yy_rsc_4_0_i_wea_d;
  yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_4_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_4_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_5_0_i_adra_d <= hybrid_core_inst_yy_rsc_5_0_i_adra_d;
  hybrid_core_inst_yy_rsc_5_0_i_qa_d <= yy_rsc_5_0_i_qa_d;
  yy_rsc_5_0_i_wea_d <= hybrid_core_inst_yy_rsc_5_0_i_wea_d;
  yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_5_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_5_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_6_0_i_adra_d <= hybrid_core_inst_yy_rsc_6_0_i_adra_d;
  hybrid_core_inst_yy_rsc_6_0_i_qa_d <= yy_rsc_6_0_i_qa_d;
  yy_rsc_6_0_i_wea_d <= hybrid_core_inst_yy_rsc_6_0_i_wea_d;
  yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_6_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_6_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_7_0_i_adra_d <= hybrid_core_inst_yy_rsc_7_0_i_adra_d;
  hybrid_core_inst_yy_rsc_7_0_i_qa_d <= yy_rsc_7_0_i_qa_d;
  yy_rsc_7_0_i_wea_d <= hybrid_core_inst_yy_rsc_7_0_i_wea_d;
  yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_7_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_7_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_8_0_i_adra_d <= hybrid_core_inst_yy_rsc_8_0_i_adra_d;
  hybrid_core_inst_yy_rsc_8_0_i_qa_d <= yy_rsc_8_0_i_qa_d;
  yy_rsc_8_0_i_wea_d <= hybrid_core_inst_yy_rsc_8_0_i_wea_d;
  yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_8_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_8_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_9_0_i_adra_d <= hybrid_core_inst_yy_rsc_9_0_i_adra_d;
  hybrid_core_inst_yy_rsc_9_0_i_qa_d <= yy_rsc_9_0_i_qa_d;
  yy_rsc_9_0_i_wea_d <= hybrid_core_inst_yy_rsc_9_0_i_wea_d;
  yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_9_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_9_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_10_0_i_adra_d <= hybrid_core_inst_yy_rsc_10_0_i_adra_d;
  hybrid_core_inst_yy_rsc_10_0_i_qa_d <= yy_rsc_10_0_i_qa_d;
  yy_rsc_10_0_i_wea_d <= hybrid_core_inst_yy_rsc_10_0_i_wea_d;
  yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_10_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_10_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_11_0_i_adra_d <= hybrid_core_inst_yy_rsc_11_0_i_adra_d;
  hybrid_core_inst_yy_rsc_11_0_i_qa_d <= yy_rsc_11_0_i_qa_d;
  yy_rsc_11_0_i_wea_d <= hybrid_core_inst_yy_rsc_11_0_i_wea_d;
  yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_11_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_11_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_12_0_i_adra_d <= hybrid_core_inst_yy_rsc_12_0_i_adra_d;
  hybrid_core_inst_yy_rsc_12_0_i_qa_d <= yy_rsc_12_0_i_qa_d;
  yy_rsc_12_0_i_wea_d <= hybrid_core_inst_yy_rsc_12_0_i_wea_d;
  yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_12_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_12_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_13_0_i_adra_d <= hybrid_core_inst_yy_rsc_13_0_i_adra_d;
  hybrid_core_inst_yy_rsc_13_0_i_qa_d <= yy_rsc_13_0_i_qa_d;
  yy_rsc_13_0_i_wea_d <= hybrid_core_inst_yy_rsc_13_0_i_wea_d;
  yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_13_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_13_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_14_0_i_adra_d <= hybrid_core_inst_yy_rsc_14_0_i_adra_d;
  hybrid_core_inst_yy_rsc_14_0_i_qa_d <= yy_rsc_14_0_i_qa_d;
  yy_rsc_14_0_i_wea_d <= hybrid_core_inst_yy_rsc_14_0_i_wea_d;
  yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_14_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_14_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_15_0_i_adra_d <= hybrid_core_inst_yy_rsc_15_0_i_adra_d;
  hybrid_core_inst_yy_rsc_15_0_i_qa_d <= yy_rsc_15_0_i_qa_d;
  yy_rsc_15_0_i_wea_d <= hybrid_core_inst_yy_rsc_15_0_i_wea_d;
  yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_15_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_15_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_16_0_i_adra_d <= hybrid_core_inst_yy_rsc_16_0_i_adra_d;
  hybrid_core_inst_yy_rsc_16_0_i_qa_d <= yy_rsc_16_0_i_qa_d;
  yy_rsc_16_0_i_wea_d <= hybrid_core_inst_yy_rsc_16_0_i_wea_d;
  yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_16_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_16_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_17_0_i_adra_d <= hybrid_core_inst_yy_rsc_17_0_i_adra_d;
  hybrid_core_inst_yy_rsc_17_0_i_qa_d <= yy_rsc_17_0_i_qa_d;
  yy_rsc_17_0_i_wea_d <= hybrid_core_inst_yy_rsc_17_0_i_wea_d;
  yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_17_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_17_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_18_0_i_adra_d <= hybrid_core_inst_yy_rsc_18_0_i_adra_d;
  hybrid_core_inst_yy_rsc_18_0_i_qa_d <= yy_rsc_18_0_i_qa_d;
  yy_rsc_18_0_i_wea_d <= hybrid_core_inst_yy_rsc_18_0_i_wea_d;
  yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_18_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_18_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_19_0_i_adra_d <= hybrid_core_inst_yy_rsc_19_0_i_adra_d;
  hybrid_core_inst_yy_rsc_19_0_i_qa_d <= yy_rsc_19_0_i_qa_d;
  yy_rsc_19_0_i_wea_d <= hybrid_core_inst_yy_rsc_19_0_i_wea_d;
  yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_19_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_19_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_20_0_i_adra_d <= hybrid_core_inst_yy_rsc_20_0_i_adra_d;
  hybrid_core_inst_yy_rsc_20_0_i_qa_d <= yy_rsc_20_0_i_qa_d;
  yy_rsc_20_0_i_wea_d <= hybrid_core_inst_yy_rsc_20_0_i_wea_d;
  yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_20_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_20_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_21_0_i_adra_d <= hybrid_core_inst_yy_rsc_21_0_i_adra_d;
  hybrid_core_inst_yy_rsc_21_0_i_qa_d <= yy_rsc_21_0_i_qa_d;
  yy_rsc_21_0_i_wea_d <= hybrid_core_inst_yy_rsc_21_0_i_wea_d;
  yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_21_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_21_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_22_0_i_adra_d <= hybrid_core_inst_yy_rsc_22_0_i_adra_d;
  hybrid_core_inst_yy_rsc_22_0_i_qa_d <= yy_rsc_22_0_i_qa_d;
  yy_rsc_22_0_i_wea_d <= hybrid_core_inst_yy_rsc_22_0_i_wea_d;
  yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_22_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_22_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_23_0_i_adra_d <= hybrid_core_inst_yy_rsc_23_0_i_adra_d;
  hybrid_core_inst_yy_rsc_23_0_i_qa_d <= yy_rsc_23_0_i_qa_d;
  yy_rsc_23_0_i_wea_d <= hybrid_core_inst_yy_rsc_23_0_i_wea_d;
  yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_23_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_23_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_24_0_i_adra_d <= hybrid_core_inst_yy_rsc_24_0_i_adra_d;
  hybrid_core_inst_yy_rsc_24_0_i_qa_d <= yy_rsc_24_0_i_qa_d;
  yy_rsc_24_0_i_wea_d <= hybrid_core_inst_yy_rsc_24_0_i_wea_d;
  yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_24_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_24_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_25_0_i_adra_d <= hybrid_core_inst_yy_rsc_25_0_i_adra_d;
  hybrid_core_inst_yy_rsc_25_0_i_qa_d <= yy_rsc_25_0_i_qa_d;
  yy_rsc_25_0_i_wea_d <= hybrid_core_inst_yy_rsc_25_0_i_wea_d;
  yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_25_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_25_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_26_0_i_adra_d <= hybrid_core_inst_yy_rsc_26_0_i_adra_d;
  hybrid_core_inst_yy_rsc_26_0_i_qa_d <= yy_rsc_26_0_i_qa_d;
  yy_rsc_26_0_i_wea_d <= hybrid_core_inst_yy_rsc_26_0_i_wea_d;
  yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_26_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_26_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_27_0_i_adra_d <= hybrid_core_inst_yy_rsc_27_0_i_adra_d;
  hybrid_core_inst_yy_rsc_27_0_i_qa_d <= yy_rsc_27_0_i_qa_d;
  yy_rsc_27_0_i_wea_d <= hybrid_core_inst_yy_rsc_27_0_i_wea_d;
  yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_27_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_27_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_28_0_i_adra_d <= hybrid_core_inst_yy_rsc_28_0_i_adra_d;
  hybrid_core_inst_yy_rsc_28_0_i_qa_d <= yy_rsc_28_0_i_qa_d;
  yy_rsc_28_0_i_wea_d <= hybrid_core_inst_yy_rsc_28_0_i_wea_d;
  yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_28_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_28_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_29_0_i_adra_d <= hybrid_core_inst_yy_rsc_29_0_i_adra_d;
  hybrid_core_inst_yy_rsc_29_0_i_qa_d <= yy_rsc_29_0_i_qa_d;
  yy_rsc_29_0_i_wea_d <= hybrid_core_inst_yy_rsc_29_0_i_wea_d;
  yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_29_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_29_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_30_0_i_adra_d <= hybrid_core_inst_yy_rsc_30_0_i_adra_d;
  hybrid_core_inst_yy_rsc_30_0_i_qa_d <= yy_rsc_30_0_i_qa_d;
  yy_rsc_30_0_i_wea_d <= hybrid_core_inst_yy_rsc_30_0_i_wea_d;
  yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_30_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_30_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  yy_rsc_31_0_i_adra_d <= hybrid_core_inst_yy_rsc_31_0_i_adra_d;
  hybrid_core_inst_yy_rsc_31_0_i_qa_d <= yy_rsc_31_0_i_qa_d;
  yy_rsc_31_0_i_wea_d <= hybrid_core_inst_yy_rsc_31_0_i_wea_d;
  yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= hybrid_core_inst_yy_rsc_31_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d <= hybrid_core_inst_yy_rsc_31_0_i_rwA_rw_ram_ir_internal_WMASK_B_d;
  S34_OUTER_LOOP_for_tf_mul_cmp_a <= hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_a;
  S34_OUTER_LOOP_for_tf_mul_cmp_b <= hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_b;
  hybrid_core_inst_S34_OUTER_LOOP_for_tf_mul_cmp_z <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'(
      UNSIGNED(S34_OUTER_LOOP_for_tf_mul_cmp_a) * UNSIGNED(S34_OUTER_LOOP_for_tf_mul_cmp_b)),
      10));
  xx_rsc_0_0_i_da_d_iff <= hybrid_core_inst_xx_rsc_0_0_i_da_d_pff;
  xx_rsc_1_0_i_da_d_iff <= hybrid_core_inst_xx_rsc_1_0_i_da_d_pff;
  xx_rsc_2_0_i_da_d_iff <= hybrid_core_inst_xx_rsc_2_0_i_da_d_pff;
  xx_rsc_3_0_i_da_d_iff <= hybrid_core_inst_xx_rsc_3_0_i_da_d_pff;
  yy_rsc_0_0_i_da_d_iff <= hybrid_core_inst_yy_rsc_0_0_i_da_d_pff;
  yy_rsc_1_0_i_da_d_iff <= hybrid_core_inst_yy_rsc_1_0_i_da_d_pff;
  yy_rsc_2_0_i_da_d_iff <= hybrid_core_inst_yy_rsc_2_0_i_da_d_pff;
  yy_rsc_3_0_i_da_d_iff <= hybrid_core_inst_yy_rsc_3_0_i_da_d_pff;

END v14;



