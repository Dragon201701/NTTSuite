// check_properties -prop -list spec.prop_ovf_spec_wrapper_ln65_1 ; # ( ovf ) (l1=1, l2=0)
module GOTH_58 ( M1TU__P_18_14 , M1TU__P_36_15 , M1TU__clk , M1TU__asm_sym_data_21
 , M1TU__asm_sym_data_17 , M1TU__OOB_X_1 , M1TU__asm_sym_data_16 , M1TU__OOB_X_2
 , M1TU__asm_sym_data_11 , M1TU__asm_sym_data_8 , M1TU__asm_sym_data_9 , M1TU__asm_sym_data_10
 , M1TU__OOB_X_3 , M1TU__asm_sym_data_3 , M1TU__asm_sym_data_0 , M1TU__asm_sym_data_1
 , M1TU__asm_sym_data_2 , M1TU__OOB_X_4 , M1TU__P_56 , M1TU__OOB_X_6 , M1TU__asm_sym_data_20
 , M1TU__OOB_X_7 , M1TU__OOB_X_8 , M1TU__OOB_X_9 ) ;
 input wire  M1TU__clk ; 
 input wire  [31:0]  M1TU__asm_sym_data_21 ; 
 input wire  [31:0]  M1TU__asm_sym_data_17 ; 
 input wire  [31:0]  M1TU__OOB_X_1 ; 
 input wire  [31:0]  M1TU__asm_sym_data_16 ; 
 input wire  [31:0]  M1TU__OOB_X_2 ; 
 input wire  [31:0]  M1TU__asm_sym_data_11 ; 
 input wire  [31:0]  M1TU__asm_sym_data_8 ; 
 input wire  [31:0]  M1TU__asm_sym_data_9 ; 
 input wire  [31:0]  M1TU__asm_sym_data_10 ; 
 input wire  [31:0]  M1TU__OOB_X_3 ; 
 input wire  [31:0]  M1TU__asm_sym_data_3 ; 
 input wire  [31:0]  M1TU__asm_sym_data_0 ; 
 input wire  [31:0]  M1TU__asm_sym_data_1 ; 
 input wire  [31:0]  M1TU__asm_sym_data_2 ; 
 input wire  [31:0]  M1TU__OOB_X_4 ; 
 input wire  [31:0]  M1TU__P_56 ; 
 input wire  [31:0]  M1TU__OOB_X_6 ; 
 input wire  [31:0]  M1TU__asm_sym_data_20 ; 
 input wire  [31:0]  M1TU__OOB_X_7 ; 
 input wire  [31:0]  M1TU__OOB_X_8 ; 
 input wire  [31:0]  M1TU__OOB_X_9 ; 
 output wire  M1TU__P_18_14 ; 
 output wire  [0:0]  M1TU__P_36_15 ; 
 wire  [0:0] E_48092 ; 
assign M1TU__P_36_15 = E_48092 ;
 wire  [0:0] E_48220 ; 
assign M1TU__P_18_14 = E_48220 ;
 wire  [0:0] E_47863 ; 
 wire  [0:0] E_47862 ; 
 wire  [0:0] E_47861 ; 
 wire  [32:0] E_48018 ; 
 wire  [31:0] E_48055 ; 
 wire  [0:0] E_48412 ; 
 wire  [19:0] E_51353 ; 
 wire  [19:0] E_48053 ; 
 wire  [18:0] E_48052 ; 
 wire  [19:0] E_48016 ; 
 wire  [0:0] E_48170 ; 
 wire  [0:0] E_48169 ; 
 wire  [0:0] E_48168 ; 
 wire  [19:0] E_48167 ; 
 wire  [19:0] E_48068 ; 
 wire  [0:0] E_48165 ; 
 wire  [0:0] E_48164 ; 
 wire  [2:0] E_48189 ; 
 wire  [2:0] E_48205 ; 
 wire  [0:0] E_48203 ; 
 wire  [0:0] E_48202 ; 
 wire  [0:0] E_48201 ; 
 wire  [0:0] E_48200 ; 
 wire  [0:0] E_48199 ; 
 wire  [19:0] E_48198 ; 
 wire  [19:0] E_48197 ; 
 wire  [0:0] E_48196 ; 
 wire  [0:0] E_48195 ; 
 wire  [0:0] E_48194 ; 
 wire  [19:0] E_48193 ; 
 wire  [19:0] E_47976 ; 
 wire  [0:0] E_48191 ; 
 wire  [0:0] E_48190 ; 
 wire  [2:0] E_48188 ; 
 wire  [0:0] E_48187 ; 
 wire  [0:0] E_48186 ; 
 wire  [0:0] E_48185 ; 
 wire  [0:0] E_48184 ; 
 wire  [19:0] E_48183 ; 
 wire  signed  [20:0] E_48036 ; 
 wire  [19:0] E_48182 ; 
 wire  [0:0] E_48181 ; 
 wire  [0:0] E_48115 ; 
 wire  [19:0] E_48179 ; 
 wire  [19:0] E_48206 ; 
 wire  [19:0] E_48141 ; 
 wire  [0:0] E_48175 ; 
 wire  [0:0] E_48174 ; 
 wire  [0:0] E_48173 ; 
 wire  [19:0] E_48172 ; 
 wire  [9:0] E_48075 ; 
 wire  [0:0] E_48156 ; 
 wire  [0:0] E_48155 ; 
 wire  [1:0] E_47804 ; 
 wire  [19:0] E_48142 ; 
 wire  signed  [20:0] E_47957 ; 
 wire  [1:0] E_47806 ; 
 wire clk ; 
assign clk = M1TU__clk ;
 wire  [19:0] E_48253 ; 
 wire  [19:0] E_48178_68655 ; 
 wire  [3:0] E_48178 ; 
 wire  [2:0] E_48176 ; 
 wire  [0:0] E_48152 ; 
 wire  [19:0] E_48151 ; 
 wire  [19:0] E_48209 ; 
 wire  [0:0] E_48150 ; 
 wire  [0:0] E_48149 ; 
 wire  [2:0] E_48148 ; 
 wire  [19:0] E_48256 ; 
 wire  [19:0] E_48092_68651 ; 
 wire  [19:0] E_48147 ; 
 wire  [19:0] E_48210 ; 
 wire  [0:0] E_48146 ; 
 wire  [0:0] E_48145 ; 
 wire  [19:0] E_48257 ; 
 wire  [0:0] E_48144 ; 
 wire  [0:0] E_48143 ; 
 wire  [0:0] E_48140 ; 
 wire  [0:0] E_48139 ; 
 wire  [2:0] E_47813 ; 
 wire  [2:0] E_47812 ; 
 wire  [2:0] E_47811 ; 
 wire  [2:0] E_47810 ; 
 wire  [0:0] E_48159 ; 
 wire  [0:0] E_48158 ; 
 wire  [2:0] E_47809 ; 
 wire  [0:0] E_48136 ; 
 wire  [2:0] E_48115_68642 ; 
 wire  [2:0] E_47807 ; 
 wire  [2:0] E_47806_68640 ; 
 wire  [2:0] E_47805 ; 
 wire  [2:0] E_47804_68639 ; 
 wire  [2:0] E_47803 ; 
 wire  [2:0] E_48163 ; 
 wire  [2:0] E_47802 ; 
 wire  [2:0] E_47801 ; 
 wire  [2:0] E_47800 ; 
 wire  [2:0] E_60005 ; 
 wire  [19:0] E_48162 ; 
 wire  [19:0] E_48207 ; 
 wire  [19:0] E_48254 ; 
 wire  [19:0] E_48157 ; 
 wire  [19:0] E_48208 ; 
 wire  [19:0] E_48255 ; 
 wire  [9:0] E_51065 ; 
 wire  [31:0] E_48055_clone_48407 ; 
 wire  [31:0] asm_sym_data_21 ; 
assign asm_sym_data_21 = M1TU__asm_sym_data_21 ;
 wire  [31:0] E_49059 ; 
 wire  [0:0] E_49046 ; 
 wire  [20:0] E_48076 ; 
 wire  [31:0] E_49057 ; 
 wire  [0:0] E_51058 ; 
 wire  [31:0] E_48073 ; 
 wire  [0:0] E_48072 ; 
 wire  [31:0] E_48071 ; 
 wire  [31:0] E_48120 ; 
 wire  [0:0] E_48347 ; 
 wire  [19:0] E_51359 ; 
 wire  [19:0] E_48117 ; 
 wire  [18:0] E_48116 ; 
 wire  [31:0] E_48120_clone_48342 ; 
assign E_48120_clone_48342 = M1TU__asm_sym_data_17 ;
 wire  [31:0] OOB_X_1 ; 
assign OOB_X_1 = M1TU__OOB_X_1 ;
 wire  [31:0] E_48114 ; 
 wire  [0:0] E_48113 ; 
 wire  [31:0] E_48112 ; 
 wire  [31:0] E_48110 ; 
 wire  [31:0] E_48108 ; 
 wire  [31:0] E_48108_clone_48355 ; 
assign E_48108_clone_48355 = M1TU__asm_sym_data_16 ;
 wire  [31:0] OOB_X_2 ; 
assign OOB_X_2 = M1TU__OOB_X_2 ;
 wire  [31:0] E_48106 ; 
 wire  [0:0] E_48373 ; 
 wire  [19:0] E_51357 ; 
 wire  [19:0] E_48102 ; 
 wire  [19:0] E_48101 ; 
 wire  [19:0] E_48040 ; 
 wire  [19:0] E_48039 ; 
 wire  signed  [31:0] E_48038 ; 
 wire  [0:0] E_48037 ; 
 wire  [5:0] E_48096 ; 
 wire  signed  [31:0] E_48035_68647 ; 
 wire  [31:0] E_48035 ; 
 wire  signed  [0:0] E_48093 ; 
 wire  signed  [31:0] E_48092_68644 ; 
 wire  [19:0] E_48258 ; 
 wire  [19:0] E_48100 ; 
 wire  [0:0] E_48098 ; 
 wire  signed  [20:0] E_48097 ; 
 wire  [19:0] E_48095 ; 
 wire  [31:0] E_48106_clone_48368 ; 
 wire  [0:0] E_51002 ; 
 wire  [19:0] E_51351 ; 
 wire  [31:0] E_50825 ; 
 wire  [0:0] E_51018 ; 
 wire  [19:0] E_51345 ; 
 wire  [19:0] E_48001 ; 
 wire  [19:0] E_48000 ; 
 wire  [19:0] E_47961 ; 
 wire  [19:0] E_47960 ; 
 wire  signed  [31:0] E_47959 ; 
 wire  [0:0] E_47958 ; 
 wire  signed  [31:0] E_47956_68643 ; 
 wire  [31:0] E_47956 ; 
 wire  [19:0] E_48260 ; 
 wire  [19:0] E_47999 ; 
 wire  signed  [31:0] E_47998 ; 
 wire  [0:0] E_47997 ; 
 wire  signed  [20:0] E_47996 ; 
 wire  signed  [31:0] E_47995_68645 ; 
 wire  [31:0] E_47995 ; 
 wire  [31:0] E_50829 ; 
 wire  [0:0] E_51038 ; 
 wire  [19:0] E_51339 ; 
 wire  [31:0] asm_sym_data_11 ; 
assign asm_sym_data_11 = M1TU__asm_sym_data_11 ;
 wire  [31:0] asm_sym_data_8 ; 
assign asm_sym_data_8 = M1TU__asm_sym_data_8 ;
 wire  [31:0] E_50905 ; 
 wire  [0:0] E_51014 ; 
 wire  [31:0] asm_sym_data_9 ; 
assign asm_sym_data_9 = M1TU__asm_sym_data_9 ;
 wire  [31:0] E_50865 ; 
 wire  [0:0] E_50994 ; 
 wire  [31:0] E_50869 ; 
 wire  [0:0] E_50998 ; 
 wire  [31:0] asm_sym_data_10 ; 
assign asm_sym_data_10 = M1TU__asm_sym_data_10 ;
 wire  [31:0] OOB_X_3 ; 
assign OOB_X_3 = M1TU__OOB_X_3 ;
 wire  [31:0] E_48091 ; 
 wire  [31:0] E_48089 ; 
 wire  [51:0] E_48087 ; 
 wire  [31:0] E_48086 ; 
 wire  [31:0] E_48086_clone_48381 ; 
 wire  [31:0] E_51037 ; 
 wire  [31:0] E_51041 ; 
 wire  [31:0] asm_sym_data_3 ; 
assign asm_sym_data_3 = M1TU__asm_sym_data_3 ;
 wire  [31:0] E_47949_clone_48524 ; 
assign E_47949_clone_48524 = M1TU__asm_sym_data_0 ;
 wire  [31:0] E_51053 ; 
 wire  [31:0] asm_sym_data_1 ; 
assign asm_sym_data_1 = M1TU__asm_sym_data_1 ;
 wire  [31:0] E_48028_clone_48446 ; 
 wire  [31:0] E_51049 ; 
 wire  [31:0] asm_sym_data_2 ; 
assign asm_sym_data_2 = M1TU__asm_sym_data_2 ;
 wire  [31:0] OOB_X_4 ; 
assign OOB_X_4 = M1TU__OOB_X_4 ;
 wire  [4:0] E_48084 ; 
 wire  [31:0] E_48083 ; 
 wire  [31:0] E_48082 ; 
 wire  [31:0] E_48259 ; 
 wire  [31:0] E_48081 ; 
assign E_48081 = M1TU__P_56 ;
 wire  [31:0] E_48080 ; 
 wire  signed  [32:0] E_48079 ; 
 wire  [31:0] E_48069 ; 
 wire  [31:0] E_48124 ; 
 wire  [0:0] E_48123 ; 
 wire  signed  [31:0] E_48122 ; 
 wire  [31:0] E_48122_68652 ; 
 wire  [31:0] E_48077 ; 
 wire  [31:0] OOB_X_6 ; 
assign OOB_X_6 = M1TU__OOB_X_6 ;
 wire  [31:0] E_48051 ; 
 wire  [0:0] E_48050 ; 
 wire  [31:0] E_48049 ; 
 wire  signed  [32:0] E_48048 ; 
 wire  [31:0] E_48047 ; 
 wire  [63:0] E_48046 ; 
 wire  [31:0] E_48045 ; 
 wire  [31:0] E_48045_clone_48420 ; 
 wire  [31:0] asm_sym_data_20 ; 
assign asm_sym_data_20 = M1TU__asm_sym_data_20 ;
 wire  [31:0] E_49053 ; 
 wire  [0:0] E_49037 ; 
 wire  [31:0] E_49051 ; 
 wire  [0:0] E_51057 ; 
 wire  [31:0] OOB_X_7 ; 
assign OOB_X_7 = M1TU__OOB_X_7 ;
 wire  [31:0] E_48043 ; 
 wire  [0:0] E_48438 ; 
 wire  [31:0] E_48043_clone_48433 ; 
 wire  [31:0] E_50681 ; 
 wire  [31:0] E_47964_clone_48511 ; 
 wire  [31:0] E_50781 ; 
 wire  [31:0] E_48004_clone_48472 ; 
 wire  [31:0] E_50733 ; 
 wire  [31:0] OOB_X_8 ; 
assign OOB_X_8 = M1TU__OOB_X_8 ;
 wire  [31:0] E_48033 ; 
 wire  [63:0] E_48032 ; 
 wire  [31:0] E_48031 ; 
 wire  [43:0] E_48030 ; 
 wire  [63:0] E_48029 ; 
 wire  [31:0] E_48028 ; 
 wire  [31:0] OOB_X_9 ; 
assign OOB_X_9 = M1TU__OOB_X_9 ;
 wire  [31:0] E_48027 ; 
 wire  signed  [32:0] E_48026 ; 
 wire  [31:0] E_47937 ; 
 wire  [0:0] E_47860 ; 
  assign /* unsigned  1-bit */  E_48092 = 1'h0;
  assign /* unsigned  1-bit */  E_48220 = ( E_47863 ? E_48115 : E_47860 ) ;
  assign /* unsigned  1-bit */  E_47863 = (E_47862 && E_48156) ;
  assign /* unsigned  1-bit */  E_47862 = ( !E_47861 ) ;
  assign /* unsigned  1-bit */  E_47861 = (E_48018 <= E_47937) ;
  assign /* unsigned 33-bit */  E_48018 = (E_48055 + E_48051) ;
  assign /* unsigned 32-bit */  E_48055 = ( E_48412 ? OOB_X_6 : E_48055_clone_48407 ) ;
  assign /* unsigned  1-bit */  E_48412 = (E_51353 > E_51065) ;
  assign /* unsigned 20-bit */  E_51353 = (E_48053 + E_48115) ;
  assign /* unsigned 20-bit */  E_48053 = (E_48052 <<< E_48115) ;
  assign /* unsigned 19-bit */  E_48052 = ( E_48016 ) ;
  assign /* unsigned 20-bit */  E_48016 = ( E_48170 ? E_48092_68651 : E_48157 ) ;
  assign /* unsigned  1-bit */  E_48170 = (E_48169 && E_48159) ;
  assign /* unsigned  1-bit */  E_48169 = ( !E_48168 ) ;
  assign /* unsigned  1-bit */  E_48168 = (E_48167 < E_48075) ;
  assign /* unsigned 20-bit */  E_48167 = (E_48068 + E_48115) ;
  assign /* unsigned 20-bit */  E_48068 = ( E_48165 ? E_48092_68651 : E_48162 ) ;
  assign /* unsigned  1-bit */  E_48165 = (E_48164 || E_48181) ;
  assign /* unsigned  1-bit */  E_48164 = (E_48189 == E_48163) ;
  CPL_FF#3  I_48047_reg ( .q ( E_48189 )  , .qbar (  )  , .d ( E_48205 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_60005 )  );
  assign /* unsigned  3-bit */  E_48205 = ( E_48203 ? E_48115_68642 : E_47813 ) ;
  assign /* unsigned  1-bit */  E_48203 = (E_48202 || E_48140) ;
  assign /* unsigned  1-bit */  E_48202 = ( E_48201 ? E_48144 : E_48092 ) ;
  assign /* unsigned  1-bit */  E_48201 = (E_48200 && E_48146) ;
  assign /* unsigned  1-bit */  E_48200 = ( !E_48199 ) ;
  assign /* unsigned  1-bit */  E_48199 = (E_48198 < E_48075) ;
  assign /* unsigned 20-bit */  E_48198 = (E_48197 + E_48115) ;
  assign /* unsigned 20-bit */  E_48197 = ( E_48196 ? E_48092_68651 : E_48147 ) ;
  assign /* unsigned  1-bit */  E_48196 = (E_48195 && E_48150) ;
  assign /* unsigned  1-bit */  E_48195 = ( !E_48194 ) ;
  assign /* unsigned  1-bit */  E_48194 = (E_48193 < E_48075) ;
  assign /* unsigned 20-bit */  E_48193 = (E_47976 + E_48115) ;
  assign /* unsigned 20-bit */  E_47976 = ( E_48191 ? E_48092_68651 : E_48151 ) ;
  assign /* unsigned  1-bit */  E_48191 = (E_48190 || E_48187) ;
  assign /* unsigned  1-bit */  E_48190 = (E_48189 == E_48188) ;
  assign /* unsigned  3-bit */  E_48188 = 3'h7;
  assign /* unsigned  1-bit */  E_48187 = ( E_48186 ? E_48152 : E_48092 ) ;
  assign /* unsigned  1-bit */  E_48186 = (E_48185 && E_48175) ;
  assign /* unsigned  1-bit */  E_48185 = ( !E_48184 ) ;
  assign /* unsigned  1-bit */  E_48184 = (E_48183 >= E_48176) ;
  assign /* unsigned 20-bit */  E_48183 = ( E_48036 ) ;
  assign /*   signed 21-bit */  E_48036 = (E_48182 - E_47806) ;
  assign /* unsigned 20-bit */  E_48182 = ( E_48181 ? E_48178_68655 : E_48179 ) ;
wire  [2:0]  E_48115_89764 = { {2{1'b0}}, E_48115 }; /* zero-padding */ 
  assign /* unsigned  1-bit */  E_48181 = (E_48189 == E_48115_89764) ;
  assign /* unsigned  1-bit */  E_48115 = 1'h1;
  CPL_FF#20  I_48049_reg ( .q ( E_48179 )  , .qbar (  )  , .d ( E_48206 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48253 )  );
  assign /* unsigned 20-bit */  E_48206 = ( E_48201 ? E_48142 : E_48141 ) ;
  assign /* unsigned 20-bit */  E_48141 = ( E_48175 ? E_48183 : E_48182 ) ;
  assign /* unsigned  1-bit */  E_48175 = (E_48174 && E_48156) ;
  assign /* unsigned  1-bit */  E_48174 = ( !E_48173 ) ;
  assign /* unsigned  1-bit */  E_48173 = (E_48172 < E_48075) ;
  assign /* unsigned 20-bit */  E_48172 = (E_48016 + E_48115) ;
  assign /* unsigned 10-bit */  E_48075 = 10'h200;
  assign /* unsigned  1-bit */  E_48156 = (E_48155 || E_48170) ;
wire  [2:0]  E_47804_89765 = { {1{1'b0}}, E_47804 }; /* zero-padding */ 
  assign /* unsigned  1-bit */  E_48155 = (E_48189 == E_47804_89765) ;
  assign /* unsigned  2-bit */  E_47804 = 2'h3;
  assign /* unsigned 20-bit */  E_48142 = ( E_47957 ) ;
  assign /*   signed 21-bit */  E_47957 = (E_48141 - E_47806) ;
  assign /* unsigned  2-bit */  E_47806 = 2'h2;
  assign /* unsigned 20-bit */  E_48253 = 20'hX; /*CDBImplicitXNone*/
  assign /* unsigned 20-bit */  E_48178_68655 = ( E_48178 ) ;
  assign /* unsigned  4-bit */  E_48178 = 4'ha;
  assign /* unsigned  3-bit */  E_48176 = 3'h6;
  assign /* unsigned  1-bit */  E_48152 = (E_48183 >= E_47806) ;
  CPL_FF#20  I_48054_reg ( .q ( E_48151 )  , .qbar (  )  , .d ( E_48209 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48256 )  );
  assign /* unsigned 20-bit */  E_48209 = ( E_48150 ? E_48193 : E_47976 ) ;
  assign /* unsigned  1-bit */  E_48150 = (E_48149 || E_48191) ;
  assign /* unsigned  1-bit */  E_48149 = (E_48189 == E_48148) ;
  assign /* unsigned  3-bit */  E_48148 = 3'h5;
  assign /* unsigned 20-bit */  E_48256 = 20'hX; /*CDBImplicitXNone*/
  assign /* unsigned 20-bit */  E_48092_68651 = ( E_48092 ) ;
  CPL_FF#20  I_48056_reg ( .q ( E_48147 )  , .qbar (  )  , .d ( E_48210 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48257 )  );
  assign /* unsigned 20-bit */  E_48210 = ( E_48146 ? E_48198 : E_48197 ) ;
  assign /* unsigned  1-bit */  E_48146 = (E_48145 || E_48196) ;
  assign /* unsigned  1-bit */  E_48145 = (E_48189 == E_48176) ;
  assign /* unsigned 20-bit */  E_48257 = 20'hX; /*CDBImplicitXNone*/
  assign /* unsigned  1-bit */  E_48144 = ( !E_48143 ) ;
  assign /* unsigned  1-bit */  E_48143 = (E_48142 >= E_47806) ;
  assign /* unsigned  1-bit */  E_48140 = ( E_48186 ? E_48139 : E_48092 ) ;
  assign /* unsigned  1-bit */  E_48139 = ( !E_48152 ) ;
  assign /* unsigned  3-bit */  E_47813 = ( E_48146 ? E_47801 : E_47812 ) ;
  assign /* unsigned  3-bit */  E_47812 = ( E_48150 ? E_47802 : E_47811 ) ;
  assign /* unsigned  3-bit */  E_47811 = ( E_48156 ? E_47805 : E_47810 ) ;
  assign /* unsigned  3-bit */  E_47810 = ( E_48159 ? E_47807 : E_47809 ) ;
  assign /* unsigned  1-bit */  E_48159 = (E_48158 || E_48165) ;
wire  [2:0]  E_47806_89766 = { {1{1'b0}}, E_47806 }; /* zero-padding */ 
  assign /* unsigned  1-bit */  E_48158 = (E_48189 == E_47806_89766) ;
  assign /* unsigned  3-bit */  E_47809 = ( E_48136 ? E_48115_68642 : E_48189 ) ;
wire  [2:0]  E_48092_89767 = { {2{1'b0}}, E_48092 }; /* zero-padding */ 
  assign /* unsigned  1-bit */  E_48136 = (E_48189 == E_48092_89767) ;
  assign /* unsigned  3-bit */  E_48115_68642 = ( E_48115 ) ;
  assign /* unsigned  3-bit */  E_47807 = ( E_48169 ? E_47809 : E_47806_68640 ) ;
  assign /* unsigned  3-bit */  E_47806_68640 = ( E_47806 ) ;
  assign /* unsigned  3-bit */  E_47805 = ( E_48174 ? E_47803 : E_47804_68639 ) ;
  assign /* unsigned  3-bit */  E_47804_68639 = ( E_47804 ) ;
  assign /* unsigned  3-bit */  E_47803 = ( E_48185 ? E_47810 : E_48163 ) ;
  assign /* unsigned  3-bit */  E_48163 = 3'h4;
  assign /* unsigned  3-bit */  E_47802 = ( E_48195 ? E_47811 : E_48148 ) ;
  assign /* unsigned  3-bit */  E_47801 = ( E_48200 ? E_47800 : E_48176 ) ;
  assign /* unsigned  3-bit */  E_47800 = ( E_48144 ? E_47812 : E_48188 ) ;
  assign /* unsigned  3-bit */  E_60005 = 3'h1;
  CPL_FF#20  I_48050_reg ( .q ( E_48162 )  , .qbar (  )  , .d ( E_48207 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48254 )  );
  assign /* unsigned 20-bit */  E_48207 = ( E_48159 ? E_48167 : E_48068 ) ;
  assign /* unsigned 20-bit */  E_48254 = 20'hX; /*CDBImplicitXNone*/
  CPL_FF#20  I_48052_reg ( .q ( E_48157 )  , .qbar (  )  , .d ( E_48208 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48255 )  );
  assign /* unsigned 20-bit */  E_48208 = ( E_48156 ? E_48172 : E_48016 ) ;
  assign /* unsigned 20-bit */  E_48255 = 20'hX; /*CDBImplicitXNone*/
  assign /* unsigned 10-bit */  E_51065 = 10'h3ff;
  assign /* unsigned 32-bit */  E_48055_clone_48407 = ( E_48159 ? E_49059 : asm_sym_data_21 ) ;
  assign /* unsigned 32-bit */  E_49059 = ( E_49046 ? E_48124 : E_49057 ) ;
wire  [20:0]  E_48053_89768 = { {1{1'b0}}, E_48053 }; /* zero-padding */ 
  assign /* unsigned  1-bit */  E_49046 = (E_48076 == E_48053_89768) ;
  assign /* unsigned 21-bit */  E_48076 = (E_48068 + E_48075) ;
  assign /* unsigned 32-bit */  E_49057 = ( E_51058 ? E_48073 : asm_sym_data_21 ) ;
  assign /* unsigned  1-bit */  E_51058 = (E_48068 == E_48053) ;
  assign /* unsigned 32-bit */  E_48073 = ( E_48072 ? E_48069 : E_48071 ) ;
  assign /* unsigned  1-bit */  E_48072 = (E_48071 > E_48083) ;
  assign /* unsigned 32-bit */  E_48071 = (E_48120 + E_48114) ;
  assign /* unsigned 32-bit */  E_48120 = ( E_48347 ? OOB_X_1 : E_48120_clone_48342 ) ;
  assign /* unsigned  1-bit */  E_48347 = (E_51359 > E_51065) ;
  assign /* unsigned 20-bit */  E_51359 = (E_48117 + E_48115) ;
  assign /* unsigned 20-bit */  E_48117 = (E_48116 <<< E_48115) ;
  assign /* unsigned 19-bit */  E_48116 = ( E_48068 ) ;
  assign /* unsigned 32-bit */  E_48114 = ( E_48113 ? E_48080 : E_48112 ) ;
  assign /* unsigned  1-bit */  E_48113 = (E_48112 >= E_48083) ;
  assign /* unsigned 32-bit */  E_48112 = (E_48110 - E_48091) ;
  assign /* unsigned 32-bit */  E_48110 = (E_48108 * E_48106) ;
  assign /* unsigned 32-bit */  E_48108 = ( E_48347 ? OOB_X_2 : E_48108_clone_48355 ) ;
  assign /* unsigned 32-bit */  E_48106 = ( E_48373 ? OOB_X_3 : E_48106_clone_48368 ) ;
  assign /* unsigned  1-bit */  E_48373 = (E_51357 > E_51065) ;
  assign /* unsigned 20-bit */  E_51357 = (E_48102 & E_48068) ;
  assign /* unsigned 20-bit */  E_48102 = ( E_48165 ? E_48100 : E_48101 ) ;
  CPL_FF#20  I_48058_reg ( .q ( E_48101 )  , .qbar (  )  , .d ( E_48040 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48258 )  );
  assign /* unsigned 20-bit */  E_48040 = ( E_48170 ? E_48039 : E_48102 ) ;
  assign /* unsigned 20-bit */  E_48039 = ( E_48038 ) ;
  assign /*   signed 32-bit */  E_48038 = ( E_48037 ? E_48092_68644 : E_48035_68647 ) ;
wire signed  [7:0]  E_48096_89769 = E_48096; /* unsign->sign */ 
  assign /* unsigned  1-bit */  E_48037 = (E_48036 > E_48096_89769) ;
  assign /* unsigned  6-bit */  E_48096 = 6'h20;
  assign /*   signed 32-bit */  E_48035_68647 = ( E_48035 ) ;
  assign /* unsigned 32-bit */  E_48035 = (E_48093 <<< E_48036) ;
  assign /*   signed  1-bit */  E_48093 = 1'sh1;
  assign /*   signed 32-bit */  E_48092_68644 = ( E_48092 ) ;
  assign /* unsigned 20-bit */  E_48258 = 20'hX; /*CDBImplicitXNone*/
  assign /* unsigned 20-bit */  E_48100 = ( E_48098 ? E_48092_68651 : E_48095 ) ;
wire signed  [7:0]  E_48096_89770 = E_48096; /* unsign->sign */ 
  assign /* unsigned  1-bit */  E_48098 = (E_48097 > E_48096_89770) ;
  assign /*   signed 21-bit */  E_48097 = (E_48182 - E_48115) ;
  assign /* unsigned 20-bit */  E_48095 = (E_48093 <<< E_48097) ;
  assign /* unsigned 32-bit */  E_48106_clone_48368 = ( E_51002 ? E_50865 : E_50825 ) ;
  assign /* unsigned  1-bit */  E_51002 = (E_51351 == E_51357) ;
  assign /* unsigned 20-bit */  E_51351 = (E_48040 & E_48016) ;
  assign /* unsigned 32-bit */  E_50825 = ( E_51018 ? E_50905 : E_50829 ) ;
  assign /* unsigned  1-bit */  E_51018 = (E_51345 == E_51357) ;
  assign /* unsigned 20-bit */  E_51345 = (E_48001 & E_47976) ;
  assign /* unsigned 20-bit */  E_48001 = ( E_48191 ? E_47999 : E_48000 ) ;
  CPL_FF#20  I_48062_reg ( .q ( E_48000 )  , .qbar (  )  , .d ( E_47961 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48260 )  );
  assign /* unsigned 20-bit */  E_47961 = ( E_48196 ? E_47960 : E_48001 ) ;
  assign /* unsigned 20-bit */  E_47960 = ( E_47959 ) ;
  assign /*   signed 32-bit */  E_47959 = ( E_47958 ? E_48092_68644 : E_47956_68643 ) ;
wire signed  [7:0]  E_48096_89771 = E_48096; /* unsign->sign */ 
  assign /* unsigned  1-bit */  E_47958 = (E_47957 > E_48096_89771) ;
  assign /*   signed 32-bit */  E_47956_68643 = ( E_47956 ) ;
  assign /* unsigned 32-bit */  E_47956 = (E_48093 <<< E_47957) ;
  assign /* unsigned 20-bit */  E_48260 = 20'hX; /*CDBImplicitXNone*/
  assign /* unsigned 20-bit */  E_47999 = ( E_47998 ) ;
  assign /*   signed 32-bit */  E_47998 = ( E_47997 ? E_48092_68644 : E_47995_68645 ) ;
wire signed  [7:0]  E_48096_89772 = E_48096; /* unsign->sign */ 
  assign /* unsigned  1-bit */  E_47997 = (E_47996 > E_48096_89772) ;
  assign /*   signed 21-bit */  E_47996 = (E_48141 - E_48115) ;
  assign /*   signed 32-bit */  E_47995_68645 = ( E_47995 ) ;
  assign /* unsigned 32-bit */  E_47995 = (E_48093 <<< E_47996) ;
  assign /* unsigned 32-bit */  E_50829 = ( E_51038 ? asm_sym_data_8 : asm_sym_data_11 ) ;
  assign /* unsigned  1-bit */  E_51038 = (E_51357 == E_51339) ;
  assign /* unsigned 20-bit */  E_51339 = (E_47961 & E_48197) ;
  assign /* unsigned 32-bit */  E_50905 = ( E_51014 ? asm_sym_data_8 : asm_sym_data_9 ) ;
  assign /* unsigned  1-bit */  E_51014 = (E_51345 == E_51339) ;
  assign /* unsigned 32-bit */  E_50865 = ( E_50994 ? E_50905 : E_50869 ) ;
  assign /* unsigned  1-bit */  E_50994 = (E_51351 == E_51345) ;
  assign /* unsigned 32-bit */  E_50869 = ( E_50998 ? asm_sym_data_8 : asm_sym_data_10 ) ;
  assign /* unsigned  1-bit */  E_50998 = (E_51351 == E_51339) ;
  assign /* unsigned 32-bit */  E_48091 = (E_48089 * E_48083) ;
  assign /* unsigned 32-bit */  E_48089 = (E_48087 >>> E_48084) ;
  assign /* unsigned 52-bit */  E_48087 = (E_48108 * E_48086) ;
  assign /* unsigned 32-bit */  E_48086 = ( E_48373 ? OOB_X_4 : E_48086_clone_48381 ) ;
  assign /* unsigned 32-bit */  E_48086_clone_48381 = ( E_51002 ? E_48028_clone_48446 : E_51037 ) ;
  assign /* unsigned 32-bit */  E_51037 = ( E_51018 ? E_51053 : E_51041 ) ;
  assign /* unsigned 32-bit */  E_51041 = ( E_51038 ? E_47949_clone_48524 : asm_sym_data_3 ) ;
  assign /* unsigned 32-bit */  E_51053 = ( E_51014 ? E_47949_clone_48524 : asm_sym_data_1 ) ;
  assign /* unsigned 32-bit */  E_48028_clone_48446 = ( E_50994 ? E_51053 : E_51049 ) ;
  assign /* unsigned 32-bit */  E_51049 = ( E_50998 ? E_47949_clone_48524 : asm_sym_data_2 ) ;
  assign /* unsigned  5-bit */  E_48084 = 5'h14;
  assign /* unsigned 32-bit */  E_48083 = ( E_48181 ? E_48081 : E_48082 ) ;
  CPL_FF#32  I_48060_reg ( .q ( E_48082 )  , .qbar (  )  , .d ( E_48083 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48259 )  );
  assign /* unsigned 32-bit */  E_48259 = 32'hX; /*CDBImplicitXNone*/
  assign /* unsigned 32-bit */  E_48080 = ( E_48079 ) ;
  assign /*   signed 33-bit */  E_48079 = (E_48112 - E_48083) ;
  assign /* unsigned 32-bit */  E_48069 = (E_48071 - E_48083) ;
  assign /* unsigned 32-bit */  E_48124 = ( E_48123 ? E_48077 : E_48122_68652 ) ;
wire signed  [2:0]  E_48092_89773 = E_48092; /* unsign->sign */ 
  assign /* unsigned  1-bit */  E_48123 = (E_48122 < E_48092_89773) ;
  assign /*   signed 32-bit */  E_48122 = (E_48120 - E_48114) ;
  assign /* unsigned 32-bit */  E_48122_68652 = ( E_48122 ) ;
  assign /* unsigned 32-bit */  E_48077 = (E_48122 + E_48083) ;
  assign /* unsigned 32-bit */  E_48051 = ( E_48050 ? E_48027 : E_48049 ) ;
  assign /* unsigned  1-bit */  E_48050 = (E_48049 >= E_48083) ;
  assign /* unsigned 32-bit */  E_48049 = ( E_48048 ) ;
  assign /*   signed 33-bit */  E_48048 = (E_48047 - E_48033) ;
  assign /* unsigned 32-bit */  E_48047 = ( E_48046 ) ;
  assign /* unsigned 64-bit */  E_48046 = (E_48045 * E_48043) ;
  assign /* unsigned 32-bit */  E_48045 = ( E_48412 ? OOB_X_7 : E_48045_clone_48420 ) ;
  assign /* unsigned 32-bit */  E_48045_clone_48420 = ( E_48159 ? E_49053 : asm_sym_data_20 ) ;
  assign /* unsigned 32-bit */  E_49053 = ( E_49037 ? E_48124 : E_49051 ) ;
wire  [20:0]  E_51353_89774 = { {1{1'b0}}, E_51353 }; /* zero-padding */ 
  assign /* unsigned  1-bit */  E_49037 = (E_48076 == E_51353_89774) ;
  assign /* unsigned 32-bit */  E_49051 = ( E_51057 ? E_48073 : asm_sym_data_20 ) ;
  assign /* unsigned  1-bit */  E_51057 = (E_48068 == E_51353) ;
  assign /* unsigned 32-bit */  E_48043 = ( E_48438 ? OOB_X_8 : E_48043_clone_48433 ) ;
  assign /* unsigned  1-bit */  E_48438 = (E_51351 > E_51065) ;
  assign /* unsigned 32-bit */  E_48043_clone_48433 = ( E_50994 ? E_48004_clone_48472 : E_50681 ) ;
  assign /* unsigned 32-bit */  E_50681 = ( E_50998 ? E_47964_clone_48511 : E_50865 ) ;
  assign /* unsigned 32-bit */  E_47964_clone_48511 = ( E_51038 ? E_48106_clone_48368 : E_50781 ) ;
  assign /* unsigned 32-bit */  E_50781 = ( E_50998 ? E_50865 : asm_sym_data_8 ) ;
  assign /* unsigned 32-bit */  E_48004_clone_48472 = ( E_51014 ? E_47964_clone_48511 : E_50733 ) ;
  assign /* unsigned 32-bit */  E_50733 = ( E_51018 ? E_48106_clone_48368 : E_50905 ) ;
  assign /* unsigned 32-bit */  E_48033 = ( E_48032 ) ;
  assign /* unsigned 64-bit */  E_48032 = (E_48031 * E_48083) ;
  assign /* unsigned 32-bit */  E_48031 = ( E_48030 ) ;
  assign /* unsigned 44-bit */  E_48030 = (E_48029 >>> E_48084) ;
  assign /* unsigned 64-bit */  E_48029 = (E_48045 * E_48028) ;
  assign /* unsigned 32-bit */  E_48028 = ( E_48438 ? OOB_X_9 : E_48028_clone_48446 ) ;
  assign /* unsigned 32-bit */  E_48027 = ( E_48026 ) ;
  assign /*   signed 33-bit */  E_48026 = (E_48049 - E_48083) ;
  assign /* unsigned 32-bit */  E_47937 = 32'hffffffff;
  CPL_FF  I_48081_reg ( .q ( E_47860 )  , .qbar (  )  , .d ( E_48220 )  , .clk ( clk )  , 
		.arst ( E_48092 )  , .arstval ( E_48092 )  );
endmodule


 
`ifndef __CPL__

module CPL_NMACROFF(q, qbar, d, clk, wen, arst, rstval, arst2, rstval2);
    parameter WIDTH = 1;
    output [WIDTH-1:0] q, qbar;
    reg    [WIDTH-1:0] q, qbar;

    input [WIDTH-1:0] d;
    input [WIDTH-1:0] rstval, rstval2;
    input             clk, wen, arst, arst2;

    always @(negedge clk or posedge arst or posedge arst2)
    begin
        if (arst)
        begin
            q <= rstval;
            qbar <= ~rstval;
        end
        else if (arst2)
        begin
            q <= rstval2;
            qbar <= ~rstval2;
        end
        else
        begin
           if( wen )
             begin
                q <= d;
                qbar <= ~d;
             end
        end
    end
endmodule



module CPL_MACROFF(q, qbar, d, clk, wen, arst, rstval, arst2, rstval2);
    parameter WIDTH = 1;
    output [WIDTH-1:0] q, qbar;
    reg    [WIDTH-1:0] q, qbar;

    input [WIDTH-1:0] d;
    input [WIDTH-1:0] rstval, rstval2;
    input             clk, wen, arst, arst2;

    always @(posedge clk or posedge arst or posedge arst2)
    begin
        if (arst)
        begin
            q <= rstval;
            qbar <= ~rstval;
        end
        else if (arst2)
        begin
            q <= rstval2;
            qbar <= ~rstval2;
        end
        else
        begin
           if( wen )
             begin
                q <= d;
                qbar <= ~d;
             end
        end
    end
endmodule


module CPL_FF(q, qbar, d, clk, arst, arstval);
    parameter WIDTH = 1;
    output [WIDTH-1:0] q, qbar;
    reg    [WIDTH-1:0] q, qbar;

    input [WIDTH-1:0] d;
    input [WIDTH-1:0] arstval;
    input             clk, arst;

    always @(posedge clk or posedge arst)
    begin
        if (arst)
        begin
            q <= arstval;
            qbar <= ~arstval;
        end
        else
        begin
            q <= d;
            qbar <= ~d;
        end
    end
endmodule


`endif // __CPL__
