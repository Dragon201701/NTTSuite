
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> ../td_ccore_solutions/modulo_dev_d3e65941ee7586d7daaa2e36d0d005555a5b_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Aug 26 01:37:26 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    modulo_dev_core
// ------------------------------------------------------------------


module modulo_dev_core (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;


  // Interconnect Declarations
  wire [63:0] base_rsci_idat;
  wire [63:0] m_rsci_idat;
  reg [63:0] return_rsci_d;
  wire ccs_ccore_start_rsci_idat;
  reg [63:0] result_rem_12_cmp_a;
  reg [63:0] result_rem_12_cmp_b;
  wire [63:0] result_rem_12_cmp_z;
  reg [63:0] result_rem_12_cmp_1_a;
  reg [63:0] result_rem_12_cmp_1_b;
  wire [63:0] result_rem_12_cmp_1_z;
  reg [63:0] result_rem_12_cmp_2_a;
  reg [63:0] result_rem_12_cmp_2_b;
  wire [63:0] result_rem_12_cmp_2_z;
  reg [63:0] result_rem_12_cmp_3_a;
  reg [63:0] result_rem_12_cmp_3_b;
  wire [63:0] result_rem_12_cmp_3_z;
  reg [63:0] result_rem_12_cmp_4_a;
  reg [63:0] result_rem_12_cmp_4_b;
  wire [63:0] result_rem_12_cmp_4_z;
  reg [63:0] result_rem_12_cmp_5_a;
  reg [63:0] result_rem_12_cmp_5_b;
  wire [63:0] result_rem_12_cmp_5_z;
  reg [63:0] result_rem_12_cmp_6_a;
  reg [63:0] result_rem_12_cmp_6_b;
  wire [63:0] result_rem_12_cmp_6_z;
  reg [63:0] result_rem_12_cmp_7_a;
  reg [63:0] result_rem_12_cmp_7_b;
  wire [63:0] result_rem_12_cmp_7_z;
  reg [63:0] result_rem_12_cmp_8_a;
  reg [63:0] result_rem_12_cmp_8_b;
  wire [63:0] result_rem_12_cmp_8_z;
  reg [63:0] result_rem_12_cmp_9_a;
  reg [63:0] result_rem_12_cmp_9_b;
  wire [63:0] result_rem_12_cmp_9_z;
  reg [63:0] result_rem_12_cmp_10_a;
  reg [63:0] result_rem_12_cmp_10_b;
  wire [63:0] result_rem_12_cmp_10_z;
  wire [3:0] result_result_acc_tmp;
  wire [4:0] nl_result_result_acc_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_3;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_11;
  wire and_dcpl_13;
  wire and_dcpl_18;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_28;
  wire and_dcpl_29;
  wire and_dcpl_30;
  wire and_dcpl_31;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_37;
  wire and_dcpl_38;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_41;
  wire and_dcpl_42;
  wire and_dcpl_43;
  wire and_dcpl_45;
  wire and_dcpl_47;
  wire and_dcpl_50;
  wire and_dcpl_51;
  wire and_dcpl_52;
  wire and_dcpl_53;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_63;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_68;
  wire and_dcpl_70;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_88;
  wire and_dcpl_89;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_96;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_117;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire and_dcpl_120;
  wire and_dcpl_122;
  wire and_dcpl_125;
  wire and_dcpl_127;
  wire and_dcpl_128;
  wire and_dcpl_129;
  wire and_dcpl_130;
  wire and_dcpl_131;
  wire and_dcpl_132;
  wire and_dcpl_133;
  wire and_dcpl_134;
  wire and_dcpl_135;
  wire and_dcpl_136;
  wire and_dcpl_137;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_142;
  wire and_dcpl_143;
  wire and_dcpl_145;
  wire and_dcpl_147;
  wire and_dcpl_149;
  wire and_dcpl_150;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_168;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_194;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_199;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire and_dcpl_214;
  wire and_dcpl_218;
  wire and_dcpl_221;
  wire and_dcpl_228;
  wire and_dcpl_232;
  wire and_dcpl_233;
  wire and_dcpl_234;
  wire and_dcpl_235;
  wire and_dcpl_237;
  wire and_dcpl_239;
  wire and_dcpl_240;
  wire and_dcpl_244;
  wire and_dcpl_249;
  wire and_dcpl_254;
  wire and_dcpl_260;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire or_tmp_2;
  wire and_dcpl_269;
  wire mux_tmp_1;
  wire and_dcpl_275;
  wire mux_tmp_3;
  wire mux_tmp_4;
  wire and_dcpl_281;
  wire mux_tmp_6;
  wire mux_tmp_7;
  wire mux_tmp_8;
  wire and_dcpl_287;
  wire mux_tmp_10;
  wire mux_tmp_11;
  wire mux_tmp_12;
  wire mux_tmp_13;
  wire and_dcpl_293;
  wire mux_tmp_15;
  wire mux_tmp_16;
  wire mux_tmp_17;
  wire mux_tmp_18;
  wire mux_tmp_19;
  wire and_dcpl_299;
  wire mux_tmp_21;
  wire mux_tmp_22;
  wire mux_tmp_23;
  wire mux_tmp_24;
  wire mux_tmp_25;
  wire mux_tmp_26;
  wire and_dcpl_305;
  wire mux_tmp_28;
  wire mux_tmp_29;
  wire mux_tmp_30;
  wire mux_tmp_31;
  wire mux_tmp_32;
  wire mux_tmp_33;
  wire mux_tmp_34;
  wire and_dcpl_311;
  wire and_tmp_6;
  wire mux_tmp_36;
  wire mux_tmp_37;
  wire and_dcpl_318;
  wire and_dcpl_319;
  wire or_tmp_102;
  wire and_dcpl_322;
  wire mux_tmp_39;
  wire and_dcpl_325;
  wire mux_tmp_41;
  wire mux_tmp_42;
  wire and_dcpl_329;
  wire mux_tmp_44;
  wire mux_tmp_45;
  wire mux_tmp_46;
  wire and_dcpl_333;
  wire mux_tmp_48;
  wire mux_tmp_49;
  wire mux_tmp_50;
  wire mux_tmp_51;
  wire and_dcpl_337;
  wire mux_tmp_53;
  wire mux_tmp_54;
  wire mux_tmp_55;
  wire mux_tmp_56;
  wire mux_tmp_57;
  wire and_dcpl_341;
  wire mux_tmp_59;
  wire mux_tmp_60;
  wire mux_tmp_61;
  wire mux_tmp_62;
  wire mux_tmp_63;
  wire mux_tmp_64;
  wire and_dcpl_344;
  wire mux_tmp_66;
  wire mux_tmp_67;
  wire mux_tmp_68;
  wire mux_tmp_69;
  wire mux_tmp_70;
  wire mux_tmp_71;
  wire mux_tmp_72;
  wire and_dcpl_347;
  wire and_tmp_13;
  wire mux_tmp_74;
  wire mux_tmp_75;
  wire and_dcpl_352;
  wire and_dcpl_353;
  wire or_tmp_202;
  wire and_dcpl_357;
  wire mux_tmp_77;
  wire and_dcpl_361;
  wire mux_tmp_79;
  wire mux_tmp_80;
  wire and_dcpl_364;
  wire mux_tmp_82;
  wire mux_tmp_83;
  wire mux_tmp_84;
  wire and_dcpl_367;
  wire mux_tmp_86;
  wire mux_tmp_87;
  wire mux_tmp_88;
  wire mux_tmp_89;
  wire and_dcpl_370;
  wire mux_tmp_91;
  wire mux_tmp_92;
  wire mux_tmp_93;
  wire mux_tmp_94;
  wire mux_tmp_95;
  wire and_dcpl_373;
  wire mux_tmp_97;
  wire mux_tmp_98;
  wire mux_tmp_99;
  wire mux_tmp_100;
  wire mux_tmp_101;
  wire mux_tmp_102;
  wire and_dcpl_377;
  wire mux_tmp_104;
  wire mux_tmp_105;
  wire mux_tmp_106;
  wire mux_tmp_107;
  wire mux_tmp_108;
  wire mux_tmp_109;
  wire mux_tmp_110;
  wire and_dcpl_381;
  wire and_tmp_20;
  wire mux_tmp_112;
  wire mux_tmp_113;
  wire and_dcpl_386;
  wire and_dcpl_387;
  wire or_tmp_302;
  wire and_dcpl_390;
  wire mux_tmp_115;
  wire and_dcpl_393;
  wire mux_tmp_117;
  wire mux_tmp_118;
  wire and_dcpl_396;
  wire mux_tmp_120;
  wire mux_tmp_121;
  wire mux_tmp_122;
  wire and_dcpl_399;
  wire mux_tmp_124;
  wire mux_tmp_125;
  wire mux_tmp_126;
  wire mux_tmp_127;
  wire and_dcpl_402;
  wire mux_tmp_129;
  wire mux_tmp_130;
  wire mux_tmp_131;
  wire mux_tmp_132;
  wire mux_tmp_133;
  wire and_dcpl_405;
  wire mux_tmp_135;
  wire mux_tmp_136;
  wire mux_tmp_137;
  wire mux_tmp_138;
  wire mux_tmp_139;
  wire mux_tmp_140;
  wire and_dcpl_408;
  wire mux_tmp_142;
  wire mux_tmp_143;
  wire mux_tmp_144;
  wire mux_tmp_145;
  wire mux_tmp_146;
  wire mux_tmp_147;
  wire mux_tmp_148;
  wire and_dcpl_411;
  wire and_tmp_27;
  wire mux_tmp_150;
  wire mux_tmp_151;
  wire and_dcpl_417;
  wire and_dcpl_418;
  wire or_tmp_402;
  wire and_dcpl_422;
  wire mux_tmp_153;
  wire and_dcpl_426;
  wire mux_tmp_155;
  wire mux_tmp_156;
  wire and_dcpl_430;
  wire mux_tmp_158;
  wire mux_tmp_159;
  wire mux_tmp_160;
  wire and_dcpl_433;
  wire mux_tmp_162;
  wire mux_tmp_163;
  wire mux_tmp_164;
  wire mux_tmp_165;
  wire and_dcpl_437;
  wire mux_tmp_167;
  wire mux_tmp_168;
  wire mux_tmp_169;
  wire mux_tmp_170;
  wire mux_tmp_171;
  wire and_dcpl_441;
  wire mux_tmp_173;
  wire mux_tmp_174;
  wire mux_tmp_175;
  wire mux_tmp_176;
  wire mux_tmp_177;
  wire mux_tmp_178;
  wire and_dcpl_444;
  wire mux_tmp_180;
  wire mux_tmp_181;
  wire mux_tmp_182;
  wire mux_tmp_183;
  wire mux_tmp_184;
  wire mux_tmp_185;
  wire mux_tmp_186;
  wire and_dcpl_447;
  wire and_tmp_34;
  wire mux_tmp_188;
  wire mux_tmp_189;
  wire and_dcpl_452;
  wire or_tmp_502;
  wire and_dcpl_455;
  wire mux_tmp_191;
  wire and_dcpl_458;
  wire mux_tmp_193;
  wire mux_tmp_194;
  wire and_dcpl_462;
  wire mux_tmp_196;
  wire mux_tmp_197;
  wire mux_tmp_198;
  wire and_dcpl_464;
  wire mux_tmp_200;
  wire mux_tmp_201;
  wire mux_tmp_202;
  wire mux_tmp_203;
  wire and_dcpl_468;
  wire mux_tmp_205;
  wire mux_tmp_206;
  wire mux_tmp_207;
  wire mux_tmp_208;
  wire mux_tmp_209;
  wire and_dcpl_472;
  wire mux_tmp_211;
  wire mux_tmp_212;
  wire mux_tmp_213;
  wire mux_tmp_214;
  wire mux_tmp_215;
  wire mux_tmp_216;
  wire and_dcpl_474;
  wire mux_tmp_218;
  wire mux_tmp_219;
  wire mux_tmp_220;
  wire mux_tmp_221;
  wire mux_tmp_222;
  wire mux_tmp_223;
  wire mux_tmp_224;
  wire and_dcpl_476;
  wire and_tmp_41;
  wire mux_tmp_226;
  wire mux_tmp_227;
  wire and_dcpl_480;
  wire or_tmp_602;
  wire and_dcpl_484;
  wire mux_tmp_229;
  wire and_dcpl_488;
  wire mux_tmp_231;
  wire mux_tmp_232;
  wire and_dcpl_491;
  wire mux_tmp_234;
  wire mux_tmp_235;
  wire mux_tmp_236;
  wire and_dcpl_493;
  wire mux_tmp_238;
  wire mux_tmp_239;
  wire mux_tmp_240;
  wire mux_tmp_241;
  wire and_dcpl_496;
  wire mux_tmp_243;
  wire mux_tmp_244;
  wire mux_tmp_245;
  wire mux_tmp_246;
  wire mux_tmp_247;
  wire and_dcpl_499;
  wire mux_tmp_249;
  wire mux_tmp_250;
  wire mux_tmp_251;
  wire mux_tmp_252;
  wire mux_tmp_253;
  wire mux_tmp_254;
  wire and_dcpl_501;
  wire mux_tmp_256;
  wire mux_tmp_257;
  wire mux_tmp_258;
  wire mux_tmp_259;
  wire mux_tmp_260;
  wire mux_tmp_261;
  wire mux_tmp_262;
  wire and_dcpl_503;
  wire and_tmp_48;
  wire mux_tmp_264;
  wire mux_tmp_265;
  wire and_dcpl_507;
  wire or_tmp_702;
  wire and_dcpl_510;
  wire mux_tmp_267;
  wire and_dcpl_513;
  wire mux_tmp_269;
  wire mux_tmp_270;
  wire and_dcpl_516;
  wire mux_tmp_272;
  wire mux_tmp_273;
  wire mux_tmp_274;
  wire and_dcpl_518;
  wire mux_tmp_276;
  wire mux_tmp_277;
  wire mux_tmp_278;
  wire mux_tmp_279;
  wire and_dcpl_521;
  wire mux_tmp_281;
  wire mux_tmp_282;
  wire mux_tmp_283;
  wire mux_tmp_284;
  wire mux_tmp_285;
  wire and_dcpl_524;
  wire mux_tmp_287;
  wire mux_tmp_288;
  wire mux_tmp_289;
  wire mux_tmp_290;
  wire mux_tmp_291;
  wire mux_tmp_292;
  wire and_dcpl_526;
  wire mux_tmp_294;
  wire mux_tmp_295;
  wire mux_tmp_296;
  wire mux_tmp_297;
  wire mux_tmp_298;
  wire mux_tmp_299;
  wire mux_tmp_300;
  wire and_dcpl_528;
  wire and_tmp_55;
  wire mux_tmp_302;
  wire mux_tmp_303;
  wire and_dcpl_532;
  wire and_dcpl_533;
  wire not_tmp_645;
  wire or_tmp_801;
  wire and_dcpl_536;
  wire mux_tmp_305;
  wire and_dcpl_539;
  wire mux_tmp_307;
  wire mux_tmp_308;
  wire and_dcpl_542;
  wire mux_tmp_310;
  wire mux_tmp_311;
  wire mux_tmp_312;
  wire and_dcpl_546;
  wire mux_tmp_314;
  wire mux_tmp_315;
  wire mux_tmp_316;
  wire mux_tmp_317;
  wire and_dcpl_549;
  wire mux_tmp_319;
  wire mux_tmp_320;
  wire mux_tmp_321;
  wire mux_tmp_322;
  wire mux_tmp_323;
  wire and_dcpl_552;
  wire mux_tmp_325;
  wire mux_tmp_326;
  wire mux_tmp_327;
  wire mux_tmp_328;
  wire mux_tmp_329;
  wire mux_tmp_330;
  wire and_dcpl_556;
  wire mux_tmp_332;
  wire mux_tmp_333;
  wire mux_tmp_334;
  wire mux_tmp_335;
  wire mux_tmp_336;
  wire mux_tmp_337;
  wire mux_tmp_338;
  wire and_dcpl_560;
  wire or_tmp_897;
  wire mux_tmp_340;
  wire mux_tmp_341;
  wire mux_tmp_342;
  wire mux_tmp_343;
  wire mux_tmp_344;
  wire mux_tmp_345;
  wire mux_tmp_346;
  wire mux_tmp_347;
  wire mux_tmp_348;
  wire and_dcpl_566;
  wire or_tmp_909;
  wire and_dcpl_568;
  wire mux_tmp_350;
  wire and_dcpl_570;
  wire mux_tmp_352;
  wire mux_tmp_353;
  wire and_dcpl_572;
  wire mux_tmp_355;
  wire mux_tmp_356;
  wire mux_tmp_357;
  wire and_dcpl_576;
  wire mux_tmp_359;
  wire mux_tmp_360;
  wire mux_tmp_361;
  wire mux_tmp_362;
  wire and_dcpl_578;
  wire mux_tmp_364;
  wire mux_tmp_365;
  wire mux_tmp_366;
  wire mux_tmp_367;
  wire mux_tmp_368;
  wire and_dcpl_580;
  wire mux_tmp_370;
  wire mux_tmp_371;
  wire mux_tmp_372;
  wire mux_tmp_373;
  wire mux_tmp_374;
  wire mux_tmp_375;
  wire and_dcpl_583;
  wire mux_tmp_377;
  wire mux_tmp_378;
  wire mux_tmp_379;
  wire mux_tmp_380;
  wire mux_tmp_381;
  wire mux_tmp_382;
  wire mux_tmp_383;
  wire and_dcpl_586;
  wire or_tmp_1005;
  wire mux_tmp_385;
  wire mux_tmp_386;
  wire mux_tmp_387;
  wire mux_tmp_388;
  wire mux_tmp_389;
  wire mux_tmp_390;
  wire mux_tmp_391;
  wire mux_tmp_392;
  wire mux_tmp_393;
  wire and_dcpl_590;
  wire or_tmp_1017;
  wire and_dcpl_592;
  wire mux_tmp_395;
  wire and_dcpl_594;
  wire mux_tmp_397;
  wire mux_tmp_398;
  wire and_dcpl_596;
  wire mux_tmp_400;
  wire mux_tmp_401;
  wire mux_tmp_402;
  wire and_dcpl_599;
  wire mux_tmp_404;
  wire mux_tmp_405;
  wire mux_tmp_406;
  wire mux_tmp_407;
  wire and_dcpl_601;
  wire mux_tmp_409;
  wire mux_tmp_410;
  wire mux_tmp_411;
  wire mux_tmp_412;
  wire mux_tmp_413;
  wire and_dcpl_603;
  wire mux_tmp_415;
  wire mux_tmp_416;
  wire mux_tmp_417;
  wire mux_tmp_418;
  wire mux_tmp_419;
  wire mux_tmp_420;
  wire and_dcpl_607;
  wire mux_tmp_422;
  wire mux_tmp_423;
  wire mux_tmp_424;
  wire mux_tmp_425;
  wire mux_tmp_426;
  wire mux_tmp_427;
  wire mux_tmp_428;
  wire and_dcpl_611;
  wire or_tmp_1113;
  wire mux_tmp_430;
  wire mux_tmp_431;
  wire mux_tmp_432;
  wire mux_tmp_433;
  wire mux_tmp_434;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire mux_tmp_437;
  wire mux_tmp_438;
  reg main_stage_0_11;
  reg asn_itm_10;
  reg [3:0] result_rem_11cyc_st_9;
  reg [3:0] result_rem_11cyc_st_8;
  reg [3:0] result_rem_11cyc_st_7;
  reg [3:0] result_rem_11cyc_st_6;
  reg [3:0] result_rem_11cyc_st_5;
  reg [3:0] result_rem_11cyc_st_4;
  reg [3:0] result_rem_11cyc_st_3;
  reg [3:0] result_rem_11cyc_st_2;
  reg [3:0] result_rem_11cyc;
  reg [3:0] result_rem_11cyc_st_11;
  reg asn_itm_11;
  reg main_stage_0_12;
  reg main_stage_0_3;
  reg asn_itm_2;
  reg main_stage_0_4;
  reg asn_itm_3;
  reg main_stage_0_5;
  reg asn_itm_4;
  reg main_stage_0_6;
  reg asn_itm_5;
  reg main_stage_0_7;
  reg asn_itm_6;
  reg main_stage_0_8;
  reg asn_itm_7;
  reg main_stage_0_9;
  reg asn_itm_8;
  reg main_stage_0_10;
  reg asn_itm_9;
  reg main_stage_0_2;
  reg asn_itm_1;
  wire result_and_1_cse;
  wire result_and_3_cse;
  wire result_and_5_cse;
  wire result_and_7_cse;
  wire result_and_9_cse;
  wire result_and_11_cse;
  wire result_and_13_cse;
  wire result_and_15_cse;
  wire result_and_17_cse;
  wire result_and_19_cse;
  wire result_and_21_cse;
  wire or_3_cse;
  wire or_8_cse;
  wire or_15_cse;
  wire or_24_cse;
  wire or_35_cse;
  wire or_48_cse;
  wire or_63_cse;
  wire or_107_cse;
  wire or_112_cse;
  wire or_119_cse;
  wire or_128_cse;
  wire or_139_cse;
  wire or_152_cse;
  wire or_167_cse;
  wire or_209_cse;
  wire or_214_cse;
  wire or_221_cse;
  wire or_230_cse;
  wire or_241_cse;
  wire or_254_cse;
  wire or_269_cse;
  wire or_311_cse;
  wire or_316_cse;
  wire or_323_cse;
  wire or_332_cse;
  wire or_343_cse;
  wire or_356_cse;
  wire or_371_cse;
  wire nand_144_cse;
  wire or_413_cse;
  wire or_418_cse;
  wire or_425_cse;
  wire or_434_cse;
  wire or_445_cse;
  wire or_458_cse;
  wire or_473_cse;
  wire nand_138_cse;
  wire or_516_cse;
  wire or_521_cse;
  wire or_528_cse;
  wire or_537_cse;
  wire and_790_cse;
  wire or_548_cse;
  wire or_561_cse;
  wire or_576_cse;
  wire nand_146_cse;
  wire or_617_cse;
  wire or_622_cse;
  wire or_629_cse;
  wire or_638_cse;
  wire or_649_cse;
  wire or_662_cse;
  wire or_677_cse;
  wire or_718_cse;
  wire nand_112_cse;
  wire nand_108_cse;
  wire nand_103_cse;
  wire nand_97_cse;
  wire or_763_cse;
  wire nand_83_cse;
  wire or_818_cse;
  wire or_823_cse;
  wire or_830_cse;
  wire or_839_cse;
  wire nand_58_cse;
  wire or_850_cse;
  wire nand_55_cse;
  wire or_863_cse;
  wire nand_51_cse;
  wire or_878_cse;
  wire and_749_cse;
  wire or_928_cse;
  wire and_747_cse;
  wire or_933_cse;
  wire and_744_cse;
  wire or_940_cse;
  wire and_740_cse;
  wire or_949_cse;
  wire or_960_cse;
  wire and_731_cse;
  wire or_973_cse;
  wire and_725_cse;
  wire nand_42_cse;
  wire or_988_cse;
  wire or_1037_cse;
  wire or_1042_cse;
  wire or_1049_cse;
  wire or_1058_cse;
  wire or_1069_cse;
  wire or_1082_cse;
  wire or_1097_cse;
  reg [63:0] base_buf_sva_mut_2;
  reg [63:0] base_buf_sva_mut_3;
  reg [63:0] base_buf_sva_mut_4;
  reg [63:0] base_buf_sva_mut_5;
  reg [63:0] base_buf_sva_mut_6;
  reg [63:0] base_buf_sva_mut_7;
  reg [63:0] base_buf_sva_mut_8;
  reg [63:0] base_buf_sva_mut_9;
  reg [63:0] base_buf_sva_mut_10;
  reg [63:0] m_buf_sva_mut_2;
  reg [63:0] m_buf_sva_mut_3;
  reg [63:0] m_buf_sva_mut_4;
  reg [63:0] m_buf_sva_mut_5;
  reg [63:0] m_buf_sva_mut_6;
  reg [63:0] m_buf_sva_mut_7;
  reg [63:0] m_buf_sva_mut_8;
  reg [63:0] m_buf_sva_mut_9;
  reg [63:0] m_buf_sva_mut_10;
  reg [63:0] base_buf_sva_mut_1_2;
  reg [63:0] base_buf_sva_mut_1_3;
  reg [63:0] base_buf_sva_mut_1_4;
  reg [63:0] base_buf_sva_mut_1_5;
  reg [63:0] base_buf_sva_mut_1_6;
  reg [63:0] base_buf_sva_mut_1_7;
  reg [63:0] base_buf_sva_mut_1_8;
  reg [63:0] base_buf_sva_mut_1_9;
  reg [63:0] base_buf_sva_mut_1_10;
  reg [63:0] m_buf_sva_mut_1_2;
  reg [63:0] m_buf_sva_mut_1_3;
  reg [63:0] m_buf_sva_mut_1_4;
  reg [63:0] m_buf_sva_mut_1_5;
  reg [63:0] m_buf_sva_mut_1_6;
  reg [63:0] m_buf_sva_mut_1_7;
  reg [63:0] m_buf_sva_mut_1_8;
  reg [63:0] m_buf_sva_mut_1_9;
  reg [63:0] m_buf_sva_mut_1_10;
  reg [63:0] base_buf_sva_mut_2_2;
  reg [63:0] base_buf_sva_mut_2_3;
  reg [63:0] base_buf_sva_mut_2_4;
  reg [63:0] base_buf_sva_mut_2_5;
  reg [63:0] base_buf_sva_mut_2_6;
  reg [63:0] base_buf_sva_mut_2_7;
  reg [63:0] base_buf_sva_mut_2_8;
  reg [63:0] base_buf_sva_mut_2_9;
  reg [63:0] base_buf_sva_mut_2_10;
  reg [63:0] m_buf_sva_mut_2_2;
  reg [63:0] m_buf_sva_mut_2_3;
  reg [63:0] m_buf_sva_mut_2_4;
  reg [63:0] m_buf_sva_mut_2_5;
  reg [63:0] m_buf_sva_mut_2_6;
  reg [63:0] m_buf_sva_mut_2_7;
  reg [63:0] m_buf_sva_mut_2_8;
  reg [63:0] m_buf_sva_mut_2_9;
  reg [63:0] m_buf_sva_mut_2_10;
  reg [63:0] base_buf_sva_mut_3_2;
  reg [63:0] base_buf_sva_mut_3_3;
  reg [63:0] base_buf_sva_mut_3_4;
  reg [63:0] base_buf_sva_mut_3_5;
  reg [63:0] base_buf_sva_mut_3_6;
  reg [63:0] base_buf_sva_mut_3_7;
  reg [63:0] base_buf_sva_mut_3_8;
  reg [63:0] base_buf_sva_mut_3_9;
  reg [63:0] base_buf_sva_mut_3_10;
  reg [63:0] m_buf_sva_mut_3_2;
  reg [63:0] m_buf_sva_mut_3_3;
  reg [63:0] m_buf_sva_mut_3_4;
  reg [63:0] m_buf_sva_mut_3_5;
  reg [63:0] m_buf_sva_mut_3_6;
  reg [63:0] m_buf_sva_mut_3_7;
  reg [63:0] m_buf_sva_mut_3_8;
  reg [63:0] m_buf_sva_mut_3_9;
  reg [63:0] m_buf_sva_mut_3_10;
  reg [63:0] base_buf_sva_mut_4_2;
  reg [63:0] base_buf_sva_mut_4_3;
  reg [63:0] base_buf_sva_mut_4_4;
  reg [63:0] base_buf_sva_mut_4_5;
  reg [63:0] base_buf_sva_mut_4_6;
  reg [63:0] base_buf_sva_mut_4_7;
  reg [63:0] base_buf_sva_mut_4_8;
  reg [63:0] base_buf_sva_mut_4_9;
  reg [63:0] base_buf_sva_mut_4_10;
  reg [63:0] m_buf_sva_mut_4_2;
  reg [63:0] m_buf_sva_mut_4_3;
  reg [63:0] m_buf_sva_mut_4_4;
  reg [63:0] m_buf_sva_mut_4_5;
  reg [63:0] m_buf_sva_mut_4_6;
  reg [63:0] m_buf_sva_mut_4_7;
  reg [63:0] m_buf_sva_mut_4_8;
  reg [63:0] m_buf_sva_mut_4_9;
  reg [63:0] m_buf_sva_mut_4_10;
  reg [63:0] base_buf_sva_mut_5_2;
  reg [63:0] base_buf_sva_mut_5_3;
  reg [63:0] base_buf_sva_mut_5_4;
  reg [63:0] base_buf_sva_mut_5_5;
  reg [63:0] base_buf_sva_mut_5_6;
  reg [63:0] base_buf_sva_mut_5_7;
  reg [63:0] base_buf_sva_mut_5_8;
  reg [63:0] base_buf_sva_mut_5_9;
  reg [63:0] base_buf_sva_mut_5_10;
  reg [63:0] m_buf_sva_mut_5_2;
  reg [63:0] m_buf_sva_mut_5_3;
  reg [63:0] m_buf_sva_mut_5_4;
  reg [63:0] m_buf_sva_mut_5_5;
  reg [63:0] m_buf_sva_mut_5_6;
  reg [63:0] m_buf_sva_mut_5_7;
  reg [63:0] m_buf_sva_mut_5_8;
  reg [63:0] m_buf_sva_mut_5_9;
  reg [63:0] m_buf_sva_mut_5_10;
  reg [63:0] base_buf_sva_mut_6_2;
  reg [63:0] base_buf_sva_mut_6_3;
  reg [63:0] base_buf_sva_mut_6_4;
  reg [63:0] base_buf_sva_mut_6_5;
  reg [63:0] base_buf_sva_mut_6_6;
  reg [63:0] base_buf_sva_mut_6_7;
  reg [63:0] base_buf_sva_mut_6_8;
  reg [63:0] base_buf_sva_mut_6_9;
  reg [63:0] base_buf_sva_mut_6_10;
  reg [63:0] m_buf_sva_mut_6_2;
  reg [63:0] m_buf_sva_mut_6_3;
  reg [63:0] m_buf_sva_mut_6_4;
  reg [63:0] m_buf_sva_mut_6_5;
  reg [63:0] m_buf_sva_mut_6_6;
  reg [63:0] m_buf_sva_mut_6_7;
  reg [63:0] m_buf_sva_mut_6_8;
  reg [63:0] m_buf_sva_mut_6_9;
  reg [63:0] m_buf_sva_mut_6_10;
  reg [63:0] base_buf_sva_mut_7_2;
  reg [63:0] base_buf_sva_mut_7_3;
  reg [63:0] base_buf_sva_mut_7_4;
  reg [63:0] base_buf_sva_mut_7_5;
  reg [63:0] base_buf_sva_mut_7_6;
  reg [63:0] base_buf_sva_mut_7_7;
  reg [63:0] base_buf_sva_mut_7_8;
  reg [63:0] base_buf_sva_mut_7_9;
  reg [63:0] base_buf_sva_mut_7_10;
  reg [63:0] m_buf_sva_mut_7_2;
  reg [63:0] m_buf_sva_mut_7_3;
  reg [63:0] m_buf_sva_mut_7_4;
  reg [63:0] m_buf_sva_mut_7_5;
  reg [63:0] m_buf_sva_mut_7_6;
  reg [63:0] m_buf_sva_mut_7_7;
  reg [63:0] m_buf_sva_mut_7_8;
  reg [63:0] m_buf_sva_mut_7_9;
  reg [63:0] m_buf_sva_mut_7_10;
  reg [63:0] base_buf_sva_mut_8_2;
  reg [63:0] base_buf_sva_mut_8_3;
  reg [63:0] base_buf_sva_mut_8_4;
  reg [63:0] base_buf_sva_mut_8_5;
  reg [63:0] base_buf_sva_mut_8_6;
  reg [63:0] base_buf_sva_mut_8_7;
  reg [63:0] base_buf_sva_mut_8_8;
  reg [63:0] base_buf_sva_mut_8_9;
  reg [63:0] base_buf_sva_mut_8_10;
  reg [63:0] m_buf_sva_mut_8_2;
  reg [63:0] m_buf_sva_mut_8_3;
  reg [63:0] m_buf_sva_mut_8_4;
  reg [63:0] m_buf_sva_mut_8_5;
  reg [63:0] m_buf_sva_mut_8_6;
  reg [63:0] m_buf_sva_mut_8_7;
  reg [63:0] m_buf_sva_mut_8_8;
  reg [63:0] m_buf_sva_mut_8_9;
  reg [63:0] m_buf_sva_mut_8_10;
  reg [63:0] base_buf_sva_mut_9_2;
  reg [63:0] base_buf_sva_mut_9_3;
  reg [63:0] base_buf_sva_mut_9_4;
  reg [63:0] base_buf_sva_mut_9_5;
  reg [63:0] base_buf_sva_mut_9_6;
  reg [63:0] base_buf_sva_mut_9_7;
  reg [63:0] base_buf_sva_mut_9_8;
  reg [63:0] base_buf_sva_mut_9_9;
  reg [63:0] base_buf_sva_mut_9_10;
  reg [63:0] m_buf_sva_mut_9_2;
  reg [63:0] m_buf_sva_mut_9_3;
  reg [63:0] m_buf_sva_mut_9_4;
  reg [63:0] m_buf_sva_mut_9_5;
  reg [63:0] m_buf_sva_mut_9_6;
  reg [63:0] m_buf_sva_mut_9_7;
  reg [63:0] m_buf_sva_mut_9_8;
  reg [63:0] m_buf_sva_mut_9_9;
  reg [63:0] m_buf_sva_mut_9_10;
  reg [63:0] base_buf_sva_mut_10_2;
  reg [63:0] base_buf_sva_mut_10_3;
  reg [63:0] base_buf_sva_mut_10_4;
  reg [63:0] base_buf_sva_mut_10_5;
  reg [63:0] base_buf_sva_mut_10_6;
  reg [63:0] base_buf_sva_mut_10_7;
  reg [63:0] base_buf_sva_mut_10_8;
  reg [63:0] base_buf_sva_mut_10_9;
  reg [63:0] base_buf_sva_mut_10_10;
  reg [63:0] m_buf_sva_mut_10_2;
  reg [63:0] m_buf_sva_mut_10_3;
  reg [63:0] m_buf_sva_mut_10_4;
  reg [63:0] m_buf_sva_mut_10_5;
  reg [63:0] m_buf_sva_mut_10_6;
  reg [63:0] m_buf_sva_mut_10_7;
  reg [63:0] m_buf_sva_mut_10_8;
  reg [63:0] m_buf_sva_mut_10_9;
  reg [63:0] m_buf_sva_mut_10_10;
  reg [3:0] result_rem_11cyc_st_10;
  wire return_rsci_d_mx0c0;
  wire return_rsci_d_mx0c1;
  wire return_rsci_d_mx0c2;
  wire return_rsci_d_mx0c3;
  wire return_rsci_d_mx0c4;
  wire return_rsci_d_mx0c5;
  wire return_rsci_d_mx0c6;
  wire return_rsci_d_mx0c7;
  wire return_rsci_d_mx0c8;
  wire return_rsci_d_mx0c9;
  wire return_rsci_d_mx0c10;
  wire [3:0] result_acc_imod_1;
  wire [5:0] nl_result_acc_imod_1;
  wire [3:0] result_acc_idiv_1;
  wire [4:0] nl_result_acc_idiv_1;
  wire m_and_cse;
  wire m_and_1_cse;
  wire m_and_2_cse;
  wire m_and_3_cse;
  wire m_and_4_cse;
  wire m_and_5_cse;
  wire m_and_6_cse;
  wire m_and_7_cse;
  wire m_and_8_cse;
  wire m_and_9_cse;
  wire m_and_10_cse;
  wire m_and_11_cse;
  wire m_and_12_cse;
  wire m_and_13_cse;
  wire m_and_14_cse;
  wire m_and_15_cse;
  wire m_and_16_cse;
  wire m_and_17_cse;
  wire m_and_18_cse;
  wire m_and_19_cse;
  wire m_and_20_cse;
  wire m_and_21_cse;
  wire m_and_22_cse;
  wire m_and_23_cse;
  wire m_and_24_cse;
  wire m_and_25_cse;
  wire m_and_26_cse;
  wire m_and_27_cse;
  wire m_and_28_cse;
  wire m_and_29_cse;
  wire m_and_30_cse;
  wire m_and_31_cse;
  wire m_and_32_cse;
  wire m_and_33_cse;
  wire m_and_34_cse;
  wire m_and_35_cse;
  wire m_and_36_cse;
  wire m_and_37_cse;
  wire m_and_38_cse;
  wire m_and_39_cse;
  wire m_and_40_cse;
  wire m_and_41_cse;
  wire m_and_42_cse;
  wire m_and_43_cse;
  wire m_and_44_cse;
  wire m_and_45_cse;
  wire m_and_46_cse;
  wire m_and_47_cse;
  wire m_and_48_cse;
  wire m_and_49_cse;
  wire m_and_50_cse;
  wire m_and_51_cse;
  wire m_and_52_cse;
  wire m_and_53_cse;
  wire m_and_54_cse;
  wire m_and_55_cse;
  wire m_and_56_cse;
  wire m_and_57_cse;
  wire m_and_58_cse;
  wire m_and_59_cse;
  wire m_and_60_cse;
  wire m_and_61_cse;
  wire m_and_62_cse;
  wire m_and_63_cse;
  wire m_and_64_cse;
  wire m_and_65_cse;
  wire m_and_66_cse;
  wire m_and_67_cse;
  wire m_and_68_cse;
  wire m_and_69_cse;
  wire m_and_70_cse;
  wire m_and_71_cse;
  wire m_and_72_cse;
  wire m_and_73_cse;
  wire m_and_74_cse;
  wire m_and_75_cse;
  wire m_and_76_cse;
  wire m_and_77_cse;
  wire m_and_78_cse;
  wire m_and_79_cse;
  wire m_and_80_cse;
  wire m_and_81_cse;
  wire m_and_82_cse;
  wire m_and_83_cse;
  wire m_and_84_cse;
  wire m_and_85_cse;
  wire m_and_86_cse;
  wire m_and_87_cse;
  wire m_and_88_cse;
  wire m_and_89_cse;
  wire m_and_90_cse;
  wire m_and_91_cse;
  wire m_and_92_cse;
  wire m_and_93_cse;
  wire m_and_94_cse;
  wire m_and_95_cse;
  wire m_and_96_cse;
  wire m_and_97_cse;
  wire m_and_98_cse;

  wire[0:0] mux_nl;
  wire[0:0] nor_691_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] or_10_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] or_17_nl;
  wire[0:0] nor_688_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] or_26_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] or_37_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_677_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] or_50_nl;
  wire[0:0] nor_673_nl;
  wire[0:0] nor_674_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] nor_676_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] or_65_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] nor_667_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] nor_670_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] or_82_nl;
  wire[0:0] or_80_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] nor_660_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nor_654_nl;
  wire[0:0] nor_655_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] or_114_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] or_121_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] or_130_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] or_141_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] or_154_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] nor_627_nl;
  wire[0:0] or_169_nl;
  wire[0:0] nor_628_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] nor_630_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] or_186_nl;
  wire[0:0] or_184_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] nor_624_nl;
  wire[0:0] mux_73_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] nor_617_nl;
  wire[0:0] and_797_nl;
  wire[0:0] or_195_nl;
  wire[0:0] mux_76_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] or_216_nl;
  wire[0:0] mux_78_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] or_223_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] mux_81_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] or_232_nl;
  wire[0:0] nor_609_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] mux_85_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] or_243_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] mux_90_nl;
  wire[0:0] nor_602_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] or_256_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] mux_96_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] or_271_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] mux_103_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] or_288_nl;
  wire[0:0] or_286_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] mux_111_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] mux_114_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] or_318_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] nor_576_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] or_325_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] mux_119_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] or_334_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] nor_565_nl;
  wire[0:0] or_345_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] or_358_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_134_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] or_373_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] mux_141_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] nor_543_nl;
  wire[0:0] or_390_nl;
  wire[0:0] or_388_nl;
  wire[0:0] nor_544_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] mux_149_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] and_796_nl;
  wire[0:0] or_399_nl;
  wire[0:0] mux_152_nl;
  wire[0:0] and_795_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] or_420_nl;
  wire[0:0] mux_154_nl;
  wire[0:0] and_794_nl;
  wire[0:0] nor_539_nl;
  wire[0:0] or_427_nl;
  wire[0:0] nor_540_nl;
  wire[0:0] mux_157_nl;
  wire[0:0] and_793_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] or_436_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] mux_161_nl;
  wire[0:0] and_792_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] or_447_nl;
  wire[0:0] nor_533_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] nor_535_nl;
  wire[0:0] mux_166_nl;
  wire[0:0] and_791_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] or_460_nl;
  wire[0:0] nor_528_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] mux_172_nl;
  wire[0:0] and_789_nl;
  wire[0:0] nor_522_nl;
  wire[0:0] or_475_nl;
  wire[0:0] and_788_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] nor_524_nl;
  wire[0:0] nor_525_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] mux_179_nl;
  wire[0:0] and_787_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] or_492_nl;
  wire[0:0] or_490_nl;
  wire[0:0] nor_517_nl;
  wire[0:0] and_785_nl;
  wire[0:0] nor_518_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] nor_521_nl;
  wire[0:0] mux_187_nl;
  wire[0:0] and_786_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] or_501_nl;
  wire[0:0] mux_190_nl;
  wire[0:0] and_784_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] or_523_nl;
  wire[0:0] mux_192_nl;
  wire[0:0] and_783_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] or_530_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] mux_195_nl;
  wire[0:0] and_782_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] or_539_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_199_nl;
  wire[0:0] and_781_nl;
  wire[0:0] nor_504_nl;
  wire[0:0] or_550_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] nor_506_nl;
  wire[0:0] nor_507_nl;
  wire[0:0] mux_204_nl;
  wire[0:0] and_780_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] or_563_nl;
  wire[0:0] nor_500_nl;
  wire[0:0] nor_501_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] nor_503_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] and_778_nl;
  wire[0:0] nor_494_nl;
  wire[0:0] or_578_nl;
  wire[0:0] and_777_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] and_776_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] or_595_nl;
  wire[0:0] or_593_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] and_774_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] nor_492_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] and_775_nl;
  wire[0:0] nor_487_nl;
  wire[0:0] and_773_nl;
  wire[0:0] or_604_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] and_772_nl;
  wire[0:0] nor_486_nl;
  wire[0:0] or_624_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] and_771_nl;
  wire[0:0] nor_484_nl;
  wire[0:0] or_631_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] and_770_nl;
  wire[0:0] nor_481_nl;
  wire[0:0] or_640_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] nor_483_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] and_769_nl;
  wire[0:0] nor_477_nl;
  wire[0:0] or_651_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] nor_480_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] and_768_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] or_664_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] nor_476_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] and_766_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] or_679_nl;
  wire[0:0] and_765_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] and_764_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] or_696_nl;
  wire[0:0] or_694_nl;
  wire[0:0] nor_462_nl;
  wire[0:0] and_762_nl;
  wire[0:0] nor_463_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] nor_465_nl;
  wire[0:0] nor_466_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] and_763_nl;
  wire[0:0] nor_459_nl;
  wire[0:0] nor_460_nl;
  wire[0:0] or_705_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] and_761_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] nand_153_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] and_760_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] nand_152_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] and_759_nl;
  wire[0:0] nor_453_nl;
  wire[0:0] nand_151_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] and_758_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] nand_96_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] nor_451_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] and_757_nl;
  wire[0:0] nor_444_nl;
  wire[0:0] nand_150_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] nor_446_nl;
  wire[0:0] nor_447_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] and_755_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] and_754_nl;
  wire[0:0] nor_440_nl;
  wire[0:0] nor_441_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] nor_443_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] and_753_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] nand_72_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] and_751_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] and_752_nl;
  wire[0:0] nor_432_nl;
  wire[0:0] and_750_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_431_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] or_825_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] nor_428_nl;
  wire[0:0] or_832_nl;
  wire[0:0] and_748_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] nor_426_nl;
  wire[0:0] or_841_nl;
  wire[0:0] and_745_nl;
  wire[0:0] and_746_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] nor_424_nl;
  wire[0:0] or_852_nl;
  wire[0:0] and_741_nl;
  wire[0:0] and_742_nl;
  wire[0:0] and_743_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] nor_423_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] or_865_nl;
  wire[0:0] and_736_nl;
  wire[0:0] and_737_nl;
  wire[0:0] and_738_nl;
  wire[0:0] and_739_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] nor_421_nl;
  wire[0:0] nor_419_nl;
  wire[0:0] or_880_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] and_732_nl;
  wire[0:0] and_733_nl;
  wire[0:0] and_734_nl;
  wire[0:0] and_735_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] nor_415_nl;
  wire[0:0] or_897_nl;
  wire[0:0] or_895_nl;
  wire[0:0] and_726_nl;
  wire[0:0] nor_416_nl;
  wire[0:0] and_727_nl;
  wire[0:0] and_728_nl;
  wire[0:0] and_729_nl;
  wire[0:0] and_730_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] nor_417_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] or_914_nl;
  wire[0:0] nor_408_nl;
  wire[0:0] or_913_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] or_912_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] or_911_nl;
  wire[0:0] nor_411_nl;
  wire[0:0] or_910_nl;
  wire[0:0] nor_412_nl;
  wire[0:0] or_909_nl;
  wire[0:0] nor_413_nl;
  wire[0:0] or_908_nl;
  wire[0:0] and_724_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] nor_406_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] or_935_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] nor_404_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] or_942_nl;
  wire[0:0] and_722_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] nor_402_nl;
  wire[0:0] nor_401_nl;
  wire[0:0] or_951_nl;
  wire[0:0] and_719_nl;
  wire[0:0] and_720_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] nor_399_nl;
  wire[0:0] or_962_nl;
  wire[0:0] and_715_nl;
  wire[0:0] and_716_nl;
  wire[0:0] and_717_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] nor_398_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] or_975_nl;
  wire[0:0] and_710_nl;
  wire[0:0] and_711_nl;
  wire[0:0] and_712_nl;
  wire[0:0] and_713_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] nor_396_nl;
  wire[0:0] nor_394_nl;
  wire[0:0] or_990_nl;
  wire[0:0] nor_395_nl;
  wire[0:0] and_706_nl;
  wire[0:0] and_707_nl;
  wire[0:0] and_708_nl;
  wire[0:0] and_709_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_393_nl;
  wire[0:0] nor_390_nl;
  wire[0:0] or_1007_nl;
  wire[0:0] or_1005_nl;
  wire[0:0] and_700_nl;
  wire[0:0] nor_391_nl;
  wire[0:0] and_701_nl;
  wire[0:0] and_702_nl;
  wire[0:0] and_703_nl;
  wire[0:0] and_704_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] nor_392_nl;
  wire[0:0] nor_383_nl;
  wire[0:0] or_1024_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] nor_385_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] nor_387_nl;
  wire[0:0] or_1020_nl;
  wire[0:0] nor_388_nl;
  wire[0:0] or_1019_nl;
  wire[0:0] nor_389_nl;
  wire[0:0] or_1018_nl;
  wire[0:0] and_697_nl;
  wire[0:0] and_698_nl;
  wire[0:0] or_1016_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_382_nl;
  wire[0:0] nor_381_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] nor_380_nl;
  wire[0:0] nor_379_nl;
  wire[0:0] or_1051_nl;
  wire[0:0] and_695_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] nor_378_nl;
  wire[0:0] nor_377_nl;
  wire[0:0] or_1060_nl;
  wire[0:0] and_692_nl;
  wire[0:0] and_693_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] nor_376_nl;
  wire[0:0] nor_375_nl;
  wire[0:0] or_1071_nl;
  wire[0:0] and_688_nl;
  wire[0:0] and_689_nl;
  wire[0:0] and_690_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] nor_374_nl;
  wire[0:0] nor_373_nl;
  wire[0:0] or_1084_nl;
  wire[0:0] and_683_nl;
  wire[0:0] and_684_nl;
  wire[0:0] and_685_nl;
  wire[0:0] and_686_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] nor_372_nl;
  wire[0:0] nor_370_nl;
  wire[0:0] or_1099_nl;
  wire[0:0] nor_371_nl;
  wire[0:0] and_679_nl;
  wire[0:0] and_680_nl;
  wire[0:0] and_681_nl;
  wire[0:0] and_682_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] nor_369_nl;
  wire[0:0] nor_366_nl;
  wire[0:0] or_1116_nl;
  wire[0:0] or_1114_nl;
  wire[0:0] and_673_nl;
  wire[0:0] nor_367_nl;
  wire[0:0] and_674_nl;
  wire[0:0] and_675_nl;
  wire[0:0] and_676_nl;
  wire[0:0] and_677_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_368_nl;
  wire[0:0] nor_358_nl;
  wire[0:0] or_1133_nl;
  wire[0:0] nor_359_nl;
  wire[0:0] or_1132_nl;
  wire[0:0] nor_360_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] nor_361_nl;
  wire[0:0] or_1130_nl;
  wire[0:0] nor_362_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] nor_363_nl;
  wire[0:0] or_1128_nl;
  wire[0:0] nor_364_nl;
  wire[0:0] or_1127_nl;
  wire[0:0] and_671_nl;
  wire[0:0] nor_365_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd64)) base_rsci (
      .dat(base_rsc_dat),
      .idat(base_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd64)) return_rsci (
      .d(return_rsci_d),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp (
      .a(result_rem_12_cmp_a),
      .b(result_rem_12_cmp_b),
      .z(result_rem_12_cmp_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_1 (
      .a(result_rem_12_cmp_1_a),
      .b(result_rem_12_cmp_1_b),
      .z(result_rem_12_cmp_1_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_2 (
      .a(result_rem_12_cmp_2_a),
      .b(result_rem_12_cmp_2_b),
      .z(result_rem_12_cmp_2_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_3 (
      .a(result_rem_12_cmp_3_a),
      .b(result_rem_12_cmp_3_b),
      .z(result_rem_12_cmp_3_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_4 (
      .a(result_rem_12_cmp_4_a),
      .b(result_rem_12_cmp_4_b),
      .z(result_rem_12_cmp_4_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_5 (
      .a(result_rem_12_cmp_5_a),
      .b(result_rem_12_cmp_5_b),
      .z(result_rem_12_cmp_5_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_6 (
      .a(result_rem_12_cmp_6_a),
      .b(result_rem_12_cmp_6_b),
      .z(result_rem_12_cmp_6_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_7 (
      .a(result_rem_12_cmp_7_a),
      .b(result_rem_12_cmp_7_b),
      .z(result_rem_12_cmp_7_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_8 (
      .a(result_rem_12_cmp_8_a),
      .b(result_rem_12_cmp_8_b),
      .z(result_rem_12_cmp_8_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_9 (
      .a(result_rem_12_cmp_9_a),
      .b(result_rem_12_cmp_9_b),
      .z(result_rem_12_cmp_9_z)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd0)) result_rem_12_cmp_10 (
      .a(result_rem_12_cmp_10_a),
      .b(result_rem_12_cmp_10_b),
      .z(result_rem_12_cmp_10_z)
    );
  assign result_and_1_cse = ccs_ccore_en & (and_dcpl_263 | and_dcpl_269 | and_dcpl_275
      | and_dcpl_281 | and_dcpl_287 | and_dcpl_293 | and_dcpl_299 | and_dcpl_305
      | and_dcpl_311 | mux_tmp_37);
  assign result_and_3_cse = ccs_ccore_en & (and_dcpl_319 | and_dcpl_322 | and_dcpl_325
      | and_dcpl_329 | and_dcpl_333 | and_dcpl_337 | and_dcpl_341 | and_dcpl_344
      | and_dcpl_347 | mux_tmp_75);
  assign result_and_5_cse = ccs_ccore_en & (and_dcpl_353 | and_dcpl_357 | and_dcpl_361
      | and_dcpl_364 | and_dcpl_367 | and_dcpl_370 | and_dcpl_373 | and_dcpl_377
      | and_dcpl_381 | mux_tmp_113);
  assign result_and_7_cse = ccs_ccore_en & (and_dcpl_387 | and_dcpl_390 | and_dcpl_393
      | and_dcpl_396 | and_dcpl_399 | and_dcpl_402 | and_dcpl_405 | and_dcpl_408
      | and_dcpl_411 | mux_tmp_151);
  assign result_and_9_cse = ccs_ccore_en & (and_dcpl_418 | and_dcpl_422 | and_dcpl_426
      | and_dcpl_430 | and_dcpl_433 | and_dcpl_437 | and_dcpl_441 | and_dcpl_444
      | and_dcpl_447 | mux_tmp_189);
  assign result_and_11_cse = ccs_ccore_en & (and_dcpl_452 | and_dcpl_455 | and_dcpl_458
      | and_dcpl_462 | and_dcpl_464 | and_dcpl_468 | and_dcpl_472 | and_dcpl_474
      | and_dcpl_476 | mux_tmp_227);
  assign result_and_13_cse = ccs_ccore_en & (and_dcpl_480 | and_dcpl_484 | and_dcpl_488
      | and_dcpl_491 | and_dcpl_493 | and_dcpl_496 | and_dcpl_499 | and_dcpl_501
      | and_dcpl_503 | mux_tmp_265);
  assign result_and_15_cse = ccs_ccore_en & (and_dcpl_507 | and_dcpl_510 | and_dcpl_513
      | and_dcpl_516 | and_dcpl_518 | and_dcpl_521 | and_dcpl_524 | and_dcpl_526
      | and_dcpl_528 | mux_tmp_303);
  assign result_and_17_cse = ccs_ccore_en & (and_dcpl_533 | and_dcpl_536 | and_dcpl_539
      | and_dcpl_542 | and_dcpl_546 | and_dcpl_549 | and_dcpl_552 | and_dcpl_556
      | and_dcpl_560 | mux_tmp_348);
  assign result_and_19_cse = ccs_ccore_en & (and_dcpl_566 | and_dcpl_568 | and_dcpl_570
      | and_dcpl_572 | and_dcpl_576 | and_dcpl_578 | and_dcpl_580 | and_dcpl_583
      | and_dcpl_586 | mux_tmp_393);
  assign result_and_21_cse = ccs_ccore_en & (and_dcpl_590 | and_dcpl_592 | and_dcpl_594
      | and_dcpl_596 | and_dcpl_599 | and_dcpl_601 | and_dcpl_603 | and_dcpl_607
      | and_dcpl_611 | mux_tmp_438);
  assign m_and_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_2;
  assign m_and_1_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_6;
  assign m_and_2_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_9;
  assign m_and_3_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_11;
  assign m_and_4_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_2;
  assign m_and_5_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_6;
  assign m_and_6_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_9;
  assign m_and_7_cse = ccs_ccore_en & and_dcpl_13 & and_dcpl_11;
  assign m_and_8_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (~ (result_rem_11cyc_st_9[0]));
  assign m_and_9_cse = ccs_ccore_en & and_dcpl_4 & and_dcpl_18 & (result_rem_11cyc_st_9[0]);
  assign m_and_10_cse = ccs_ccore_en & and_dcpl_4 & (result_rem_11cyc_st_9[3]) &
      (result_rem_11cyc_st_9[1]) & (~ (result_rem_11cyc_st_9[0]));
  assign m_and_11_cse = ccs_ccore_en & and_dcpl_30;
  assign m_and_12_cse = ccs_ccore_en & and_dcpl_32;
  assign m_and_13_cse = ccs_ccore_en & and_dcpl_35;
  assign m_and_14_cse = ccs_ccore_en & and_dcpl_37;
  assign m_and_15_cse = ccs_ccore_en & and_dcpl_39;
  assign m_and_16_cse = ccs_ccore_en & and_dcpl_40;
  assign m_and_17_cse = ccs_ccore_en & and_dcpl_41;
  assign m_and_18_cse = ccs_ccore_en & and_dcpl_42;
  assign m_and_19_cse = ccs_ccore_en & and_dcpl_45;
  assign m_and_20_cse = ccs_ccore_en & and_dcpl_47;
  assign m_and_21_cse = ccs_ccore_en & and_dcpl_50;
  assign m_and_22_cse = ccs_ccore_en & and_dcpl_55;
  assign m_and_23_cse = ccs_ccore_en & and_dcpl_58;
  assign m_and_24_cse = ccs_ccore_en & and_dcpl_60;
  assign m_and_25_cse = ccs_ccore_en & and_dcpl_62;
  assign m_and_26_cse = ccs_ccore_en & and_dcpl_65;
  assign m_and_27_cse = ccs_ccore_en & and_dcpl_68;
  assign m_and_28_cse = ccs_ccore_en & and_dcpl_70;
  assign m_and_29_cse = ccs_ccore_en & and_dcpl_72;
  assign m_and_30_cse = ccs_ccore_en & and_dcpl_74;
  assign m_and_31_cse = ccs_ccore_en & and_dcpl_75;
  assign m_and_32_cse = ccs_ccore_en & and_dcpl_76;
  assign m_and_33_cse = ccs_ccore_en & and_dcpl_81;
  assign m_and_34_cse = ccs_ccore_en & and_dcpl_84;
  assign m_and_35_cse = ccs_ccore_en & and_dcpl_86;
  assign m_and_36_cse = ccs_ccore_en & and_dcpl_88;
  assign m_and_37_cse = ccs_ccore_en & and_dcpl_91;
  assign m_and_38_cse = ccs_ccore_en & and_dcpl_94;
  assign m_and_39_cse = ccs_ccore_en & and_dcpl_96;
  assign m_and_40_cse = ccs_ccore_en & and_dcpl_98;
  assign m_and_41_cse = ccs_ccore_en & and_dcpl_100;
  assign m_and_42_cse = ccs_ccore_en & and_dcpl_101;
  assign m_and_43_cse = ccs_ccore_en & and_dcpl_102;
  assign m_and_44_cse = ccs_ccore_en & and_dcpl_107;
  assign m_and_45_cse = ccs_ccore_en & and_dcpl_110;
  assign m_and_46_cse = ccs_ccore_en & and_dcpl_112;
  assign m_and_47_cse = ccs_ccore_en & and_dcpl_114;
  assign m_and_48_cse = ccs_ccore_en & and_dcpl_116;
  assign m_and_49_cse = ccs_ccore_en & and_dcpl_117;
  assign m_and_50_cse = ccs_ccore_en & and_dcpl_118;
  assign m_and_51_cse = ccs_ccore_en & and_dcpl_119;
  assign m_and_52_cse = ccs_ccore_en & and_dcpl_122;
  assign m_and_53_cse = ccs_ccore_en & and_dcpl_125;
  assign m_and_54_cse = ccs_ccore_en & and_dcpl_127;
  assign m_and_55_cse = ccs_ccore_en & and_dcpl_132;
  assign m_and_56_cse = ccs_ccore_en & and_dcpl_135;
  assign m_and_57_cse = ccs_ccore_en & and_dcpl_137;
  assign m_and_58_cse = ccs_ccore_en & and_dcpl_139;
  assign m_and_59_cse = ccs_ccore_en & and_dcpl_142;
  assign m_and_60_cse = ccs_ccore_en & and_dcpl_145;
  assign m_and_61_cse = ccs_ccore_en & and_dcpl_147;
  assign m_and_62_cse = ccs_ccore_en & and_dcpl_149;
  assign m_and_63_cse = ccs_ccore_en & and_dcpl_151;
  assign m_and_64_cse = ccs_ccore_en & and_dcpl_152;
  assign m_and_65_cse = ccs_ccore_en & and_dcpl_153;
  assign m_and_66_cse = ccs_ccore_en & and_dcpl_158;
  assign m_and_67_cse = ccs_ccore_en & and_dcpl_160;
  assign m_and_68_cse = ccs_ccore_en & and_dcpl_163;
  assign m_and_69_cse = ccs_ccore_en & and_dcpl_165;
  assign m_and_70_cse = ccs_ccore_en & and_dcpl_168;
  assign m_and_71_cse = ccs_ccore_en & and_dcpl_170;
  assign m_and_72_cse = ccs_ccore_en & and_dcpl_173;
  assign m_and_73_cse = ccs_ccore_en & and_dcpl_175;
  assign m_and_74_cse = ccs_ccore_en & and_dcpl_177;
  assign m_and_75_cse = ccs_ccore_en & and_dcpl_178;
  assign m_and_76_cse = ccs_ccore_en & and_dcpl_179;
  assign m_and_77_cse = ccs_ccore_en & and_dcpl_184;
  assign m_and_78_cse = ccs_ccore_en & and_dcpl_186;
  assign m_and_79_cse = ccs_ccore_en & and_dcpl_189;
  assign m_and_80_cse = ccs_ccore_en & and_dcpl_191;
  assign m_and_81_cse = ccs_ccore_en & and_dcpl_194;
  assign m_and_82_cse = ccs_ccore_en & and_dcpl_196;
  assign m_and_83_cse = ccs_ccore_en & and_dcpl_199;
  assign m_and_84_cse = ccs_ccore_en & and_dcpl_201;
  assign m_and_85_cse = ccs_ccore_en & and_dcpl_203;
  assign m_and_86_cse = ccs_ccore_en & and_dcpl_204;
  assign m_and_87_cse = ccs_ccore_en & and_dcpl_205;
  assign m_and_88_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_207;
  assign m_and_89_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_212;
  assign m_and_90_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_214;
  assign m_and_91_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_211 & (result_rem_11cyc[1]);
  assign m_and_92_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_218 & (~ (result_rem_11cyc[1]));
  assign m_and_93_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_221 & (~ (result_rem_11cyc[1]));
  assign m_and_94_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_218 & (result_rem_11cyc[1]);
  assign m_and_95_cse = ccs_ccore_en & and_dcpl_209 & and_dcpl_221 & (result_rem_11cyc[1]);
  assign m_and_96_cse = ccs_ccore_en & and_dcpl_228 & and_dcpl_207;
  assign m_and_97_cse = ccs_ccore_en & and_dcpl_228 & and_dcpl_212;
  assign m_and_98_cse = ccs_ccore_en & and_dcpl_228 & and_dcpl_214;
  assign nl_result_result_acc_tmp = conv_u2u_2_4(signext_2_1(result_acc_imod_1[3]))
      + conv_u2u_3_4(result_acc_imod_1[2:0]);
  assign result_result_acc_tmp = nl_result_result_acc_tmp[3:0];
  assign nl_result_acc_imod_1 = conv_u2s_3_4(result_acc_idiv_1[2:0]) + conv_u2s_3_4({(~
      (result_acc_idiv_1[3])) , 2'b00}) + conv_s2s_3_4({2'b10 , (result_acc_idiv_1[3])});
  assign result_acc_imod_1 = nl_result_acc_imod_1[3:0];
  assign nl_result_acc_idiv_1 = result_rem_11cyc + 4'b0001;
  assign result_acc_idiv_1 = nl_result_acc_idiv_1[3:0];
  assign and_dcpl_1 = ~((result_rem_11cyc_st_9[3]) | (result_rem_11cyc_st_9[1]));
  assign and_dcpl_2 = and_dcpl_1 & (~ (result_rem_11cyc_st_9[0]));
  assign and_dcpl_3 = main_stage_0_10 & asn_itm_9;
  assign and_dcpl_4 = and_dcpl_3 & (~ (result_rem_11cyc_st_9[2]));
  assign and_dcpl_6 = and_dcpl_1 & (result_rem_11cyc_st_9[0]);
  assign and_dcpl_8 = (~ (result_rem_11cyc_st_9[3])) & (result_rem_11cyc_st_9[1]);
  assign and_dcpl_9 = and_dcpl_8 & (~ (result_rem_11cyc_st_9[0]));
  assign and_dcpl_11 = and_dcpl_8 & (result_rem_11cyc_st_9[0]);
  assign and_dcpl_13 = and_dcpl_3 & (result_rem_11cyc_st_9[2]);
  assign and_dcpl_18 = (result_rem_11cyc_st_9[3]) & (~ (result_rem_11cyc_st_9[1]));
  assign and_dcpl_26 = ~((result_rem_11cyc_st_8[3]) | (result_rem_11cyc_st_8[1]));
  assign and_dcpl_27 = and_dcpl_26 & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_28 = main_stage_0_9 & asn_itm_8;
  assign and_dcpl_29 = and_dcpl_28 & (~ (result_rem_11cyc_st_8[2]));
  assign and_dcpl_30 = and_dcpl_29 & and_dcpl_27;
  assign and_dcpl_31 = and_dcpl_26 & (result_rem_11cyc_st_8[0]);
  assign and_dcpl_32 = and_dcpl_29 & and_dcpl_31;
  assign and_dcpl_33 = (~ (result_rem_11cyc_st_8[3])) & (result_rem_11cyc_st_8[1]);
  assign and_dcpl_34 = and_dcpl_33 & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_35 = and_dcpl_29 & and_dcpl_34;
  assign and_dcpl_36 = and_dcpl_33 & (result_rem_11cyc_st_8[0]);
  assign and_dcpl_37 = and_dcpl_29 & and_dcpl_36;
  assign and_dcpl_38 = and_dcpl_28 & (result_rem_11cyc_st_8[2]);
  assign and_dcpl_39 = and_dcpl_38 & and_dcpl_27;
  assign and_dcpl_40 = and_dcpl_38 & and_dcpl_31;
  assign and_dcpl_41 = and_dcpl_38 & and_dcpl_34;
  assign and_dcpl_42 = and_dcpl_38 & and_dcpl_36;
  assign and_dcpl_43 = (result_rem_11cyc_st_8[3]) & (~ (result_rem_11cyc_st_8[1]));
  assign and_dcpl_45 = and_dcpl_29 & and_dcpl_43 & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_47 = and_dcpl_29 & and_dcpl_43 & (result_rem_11cyc_st_8[0]);
  assign and_dcpl_50 = and_dcpl_29 & (result_rem_11cyc_st_8[3]) & (result_rem_11cyc_st_8[1])
      & (~ (result_rem_11cyc_st_8[0]));
  assign and_dcpl_51 = ~((result_rem_11cyc_st_7[2]) | (result_rem_11cyc_st_7[0]));
  assign and_dcpl_52 = and_dcpl_51 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_53 = main_stage_0_8 & asn_itm_7;
  assign and_dcpl_54 = and_dcpl_53 & (~ (result_rem_11cyc_st_7[3]));
  assign and_dcpl_55 = and_dcpl_54 & and_dcpl_52;
  assign and_dcpl_56 = (~ (result_rem_11cyc_st_7[2])) & (result_rem_11cyc_st_7[0]);
  assign and_dcpl_57 = and_dcpl_56 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_58 = and_dcpl_54 & and_dcpl_57;
  assign and_dcpl_59 = and_dcpl_51 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_60 = and_dcpl_54 & and_dcpl_59;
  assign and_dcpl_62 = and_dcpl_54 & and_dcpl_56 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_63 = (result_rem_11cyc_st_7[2]) & (~ (result_rem_11cyc_st_7[0]));
  assign and_dcpl_65 = and_dcpl_54 & and_dcpl_63 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_66 = (result_rem_11cyc_st_7[2]) & (result_rem_11cyc_st_7[0]);
  assign and_dcpl_68 = and_dcpl_54 & and_dcpl_66 & (~ (result_rem_11cyc_st_7[1]));
  assign and_dcpl_70 = and_dcpl_54 & and_dcpl_63 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_72 = and_dcpl_54 & and_dcpl_66 & (result_rem_11cyc_st_7[1]);
  assign and_dcpl_73 = and_dcpl_53 & (result_rem_11cyc_st_7[3]);
  assign and_dcpl_74 = and_dcpl_73 & and_dcpl_52;
  assign and_dcpl_75 = and_dcpl_73 & and_dcpl_57;
  assign and_dcpl_76 = and_dcpl_73 & and_dcpl_59;
  assign and_dcpl_77 = ~((result_rem_11cyc_st_6[2]) | (result_rem_11cyc_st_6[0]));
  assign and_dcpl_78 = and_dcpl_77 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_79 = main_stage_0_7 & asn_itm_6;
  assign and_dcpl_80 = and_dcpl_79 & (~ (result_rem_11cyc_st_6[3]));
  assign and_dcpl_81 = and_dcpl_80 & and_dcpl_78;
  assign and_dcpl_82 = (~ (result_rem_11cyc_st_6[2])) & (result_rem_11cyc_st_6[0]);
  assign and_dcpl_83 = and_dcpl_82 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_84 = and_dcpl_80 & and_dcpl_83;
  assign and_dcpl_85 = and_dcpl_77 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_86 = and_dcpl_80 & and_dcpl_85;
  assign and_dcpl_88 = and_dcpl_80 & and_dcpl_82 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_89 = (result_rem_11cyc_st_6[2]) & (~ (result_rem_11cyc_st_6[0]));
  assign and_dcpl_91 = and_dcpl_80 & and_dcpl_89 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_92 = (result_rem_11cyc_st_6[2]) & (result_rem_11cyc_st_6[0]);
  assign and_dcpl_94 = and_dcpl_80 & and_dcpl_92 & (~ (result_rem_11cyc_st_6[1]));
  assign and_dcpl_96 = and_dcpl_80 & and_dcpl_89 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_98 = and_dcpl_80 & and_dcpl_92 & (result_rem_11cyc_st_6[1]);
  assign and_dcpl_99 = and_dcpl_79 & (result_rem_11cyc_st_6[3]);
  assign and_dcpl_100 = and_dcpl_99 & and_dcpl_78;
  assign and_dcpl_101 = and_dcpl_99 & and_dcpl_83;
  assign and_dcpl_102 = and_dcpl_99 & and_dcpl_85;
  assign and_dcpl_103 = ~((result_rem_11cyc_st_5[3]) | (result_rem_11cyc_st_5[0]));
  assign and_dcpl_104 = and_dcpl_103 & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_105 = main_stage_0_6 & asn_itm_5;
  assign and_dcpl_106 = and_dcpl_105 & (~ (result_rem_11cyc_st_5[2]));
  assign and_dcpl_107 = and_dcpl_106 & and_dcpl_104;
  assign and_dcpl_108 = (~ (result_rem_11cyc_st_5[3])) & (result_rem_11cyc_st_5[0]);
  assign and_dcpl_109 = and_dcpl_108 & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_110 = and_dcpl_106 & and_dcpl_109;
  assign and_dcpl_111 = and_dcpl_103 & (result_rem_11cyc_st_5[1]);
  assign and_dcpl_112 = and_dcpl_106 & and_dcpl_111;
  assign and_dcpl_113 = and_dcpl_108 & (result_rem_11cyc_st_5[1]);
  assign and_dcpl_114 = and_dcpl_106 & and_dcpl_113;
  assign and_dcpl_115 = and_dcpl_105 & (result_rem_11cyc_st_5[2]);
  assign and_dcpl_116 = and_dcpl_115 & and_dcpl_104;
  assign and_dcpl_117 = and_dcpl_115 & and_dcpl_109;
  assign and_dcpl_118 = and_dcpl_115 & and_dcpl_111;
  assign and_dcpl_119 = and_dcpl_115 & and_dcpl_113;
  assign and_dcpl_120 = (result_rem_11cyc_st_5[3]) & (~ (result_rem_11cyc_st_5[0]));
  assign and_dcpl_122 = and_dcpl_106 & and_dcpl_120 & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_125 = and_dcpl_106 & (result_rem_11cyc_st_5[3]) & (result_rem_11cyc_st_5[0])
      & (~ (result_rem_11cyc_st_5[1]));
  assign and_dcpl_127 = and_dcpl_106 & and_dcpl_120 & (result_rem_11cyc_st_5[1]);
  assign and_dcpl_128 = ~((result_rem_11cyc_st_4[2]) | (result_rem_11cyc_st_4[0]));
  assign and_dcpl_129 = and_dcpl_128 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_130 = main_stage_0_5 & asn_itm_4;
  assign and_dcpl_131 = and_dcpl_130 & (~ (result_rem_11cyc_st_4[3]));
  assign and_dcpl_132 = and_dcpl_131 & and_dcpl_129;
  assign and_dcpl_133 = (~ (result_rem_11cyc_st_4[2])) & (result_rem_11cyc_st_4[0]);
  assign and_dcpl_134 = and_dcpl_133 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_135 = and_dcpl_131 & and_dcpl_134;
  assign and_dcpl_136 = and_dcpl_128 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_137 = and_dcpl_131 & and_dcpl_136;
  assign and_dcpl_139 = and_dcpl_131 & and_dcpl_133 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_140 = (result_rem_11cyc_st_4[2]) & (~ (result_rem_11cyc_st_4[0]));
  assign and_dcpl_142 = and_dcpl_131 & and_dcpl_140 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_143 = (result_rem_11cyc_st_4[2]) & (result_rem_11cyc_st_4[0]);
  assign and_dcpl_145 = and_dcpl_131 & and_dcpl_143 & (~ (result_rem_11cyc_st_4[1]));
  assign and_dcpl_147 = and_dcpl_131 & and_dcpl_140 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_149 = and_dcpl_131 & and_dcpl_143 & (result_rem_11cyc_st_4[1]);
  assign and_dcpl_150 = and_dcpl_130 & (result_rem_11cyc_st_4[3]);
  assign and_dcpl_151 = and_dcpl_150 & and_dcpl_129;
  assign and_dcpl_152 = and_dcpl_150 & and_dcpl_134;
  assign and_dcpl_153 = and_dcpl_150 & and_dcpl_136;
  assign and_dcpl_154 = ~((result_rem_11cyc_st_3[2:1]!=2'b00));
  assign and_dcpl_155 = and_dcpl_154 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_156 = main_stage_0_4 & asn_itm_3;
  assign and_dcpl_157 = and_dcpl_156 & (~ (result_rem_11cyc_st_3[3]));
  assign and_dcpl_158 = and_dcpl_157 & and_dcpl_155;
  assign and_dcpl_159 = and_dcpl_154 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_160 = and_dcpl_157 & and_dcpl_159;
  assign and_dcpl_161 = (result_rem_11cyc_st_3[2:1]==2'b01);
  assign and_dcpl_162 = and_dcpl_161 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_163 = and_dcpl_157 & and_dcpl_162;
  assign and_dcpl_165 = and_dcpl_157 & and_dcpl_161 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_166 = (result_rem_11cyc_st_3[2:1]==2'b10);
  assign and_dcpl_168 = and_dcpl_157 & and_dcpl_166 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_170 = and_dcpl_157 & and_dcpl_166 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_171 = (result_rem_11cyc_st_3[2:1]==2'b11);
  assign and_dcpl_173 = and_dcpl_157 & and_dcpl_171 & (~ (result_rem_11cyc_st_3[0]));
  assign and_dcpl_175 = and_dcpl_157 & and_dcpl_171 & (result_rem_11cyc_st_3[0]);
  assign and_dcpl_176 = and_dcpl_156 & (result_rem_11cyc_st_3[3]);
  assign and_dcpl_177 = and_dcpl_176 & and_dcpl_155;
  assign and_dcpl_178 = and_dcpl_176 & and_dcpl_159;
  assign and_dcpl_179 = and_dcpl_176 & and_dcpl_162;
  assign and_dcpl_180 = ~((result_rem_11cyc_st_2[2:1]!=2'b00));
  assign and_dcpl_181 = and_dcpl_180 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_182 = main_stage_0_3 & asn_itm_2;
  assign and_dcpl_183 = and_dcpl_182 & (~ (result_rem_11cyc_st_2[3]));
  assign and_dcpl_184 = and_dcpl_183 & and_dcpl_181;
  assign and_dcpl_185 = and_dcpl_180 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_186 = and_dcpl_183 & and_dcpl_185;
  assign and_dcpl_187 = (result_rem_11cyc_st_2[2:1]==2'b01);
  assign and_dcpl_188 = and_dcpl_187 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_189 = and_dcpl_183 & and_dcpl_188;
  assign and_dcpl_191 = and_dcpl_183 & and_dcpl_187 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_192 = (result_rem_11cyc_st_2[2:1]==2'b10);
  assign and_dcpl_194 = and_dcpl_183 & and_dcpl_192 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_196 = and_dcpl_183 & and_dcpl_192 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_197 = (result_rem_11cyc_st_2[2:1]==2'b11);
  assign and_dcpl_199 = and_dcpl_183 & and_dcpl_197 & (~ (result_rem_11cyc_st_2[0]));
  assign and_dcpl_201 = and_dcpl_183 & and_dcpl_197 & (result_rem_11cyc_st_2[0]);
  assign and_dcpl_202 = and_dcpl_182 & (result_rem_11cyc_st_2[3]);
  assign and_dcpl_203 = and_dcpl_202 & and_dcpl_181;
  assign and_dcpl_204 = and_dcpl_202 & and_dcpl_185;
  assign and_dcpl_205 = and_dcpl_202 & and_dcpl_188;
  assign and_dcpl_206 = ~((result_rem_11cyc[2]) | (result_rem_11cyc[0]));
  assign and_dcpl_207 = and_dcpl_206 & (~ (result_rem_11cyc[1]));
  assign and_dcpl_208 = main_stage_0_2 & asn_itm_1;
  assign and_dcpl_209 = and_dcpl_208 & (~ (result_rem_11cyc[3]));
  assign and_dcpl_211 = (~ (result_rem_11cyc[2])) & (result_rem_11cyc[0]);
  assign and_dcpl_212 = and_dcpl_211 & (~ (result_rem_11cyc[1]));
  assign and_dcpl_214 = and_dcpl_206 & (result_rem_11cyc[1]);
  assign and_dcpl_218 = (result_rem_11cyc[2]) & (~ (result_rem_11cyc[0]));
  assign and_dcpl_221 = (result_rem_11cyc[2]) & (result_rem_11cyc[0]);
  assign and_dcpl_228 = and_dcpl_208 & (result_rem_11cyc[3]);
  assign and_dcpl_232 = ~((result_rem_11cyc_st_11[2:1]!=2'b00));
  assign and_dcpl_233 = and_dcpl_232 & (~ (result_rem_11cyc_st_11[0]));
  assign and_dcpl_234 = main_stage_0_12 & asn_itm_11;
  assign and_dcpl_235 = and_dcpl_234 & (~ (result_rem_11cyc_st_11[3]));
  assign and_dcpl_237 = and_dcpl_232 & (result_rem_11cyc_st_11[0]);
  assign and_dcpl_239 = (result_rem_11cyc_st_11[2:1]==2'b01);
  assign and_dcpl_240 = and_dcpl_239 & (~ (result_rem_11cyc_st_11[0]));
  assign and_dcpl_244 = (result_rem_11cyc_st_11[2:1]==2'b10);
  assign and_dcpl_249 = (result_rem_11cyc_st_11[2:1]==2'b11);
  assign and_dcpl_254 = and_dcpl_234 & (result_rem_11cyc_st_11[3]);
  assign and_dcpl_260 = ~((result_result_acc_tmp[1:0]!=2'b00));
  assign and_dcpl_261 = ccs_ccore_start_rsci_idat & (~ (result_result_acc_tmp[2]));
  assign and_dcpl_262 = and_dcpl_261 & (~ (result_result_acc_tmp[3]));
  assign and_dcpl_263 = and_dcpl_262 & and_dcpl_260;
  assign or_tmp_2 = (result_rem_11cyc!=4'b0000) | (~ and_dcpl_208);
  assign or_3_cse = (result_result_acc_tmp!=4'b0000);
  assign nor_691_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_2));
  assign mux_nl = MUX_s_1_2_2(nor_691_nl, or_tmp_2, or_3_cse);
  assign and_dcpl_269 = mux_nl & and_dcpl_184;
  assign or_8_cse = (result_rem_11cyc!=4'b0000);
  assign nor_690_nl = ~(and_dcpl_208 | and_dcpl_184);
  assign or_10_nl = (result_rem_11cyc_st_2!=4'b0000) | (~ and_dcpl_182);
  assign mux_tmp_1 = MUX_s_1_2_2(nor_690_nl, or_10_nl, or_8_cse);
  assign nor_689_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_1));
  assign mux_2_nl = MUX_s_1_2_2(nor_689_nl, mux_tmp_1, or_3_cse);
  assign and_dcpl_275 = mux_2_nl & and_dcpl_158;
  assign or_15_cse = (result_rem_11cyc_st_2!=4'b0000);
  assign nor_687_nl = ~(and_dcpl_182 | and_dcpl_158);
  assign or_17_nl = (result_rem_11cyc_st_3!=4'b0000) | (~ and_dcpl_156);
  assign mux_tmp_3 = MUX_s_1_2_2(nor_687_nl, or_17_nl, or_15_cse);
  assign nor_688_nl = ~(and_dcpl_208 | (~ mux_tmp_3));
  assign mux_tmp_4 = MUX_s_1_2_2(nor_688_nl, mux_tmp_3, or_8_cse);
  assign nor_686_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_4));
  assign mux_5_nl = MUX_s_1_2_2(nor_686_nl, mux_tmp_4, or_3_cse);
  assign and_dcpl_281 = mux_5_nl & and_dcpl_132;
  assign or_24_cse = (result_rem_11cyc_st_3!=4'b0000);
  assign nor_683_nl = ~(and_dcpl_156 | and_dcpl_132);
  assign or_26_nl = (result_rem_11cyc_st_4!=4'b0000) | (~ and_dcpl_130);
  assign mux_tmp_6 = MUX_s_1_2_2(nor_683_nl, or_26_nl, or_24_cse);
  assign nor_684_nl = ~(and_dcpl_182 | (~ mux_tmp_6));
  assign mux_tmp_7 = MUX_s_1_2_2(nor_684_nl, mux_tmp_6, or_15_cse);
  assign nor_685_nl = ~(and_dcpl_208 | (~ mux_tmp_7));
  assign mux_tmp_8 = MUX_s_1_2_2(nor_685_nl, mux_tmp_7, or_8_cse);
  assign nor_682_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_8));
  assign mux_9_nl = MUX_s_1_2_2(nor_682_nl, mux_tmp_8, or_3_cse);
  assign and_dcpl_287 = mux_9_nl & and_dcpl_107;
  assign or_35_cse = (result_rem_11cyc_st_4!=4'b0000);
  assign nor_678_nl = ~(and_dcpl_130 | and_dcpl_107);
  assign or_37_nl = (result_rem_11cyc_st_5!=4'b0000) | (~ and_dcpl_105);
  assign mux_tmp_10 = MUX_s_1_2_2(nor_678_nl, or_37_nl, or_35_cse);
  assign nor_679_nl = ~(and_dcpl_156 | (~ mux_tmp_10));
  assign mux_tmp_11 = MUX_s_1_2_2(nor_679_nl, mux_tmp_10, or_24_cse);
  assign nor_680_nl = ~(and_dcpl_182 | (~ mux_tmp_11));
  assign mux_tmp_12 = MUX_s_1_2_2(nor_680_nl, mux_tmp_11, or_15_cse);
  assign nor_681_nl = ~(and_dcpl_208 | (~ mux_tmp_12));
  assign mux_tmp_13 = MUX_s_1_2_2(nor_681_nl, mux_tmp_12, or_8_cse);
  assign nor_677_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_13));
  assign mux_14_nl = MUX_s_1_2_2(nor_677_nl, mux_tmp_13, or_3_cse);
  assign and_dcpl_293 = mux_14_nl & and_dcpl_81;
  assign or_48_cse = (result_rem_11cyc_st_5!=4'b0000);
  assign nor_672_nl = ~(and_dcpl_105 | and_dcpl_81);
  assign or_50_nl = (result_rem_11cyc_st_6!=4'b0000) | (~ and_dcpl_79);
  assign mux_tmp_15 = MUX_s_1_2_2(nor_672_nl, or_50_nl, or_48_cse);
  assign nor_673_nl = ~(and_dcpl_130 | (~ mux_tmp_15));
  assign mux_tmp_16 = MUX_s_1_2_2(nor_673_nl, mux_tmp_15, or_35_cse);
  assign nor_674_nl = ~(and_dcpl_156 | (~ mux_tmp_16));
  assign mux_tmp_17 = MUX_s_1_2_2(nor_674_nl, mux_tmp_16, or_24_cse);
  assign nor_675_nl = ~(and_dcpl_182 | (~ mux_tmp_17));
  assign mux_tmp_18 = MUX_s_1_2_2(nor_675_nl, mux_tmp_17, or_15_cse);
  assign nor_676_nl = ~(and_dcpl_208 | (~ mux_tmp_18));
  assign mux_tmp_19 = MUX_s_1_2_2(nor_676_nl, mux_tmp_18, or_8_cse);
  assign nor_671_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_19));
  assign mux_20_nl = MUX_s_1_2_2(nor_671_nl, mux_tmp_19, or_3_cse);
  assign and_dcpl_299 = mux_20_nl & and_dcpl_55;
  assign or_63_cse = (result_rem_11cyc_st_6!=4'b0000);
  assign nor_665_nl = ~(and_dcpl_79 | and_dcpl_55);
  assign or_65_nl = (result_rem_11cyc_st_7!=4'b0000) | (~ and_dcpl_53);
  assign mux_tmp_21 = MUX_s_1_2_2(nor_665_nl, or_65_nl, or_63_cse);
  assign nor_666_nl = ~(and_dcpl_105 | (~ mux_tmp_21));
  assign mux_tmp_22 = MUX_s_1_2_2(nor_666_nl, mux_tmp_21, or_48_cse);
  assign nor_667_nl = ~(and_dcpl_130 | (~ mux_tmp_22));
  assign mux_tmp_23 = MUX_s_1_2_2(nor_667_nl, mux_tmp_22, or_35_cse);
  assign nor_668_nl = ~(and_dcpl_156 | (~ mux_tmp_23));
  assign mux_tmp_24 = MUX_s_1_2_2(nor_668_nl, mux_tmp_23, or_24_cse);
  assign nor_669_nl = ~(and_dcpl_182 | (~ mux_tmp_24));
  assign mux_tmp_25 = MUX_s_1_2_2(nor_669_nl, mux_tmp_24, or_15_cse);
  assign nor_670_nl = ~(and_dcpl_208 | (~ mux_tmp_25));
  assign mux_tmp_26 = MUX_s_1_2_2(nor_670_nl, mux_tmp_25, or_8_cse);
  assign nor_664_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_26));
  assign mux_27_nl = MUX_s_1_2_2(nor_664_nl, mux_tmp_26, or_3_cse);
  assign and_dcpl_305 = mux_27_nl & and_dcpl_30;
  assign nor_656_nl = ~(and_dcpl_53 | and_dcpl_30);
  assign or_82_nl = (result_rem_11cyc_st_8!=4'b0000) | (~ and_dcpl_28);
  assign or_80_nl = (result_rem_11cyc_st_7!=4'b0000);
  assign mux_tmp_28 = MUX_s_1_2_2(nor_656_nl, or_82_nl, or_80_nl);
  assign nor_657_nl = ~(and_dcpl_79 | (~ mux_tmp_28));
  assign mux_tmp_29 = MUX_s_1_2_2(nor_657_nl, mux_tmp_28, or_63_cse);
  assign nor_658_nl = ~(and_dcpl_105 | (~ mux_tmp_29));
  assign mux_tmp_30 = MUX_s_1_2_2(nor_658_nl, mux_tmp_29, or_48_cse);
  assign nor_659_nl = ~(and_dcpl_130 | (~ mux_tmp_30));
  assign mux_tmp_31 = MUX_s_1_2_2(nor_659_nl, mux_tmp_30, or_35_cse);
  assign nor_660_nl = ~(and_dcpl_156 | (~ mux_tmp_31));
  assign mux_tmp_32 = MUX_s_1_2_2(nor_660_nl, mux_tmp_31, or_24_cse);
  assign nor_661_nl = ~(and_dcpl_182 | (~ mux_tmp_32));
  assign mux_tmp_33 = MUX_s_1_2_2(nor_661_nl, mux_tmp_32, or_15_cse);
  assign nor_662_nl = ~(and_dcpl_208 | (~ mux_tmp_33));
  assign mux_tmp_34 = MUX_s_1_2_2(nor_662_nl, mux_tmp_33, or_8_cse);
  assign nor_663_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_34));
  assign mux_35_nl = MUX_s_1_2_2(nor_663_nl, mux_tmp_34, or_3_cse);
  assign and_dcpl_311 = mux_35_nl & and_dcpl_4 & and_dcpl_2;
  assign and_tmp_6 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0000))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0000)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0000)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0000)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0000)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0000)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0000)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0000));
  assign nor_654_nl = ~(and_dcpl_208 | (~ and_tmp_6));
  assign mux_tmp_36 = MUX_s_1_2_2(nor_654_nl, and_tmp_6, or_8_cse);
  assign nor_655_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_36));
  assign mux_tmp_37 = MUX_s_1_2_2(nor_655_nl, mux_tmp_36, or_3_cse);
  assign and_dcpl_318 = (result_result_acc_tmp[1:0]==2'b01);
  assign and_dcpl_319 = and_dcpl_262 & and_dcpl_318;
  assign or_tmp_102 = (result_rem_11cyc!=4'b0001) | (~ and_dcpl_208);
  assign or_107_cse = (result_result_acc_tmp!=4'b0001);
  assign nor_653_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_102));
  assign mux_38_nl = MUX_s_1_2_2(nor_653_nl, or_tmp_102, or_107_cse);
  assign and_dcpl_322 = mux_38_nl & and_dcpl_186;
  assign or_112_cse = (result_rem_11cyc!=4'b0001);
  assign nor_652_nl = ~(and_dcpl_208 | and_dcpl_186);
  assign or_114_nl = (result_rem_11cyc_st_2!=4'b0001) | (~ and_dcpl_182);
  assign mux_tmp_39 = MUX_s_1_2_2(nor_652_nl, or_114_nl, or_112_cse);
  assign nor_651_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_39));
  assign mux_40_nl = MUX_s_1_2_2(nor_651_nl, mux_tmp_39, or_107_cse);
  assign and_dcpl_325 = mux_40_nl & and_dcpl_160;
  assign or_119_cse = (result_rem_11cyc_st_2!=4'b0001);
  assign nor_649_nl = ~(and_dcpl_182 | and_dcpl_160);
  assign or_121_nl = (result_rem_11cyc_st_3!=4'b0001) | (~ and_dcpl_156);
  assign mux_tmp_41 = MUX_s_1_2_2(nor_649_nl, or_121_nl, or_119_cse);
  assign nor_650_nl = ~(and_dcpl_208 | (~ mux_tmp_41));
  assign mux_tmp_42 = MUX_s_1_2_2(nor_650_nl, mux_tmp_41, or_112_cse);
  assign nor_648_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_42));
  assign mux_43_nl = MUX_s_1_2_2(nor_648_nl, mux_tmp_42, or_107_cse);
  assign and_dcpl_329 = mux_43_nl & and_dcpl_135;
  assign or_128_cse = (result_rem_11cyc_st_3!=4'b0001);
  assign nor_645_nl = ~(and_dcpl_156 | and_dcpl_135);
  assign or_130_nl = (result_rem_11cyc_st_4!=4'b0001) | (~ and_dcpl_130);
  assign mux_tmp_44 = MUX_s_1_2_2(nor_645_nl, or_130_nl, or_128_cse);
  assign nor_646_nl = ~(and_dcpl_182 | (~ mux_tmp_44));
  assign mux_tmp_45 = MUX_s_1_2_2(nor_646_nl, mux_tmp_44, or_119_cse);
  assign nor_647_nl = ~(and_dcpl_208 | (~ mux_tmp_45));
  assign mux_tmp_46 = MUX_s_1_2_2(nor_647_nl, mux_tmp_45, or_112_cse);
  assign nor_644_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_46));
  assign mux_47_nl = MUX_s_1_2_2(nor_644_nl, mux_tmp_46, or_107_cse);
  assign and_dcpl_333 = mux_47_nl & and_dcpl_110;
  assign or_139_cse = (result_rem_11cyc_st_4!=4'b0001);
  assign nor_640_nl = ~(and_dcpl_130 | and_dcpl_110);
  assign or_141_nl = (result_rem_11cyc_st_5!=4'b0001) | (~ and_dcpl_105);
  assign mux_tmp_48 = MUX_s_1_2_2(nor_640_nl, or_141_nl, or_139_cse);
  assign nor_641_nl = ~(and_dcpl_156 | (~ mux_tmp_48));
  assign mux_tmp_49 = MUX_s_1_2_2(nor_641_nl, mux_tmp_48, or_128_cse);
  assign nor_642_nl = ~(and_dcpl_182 | (~ mux_tmp_49));
  assign mux_tmp_50 = MUX_s_1_2_2(nor_642_nl, mux_tmp_49, or_119_cse);
  assign nor_643_nl = ~(and_dcpl_208 | (~ mux_tmp_50));
  assign mux_tmp_51 = MUX_s_1_2_2(nor_643_nl, mux_tmp_50, or_112_cse);
  assign nor_639_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_51));
  assign mux_52_nl = MUX_s_1_2_2(nor_639_nl, mux_tmp_51, or_107_cse);
  assign and_dcpl_337 = mux_52_nl & and_dcpl_84;
  assign or_152_cse = (result_rem_11cyc_st_5!=4'b0001);
  assign nor_634_nl = ~(and_dcpl_105 | and_dcpl_84);
  assign or_154_nl = (result_rem_11cyc_st_6!=4'b0001) | (~ and_dcpl_79);
  assign mux_tmp_53 = MUX_s_1_2_2(nor_634_nl, or_154_nl, or_152_cse);
  assign nor_635_nl = ~(and_dcpl_130 | (~ mux_tmp_53));
  assign mux_tmp_54 = MUX_s_1_2_2(nor_635_nl, mux_tmp_53, or_139_cse);
  assign nor_636_nl = ~(and_dcpl_156 | (~ mux_tmp_54));
  assign mux_tmp_55 = MUX_s_1_2_2(nor_636_nl, mux_tmp_54, or_128_cse);
  assign nor_637_nl = ~(and_dcpl_182 | (~ mux_tmp_55));
  assign mux_tmp_56 = MUX_s_1_2_2(nor_637_nl, mux_tmp_55, or_119_cse);
  assign nor_638_nl = ~(and_dcpl_208 | (~ mux_tmp_56));
  assign mux_tmp_57 = MUX_s_1_2_2(nor_638_nl, mux_tmp_56, or_112_cse);
  assign nor_633_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_57));
  assign mux_58_nl = MUX_s_1_2_2(nor_633_nl, mux_tmp_57, or_107_cse);
  assign and_dcpl_341 = mux_58_nl & and_dcpl_58;
  assign or_167_cse = (result_rem_11cyc_st_6!=4'b0001);
  assign nor_627_nl = ~(and_dcpl_79 | and_dcpl_58);
  assign or_169_nl = (result_rem_11cyc_st_7!=4'b0001) | (~ and_dcpl_53);
  assign mux_tmp_59 = MUX_s_1_2_2(nor_627_nl, or_169_nl, or_167_cse);
  assign nor_628_nl = ~(and_dcpl_105 | (~ mux_tmp_59));
  assign mux_tmp_60 = MUX_s_1_2_2(nor_628_nl, mux_tmp_59, or_152_cse);
  assign nor_629_nl = ~(and_dcpl_130 | (~ mux_tmp_60));
  assign mux_tmp_61 = MUX_s_1_2_2(nor_629_nl, mux_tmp_60, or_139_cse);
  assign nor_630_nl = ~(and_dcpl_156 | (~ mux_tmp_61));
  assign mux_tmp_62 = MUX_s_1_2_2(nor_630_nl, mux_tmp_61, or_128_cse);
  assign nor_631_nl = ~(and_dcpl_182 | (~ mux_tmp_62));
  assign mux_tmp_63 = MUX_s_1_2_2(nor_631_nl, mux_tmp_62, or_119_cse);
  assign nor_632_nl = ~(and_dcpl_208 | (~ mux_tmp_63));
  assign mux_tmp_64 = MUX_s_1_2_2(nor_632_nl, mux_tmp_63, or_112_cse);
  assign nor_626_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_64));
  assign mux_65_nl = MUX_s_1_2_2(nor_626_nl, mux_tmp_64, or_107_cse);
  assign and_dcpl_344 = mux_65_nl & and_dcpl_32;
  assign nor_618_nl = ~(and_dcpl_53 | and_dcpl_32);
  assign or_186_nl = (result_rem_11cyc_st_8!=4'b0001) | (~ and_dcpl_28);
  assign or_184_nl = (result_rem_11cyc_st_7!=4'b0001);
  assign mux_tmp_66 = MUX_s_1_2_2(nor_618_nl, or_186_nl, or_184_nl);
  assign nor_619_nl = ~(and_dcpl_79 | (~ mux_tmp_66));
  assign mux_tmp_67 = MUX_s_1_2_2(nor_619_nl, mux_tmp_66, or_167_cse);
  assign nor_620_nl = ~(and_dcpl_105 | (~ mux_tmp_67));
  assign mux_tmp_68 = MUX_s_1_2_2(nor_620_nl, mux_tmp_67, or_152_cse);
  assign nor_621_nl = ~(and_dcpl_130 | (~ mux_tmp_68));
  assign mux_tmp_69 = MUX_s_1_2_2(nor_621_nl, mux_tmp_68, or_139_cse);
  assign nor_622_nl = ~(and_dcpl_156 | (~ mux_tmp_69));
  assign mux_tmp_70 = MUX_s_1_2_2(nor_622_nl, mux_tmp_69, or_128_cse);
  assign nor_623_nl = ~(and_dcpl_182 | (~ mux_tmp_70));
  assign mux_tmp_71 = MUX_s_1_2_2(nor_623_nl, mux_tmp_70, or_119_cse);
  assign nor_624_nl = ~(and_dcpl_208 | (~ mux_tmp_71));
  assign mux_tmp_72 = MUX_s_1_2_2(nor_624_nl, mux_tmp_71, or_112_cse);
  assign nor_625_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_72));
  assign mux_73_nl = MUX_s_1_2_2(nor_625_nl, mux_tmp_72, or_107_cse);
  assign and_dcpl_347 = mux_73_nl & and_dcpl_4 & and_dcpl_6;
  assign and_tmp_13 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0001))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0001)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0001)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0001)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0001)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0001)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0001)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0001));
  assign nor_617_nl = ~(and_dcpl_208 | (~ and_tmp_13));
  assign mux_tmp_74 = MUX_s_1_2_2(nor_617_nl, and_tmp_13, or_112_cse);
  assign nand_146_cse = ~((result_result_acc_tmp[0]) & ccs_ccore_start_rsci_idat);
  assign and_797_nl = nand_146_cse & mux_tmp_74;
  assign or_195_nl = (result_result_acc_tmp[3:1]!=3'b000);
  assign mux_tmp_75 = MUX_s_1_2_2(and_797_nl, mux_tmp_74, or_195_nl);
  assign and_dcpl_352 = (result_result_acc_tmp[1:0]==2'b10);
  assign and_dcpl_353 = and_dcpl_262 & and_dcpl_352;
  assign or_tmp_202 = (result_rem_11cyc!=4'b0010) | (~ and_dcpl_208);
  assign or_209_cse = (result_result_acc_tmp!=4'b0010);
  assign nor_616_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_202));
  assign mux_76_nl = MUX_s_1_2_2(nor_616_nl, or_tmp_202, or_209_cse);
  assign and_dcpl_357 = mux_76_nl & and_dcpl_189;
  assign or_214_cse = (result_rem_11cyc!=4'b0010);
  assign nor_615_nl = ~(and_dcpl_208 | and_dcpl_189);
  assign or_216_nl = (result_rem_11cyc_st_2!=4'b0010) | (~ and_dcpl_182);
  assign mux_tmp_77 = MUX_s_1_2_2(nor_615_nl, or_216_nl, or_214_cse);
  assign nor_614_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_77));
  assign mux_78_nl = MUX_s_1_2_2(nor_614_nl, mux_tmp_77, or_209_cse);
  assign and_dcpl_361 = mux_78_nl & and_dcpl_163;
  assign or_221_cse = (result_rem_11cyc_st_2!=4'b0010);
  assign nor_612_nl = ~(and_dcpl_182 | and_dcpl_163);
  assign or_223_nl = (result_rem_11cyc_st_3!=4'b0010) | (~ and_dcpl_156);
  assign mux_tmp_79 = MUX_s_1_2_2(nor_612_nl, or_223_nl, or_221_cse);
  assign nor_613_nl = ~(and_dcpl_208 | (~ mux_tmp_79));
  assign mux_tmp_80 = MUX_s_1_2_2(nor_613_nl, mux_tmp_79, or_214_cse);
  assign nor_611_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_80));
  assign mux_81_nl = MUX_s_1_2_2(nor_611_nl, mux_tmp_80, or_209_cse);
  assign and_dcpl_364 = mux_81_nl & and_dcpl_137;
  assign or_230_cse = (result_rem_11cyc_st_3!=4'b0010);
  assign nor_608_nl = ~(and_dcpl_156 | and_dcpl_137);
  assign or_232_nl = (result_rem_11cyc_st_4!=4'b0010) | (~ and_dcpl_130);
  assign mux_tmp_82 = MUX_s_1_2_2(nor_608_nl, or_232_nl, or_230_cse);
  assign nor_609_nl = ~(and_dcpl_182 | (~ mux_tmp_82));
  assign mux_tmp_83 = MUX_s_1_2_2(nor_609_nl, mux_tmp_82, or_221_cse);
  assign nor_610_nl = ~(and_dcpl_208 | (~ mux_tmp_83));
  assign mux_tmp_84 = MUX_s_1_2_2(nor_610_nl, mux_tmp_83, or_214_cse);
  assign nor_607_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_84));
  assign mux_85_nl = MUX_s_1_2_2(nor_607_nl, mux_tmp_84, or_209_cse);
  assign and_dcpl_367 = mux_85_nl & and_dcpl_112;
  assign or_241_cse = (result_rem_11cyc_st_4!=4'b0010);
  assign nor_603_nl = ~(and_dcpl_130 | and_dcpl_112);
  assign or_243_nl = (result_rem_11cyc_st_5!=4'b0010) | (~ and_dcpl_105);
  assign mux_tmp_86 = MUX_s_1_2_2(nor_603_nl, or_243_nl, or_241_cse);
  assign nor_604_nl = ~(and_dcpl_156 | (~ mux_tmp_86));
  assign mux_tmp_87 = MUX_s_1_2_2(nor_604_nl, mux_tmp_86, or_230_cse);
  assign nor_605_nl = ~(and_dcpl_182 | (~ mux_tmp_87));
  assign mux_tmp_88 = MUX_s_1_2_2(nor_605_nl, mux_tmp_87, or_221_cse);
  assign nor_606_nl = ~(and_dcpl_208 | (~ mux_tmp_88));
  assign mux_tmp_89 = MUX_s_1_2_2(nor_606_nl, mux_tmp_88, or_214_cse);
  assign nor_602_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_89));
  assign mux_90_nl = MUX_s_1_2_2(nor_602_nl, mux_tmp_89, or_209_cse);
  assign and_dcpl_370 = mux_90_nl & and_dcpl_86;
  assign or_254_cse = (result_rem_11cyc_st_5!=4'b0010);
  assign nor_597_nl = ~(and_dcpl_105 | and_dcpl_86);
  assign or_256_nl = (result_rem_11cyc_st_6!=4'b0010) | (~ and_dcpl_79);
  assign mux_tmp_91 = MUX_s_1_2_2(nor_597_nl, or_256_nl, or_254_cse);
  assign nor_598_nl = ~(and_dcpl_130 | (~ mux_tmp_91));
  assign mux_tmp_92 = MUX_s_1_2_2(nor_598_nl, mux_tmp_91, or_241_cse);
  assign nor_599_nl = ~(and_dcpl_156 | (~ mux_tmp_92));
  assign mux_tmp_93 = MUX_s_1_2_2(nor_599_nl, mux_tmp_92, or_230_cse);
  assign nor_600_nl = ~(and_dcpl_182 | (~ mux_tmp_93));
  assign mux_tmp_94 = MUX_s_1_2_2(nor_600_nl, mux_tmp_93, or_221_cse);
  assign nor_601_nl = ~(and_dcpl_208 | (~ mux_tmp_94));
  assign mux_tmp_95 = MUX_s_1_2_2(nor_601_nl, mux_tmp_94, or_214_cse);
  assign nor_596_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_95));
  assign mux_96_nl = MUX_s_1_2_2(nor_596_nl, mux_tmp_95, or_209_cse);
  assign and_dcpl_373 = mux_96_nl & and_dcpl_60;
  assign or_269_cse = (result_rem_11cyc_st_6!=4'b0010);
  assign nor_590_nl = ~(and_dcpl_79 | and_dcpl_60);
  assign or_271_nl = (result_rem_11cyc_st_7!=4'b0010) | (~ and_dcpl_53);
  assign mux_tmp_97 = MUX_s_1_2_2(nor_590_nl, or_271_nl, or_269_cse);
  assign nor_591_nl = ~(and_dcpl_105 | (~ mux_tmp_97));
  assign mux_tmp_98 = MUX_s_1_2_2(nor_591_nl, mux_tmp_97, or_254_cse);
  assign nor_592_nl = ~(and_dcpl_130 | (~ mux_tmp_98));
  assign mux_tmp_99 = MUX_s_1_2_2(nor_592_nl, mux_tmp_98, or_241_cse);
  assign nor_593_nl = ~(and_dcpl_156 | (~ mux_tmp_99));
  assign mux_tmp_100 = MUX_s_1_2_2(nor_593_nl, mux_tmp_99, or_230_cse);
  assign nor_594_nl = ~(and_dcpl_182 | (~ mux_tmp_100));
  assign mux_tmp_101 = MUX_s_1_2_2(nor_594_nl, mux_tmp_100, or_221_cse);
  assign nor_595_nl = ~(and_dcpl_208 | (~ mux_tmp_101));
  assign mux_tmp_102 = MUX_s_1_2_2(nor_595_nl, mux_tmp_101, or_214_cse);
  assign nor_589_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_102));
  assign mux_103_nl = MUX_s_1_2_2(nor_589_nl, mux_tmp_102, or_209_cse);
  assign and_dcpl_377 = mux_103_nl & and_dcpl_35;
  assign nor_581_nl = ~(and_dcpl_53 | and_dcpl_35);
  assign or_288_nl = (result_rem_11cyc_st_8!=4'b0010) | (~ and_dcpl_28);
  assign or_286_nl = (result_rem_11cyc_st_7!=4'b0010);
  assign mux_tmp_104 = MUX_s_1_2_2(nor_581_nl, or_288_nl, or_286_nl);
  assign nor_582_nl = ~(and_dcpl_79 | (~ mux_tmp_104));
  assign mux_tmp_105 = MUX_s_1_2_2(nor_582_nl, mux_tmp_104, or_269_cse);
  assign nor_583_nl = ~(and_dcpl_105 | (~ mux_tmp_105));
  assign mux_tmp_106 = MUX_s_1_2_2(nor_583_nl, mux_tmp_105, or_254_cse);
  assign nor_584_nl = ~(and_dcpl_130 | (~ mux_tmp_106));
  assign mux_tmp_107 = MUX_s_1_2_2(nor_584_nl, mux_tmp_106, or_241_cse);
  assign nor_585_nl = ~(and_dcpl_156 | (~ mux_tmp_107));
  assign mux_tmp_108 = MUX_s_1_2_2(nor_585_nl, mux_tmp_107, or_230_cse);
  assign nor_586_nl = ~(and_dcpl_182 | (~ mux_tmp_108));
  assign mux_tmp_109 = MUX_s_1_2_2(nor_586_nl, mux_tmp_108, or_221_cse);
  assign nor_587_nl = ~(and_dcpl_208 | (~ mux_tmp_109));
  assign mux_tmp_110 = MUX_s_1_2_2(nor_587_nl, mux_tmp_109, or_214_cse);
  assign nor_588_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_110));
  assign mux_111_nl = MUX_s_1_2_2(nor_588_nl, mux_tmp_110, or_209_cse);
  assign and_dcpl_381 = mux_111_nl & and_dcpl_4 & and_dcpl_9;
  assign and_tmp_20 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0010))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0010)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0010)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0010)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0010)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0010)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0010)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0010));
  assign nor_579_nl = ~(and_dcpl_208 | (~ and_tmp_20));
  assign mux_tmp_112 = MUX_s_1_2_2(nor_579_nl, and_tmp_20, or_214_cse);
  assign nor_580_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_112));
  assign mux_tmp_113 = MUX_s_1_2_2(nor_580_nl, mux_tmp_112, or_209_cse);
  assign and_dcpl_386 = (result_result_acc_tmp[1:0]==2'b11);
  assign and_dcpl_387 = and_dcpl_262 & and_dcpl_386;
  assign or_tmp_302 = (result_rem_11cyc!=4'b0011) | (~ and_dcpl_208);
  assign or_311_cse = (result_result_acc_tmp!=4'b0011);
  assign nor_578_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_302));
  assign mux_114_nl = MUX_s_1_2_2(nor_578_nl, or_tmp_302, or_311_cse);
  assign and_dcpl_390 = mux_114_nl & and_dcpl_191;
  assign or_316_cse = (result_rem_11cyc!=4'b0011);
  assign nor_577_nl = ~(and_dcpl_208 | and_dcpl_191);
  assign or_318_nl = (result_rem_11cyc_st_2!=4'b0011) | (~ and_dcpl_182);
  assign mux_tmp_115 = MUX_s_1_2_2(nor_577_nl, or_318_nl, or_316_cse);
  assign nor_576_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_115));
  assign mux_116_nl = MUX_s_1_2_2(nor_576_nl, mux_tmp_115, or_311_cse);
  assign and_dcpl_393 = mux_116_nl & and_dcpl_165;
  assign or_323_cse = (result_rem_11cyc_st_2!=4'b0011);
  assign nor_574_nl = ~(and_dcpl_182 | and_dcpl_165);
  assign or_325_nl = (result_rem_11cyc_st_3!=4'b0011) | (~ and_dcpl_156);
  assign mux_tmp_117 = MUX_s_1_2_2(nor_574_nl, or_325_nl, or_323_cse);
  assign nor_575_nl = ~(and_dcpl_208 | (~ mux_tmp_117));
  assign mux_tmp_118 = MUX_s_1_2_2(nor_575_nl, mux_tmp_117, or_316_cse);
  assign nor_573_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_118));
  assign mux_119_nl = MUX_s_1_2_2(nor_573_nl, mux_tmp_118, or_311_cse);
  assign and_dcpl_396 = mux_119_nl & and_dcpl_139;
  assign or_332_cse = (result_rem_11cyc_st_3!=4'b0011);
  assign nor_570_nl = ~(and_dcpl_156 | and_dcpl_139);
  assign or_334_nl = (result_rem_11cyc_st_4!=4'b0011) | (~ and_dcpl_130);
  assign mux_tmp_120 = MUX_s_1_2_2(nor_570_nl, or_334_nl, or_332_cse);
  assign nor_571_nl = ~(and_dcpl_182 | (~ mux_tmp_120));
  assign mux_tmp_121 = MUX_s_1_2_2(nor_571_nl, mux_tmp_120, or_323_cse);
  assign nor_572_nl = ~(and_dcpl_208 | (~ mux_tmp_121));
  assign mux_tmp_122 = MUX_s_1_2_2(nor_572_nl, mux_tmp_121, or_316_cse);
  assign nor_569_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_122));
  assign mux_123_nl = MUX_s_1_2_2(nor_569_nl, mux_tmp_122, or_311_cse);
  assign and_dcpl_399 = mux_123_nl & and_dcpl_114;
  assign or_343_cse = (result_rem_11cyc_st_4!=4'b0011);
  assign nor_565_nl = ~(and_dcpl_130 | and_dcpl_114);
  assign or_345_nl = (result_rem_11cyc_st_5!=4'b0011) | (~ and_dcpl_105);
  assign mux_tmp_124 = MUX_s_1_2_2(nor_565_nl, or_345_nl, or_343_cse);
  assign nor_566_nl = ~(and_dcpl_156 | (~ mux_tmp_124));
  assign mux_tmp_125 = MUX_s_1_2_2(nor_566_nl, mux_tmp_124, or_332_cse);
  assign nor_567_nl = ~(and_dcpl_182 | (~ mux_tmp_125));
  assign mux_tmp_126 = MUX_s_1_2_2(nor_567_nl, mux_tmp_125, or_323_cse);
  assign nor_568_nl = ~(and_dcpl_208 | (~ mux_tmp_126));
  assign mux_tmp_127 = MUX_s_1_2_2(nor_568_nl, mux_tmp_126, or_316_cse);
  assign nor_564_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_127));
  assign mux_128_nl = MUX_s_1_2_2(nor_564_nl, mux_tmp_127, or_311_cse);
  assign and_dcpl_402 = mux_128_nl & and_dcpl_88;
  assign or_356_cse = (result_rem_11cyc_st_5!=4'b0011);
  assign nor_559_nl = ~(and_dcpl_105 | and_dcpl_88);
  assign or_358_nl = (result_rem_11cyc_st_6!=4'b0011) | (~ and_dcpl_79);
  assign mux_tmp_129 = MUX_s_1_2_2(nor_559_nl, or_358_nl, or_356_cse);
  assign nor_560_nl = ~(and_dcpl_130 | (~ mux_tmp_129));
  assign mux_tmp_130 = MUX_s_1_2_2(nor_560_nl, mux_tmp_129, or_343_cse);
  assign nor_561_nl = ~(and_dcpl_156 | (~ mux_tmp_130));
  assign mux_tmp_131 = MUX_s_1_2_2(nor_561_nl, mux_tmp_130, or_332_cse);
  assign nor_562_nl = ~(and_dcpl_182 | (~ mux_tmp_131));
  assign mux_tmp_132 = MUX_s_1_2_2(nor_562_nl, mux_tmp_131, or_323_cse);
  assign nor_563_nl = ~(and_dcpl_208 | (~ mux_tmp_132));
  assign mux_tmp_133 = MUX_s_1_2_2(nor_563_nl, mux_tmp_132, or_316_cse);
  assign nor_558_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_133));
  assign mux_134_nl = MUX_s_1_2_2(nor_558_nl, mux_tmp_133, or_311_cse);
  assign and_dcpl_405 = mux_134_nl & and_dcpl_62;
  assign or_371_cse = (result_rem_11cyc_st_6!=4'b0011);
  assign nor_552_nl = ~(and_dcpl_79 | and_dcpl_62);
  assign or_373_nl = (result_rem_11cyc_st_7!=4'b0011) | (~ and_dcpl_53);
  assign mux_tmp_135 = MUX_s_1_2_2(nor_552_nl, or_373_nl, or_371_cse);
  assign nor_553_nl = ~(and_dcpl_105 | (~ mux_tmp_135));
  assign mux_tmp_136 = MUX_s_1_2_2(nor_553_nl, mux_tmp_135, or_356_cse);
  assign nor_554_nl = ~(and_dcpl_130 | (~ mux_tmp_136));
  assign mux_tmp_137 = MUX_s_1_2_2(nor_554_nl, mux_tmp_136, or_343_cse);
  assign nor_555_nl = ~(and_dcpl_156 | (~ mux_tmp_137));
  assign mux_tmp_138 = MUX_s_1_2_2(nor_555_nl, mux_tmp_137, or_332_cse);
  assign nor_556_nl = ~(and_dcpl_182 | (~ mux_tmp_138));
  assign mux_tmp_139 = MUX_s_1_2_2(nor_556_nl, mux_tmp_138, or_323_cse);
  assign nor_557_nl = ~(and_dcpl_208 | (~ mux_tmp_139));
  assign mux_tmp_140 = MUX_s_1_2_2(nor_557_nl, mux_tmp_139, or_316_cse);
  assign nor_551_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_140));
  assign mux_141_nl = MUX_s_1_2_2(nor_551_nl, mux_tmp_140, or_311_cse);
  assign and_dcpl_408 = mux_141_nl & and_dcpl_37;
  assign nor_543_nl = ~(and_dcpl_53 | and_dcpl_37);
  assign or_390_nl = (result_rem_11cyc_st_8!=4'b0011) | (~ and_dcpl_28);
  assign or_388_nl = (result_rem_11cyc_st_7!=4'b0011);
  assign mux_tmp_142 = MUX_s_1_2_2(nor_543_nl, or_390_nl, or_388_nl);
  assign nor_544_nl = ~(and_dcpl_79 | (~ mux_tmp_142));
  assign mux_tmp_143 = MUX_s_1_2_2(nor_544_nl, mux_tmp_142, or_371_cse);
  assign nor_545_nl = ~(and_dcpl_105 | (~ mux_tmp_143));
  assign mux_tmp_144 = MUX_s_1_2_2(nor_545_nl, mux_tmp_143, or_356_cse);
  assign nor_546_nl = ~(and_dcpl_130 | (~ mux_tmp_144));
  assign mux_tmp_145 = MUX_s_1_2_2(nor_546_nl, mux_tmp_144, or_343_cse);
  assign nor_547_nl = ~(and_dcpl_156 | (~ mux_tmp_145));
  assign mux_tmp_146 = MUX_s_1_2_2(nor_547_nl, mux_tmp_145, or_332_cse);
  assign nor_548_nl = ~(and_dcpl_182 | (~ mux_tmp_146));
  assign mux_tmp_147 = MUX_s_1_2_2(nor_548_nl, mux_tmp_146, or_323_cse);
  assign nor_549_nl = ~(and_dcpl_208 | (~ mux_tmp_147));
  assign mux_tmp_148 = MUX_s_1_2_2(nor_549_nl, mux_tmp_147, or_316_cse);
  assign nor_550_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_148));
  assign mux_149_nl = MUX_s_1_2_2(nor_550_nl, mux_tmp_148, or_311_cse);
  assign and_dcpl_411 = mux_149_nl & and_dcpl_4 & and_dcpl_11;
  assign and_tmp_27 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0011))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0011)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0011)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0011)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0011)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0011)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0011)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0011));
  assign nor_542_nl = ~(and_dcpl_208 | (~ and_tmp_27));
  assign mux_tmp_150 = MUX_s_1_2_2(nor_542_nl, and_tmp_27, or_316_cse);
  assign and_796_nl = (~((result_result_acc_tmp[1:0]==2'b11) & ccs_ccore_start_rsci_idat))
      & mux_tmp_150;
  assign or_399_nl = (result_result_acc_tmp[3:2]!=2'b00);
  assign mux_tmp_151 = MUX_s_1_2_2(and_796_nl, mux_tmp_150, or_399_nl);
  assign and_dcpl_417 = ccs_ccore_start_rsci_idat & (result_result_acc_tmp[3:2]==2'b01);
  assign and_dcpl_418 = and_dcpl_417 & and_dcpl_260;
  assign or_tmp_402 = (result_rem_11cyc!=4'b0100) | (~ and_dcpl_208);
  assign nand_144_cse = ~((result_result_acc_tmp[2]) & ccs_ccore_start_rsci_idat);
  assign or_413_cse = (result_result_acc_tmp[1]) | (result_result_acc_tmp[0]) | (result_result_acc_tmp[3]);
  assign and_795_nl = nand_144_cse & or_tmp_402;
  assign mux_152_nl = MUX_s_1_2_2(and_795_nl, or_tmp_402, or_413_cse);
  assign and_dcpl_422 = mux_152_nl & and_dcpl_194;
  assign or_418_cse = (result_rem_11cyc!=4'b0100);
  assign nor_541_nl = ~(and_dcpl_208 | and_dcpl_194);
  assign or_420_nl = (result_rem_11cyc_st_2!=4'b0100) | (~ and_dcpl_182);
  assign mux_tmp_153 = MUX_s_1_2_2(nor_541_nl, or_420_nl, or_418_cse);
  assign and_794_nl = nand_144_cse & mux_tmp_153;
  assign mux_154_nl = MUX_s_1_2_2(and_794_nl, mux_tmp_153, or_413_cse);
  assign and_dcpl_426 = mux_154_nl & and_dcpl_168;
  assign or_425_cse = (result_rem_11cyc_st_2!=4'b0100);
  assign nor_539_nl = ~(and_dcpl_182 | and_dcpl_168);
  assign or_427_nl = (result_rem_11cyc_st_3!=4'b0100) | (~ and_dcpl_156);
  assign mux_tmp_155 = MUX_s_1_2_2(nor_539_nl, or_427_nl, or_425_cse);
  assign nor_540_nl = ~(and_dcpl_208 | (~ mux_tmp_155));
  assign mux_tmp_156 = MUX_s_1_2_2(nor_540_nl, mux_tmp_155, or_418_cse);
  assign and_793_nl = nand_144_cse & mux_tmp_156;
  assign mux_157_nl = MUX_s_1_2_2(and_793_nl, mux_tmp_156, or_413_cse);
  assign and_dcpl_430 = mux_157_nl & and_dcpl_142;
  assign or_434_cse = (result_rem_11cyc_st_3!=4'b0100);
  assign nor_536_nl = ~(and_dcpl_156 | and_dcpl_142);
  assign or_436_nl = (result_rem_11cyc_st_4!=4'b0100) | (~ and_dcpl_130);
  assign mux_tmp_158 = MUX_s_1_2_2(nor_536_nl, or_436_nl, or_434_cse);
  assign nor_537_nl = ~(and_dcpl_182 | (~ mux_tmp_158));
  assign mux_tmp_159 = MUX_s_1_2_2(nor_537_nl, mux_tmp_158, or_425_cse);
  assign nor_538_nl = ~(and_dcpl_208 | (~ mux_tmp_159));
  assign mux_tmp_160 = MUX_s_1_2_2(nor_538_nl, mux_tmp_159, or_418_cse);
  assign and_792_nl = nand_144_cse & mux_tmp_160;
  assign mux_161_nl = MUX_s_1_2_2(and_792_nl, mux_tmp_160, or_413_cse);
  assign and_dcpl_433 = mux_161_nl & and_dcpl_116;
  assign or_445_cse = (result_rem_11cyc_st_4!=4'b0100);
  assign nor_532_nl = ~(and_dcpl_130 | and_dcpl_116);
  assign or_447_nl = (result_rem_11cyc_st_5[1]) | (result_rem_11cyc_st_5[0]) | (result_rem_11cyc_st_5[3])
      | (~ and_dcpl_115);
  assign mux_tmp_162 = MUX_s_1_2_2(nor_532_nl, or_447_nl, or_445_cse);
  assign nor_533_nl = ~(and_dcpl_156 | (~ mux_tmp_162));
  assign mux_tmp_163 = MUX_s_1_2_2(nor_533_nl, mux_tmp_162, or_434_cse);
  assign nor_534_nl = ~(and_dcpl_182 | (~ mux_tmp_163));
  assign mux_tmp_164 = MUX_s_1_2_2(nor_534_nl, mux_tmp_163, or_425_cse);
  assign nor_535_nl = ~(and_dcpl_208 | (~ mux_tmp_164));
  assign mux_tmp_165 = MUX_s_1_2_2(nor_535_nl, mux_tmp_164, or_418_cse);
  assign and_791_nl = nand_144_cse & mux_tmp_165;
  assign mux_166_nl = MUX_s_1_2_2(and_791_nl, mux_tmp_165, or_413_cse);
  assign and_dcpl_437 = mux_166_nl & and_dcpl_91;
  assign or_458_cse = (result_rem_11cyc_st_5[1]) | (result_rem_11cyc_st_5[0]) | (result_rem_11cyc_st_5[3]);
  assign and_790_cse = (result_rem_11cyc_st_5[2]) & asn_itm_5 & main_stage_0_6;
  assign nor_527_nl = ~(and_790_cse | and_dcpl_91);
  assign or_460_nl = (result_rem_11cyc_st_6!=4'b0100) | (~ and_dcpl_79);
  assign mux_tmp_167 = MUX_s_1_2_2(nor_527_nl, or_460_nl, or_458_cse);
  assign nor_528_nl = ~(and_dcpl_130 | (~ mux_tmp_167));
  assign mux_tmp_168 = MUX_s_1_2_2(nor_528_nl, mux_tmp_167, or_445_cse);
  assign nor_529_nl = ~(and_dcpl_156 | (~ mux_tmp_168));
  assign mux_tmp_169 = MUX_s_1_2_2(nor_529_nl, mux_tmp_168, or_434_cse);
  assign nor_530_nl = ~(and_dcpl_182 | (~ mux_tmp_169));
  assign mux_tmp_170 = MUX_s_1_2_2(nor_530_nl, mux_tmp_169, or_425_cse);
  assign nor_531_nl = ~(and_dcpl_208 | (~ mux_tmp_170));
  assign mux_tmp_171 = MUX_s_1_2_2(nor_531_nl, mux_tmp_170, or_418_cse);
  assign and_789_nl = nand_144_cse & mux_tmp_171;
  assign mux_172_nl = MUX_s_1_2_2(and_789_nl, mux_tmp_171, or_413_cse);
  assign and_dcpl_441 = mux_172_nl & and_dcpl_65;
  assign or_473_cse = (result_rem_11cyc_st_6!=4'b0100);
  assign nor_522_nl = ~(and_dcpl_79 | and_dcpl_65);
  assign or_475_nl = (result_rem_11cyc_st_7!=4'b0100) | (~ and_dcpl_53);
  assign mux_tmp_173 = MUX_s_1_2_2(nor_522_nl, or_475_nl, or_473_cse);
  assign nand_138_cse = ~((result_rem_11cyc_st_5[2]) & asn_itm_5 & main_stage_0_6);
  assign and_788_nl = nand_138_cse & mux_tmp_173;
  assign mux_tmp_174 = MUX_s_1_2_2(and_788_nl, mux_tmp_173, or_458_cse);
  assign nor_523_nl = ~(and_dcpl_130 | (~ mux_tmp_174));
  assign mux_tmp_175 = MUX_s_1_2_2(nor_523_nl, mux_tmp_174, or_445_cse);
  assign nor_524_nl = ~(and_dcpl_156 | (~ mux_tmp_175));
  assign mux_tmp_176 = MUX_s_1_2_2(nor_524_nl, mux_tmp_175, or_434_cse);
  assign nor_525_nl = ~(and_dcpl_182 | (~ mux_tmp_176));
  assign mux_tmp_177 = MUX_s_1_2_2(nor_525_nl, mux_tmp_176, or_425_cse);
  assign nor_526_nl = ~(and_dcpl_208 | (~ mux_tmp_177));
  assign mux_tmp_178 = MUX_s_1_2_2(nor_526_nl, mux_tmp_177, or_418_cse);
  assign and_787_nl = nand_144_cse & mux_tmp_178;
  assign mux_179_nl = MUX_s_1_2_2(and_787_nl, mux_tmp_178, or_413_cse);
  assign and_dcpl_444 = mux_179_nl & and_dcpl_39;
  assign nor_516_nl = ~(and_dcpl_53 | and_dcpl_39);
  assign or_492_nl = (result_rem_11cyc_st_8[0]) | (result_rem_11cyc_st_8[1]) | (result_rem_11cyc_st_8[3])
      | (~ and_dcpl_38);
  assign or_490_nl = (result_rem_11cyc_st_7!=4'b0100);
  assign mux_tmp_180 = MUX_s_1_2_2(nor_516_nl, or_492_nl, or_490_nl);
  assign nor_517_nl = ~(and_dcpl_79 | (~ mux_tmp_180));
  assign mux_tmp_181 = MUX_s_1_2_2(nor_517_nl, mux_tmp_180, or_473_cse);
  assign and_785_nl = nand_138_cse & mux_tmp_181;
  assign mux_tmp_182 = MUX_s_1_2_2(and_785_nl, mux_tmp_181, or_458_cse);
  assign nor_518_nl = ~(and_dcpl_130 | (~ mux_tmp_182));
  assign mux_tmp_183 = MUX_s_1_2_2(nor_518_nl, mux_tmp_182, or_445_cse);
  assign nor_519_nl = ~(and_dcpl_156 | (~ mux_tmp_183));
  assign mux_tmp_184 = MUX_s_1_2_2(nor_519_nl, mux_tmp_183, or_434_cse);
  assign nor_520_nl = ~(and_dcpl_182 | (~ mux_tmp_184));
  assign mux_tmp_185 = MUX_s_1_2_2(nor_520_nl, mux_tmp_184, or_425_cse);
  assign nor_521_nl = ~(and_dcpl_208 | (~ mux_tmp_185));
  assign mux_tmp_186 = MUX_s_1_2_2(nor_521_nl, mux_tmp_185, or_418_cse);
  assign and_786_nl = nand_144_cse & mux_tmp_186;
  assign mux_187_nl = MUX_s_1_2_2(and_786_nl, mux_tmp_186, or_413_cse);
  assign and_dcpl_447 = mux_187_nl & and_dcpl_13 & and_dcpl_2;
  assign and_tmp_34 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0100))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0100)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0100)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0100)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0100)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0100)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0100)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0100));
  assign nor_514_nl = ~(and_dcpl_208 | (~ and_tmp_34));
  assign mux_tmp_188 = MUX_s_1_2_2(nor_514_nl, and_tmp_34, or_418_cse);
  assign nor_515_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_188));
  assign or_501_nl = (result_result_acc_tmp!=4'b0100);
  assign mux_tmp_189 = MUX_s_1_2_2(nor_515_nl, mux_tmp_188, or_501_nl);
  assign and_dcpl_452 = and_dcpl_417 & and_dcpl_318;
  assign or_tmp_502 = (result_rem_11cyc!=4'b0101) | (~ and_dcpl_208);
  assign or_516_cse = (result_result_acc_tmp[1]) | (~ (result_result_acc_tmp[0]))
      | (result_result_acc_tmp[3]);
  assign and_784_nl = nand_144_cse & or_tmp_502;
  assign mux_190_nl = MUX_s_1_2_2(and_784_nl, or_tmp_502, or_516_cse);
  assign and_dcpl_455 = mux_190_nl & and_dcpl_196;
  assign or_521_cse = (result_rem_11cyc!=4'b0101);
  assign nor_513_nl = ~(and_dcpl_208 | and_dcpl_196);
  assign or_523_nl = (result_rem_11cyc_st_2!=4'b0101) | (~ and_dcpl_182);
  assign mux_tmp_191 = MUX_s_1_2_2(nor_513_nl, or_523_nl, or_521_cse);
  assign and_783_nl = nand_144_cse & mux_tmp_191;
  assign mux_192_nl = MUX_s_1_2_2(and_783_nl, mux_tmp_191, or_516_cse);
  assign and_dcpl_458 = mux_192_nl & and_dcpl_170;
  assign or_528_cse = (result_rem_11cyc_st_2!=4'b0101);
  assign nor_511_nl = ~(and_dcpl_182 | and_dcpl_170);
  assign or_530_nl = (result_rem_11cyc_st_3!=4'b0101) | (~ and_dcpl_156);
  assign mux_tmp_193 = MUX_s_1_2_2(nor_511_nl, or_530_nl, or_528_cse);
  assign nor_512_nl = ~(and_dcpl_208 | (~ mux_tmp_193));
  assign mux_tmp_194 = MUX_s_1_2_2(nor_512_nl, mux_tmp_193, or_521_cse);
  assign and_782_nl = nand_144_cse & mux_tmp_194;
  assign mux_195_nl = MUX_s_1_2_2(and_782_nl, mux_tmp_194, or_516_cse);
  assign and_dcpl_462 = mux_195_nl & and_dcpl_145;
  assign or_537_cse = (result_rem_11cyc_st_3!=4'b0101);
  assign nor_508_nl = ~(and_dcpl_156 | and_dcpl_145);
  assign or_539_nl = (result_rem_11cyc_st_4!=4'b0101) | (~ and_dcpl_130);
  assign mux_tmp_196 = MUX_s_1_2_2(nor_508_nl, or_539_nl, or_537_cse);
  assign nor_509_nl = ~(and_dcpl_182 | (~ mux_tmp_196));
  assign mux_tmp_197 = MUX_s_1_2_2(nor_509_nl, mux_tmp_196, or_528_cse);
  assign nor_510_nl = ~(and_dcpl_208 | (~ mux_tmp_197));
  assign mux_tmp_198 = MUX_s_1_2_2(nor_510_nl, mux_tmp_197, or_521_cse);
  assign and_781_nl = nand_144_cse & mux_tmp_198;
  assign mux_199_nl = MUX_s_1_2_2(and_781_nl, mux_tmp_198, or_516_cse);
  assign and_dcpl_464 = mux_199_nl & and_dcpl_117;
  assign or_548_cse = (result_rem_11cyc_st_4!=4'b0101);
  assign nor_504_nl = ~(and_dcpl_130 | and_dcpl_117);
  assign or_550_nl = (result_rem_11cyc_st_5[1]) | (~ (result_rem_11cyc_st_5[0]))
      | (result_rem_11cyc_st_5[3]) | (~ and_dcpl_115);
  assign mux_tmp_200 = MUX_s_1_2_2(nor_504_nl, or_550_nl, or_548_cse);
  assign nor_505_nl = ~(and_dcpl_156 | (~ mux_tmp_200));
  assign mux_tmp_201 = MUX_s_1_2_2(nor_505_nl, mux_tmp_200, or_537_cse);
  assign nor_506_nl = ~(and_dcpl_182 | (~ mux_tmp_201));
  assign mux_tmp_202 = MUX_s_1_2_2(nor_506_nl, mux_tmp_201, or_528_cse);
  assign nor_507_nl = ~(and_dcpl_208 | (~ mux_tmp_202));
  assign mux_tmp_203 = MUX_s_1_2_2(nor_507_nl, mux_tmp_202, or_521_cse);
  assign and_780_nl = nand_144_cse & mux_tmp_203;
  assign mux_204_nl = MUX_s_1_2_2(and_780_nl, mux_tmp_203, or_516_cse);
  assign and_dcpl_468 = mux_204_nl & and_dcpl_94;
  assign or_561_cse = (result_rem_11cyc_st_5[1]) | (~ (result_rem_11cyc_st_5[0]))
      | (result_rem_11cyc_st_5[3]);
  assign nor_499_nl = ~(and_790_cse | and_dcpl_94);
  assign or_563_nl = (result_rem_11cyc_st_6!=4'b0101) | (~ and_dcpl_79);
  assign mux_tmp_205 = MUX_s_1_2_2(nor_499_nl, or_563_nl, or_561_cse);
  assign nor_500_nl = ~(and_dcpl_130 | (~ mux_tmp_205));
  assign mux_tmp_206 = MUX_s_1_2_2(nor_500_nl, mux_tmp_205, or_548_cse);
  assign nor_501_nl = ~(and_dcpl_156 | (~ mux_tmp_206));
  assign mux_tmp_207 = MUX_s_1_2_2(nor_501_nl, mux_tmp_206, or_537_cse);
  assign nor_502_nl = ~(and_dcpl_182 | (~ mux_tmp_207));
  assign mux_tmp_208 = MUX_s_1_2_2(nor_502_nl, mux_tmp_207, or_528_cse);
  assign nor_503_nl = ~(and_dcpl_208 | (~ mux_tmp_208));
  assign mux_tmp_209 = MUX_s_1_2_2(nor_503_nl, mux_tmp_208, or_521_cse);
  assign and_778_nl = nand_144_cse & mux_tmp_209;
  assign mux_210_nl = MUX_s_1_2_2(and_778_nl, mux_tmp_209, or_516_cse);
  assign and_dcpl_472 = mux_210_nl & and_dcpl_68;
  assign or_576_cse = (result_rem_11cyc_st_6!=4'b0101);
  assign nor_494_nl = ~(and_dcpl_79 | and_dcpl_68);
  assign or_578_nl = (result_rem_11cyc_st_7!=4'b0101) | (~ and_dcpl_53);
  assign mux_tmp_211 = MUX_s_1_2_2(nor_494_nl, or_578_nl, or_576_cse);
  assign and_777_nl = nand_138_cse & mux_tmp_211;
  assign mux_tmp_212 = MUX_s_1_2_2(and_777_nl, mux_tmp_211, or_561_cse);
  assign nor_495_nl = ~(and_dcpl_130 | (~ mux_tmp_212));
  assign mux_tmp_213 = MUX_s_1_2_2(nor_495_nl, mux_tmp_212, or_548_cse);
  assign nor_496_nl = ~(and_dcpl_156 | (~ mux_tmp_213));
  assign mux_tmp_214 = MUX_s_1_2_2(nor_496_nl, mux_tmp_213, or_537_cse);
  assign nor_497_nl = ~(and_dcpl_182 | (~ mux_tmp_214));
  assign mux_tmp_215 = MUX_s_1_2_2(nor_497_nl, mux_tmp_214, or_528_cse);
  assign nor_498_nl = ~(and_dcpl_208 | (~ mux_tmp_215));
  assign mux_tmp_216 = MUX_s_1_2_2(nor_498_nl, mux_tmp_215, or_521_cse);
  assign and_776_nl = nand_144_cse & mux_tmp_216;
  assign mux_217_nl = MUX_s_1_2_2(and_776_nl, mux_tmp_216, or_516_cse);
  assign and_dcpl_474 = mux_217_nl & and_dcpl_40;
  assign nor_488_nl = ~(and_dcpl_53 | and_dcpl_40);
  assign or_595_nl = (~ (result_rem_11cyc_st_8[0])) | (result_rem_11cyc_st_8[1])
      | (result_rem_11cyc_st_8[3]) | (~ and_dcpl_38);
  assign or_593_nl = (result_rem_11cyc_st_7!=4'b0101);
  assign mux_tmp_218 = MUX_s_1_2_2(nor_488_nl, or_595_nl, or_593_nl);
  assign nor_489_nl = ~(and_dcpl_79 | (~ mux_tmp_218));
  assign mux_tmp_219 = MUX_s_1_2_2(nor_489_nl, mux_tmp_218, or_576_cse);
  assign and_774_nl = nand_138_cse & mux_tmp_219;
  assign mux_tmp_220 = MUX_s_1_2_2(and_774_nl, mux_tmp_219, or_561_cse);
  assign nor_490_nl = ~(and_dcpl_130 | (~ mux_tmp_220));
  assign mux_tmp_221 = MUX_s_1_2_2(nor_490_nl, mux_tmp_220, or_548_cse);
  assign nor_491_nl = ~(and_dcpl_156 | (~ mux_tmp_221));
  assign mux_tmp_222 = MUX_s_1_2_2(nor_491_nl, mux_tmp_221, or_537_cse);
  assign nor_492_nl = ~(and_dcpl_182 | (~ mux_tmp_222));
  assign mux_tmp_223 = MUX_s_1_2_2(nor_492_nl, mux_tmp_222, or_528_cse);
  assign nor_493_nl = ~(and_dcpl_208 | (~ mux_tmp_223));
  assign mux_tmp_224 = MUX_s_1_2_2(nor_493_nl, mux_tmp_223, or_521_cse);
  assign and_775_nl = nand_144_cse & mux_tmp_224;
  assign mux_225_nl = MUX_s_1_2_2(and_775_nl, mux_tmp_224, or_516_cse);
  assign and_dcpl_476 = mux_225_nl & and_dcpl_13 & and_dcpl_6;
  assign and_tmp_41 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0101))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0101)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0101)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0101)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0101)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0101)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0101)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0101));
  assign nor_487_nl = ~(and_dcpl_208 | (~ and_tmp_41));
  assign mux_tmp_226 = MUX_s_1_2_2(nor_487_nl, and_tmp_41, or_521_cse);
  assign and_773_nl = nand_146_cse & mux_tmp_226;
  assign or_604_nl = (result_result_acc_tmp[3:1]!=3'b010);
  assign mux_tmp_227 = MUX_s_1_2_2(and_773_nl, mux_tmp_226, or_604_nl);
  assign and_dcpl_480 = and_dcpl_417 & and_dcpl_352;
  assign or_tmp_602 = (result_rem_11cyc!=4'b0110) | (~ and_dcpl_208);
  assign or_617_cse = (~ (result_result_acc_tmp[1])) | (result_result_acc_tmp[0])
      | (result_result_acc_tmp[3]);
  assign and_772_nl = nand_144_cse & or_tmp_602;
  assign mux_228_nl = MUX_s_1_2_2(and_772_nl, or_tmp_602, or_617_cse);
  assign and_dcpl_484 = mux_228_nl & and_dcpl_199;
  assign or_622_cse = (result_rem_11cyc!=4'b0110);
  assign nor_486_nl = ~(and_dcpl_208 | and_dcpl_199);
  assign or_624_nl = (result_rem_11cyc_st_2!=4'b0110) | (~ and_dcpl_182);
  assign mux_tmp_229 = MUX_s_1_2_2(nor_486_nl, or_624_nl, or_622_cse);
  assign and_771_nl = nand_144_cse & mux_tmp_229;
  assign mux_230_nl = MUX_s_1_2_2(and_771_nl, mux_tmp_229, or_617_cse);
  assign and_dcpl_488 = mux_230_nl & and_dcpl_173;
  assign or_629_cse = (result_rem_11cyc_st_2!=4'b0110);
  assign nor_484_nl = ~(and_dcpl_182 | and_dcpl_173);
  assign or_631_nl = (result_rem_11cyc_st_3!=4'b0110) | (~ and_dcpl_156);
  assign mux_tmp_231 = MUX_s_1_2_2(nor_484_nl, or_631_nl, or_629_cse);
  assign nor_485_nl = ~(and_dcpl_208 | (~ mux_tmp_231));
  assign mux_tmp_232 = MUX_s_1_2_2(nor_485_nl, mux_tmp_231, or_622_cse);
  assign and_770_nl = nand_144_cse & mux_tmp_232;
  assign mux_233_nl = MUX_s_1_2_2(and_770_nl, mux_tmp_232, or_617_cse);
  assign and_dcpl_491 = mux_233_nl & and_dcpl_147;
  assign or_638_cse = (result_rem_11cyc_st_3!=4'b0110);
  assign nor_481_nl = ~(and_dcpl_156 | and_dcpl_147);
  assign or_640_nl = (result_rem_11cyc_st_4!=4'b0110) | (~ and_dcpl_130);
  assign mux_tmp_234 = MUX_s_1_2_2(nor_481_nl, or_640_nl, or_638_cse);
  assign nor_482_nl = ~(and_dcpl_182 | (~ mux_tmp_234));
  assign mux_tmp_235 = MUX_s_1_2_2(nor_482_nl, mux_tmp_234, or_629_cse);
  assign nor_483_nl = ~(and_dcpl_208 | (~ mux_tmp_235));
  assign mux_tmp_236 = MUX_s_1_2_2(nor_483_nl, mux_tmp_235, or_622_cse);
  assign and_769_nl = nand_144_cse & mux_tmp_236;
  assign mux_237_nl = MUX_s_1_2_2(and_769_nl, mux_tmp_236, or_617_cse);
  assign and_dcpl_493 = mux_237_nl & and_dcpl_118;
  assign or_649_cse = (result_rem_11cyc_st_4!=4'b0110);
  assign nor_477_nl = ~(and_dcpl_130 | and_dcpl_118);
  assign or_651_nl = (~ (result_rem_11cyc_st_5[1])) | (result_rem_11cyc_st_5[0])
      | (result_rem_11cyc_st_5[3]) | (~ and_dcpl_115);
  assign mux_tmp_238 = MUX_s_1_2_2(nor_477_nl, or_651_nl, or_649_cse);
  assign nor_478_nl = ~(and_dcpl_156 | (~ mux_tmp_238));
  assign mux_tmp_239 = MUX_s_1_2_2(nor_478_nl, mux_tmp_238, or_638_cse);
  assign nor_479_nl = ~(and_dcpl_182 | (~ mux_tmp_239));
  assign mux_tmp_240 = MUX_s_1_2_2(nor_479_nl, mux_tmp_239, or_629_cse);
  assign nor_480_nl = ~(and_dcpl_208 | (~ mux_tmp_240));
  assign mux_tmp_241 = MUX_s_1_2_2(nor_480_nl, mux_tmp_240, or_622_cse);
  assign and_768_nl = nand_144_cse & mux_tmp_241;
  assign mux_242_nl = MUX_s_1_2_2(and_768_nl, mux_tmp_241, or_617_cse);
  assign and_dcpl_496 = mux_242_nl & and_dcpl_96;
  assign or_662_cse = (~ (result_rem_11cyc_st_5[1])) | (result_rem_11cyc_st_5[0])
      | (result_rem_11cyc_st_5[3]);
  assign nor_472_nl = ~(and_790_cse | and_dcpl_96);
  assign or_664_nl = (result_rem_11cyc_st_6!=4'b0110) | (~ and_dcpl_79);
  assign mux_tmp_243 = MUX_s_1_2_2(nor_472_nl, or_664_nl, or_662_cse);
  assign nor_473_nl = ~(and_dcpl_130 | (~ mux_tmp_243));
  assign mux_tmp_244 = MUX_s_1_2_2(nor_473_nl, mux_tmp_243, or_649_cse);
  assign nor_474_nl = ~(and_dcpl_156 | (~ mux_tmp_244));
  assign mux_tmp_245 = MUX_s_1_2_2(nor_474_nl, mux_tmp_244, or_638_cse);
  assign nor_475_nl = ~(and_dcpl_182 | (~ mux_tmp_245));
  assign mux_tmp_246 = MUX_s_1_2_2(nor_475_nl, mux_tmp_245, or_629_cse);
  assign nor_476_nl = ~(and_dcpl_208 | (~ mux_tmp_246));
  assign mux_tmp_247 = MUX_s_1_2_2(nor_476_nl, mux_tmp_246, or_622_cse);
  assign and_766_nl = nand_144_cse & mux_tmp_247;
  assign mux_248_nl = MUX_s_1_2_2(and_766_nl, mux_tmp_247, or_617_cse);
  assign and_dcpl_499 = mux_248_nl & and_dcpl_70;
  assign or_677_cse = (result_rem_11cyc_st_6!=4'b0110);
  assign nor_467_nl = ~(and_dcpl_79 | and_dcpl_70);
  assign or_679_nl = (result_rem_11cyc_st_7!=4'b0110) | (~ and_dcpl_53);
  assign mux_tmp_249 = MUX_s_1_2_2(nor_467_nl, or_679_nl, or_677_cse);
  assign and_765_nl = nand_138_cse & mux_tmp_249;
  assign mux_tmp_250 = MUX_s_1_2_2(and_765_nl, mux_tmp_249, or_662_cse);
  assign nor_468_nl = ~(and_dcpl_130 | (~ mux_tmp_250));
  assign mux_tmp_251 = MUX_s_1_2_2(nor_468_nl, mux_tmp_250, or_649_cse);
  assign nor_469_nl = ~(and_dcpl_156 | (~ mux_tmp_251));
  assign mux_tmp_252 = MUX_s_1_2_2(nor_469_nl, mux_tmp_251, or_638_cse);
  assign nor_470_nl = ~(and_dcpl_182 | (~ mux_tmp_252));
  assign mux_tmp_253 = MUX_s_1_2_2(nor_470_nl, mux_tmp_252, or_629_cse);
  assign nor_471_nl = ~(and_dcpl_208 | (~ mux_tmp_253));
  assign mux_tmp_254 = MUX_s_1_2_2(nor_471_nl, mux_tmp_253, or_622_cse);
  assign and_764_nl = nand_144_cse & mux_tmp_254;
  assign mux_255_nl = MUX_s_1_2_2(and_764_nl, mux_tmp_254, or_617_cse);
  assign and_dcpl_501 = mux_255_nl & and_dcpl_41;
  assign nor_461_nl = ~(and_dcpl_53 | and_dcpl_41);
  assign or_696_nl = (result_rem_11cyc_st_8[0]) | (~ (result_rem_11cyc_st_8[1]))
      | (result_rem_11cyc_st_8[3]) | (~ and_dcpl_38);
  assign or_694_nl = (result_rem_11cyc_st_7!=4'b0110);
  assign mux_tmp_256 = MUX_s_1_2_2(nor_461_nl, or_696_nl, or_694_nl);
  assign nor_462_nl = ~(and_dcpl_79 | (~ mux_tmp_256));
  assign mux_tmp_257 = MUX_s_1_2_2(nor_462_nl, mux_tmp_256, or_677_cse);
  assign and_762_nl = nand_138_cse & mux_tmp_257;
  assign mux_tmp_258 = MUX_s_1_2_2(and_762_nl, mux_tmp_257, or_662_cse);
  assign nor_463_nl = ~(and_dcpl_130 | (~ mux_tmp_258));
  assign mux_tmp_259 = MUX_s_1_2_2(nor_463_nl, mux_tmp_258, or_649_cse);
  assign nor_464_nl = ~(and_dcpl_156 | (~ mux_tmp_259));
  assign mux_tmp_260 = MUX_s_1_2_2(nor_464_nl, mux_tmp_259, or_638_cse);
  assign nor_465_nl = ~(and_dcpl_182 | (~ mux_tmp_260));
  assign mux_tmp_261 = MUX_s_1_2_2(nor_465_nl, mux_tmp_260, or_629_cse);
  assign nor_466_nl = ~(and_dcpl_208 | (~ mux_tmp_261));
  assign mux_tmp_262 = MUX_s_1_2_2(nor_466_nl, mux_tmp_261, or_622_cse);
  assign and_763_nl = nand_144_cse & mux_tmp_262;
  assign mux_263_nl = MUX_s_1_2_2(and_763_nl, mux_tmp_262, or_617_cse);
  assign and_dcpl_503 = mux_263_nl & and_dcpl_13 & and_dcpl_9;
  assign and_tmp_48 = ((~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2!=4'b0110))
      & ((~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3!=4'b0110)) &
      ((~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4!=4'b0110)) & ((~
      main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5!=4'b0110)) & ((~ main_stage_0_7)
      | (~ asn_itm_6) | (result_rem_11cyc_st_6!=4'b0110)) & ((~ main_stage_0_8) |
      (~ asn_itm_7) | (result_rem_11cyc_st_7!=4'b0110)) & ((~ main_stage_0_9) | (~
      asn_itm_8) | (result_rem_11cyc_st_8!=4'b0110)) & ((~ main_stage_0_10) | (~
      asn_itm_9) | (result_rem_11cyc_st_9!=4'b0110));
  assign nor_459_nl = ~(and_dcpl_208 | (~ and_tmp_48));
  assign mux_tmp_264 = MUX_s_1_2_2(nor_459_nl, and_tmp_48, or_622_cse);
  assign nor_460_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_264));
  assign or_705_nl = (result_result_acc_tmp!=4'b0110);
  assign mux_tmp_265 = MUX_s_1_2_2(nor_460_nl, mux_tmp_264, or_705_nl);
  assign and_dcpl_507 = and_dcpl_417 & and_dcpl_386;
  assign or_tmp_702 = ~((result_rem_11cyc==4'b0111) & and_dcpl_208);
  assign or_718_cse = (~ (result_result_acc_tmp[1])) | (~ (result_result_acc_tmp[0]))
      | (result_result_acc_tmp[3]);
  assign and_761_nl = nand_144_cse & or_tmp_702;
  assign mux_266_nl = MUX_s_1_2_2(and_761_nl, or_tmp_702, or_718_cse);
  assign and_dcpl_510 = mux_266_nl & and_dcpl_201;
  assign nand_112_cse = ~((result_rem_11cyc==4'b0111));
  assign nor_458_nl = ~(and_dcpl_208 | and_dcpl_201);
  assign nand_153_nl = ~((result_rem_11cyc_st_2==4'b0111) & and_dcpl_182);
  assign mux_tmp_267 = MUX_s_1_2_2(nor_458_nl, nand_153_nl, nand_112_cse);
  assign and_760_nl = nand_144_cse & mux_tmp_267;
  assign mux_268_nl = MUX_s_1_2_2(and_760_nl, mux_tmp_267, or_718_cse);
  assign and_dcpl_513 = mux_268_nl & and_dcpl_175;
  assign nand_108_cse = ~((result_rem_11cyc_st_2==4'b0111));
  assign nor_456_nl = ~(and_dcpl_182 | and_dcpl_175);
  assign nand_152_nl = ~((result_rem_11cyc_st_3==4'b0111) & and_dcpl_156);
  assign mux_tmp_269 = MUX_s_1_2_2(nor_456_nl, nand_152_nl, nand_108_cse);
  assign nor_457_nl = ~(and_dcpl_208 | (~ mux_tmp_269));
  assign mux_tmp_270 = MUX_s_1_2_2(nor_457_nl, mux_tmp_269, nand_112_cse);
  assign and_759_nl = nand_144_cse & mux_tmp_270;
  assign mux_271_nl = MUX_s_1_2_2(and_759_nl, mux_tmp_270, or_718_cse);
  assign and_dcpl_516 = mux_271_nl & and_dcpl_149;
  assign nand_103_cse = ~((result_rem_11cyc_st_3==4'b0111));
  assign nor_453_nl = ~(and_dcpl_156 | and_dcpl_149);
  assign nand_151_nl = ~((result_rem_11cyc_st_4==4'b0111) & and_dcpl_130);
  assign mux_tmp_272 = MUX_s_1_2_2(nor_453_nl, nand_151_nl, nand_103_cse);
  assign nor_454_nl = ~(and_dcpl_182 | (~ mux_tmp_272));
  assign mux_tmp_273 = MUX_s_1_2_2(nor_454_nl, mux_tmp_272, nand_108_cse);
  assign nor_455_nl = ~(and_dcpl_208 | (~ mux_tmp_273));
  assign mux_tmp_274 = MUX_s_1_2_2(nor_455_nl, mux_tmp_273, nand_112_cse);
  assign and_758_nl = nand_144_cse & mux_tmp_274;
  assign mux_275_nl = MUX_s_1_2_2(and_758_nl, mux_tmp_274, or_718_cse);
  assign and_dcpl_518 = mux_275_nl & and_dcpl_119;
  assign nand_97_cse = ~((result_rem_11cyc_st_4==4'b0111));
  assign nor_449_nl = ~(and_dcpl_130 | and_dcpl_119);
  assign nand_96_nl = ~((result_rem_11cyc_st_5[1]) & (result_rem_11cyc_st_5[0]) &
      (~ (result_rem_11cyc_st_5[3])) & and_dcpl_115);
  assign mux_tmp_276 = MUX_s_1_2_2(nor_449_nl, nand_96_nl, nand_97_cse);
  assign nor_450_nl = ~(and_dcpl_156 | (~ mux_tmp_276));
  assign mux_tmp_277 = MUX_s_1_2_2(nor_450_nl, mux_tmp_276, nand_103_cse);
  assign nor_451_nl = ~(and_dcpl_182 | (~ mux_tmp_277));
  assign mux_tmp_278 = MUX_s_1_2_2(nor_451_nl, mux_tmp_277, nand_108_cse);
  assign nor_452_nl = ~(and_dcpl_208 | (~ mux_tmp_278));
  assign mux_tmp_279 = MUX_s_1_2_2(nor_452_nl, mux_tmp_278, nand_112_cse);
  assign and_757_nl = nand_144_cse & mux_tmp_279;
  assign mux_280_nl = MUX_s_1_2_2(and_757_nl, mux_tmp_279, or_718_cse);
  assign and_dcpl_521 = mux_280_nl & and_dcpl_98;
  assign or_763_cse = (~ (result_rem_11cyc_st_5[1])) | (~ (result_rem_11cyc_st_5[0]))
      | (result_rem_11cyc_st_5[3]);
  assign nor_444_nl = ~(and_790_cse | and_dcpl_98);
  assign nand_150_nl = ~((result_rem_11cyc_st_6==4'b0111) & and_dcpl_79);
  assign mux_tmp_281 = MUX_s_1_2_2(nor_444_nl, nand_150_nl, or_763_cse);
  assign nor_445_nl = ~(and_dcpl_130 | (~ mux_tmp_281));
  assign mux_tmp_282 = MUX_s_1_2_2(nor_445_nl, mux_tmp_281, nand_97_cse);
  assign nor_446_nl = ~(and_dcpl_156 | (~ mux_tmp_282));
  assign mux_tmp_283 = MUX_s_1_2_2(nor_446_nl, mux_tmp_282, nand_103_cse);
  assign nor_447_nl = ~(and_dcpl_182 | (~ mux_tmp_283));
  assign mux_tmp_284 = MUX_s_1_2_2(nor_447_nl, mux_tmp_283, nand_108_cse);
  assign nor_448_nl = ~(and_dcpl_208 | (~ mux_tmp_284));
  assign mux_tmp_285 = MUX_s_1_2_2(nor_448_nl, mux_tmp_284, nand_112_cse);
  assign and_755_nl = nand_144_cse & mux_tmp_285;
  assign mux_286_nl = MUX_s_1_2_2(and_755_nl, mux_tmp_285, or_718_cse);
  assign and_dcpl_524 = mux_286_nl & and_dcpl_72;
  assign nand_83_cse = ~((result_rem_11cyc_st_6==4'b0111));
  assign nor_439_nl = ~(and_dcpl_79 | and_dcpl_72);
  assign nand_149_nl = ~((result_rem_11cyc_st_7==4'b0111) & and_dcpl_53);
  assign mux_tmp_287 = MUX_s_1_2_2(nor_439_nl, nand_149_nl, nand_83_cse);
  assign and_754_nl = nand_138_cse & mux_tmp_287;
  assign mux_tmp_288 = MUX_s_1_2_2(and_754_nl, mux_tmp_287, or_763_cse);
  assign nor_440_nl = ~(and_dcpl_130 | (~ mux_tmp_288));
  assign mux_tmp_289 = MUX_s_1_2_2(nor_440_nl, mux_tmp_288, nand_97_cse);
  assign nor_441_nl = ~(and_dcpl_156 | (~ mux_tmp_289));
  assign mux_tmp_290 = MUX_s_1_2_2(nor_441_nl, mux_tmp_289, nand_103_cse);
  assign nor_442_nl = ~(and_dcpl_182 | (~ mux_tmp_290));
  assign mux_tmp_291 = MUX_s_1_2_2(nor_442_nl, mux_tmp_290, nand_108_cse);
  assign nor_443_nl = ~(and_dcpl_208 | (~ mux_tmp_291));
  assign mux_tmp_292 = MUX_s_1_2_2(nor_443_nl, mux_tmp_291, nand_112_cse);
  assign and_753_nl = nand_144_cse & mux_tmp_292;
  assign mux_293_nl = MUX_s_1_2_2(and_753_nl, mux_tmp_292, or_718_cse);
  assign and_dcpl_526 = mux_293_nl & and_dcpl_42;
  assign nor_433_nl = ~(and_dcpl_53 | and_dcpl_42);
  assign nand_72_nl = ~((result_rem_11cyc_st_8[0]) & (result_rem_11cyc_st_8[1]) &
      (~ (result_rem_11cyc_st_8[3])) & and_dcpl_38);
  assign nand_73_nl = ~((result_rem_11cyc_st_7==4'b0111));
  assign mux_tmp_294 = MUX_s_1_2_2(nor_433_nl, nand_72_nl, nand_73_nl);
  assign nor_434_nl = ~(and_dcpl_79 | (~ mux_tmp_294));
  assign mux_tmp_295 = MUX_s_1_2_2(nor_434_nl, mux_tmp_294, nand_83_cse);
  assign and_751_nl = nand_138_cse & mux_tmp_295;
  assign mux_tmp_296 = MUX_s_1_2_2(and_751_nl, mux_tmp_295, or_763_cse);
  assign nor_435_nl = ~(and_dcpl_130 | (~ mux_tmp_296));
  assign mux_tmp_297 = MUX_s_1_2_2(nor_435_nl, mux_tmp_296, nand_97_cse);
  assign nor_436_nl = ~(and_dcpl_156 | (~ mux_tmp_297));
  assign mux_tmp_298 = MUX_s_1_2_2(nor_436_nl, mux_tmp_297, nand_103_cse);
  assign nor_437_nl = ~(and_dcpl_182 | (~ mux_tmp_298));
  assign mux_tmp_299 = MUX_s_1_2_2(nor_437_nl, mux_tmp_298, nand_108_cse);
  assign nor_438_nl = ~(and_dcpl_208 | (~ mux_tmp_299));
  assign mux_tmp_300 = MUX_s_1_2_2(nor_438_nl, mux_tmp_299, nand_112_cse);
  assign and_752_nl = nand_144_cse & mux_tmp_300;
  assign mux_301_nl = MUX_s_1_2_2(and_752_nl, mux_tmp_300, or_718_cse);
  assign and_dcpl_528 = mux_301_nl & and_dcpl_13 & and_dcpl_11;
  assign and_tmp_55 = (~(main_stage_0_3 & asn_itm_2 & (result_rem_11cyc_st_2==4'b0111)))
      & (~(main_stage_0_4 & asn_itm_3 & (result_rem_11cyc_st_3==4'b0111))) & (~(main_stage_0_5
      & asn_itm_4 & (result_rem_11cyc_st_4==4'b0111))) & (~(main_stage_0_6 & asn_itm_5
      & (result_rem_11cyc_st_5==4'b0111))) & (~(main_stage_0_7 & asn_itm_6 & (result_rem_11cyc_st_6==4'b0111)))
      & (~(main_stage_0_8 & asn_itm_7 & (result_rem_11cyc_st_7==4'b0111))) & (~(main_stage_0_9
      & asn_itm_8 & (result_rem_11cyc_st_8==4'b0111))) & (~(main_stage_0_10 & asn_itm_9
      & (result_rem_11cyc_st_9==4'b0111)));
  assign nor_432_nl = ~(and_dcpl_208 | (~ and_tmp_55));
  assign mux_tmp_302 = MUX_s_1_2_2(nor_432_nl, and_tmp_55, nand_112_cse);
  assign and_750_nl = (~((result_result_acc_tmp[2:0]==3'b111) & ccs_ccore_start_rsci_idat))
      & mux_tmp_302;
  assign mux_tmp_303 = MUX_s_1_2_2(and_750_nl, mux_tmp_302, result_result_acc_tmp[3]);
  assign and_dcpl_532 = and_dcpl_261 & (result_result_acc_tmp[3]);
  assign and_dcpl_533 = and_dcpl_532 & and_dcpl_260;
  assign not_tmp_645 = ~((result_rem_11cyc[3]) & asn_itm_1 & main_stage_0_2);
  assign or_tmp_801 = (result_rem_11cyc[2:0]!=3'b000) | not_tmp_645;
  assign or_818_cse = (result_result_acc_tmp!=4'b1000);
  assign nor_431_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_801));
  assign mux_304_nl = MUX_s_1_2_2(nor_431_nl, or_tmp_801, or_818_cse);
  assign and_dcpl_536 = mux_304_nl & and_dcpl_203;
  assign or_823_cse = (result_rem_11cyc[2:0]!=3'b000);
  assign and_749_cse = (result_rem_11cyc[3]) & asn_itm_1 & main_stage_0_2;
  assign nor_430_nl = ~(and_749_cse | and_dcpl_203);
  assign or_825_nl = (result_rem_11cyc_st_2[2:0]!=3'b000) | (~ and_dcpl_202);
  assign mux_tmp_305 = MUX_s_1_2_2(nor_430_nl, or_825_nl, or_823_cse);
  assign nor_429_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_305));
  assign mux_306_nl = MUX_s_1_2_2(nor_429_nl, mux_tmp_305, or_818_cse);
  assign and_dcpl_539 = mux_306_nl & and_dcpl_177;
  assign or_830_cse = (result_rem_11cyc_st_2[2:0]!=3'b000);
  assign and_747_cse = (result_rem_11cyc_st_2[3]) & asn_itm_2 & main_stage_0_3;
  assign nor_428_nl = ~(and_747_cse | and_dcpl_177);
  assign or_832_nl = (result_rem_11cyc_st_3[2:0]!=3'b000) | (~ and_dcpl_176);
  assign mux_tmp_307 = MUX_s_1_2_2(nor_428_nl, or_832_nl, or_830_cse);
  assign and_748_nl = not_tmp_645 & mux_tmp_307;
  assign mux_tmp_308 = MUX_s_1_2_2(and_748_nl, mux_tmp_307, or_823_cse);
  assign nor_427_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_308));
  assign mux_309_nl = MUX_s_1_2_2(nor_427_nl, mux_tmp_308, or_818_cse);
  assign and_dcpl_542 = mux_309_nl & and_dcpl_151;
  assign or_839_cse = (result_rem_11cyc_st_3[2:0]!=3'b000);
  assign and_744_cse = (result_rem_11cyc_st_3[3]) & asn_itm_3 & main_stage_0_4;
  assign nor_426_nl = ~(and_744_cse | and_dcpl_151);
  assign or_841_nl = (result_rem_11cyc_st_4[2:0]!=3'b000) | (~ and_dcpl_150);
  assign mux_tmp_310 = MUX_s_1_2_2(nor_426_nl, or_841_nl, or_839_cse);
  assign nand_58_cse = ~((result_rem_11cyc_st_2[3]) & asn_itm_2 & main_stage_0_3);
  assign and_745_nl = nand_58_cse & mux_tmp_310;
  assign mux_tmp_311 = MUX_s_1_2_2(and_745_nl, mux_tmp_310, or_830_cse);
  assign and_746_nl = not_tmp_645 & mux_tmp_311;
  assign mux_tmp_312 = MUX_s_1_2_2(and_746_nl, mux_tmp_311, or_823_cse);
  assign nor_425_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_312));
  assign mux_313_nl = MUX_s_1_2_2(nor_425_nl, mux_tmp_312, or_818_cse);
  assign and_dcpl_546 = mux_313_nl & and_dcpl_122;
  assign or_850_cse = (result_rem_11cyc_st_4[2:0]!=3'b000);
  assign and_740_cse = (result_rem_11cyc_st_4[3]) & asn_itm_4 & main_stage_0_5;
  assign nor_424_nl = ~(and_740_cse | and_dcpl_122);
  assign or_852_nl = (result_rem_11cyc_st_5!=4'b1000) | (~ and_dcpl_105);
  assign mux_tmp_314 = MUX_s_1_2_2(nor_424_nl, or_852_nl, or_850_cse);
  assign nand_55_cse = ~((result_rem_11cyc_st_3[3]) & asn_itm_3 & main_stage_0_4);
  assign and_741_nl = nand_55_cse & mux_tmp_314;
  assign mux_tmp_315 = MUX_s_1_2_2(and_741_nl, mux_tmp_314, or_839_cse);
  assign and_742_nl = nand_58_cse & mux_tmp_315;
  assign mux_tmp_316 = MUX_s_1_2_2(and_742_nl, mux_tmp_315, or_830_cse);
  assign and_743_nl = not_tmp_645 & mux_tmp_316;
  assign mux_tmp_317 = MUX_s_1_2_2(and_743_nl, mux_tmp_316, or_823_cse);
  assign nor_423_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_317));
  assign mux_318_nl = MUX_s_1_2_2(nor_423_nl, mux_tmp_317, or_818_cse);
  assign and_dcpl_549 = mux_318_nl & and_dcpl_100;
  assign or_863_cse = (result_rem_11cyc_st_5!=4'b1000);
  assign nor_422_nl = ~(and_dcpl_105 | and_dcpl_100);
  assign or_865_nl = (result_rem_11cyc_st_6[2:0]!=3'b000) | (~ and_dcpl_99);
  assign mux_tmp_319 = MUX_s_1_2_2(nor_422_nl, or_865_nl, or_863_cse);
  assign nand_51_cse = ~((result_rem_11cyc_st_4[3]) & asn_itm_4 & main_stage_0_5);
  assign and_736_nl = nand_51_cse & mux_tmp_319;
  assign mux_tmp_320 = MUX_s_1_2_2(and_736_nl, mux_tmp_319, or_850_cse);
  assign and_737_nl = nand_55_cse & mux_tmp_320;
  assign mux_tmp_321 = MUX_s_1_2_2(and_737_nl, mux_tmp_320, or_839_cse);
  assign and_738_nl = nand_58_cse & mux_tmp_321;
  assign mux_tmp_322 = MUX_s_1_2_2(and_738_nl, mux_tmp_321, or_830_cse);
  assign and_739_nl = not_tmp_645 & mux_tmp_322;
  assign mux_tmp_323 = MUX_s_1_2_2(and_739_nl, mux_tmp_322, or_823_cse);
  assign nor_421_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_323));
  assign mux_324_nl = MUX_s_1_2_2(nor_421_nl, mux_tmp_323, or_818_cse);
  assign and_dcpl_552 = mux_324_nl & and_dcpl_74;
  assign or_878_cse = (result_rem_11cyc_st_6[2:0]!=3'b000);
  assign and_731_cse = (result_rem_11cyc_st_6[3]) & asn_itm_6 & main_stage_0_7;
  assign nor_419_nl = ~(and_731_cse | and_dcpl_74);
  assign or_880_nl = (result_rem_11cyc_st_7[2:0]!=3'b000) | (~ and_dcpl_73);
  assign mux_tmp_325 = MUX_s_1_2_2(nor_419_nl, or_880_nl, or_878_cse);
  assign nor_420_nl = ~(and_dcpl_105 | (~ mux_tmp_325));
  assign mux_tmp_326 = MUX_s_1_2_2(nor_420_nl, mux_tmp_325, or_863_cse);
  assign and_732_nl = nand_51_cse & mux_tmp_326;
  assign mux_tmp_327 = MUX_s_1_2_2(and_732_nl, mux_tmp_326, or_850_cse);
  assign and_733_nl = nand_55_cse & mux_tmp_327;
  assign mux_tmp_328 = MUX_s_1_2_2(and_733_nl, mux_tmp_327, or_839_cse);
  assign and_734_nl = nand_58_cse & mux_tmp_328;
  assign mux_tmp_329 = MUX_s_1_2_2(and_734_nl, mux_tmp_328, or_830_cse);
  assign and_735_nl = not_tmp_645 & mux_tmp_329;
  assign mux_tmp_330 = MUX_s_1_2_2(and_735_nl, mux_tmp_329, or_823_cse);
  assign nor_418_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_330));
  assign mux_331_nl = MUX_s_1_2_2(nor_418_nl, mux_tmp_330, or_818_cse);
  assign and_dcpl_556 = mux_331_nl & and_dcpl_45;
  assign and_725_cse = (result_rem_11cyc_st_7[3]) & asn_itm_7 & main_stage_0_8;
  assign nor_415_nl = ~(and_725_cse | and_dcpl_45);
  assign or_897_nl = (result_rem_11cyc_st_8!=4'b1000) | (~ and_dcpl_28);
  assign or_895_nl = (result_rem_11cyc_st_7[2:0]!=3'b000);
  assign mux_tmp_332 = MUX_s_1_2_2(nor_415_nl, or_897_nl, or_895_nl);
  assign nand_42_cse = ~((result_rem_11cyc_st_6[3]) & asn_itm_6 & main_stage_0_7);
  assign and_726_nl = nand_42_cse & mux_tmp_332;
  assign mux_tmp_333 = MUX_s_1_2_2(and_726_nl, mux_tmp_332, or_878_cse);
  assign nor_416_nl = ~(and_dcpl_105 | (~ mux_tmp_333));
  assign mux_tmp_334 = MUX_s_1_2_2(nor_416_nl, mux_tmp_333, or_863_cse);
  assign and_727_nl = nand_51_cse & mux_tmp_334;
  assign mux_tmp_335 = MUX_s_1_2_2(and_727_nl, mux_tmp_334, or_850_cse);
  assign and_728_nl = nand_55_cse & mux_tmp_335;
  assign mux_tmp_336 = MUX_s_1_2_2(and_728_nl, mux_tmp_335, or_839_cse);
  assign and_729_nl = nand_58_cse & mux_tmp_336;
  assign mux_tmp_337 = MUX_s_1_2_2(and_729_nl, mux_tmp_336, or_830_cse);
  assign and_730_nl = not_tmp_645 & mux_tmp_337;
  assign mux_tmp_338 = MUX_s_1_2_2(and_730_nl, mux_tmp_337, or_823_cse);
  assign nor_417_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_338));
  assign mux_339_nl = MUX_s_1_2_2(nor_417_nl, mux_tmp_338, or_818_cse);
  assign and_dcpl_560 = mux_339_nl & and_dcpl_4 & and_dcpl_18 & (~ (result_rem_11cyc_st_9[0]));
  assign or_tmp_897 = (~ main_stage_0_10) | (~ asn_itm_9) | (result_rem_11cyc_st_9!=4'b1000);
  assign nor_407_nl = ~((result_rem_11cyc_st_8[3]) | (~ or_tmp_897));
  assign or_914_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (result_rem_11cyc_st_8[2:0]!=3'b000);
  assign mux_tmp_340 = MUX_s_1_2_2(nor_407_nl, or_tmp_897, or_914_nl);
  assign nor_408_nl = ~((result_rem_11cyc_st_7[3]) | (~ mux_tmp_340));
  assign or_913_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (result_rem_11cyc_st_7[2:0]!=3'b000);
  assign mux_tmp_341 = MUX_s_1_2_2(nor_408_nl, mux_tmp_340, or_913_nl);
  assign nor_409_nl = ~((result_rem_11cyc_st_6[3]) | (~ mux_tmp_341));
  assign or_912_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (result_rem_11cyc_st_6[2:0]!=3'b000);
  assign mux_tmp_342 = MUX_s_1_2_2(nor_409_nl, mux_tmp_341, or_912_nl);
  assign nor_410_nl = ~((result_rem_11cyc_st_5[3]) | (~ mux_tmp_342));
  assign or_911_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5[2:0]!=3'b000);
  assign mux_tmp_343 = MUX_s_1_2_2(nor_410_nl, mux_tmp_342, or_911_nl);
  assign nor_411_nl = ~((result_rem_11cyc_st_4[3]) | (~ mux_tmp_343));
  assign or_910_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4[2:0]!=3'b000);
  assign mux_tmp_344 = MUX_s_1_2_2(nor_411_nl, mux_tmp_343, or_910_nl);
  assign nor_412_nl = ~((result_rem_11cyc_st_3[3]) | (~ mux_tmp_344));
  assign or_909_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3[2:0]!=3'b000);
  assign mux_tmp_345 = MUX_s_1_2_2(nor_412_nl, mux_tmp_344, or_909_nl);
  assign nor_413_nl = ~((result_rem_11cyc_st_2[3]) | (~ mux_tmp_345));
  assign or_908_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2[2:0]!=3'b000);
  assign mux_tmp_346 = MUX_s_1_2_2(nor_413_nl, mux_tmp_345, or_908_nl);
  assign and_724_nl = not_tmp_645 & mux_tmp_346;
  assign mux_tmp_347 = MUX_s_1_2_2(and_724_nl, mux_tmp_346, or_823_cse);
  assign nor_414_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_347));
  assign mux_tmp_348 = MUX_s_1_2_2(nor_414_nl, mux_tmp_347, or_818_cse);
  assign and_dcpl_566 = and_dcpl_532 & and_dcpl_318;
  assign or_tmp_909 = (result_rem_11cyc[2:0]!=3'b001) | not_tmp_645;
  assign or_928_cse = (result_result_acc_tmp!=4'b1001);
  assign nor_406_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_909));
  assign mux_349_nl = MUX_s_1_2_2(nor_406_nl, or_tmp_909, or_928_cse);
  assign and_dcpl_568 = mux_349_nl & and_dcpl_204;
  assign or_933_cse = (result_rem_11cyc[2:0]!=3'b001);
  assign nor_405_nl = ~(and_749_cse | and_dcpl_204);
  assign or_935_nl = (result_rem_11cyc_st_2[2:0]!=3'b001) | (~ and_dcpl_202);
  assign mux_tmp_350 = MUX_s_1_2_2(nor_405_nl, or_935_nl, or_933_cse);
  assign nor_404_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_350));
  assign mux_351_nl = MUX_s_1_2_2(nor_404_nl, mux_tmp_350, or_928_cse);
  assign and_dcpl_570 = mux_351_nl & and_dcpl_178;
  assign or_940_cse = (result_rem_11cyc_st_2[2:0]!=3'b001);
  assign nor_403_nl = ~(and_747_cse | and_dcpl_178);
  assign or_942_nl = (result_rem_11cyc_st_3[2:0]!=3'b001) | (~ and_dcpl_176);
  assign mux_tmp_352 = MUX_s_1_2_2(nor_403_nl, or_942_nl, or_940_cse);
  assign and_722_nl = not_tmp_645 & mux_tmp_352;
  assign mux_tmp_353 = MUX_s_1_2_2(and_722_nl, mux_tmp_352, or_933_cse);
  assign nor_402_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_353));
  assign mux_354_nl = MUX_s_1_2_2(nor_402_nl, mux_tmp_353, or_928_cse);
  assign and_dcpl_572 = mux_354_nl & and_dcpl_152;
  assign or_949_cse = (result_rem_11cyc_st_3[2:0]!=3'b001);
  assign nor_401_nl = ~(and_744_cse | and_dcpl_152);
  assign or_951_nl = (result_rem_11cyc_st_4[2:0]!=3'b001) | (~ and_dcpl_150);
  assign mux_tmp_355 = MUX_s_1_2_2(nor_401_nl, or_951_nl, or_949_cse);
  assign and_719_nl = nand_58_cse & mux_tmp_355;
  assign mux_tmp_356 = MUX_s_1_2_2(and_719_nl, mux_tmp_355, or_940_cse);
  assign and_720_nl = not_tmp_645 & mux_tmp_356;
  assign mux_tmp_357 = MUX_s_1_2_2(and_720_nl, mux_tmp_356, or_933_cse);
  assign nor_400_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_357));
  assign mux_358_nl = MUX_s_1_2_2(nor_400_nl, mux_tmp_357, or_928_cse);
  assign and_dcpl_576 = mux_358_nl & and_dcpl_125;
  assign or_960_cse = (result_rem_11cyc_st_4[2:0]!=3'b001);
  assign nor_399_nl = ~(and_740_cse | and_dcpl_125);
  assign or_962_nl = (result_rem_11cyc_st_5!=4'b1001) | (~ and_dcpl_105);
  assign mux_tmp_359 = MUX_s_1_2_2(nor_399_nl, or_962_nl, or_960_cse);
  assign and_715_nl = nand_55_cse & mux_tmp_359;
  assign mux_tmp_360 = MUX_s_1_2_2(and_715_nl, mux_tmp_359, or_949_cse);
  assign and_716_nl = nand_58_cse & mux_tmp_360;
  assign mux_tmp_361 = MUX_s_1_2_2(and_716_nl, mux_tmp_360, or_940_cse);
  assign and_717_nl = not_tmp_645 & mux_tmp_361;
  assign mux_tmp_362 = MUX_s_1_2_2(and_717_nl, mux_tmp_361, or_933_cse);
  assign nor_398_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_362));
  assign mux_363_nl = MUX_s_1_2_2(nor_398_nl, mux_tmp_362, or_928_cse);
  assign and_dcpl_578 = mux_363_nl & and_dcpl_101;
  assign or_973_cse = (result_rem_11cyc_st_5!=4'b1001);
  assign nor_397_nl = ~(and_dcpl_105 | and_dcpl_101);
  assign or_975_nl = (result_rem_11cyc_st_6[2:0]!=3'b001) | (~ and_dcpl_99);
  assign mux_tmp_364 = MUX_s_1_2_2(nor_397_nl, or_975_nl, or_973_cse);
  assign and_710_nl = nand_51_cse & mux_tmp_364;
  assign mux_tmp_365 = MUX_s_1_2_2(and_710_nl, mux_tmp_364, or_960_cse);
  assign and_711_nl = nand_55_cse & mux_tmp_365;
  assign mux_tmp_366 = MUX_s_1_2_2(and_711_nl, mux_tmp_365, or_949_cse);
  assign and_712_nl = nand_58_cse & mux_tmp_366;
  assign mux_tmp_367 = MUX_s_1_2_2(and_712_nl, mux_tmp_366, or_940_cse);
  assign and_713_nl = not_tmp_645 & mux_tmp_367;
  assign mux_tmp_368 = MUX_s_1_2_2(and_713_nl, mux_tmp_367, or_933_cse);
  assign nor_396_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_368));
  assign mux_369_nl = MUX_s_1_2_2(nor_396_nl, mux_tmp_368, or_928_cse);
  assign and_dcpl_580 = mux_369_nl & and_dcpl_75;
  assign or_988_cse = (result_rem_11cyc_st_6[2:0]!=3'b001);
  assign nor_394_nl = ~(and_731_cse | and_dcpl_75);
  assign or_990_nl = (result_rem_11cyc_st_7[2:0]!=3'b001) | (~ and_dcpl_73);
  assign mux_tmp_370 = MUX_s_1_2_2(nor_394_nl, or_990_nl, or_988_cse);
  assign nor_395_nl = ~(and_dcpl_105 | (~ mux_tmp_370));
  assign mux_tmp_371 = MUX_s_1_2_2(nor_395_nl, mux_tmp_370, or_973_cse);
  assign and_706_nl = nand_51_cse & mux_tmp_371;
  assign mux_tmp_372 = MUX_s_1_2_2(and_706_nl, mux_tmp_371, or_960_cse);
  assign and_707_nl = nand_55_cse & mux_tmp_372;
  assign mux_tmp_373 = MUX_s_1_2_2(and_707_nl, mux_tmp_372, or_949_cse);
  assign and_708_nl = nand_58_cse & mux_tmp_373;
  assign mux_tmp_374 = MUX_s_1_2_2(and_708_nl, mux_tmp_373, or_940_cse);
  assign and_709_nl = not_tmp_645 & mux_tmp_374;
  assign mux_tmp_375 = MUX_s_1_2_2(and_709_nl, mux_tmp_374, or_933_cse);
  assign nor_393_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_375));
  assign mux_376_nl = MUX_s_1_2_2(nor_393_nl, mux_tmp_375, or_928_cse);
  assign and_dcpl_583 = mux_376_nl & and_dcpl_47;
  assign nor_390_nl = ~(and_725_cse | and_dcpl_47);
  assign or_1007_nl = (result_rem_11cyc_st_8!=4'b1001) | (~ and_dcpl_28);
  assign or_1005_nl = (result_rem_11cyc_st_7[2:0]!=3'b001);
  assign mux_tmp_377 = MUX_s_1_2_2(nor_390_nl, or_1007_nl, or_1005_nl);
  assign and_700_nl = nand_42_cse & mux_tmp_377;
  assign mux_tmp_378 = MUX_s_1_2_2(and_700_nl, mux_tmp_377, or_988_cse);
  assign nor_391_nl = ~(and_dcpl_105 | (~ mux_tmp_378));
  assign mux_tmp_379 = MUX_s_1_2_2(nor_391_nl, mux_tmp_378, or_973_cse);
  assign and_701_nl = nand_51_cse & mux_tmp_379;
  assign mux_tmp_380 = MUX_s_1_2_2(and_701_nl, mux_tmp_379, or_960_cse);
  assign and_702_nl = nand_55_cse & mux_tmp_380;
  assign mux_tmp_381 = MUX_s_1_2_2(and_702_nl, mux_tmp_380, or_949_cse);
  assign and_703_nl = nand_58_cse & mux_tmp_381;
  assign mux_tmp_382 = MUX_s_1_2_2(and_703_nl, mux_tmp_381, or_940_cse);
  assign and_704_nl = not_tmp_645 & mux_tmp_382;
  assign mux_tmp_383 = MUX_s_1_2_2(and_704_nl, mux_tmp_382, or_933_cse);
  assign nor_392_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_383));
  assign mux_384_nl = MUX_s_1_2_2(nor_392_nl, mux_tmp_383, or_928_cse);
  assign and_dcpl_586 = mux_384_nl & and_dcpl_4 & and_dcpl_18 & (result_rem_11cyc_st_9[0]);
  assign or_tmp_1005 = (~ main_stage_0_10) | (~ asn_itm_9) | (result_rem_11cyc_st_9!=4'b1001);
  assign nor_383_nl = ~((result_rem_11cyc_st_8[3]) | (~ or_tmp_1005));
  assign or_1024_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (result_rem_11cyc_st_8[2:0]!=3'b001);
  assign mux_tmp_385 = MUX_s_1_2_2(nor_383_nl, or_tmp_1005, or_1024_nl);
  assign nor_384_nl = ~((result_rem_11cyc_st_7[3]) | (~ mux_tmp_385));
  assign or_1023_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (result_rem_11cyc_st_7[2:0]!=3'b001);
  assign mux_tmp_386 = MUX_s_1_2_2(nor_384_nl, mux_tmp_385, or_1023_nl);
  assign nor_385_nl = ~((result_rem_11cyc_st_6[3]) | (~ mux_tmp_386));
  assign or_1022_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (result_rem_11cyc_st_6[2:0]!=3'b001);
  assign mux_tmp_387 = MUX_s_1_2_2(nor_385_nl, mux_tmp_386, or_1022_nl);
  assign nor_386_nl = ~((result_rem_11cyc_st_5[3]) | (~ mux_tmp_387));
  assign or_1021_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5[2:0]!=3'b001);
  assign mux_tmp_388 = MUX_s_1_2_2(nor_386_nl, mux_tmp_387, or_1021_nl);
  assign nor_387_nl = ~((result_rem_11cyc_st_4[3]) | (~ mux_tmp_388));
  assign or_1020_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4[2:0]!=3'b001);
  assign mux_tmp_389 = MUX_s_1_2_2(nor_387_nl, mux_tmp_388, or_1020_nl);
  assign nor_388_nl = ~((result_rem_11cyc_st_3[3]) | (~ mux_tmp_389));
  assign or_1019_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3[2:0]!=3'b001);
  assign mux_tmp_390 = MUX_s_1_2_2(nor_388_nl, mux_tmp_389, or_1019_nl);
  assign nor_389_nl = ~((result_rem_11cyc_st_2[3]) | (~ mux_tmp_390));
  assign or_1018_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2[2:0]!=3'b001);
  assign mux_tmp_391 = MUX_s_1_2_2(nor_389_nl, mux_tmp_390, or_1018_nl);
  assign and_697_nl = not_tmp_645 & mux_tmp_391;
  assign mux_tmp_392 = MUX_s_1_2_2(and_697_nl, mux_tmp_391, or_933_cse);
  assign and_698_nl = nand_146_cse & mux_tmp_392;
  assign or_1016_nl = (result_result_acc_tmp[3:1]!=3'b100);
  assign mux_tmp_393 = MUX_s_1_2_2(and_698_nl, mux_tmp_392, or_1016_nl);
  assign and_dcpl_590 = and_dcpl_532 & and_dcpl_352;
  assign or_tmp_1017 = (result_rem_11cyc[2:0]!=3'b010) | not_tmp_645;
  assign or_1037_cse = (result_result_acc_tmp!=4'b1010);
  assign nor_382_nl = ~(ccs_ccore_start_rsci_idat | (~ or_tmp_1017));
  assign mux_394_nl = MUX_s_1_2_2(nor_382_nl, or_tmp_1017, or_1037_cse);
  assign and_dcpl_592 = mux_394_nl & and_dcpl_205;
  assign or_1042_cse = (result_rem_11cyc[2:0]!=3'b010);
  assign nor_381_nl = ~(and_749_cse | and_dcpl_205);
  assign or_1044_nl = (result_rem_11cyc_st_2[2:0]!=3'b010) | (~ and_dcpl_202);
  assign mux_tmp_395 = MUX_s_1_2_2(nor_381_nl, or_1044_nl, or_1042_cse);
  assign nor_380_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_395));
  assign mux_396_nl = MUX_s_1_2_2(nor_380_nl, mux_tmp_395, or_1037_cse);
  assign and_dcpl_594 = mux_396_nl & and_dcpl_179;
  assign or_1049_cse = (result_rem_11cyc_st_2[2:0]!=3'b010);
  assign nor_379_nl = ~(and_747_cse | and_dcpl_179);
  assign or_1051_nl = (result_rem_11cyc_st_3[2:0]!=3'b010) | (~ and_dcpl_176);
  assign mux_tmp_397 = MUX_s_1_2_2(nor_379_nl, or_1051_nl, or_1049_cse);
  assign and_695_nl = not_tmp_645 & mux_tmp_397;
  assign mux_tmp_398 = MUX_s_1_2_2(and_695_nl, mux_tmp_397, or_1042_cse);
  assign nor_378_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_398));
  assign mux_399_nl = MUX_s_1_2_2(nor_378_nl, mux_tmp_398, or_1037_cse);
  assign and_dcpl_596 = mux_399_nl & and_dcpl_153;
  assign or_1058_cse = (result_rem_11cyc_st_3[2:0]!=3'b010);
  assign nor_377_nl = ~(and_744_cse | and_dcpl_153);
  assign or_1060_nl = (result_rem_11cyc_st_4[2:0]!=3'b010) | (~ and_dcpl_150);
  assign mux_tmp_400 = MUX_s_1_2_2(nor_377_nl, or_1060_nl, or_1058_cse);
  assign and_692_nl = nand_58_cse & mux_tmp_400;
  assign mux_tmp_401 = MUX_s_1_2_2(and_692_nl, mux_tmp_400, or_1049_cse);
  assign and_693_nl = not_tmp_645 & mux_tmp_401;
  assign mux_tmp_402 = MUX_s_1_2_2(and_693_nl, mux_tmp_401, or_1042_cse);
  assign nor_376_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_402));
  assign mux_403_nl = MUX_s_1_2_2(nor_376_nl, mux_tmp_402, or_1037_cse);
  assign and_dcpl_599 = mux_403_nl & and_dcpl_127;
  assign or_1069_cse = (result_rem_11cyc_st_4[2:0]!=3'b010);
  assign nor_375_nl = ~(and_740_cse | and_dcpl_127);
  assign or_1071_nl = (result_rem_11cyc_st_5!=4'b1010) | (~ and_dcpl_105);
  assign mux_tmp_404 = MUX_s_1_2_2(nor_375_nl, or_1071_nl, or_1069_cse);
  assign and_688_nl = nand_55_cse & mux_tmp_404;
  assign mux_tmp_405 = MUX_s_1_2_2(and_688_nl, mux_tmp_404, or_1058_cse);
  assign and_689_nl = nand_58_cse & mux_tmp_405;
  assign mux_tmp_406 = MUX_s_1_2_2(and_689_nl, mux_tmp_405, or_1049_cse);
  assign and_690_nl = not_tmp_645 & mux_tmp_406;
  assign mux_tmp_407 = MUX_s_1_2_2(and_690_nl, mux_tmp_406, or_1042_cse);
  assign nor_374_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_407));
  assign mux_408_nl = MUX_s_1_2_2(nor_374_nl, mux_tmp_407, or_1037_cse);
  assign and_dcpl_601 = mux_408_nl & and_dcpl_102;
  assign or_1082_cse = (result_rem_11cyc_st_5!=4'b1010);
  assign nor_373_nl = ~(and_dcpl_105 | and_dcpl_102);
  assign or_1084_nl = (result_rem_11cyc_st_6[2:0]!=3'b010) | (~ and_dcpl_99);
  assign mux_tmp_409 = MUX_s_1_2_2(nor_373_nl, or_1084_nl, or_1082_cse);
  assign and_683_nl = nand_51_cse & mux_tmp_409;
  assign mux_tmp_410 = MUX_s_1_2_2(and_683_nl, mux_tmp_409, or_1069_cse);
  assign and_684_nl = nand_55_cse & mux_tmp_410;
  assign mux_tmp_411 = MUX_s_1_2_2(and_684_nl, mux_tmp_410, or_1058_cse);
  assign and_685_nl = nand_58_cse & mux_tmp_411;
  assign mux_tmp_412 = MUX_s_1_2_2(and_685_nl, mux_tmp_411, or_1049_cse);
  assign and_686_nl = not_tmp_645 & mux_tmp_412;
  assign mux_tmp_413 = MUX_s_1_2_2(and_686_nl, mux_tmp_412, or_1042_cse);
  assign nor_372_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_413));
  assign mux_414_nl = MUX_s_1_2_2(nor_372_nl, mux_tmp_413, or_1037_cse);
  assign and_dcpl_603 = mux_414_nl & and_dcpl_76;
  assign or_1097_cse = (result_rem_11cyc_st_6[2:0]!=3'b010);
  assign nor_370_nl = ~(and_731_cse | and_dcpl_76);
  assign or_1099_nl = (result_rem_11cyc_st_7[2:0]!=3'b010) | (~ and_dcpl_73);
  assign mux_tmp_415 = MUX_s_1_2_2(nor_370_nl, or_1099_nl, or_1097_cse);
  assign nor_371_nl = ~(and_dcpl_105 | (~ mux_tmp_415));
  assign mux_tmp_416 = MUX_s_1_2_2(nor_371_nl, mux_tmp_415, or_1082_cse);
  assign and_679_nl = nand_51_cse & mux_tmp_416;
  assign mux_tmp_417 = MUX_s_1_2_2(and_679_nl, mux_tmp_416, or_1069_cse);
  assign and_680_nl = nand_55_cse & mux_tmp_417;
  assign mux_tmp_418 = MUX_s_1_2_2(and_680_nl, mux_tmp_417, or_1058_cse);
  assign and_681_nl = nand_58_cse & mux_tmp_418;
  assign mux_tmp_419 = MUX_s_1_2_2(and_681_nl, mux_tmp_418, or_1049_cse);
  assign and_682_nl = not_tmp_645 & mux_tmp_419;
  assign mux_tmp_420 = MUX_s_1_2_2(and_682_nl, mux_tmp_419, or_1042_cse);
  assign nor_369_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_420));
  assign mux_421_nl = MUX_s_1_2_2(nor_369_nl, mux_tmp_420, or_1037_cse);
  assign and_dcpl_607 = mux_421_nl & and_dcpl_50;
  assign nor_366_nl = ~(and_725_cse | and_dcpl_50);
  assign or_1116_nl = (result_rem_11cyc_st_8!=4'b1010) | (~ and_dcpl_28);
  assign or_1114_nl = (result_rem_11cyc_st_7[2:0]!=3'b010);
  assign mux_tmp_422 = MUX_s_1_2_2(nor_366_nl, or_1116_nl, or_1114_nl);
  assign and_673_nl = nand_42_cse & mux_tmp_422;
  assign mux_tmp_423 = MUX_s_1_2_2(and_673_nl, mux_tmp_422, or_1097_cse);
  assign nor_367_nl = ~(and_dcpl_105 | (~ mux_tmp_423));
  assign mux_tmp_424 = MUX_s_1_2_2(nor_367_nl, mux_tmp_423, or_1082_cse);
  assign and_674_nl = nand_51_cse & mux_tmp_424;
  assign mux_tmp_425 = MUX_s_1_2_2(and_674_nl, mux_tmp_424, or_1069_cse);
  assign and_675_nl = nand_55_cse & mux_tmp_425;
  assign mux_tmp_426 = MUX_s_1_2_2(and_675_nl, mux_tmp_425, or_1058_cse);
  assign and_676_nl = nand_58_cse & mux_tmp_426;
  assign mux_tmp_427 = MUX_s_1_2_2(and_676_nl, mux_tmp_426, or_1049_cse);
  assign and_677_nl = not_tmp_645 & mux_tmp_427;
  assign mux_tmp_428 = MUX_s_1_2_2(and_677_nl, mux_tmp_427, or_1042_cse);
  assign nor_368_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_428));
  assign mux_429_nl = MUX_s_1_2_2(nor_368_nl, mux_tmp_428, or_1037_cse);
  assign and_dcpl_611 = mux_429_nl & and_dcpl_4 & (result_rem_11cyc_st_9[3]) & (result_rem_11cyc_st_9[1])
      & (~ (result_rem_11cyc_st_9[0]));
  assign or_tmp_1113 = (~ main_stage_0_10) | (~ asn_itm_9) | (result_rem_11cyc_st_9!=4'b1010);
  assign nor_358_nl = ~((result_rem_11cyc_st_8[3]) | (~ or_tmp_1113));
  assign or_1133_nl = (~ main_stage_0_9) | (~ asn_itm_8) | (result_rem_11cyc_st_8[2:0]!=3'b010);
  assign mux_tmp_430 = MUX_s_1_2_2(nor_358_nl, or_tmp_1113, or_1133_nl);
  assign nor_359_nl = ~((result_rem_11cyc_st_7[3]) | (~ mux_tmp_430));
  assign or_1132_nl = (~ main_stage_0_8) | (~ asn_itm_7) | (result_rem_11cyc_st_7[2:0]!=3'b010);
  assign mux_tmp_431 = MUX_s_1_2_2(nor_359_nl, mux_tmp_430, or_1132_nl);
  assign nor_360_nl = ~((result_rem_11cyc_st_6[3]) | (~ mux_tmp_431));
  assign or_1131_nl = (~ main_stage_0_7) | (~ asn_itm_6) | (result_rem_11cyc_st_6[2:0]!=3'b010);
  assign mux_tmp_432 = MUX_s_1_2_2(nor_360_nl, mux_tmp_431, or_1131_nl);
  assign nor_361_nl = ~((result_rem_11cyc_st_5[3]) | (~ mux_tmp_432));
  assign or_1130_nl = (~ main_stage_0_6) | (~ asn_itm_5) | (result_rem_11cyc_st_5[2:0]!=3'b010);
  assign mux_tmp_433 = MUX_s_1_2_2(nor_361_nl, mux_tmp_432, or_1130_nl);
  assign nor_362_nl = ~((result_rem_11cyc_st_4[3]) | (~ mux_tmp_433));
  assign or_1129_nl = (~ main_stage_0_5) | (~ asn_itm_4) | (result_rem_11cyc_st_4[2:0]!=3'b010);
  assign mux_tmp_434 = MUX_s_1_2_2(nor_362_nl, mux_tmp_433, or_1129_nl);
  assign nor_363_nl = ~((result_rem_11cyc_st_3[3]) | (~ mux_tmp_434));
  assign or_1128_nl = (~ main_stage_0_4) | (~ asn_itm_3) | (result_rem_11cyc_st_3[2:0]!=3'b010);
  assign mux_tmp_435 = MUX_s_1_2_2(nor_363_nl, mux_tmp_434, or_1128_nl);
  assign nor_364_nl = ~((result_rem_11cyc_st_2[3]) | (~ mux_tmp_435));
  assign or_1127_nl = (~ main_stage_0_3) | (~ asn_itm_2) | (result_rem_11cyc_st_2[2:0]!=3'b010);
  assign mux_tmp_436 = MUX_s_1_2_2(nor_364_nl, mux_tmp_435, or_1127_nl);
  assign and_671_nl = not_tmp_645 & mux_tmp_436;
  assign mux_tmp_437 = MUX_s_1_2_2(and_671_nl, mux_tmp_436, or_1042_cse);
  assign nor_365_nl = ~(ccs_ccore_start_rsci_idat | (~ mux_tmp_437));
  assign mux_tmp_438 = MUX_s_1_2_2(nor_365_nl, mux_tmp_437, or_1037_cse);
  assign return_rsci_d_mx0c0 = and_dcpl_235 & and_dcpl_233;
  assign return_rsci_d_mx0c1 = and_dcpl_235 & and_dcpl_237;
  assign return_rsci_d_mx0c2 = and_dcpl_235 & and_dcpl_240;
  assign return_rsci_d_mx0c3 = and_dcpl_235 & and_dcpl_239 & (result_rem_11cyc_st_11[0]);
  assign return_rsci_d_mx0c4 = and_dcpl_235 & and_dcpl_244 & (~ (result_rem_11cyc_st_11[0]));
  assign return_rsci_d_mx0c5 = and_dcpl_235 & and_dcpl_244 & (result_rem_11cyc_st_11[0]);
  assign return_rsci_d_mx0c6 = and_dcpl_235 & and_dcpl_249 & (~ (result_rem_11cyc_st_11[0]));
  assign return_rsci_d_mx0c7 = and_dcpl_235 & and_dcpl_249 & (result_rem_11cyc_st_11[0]);
  assign return_rsci_d_mx0c8 = and_dcpl_254 & and_dcpl_233;
  assign return_rsci_d_mx0c9 = and_dcpl_254 & and_dcpl_237;
  assign return_rsci_d_mx0c10 = and_dcpl_254 & and_dcpl_240;
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_en & (return_rsci_d_mx0c0 | return_rsci_d_mx0c1 | return_rsci_d_mx0c2
        | return_rsci_d_mx0c3 | return_rsci_d_mx0c4 | return_rsci_d_mx0c5 | return_rsci_d_mx0c6
        | return_rsci_d_mx0c7 | return_rsci_d_mx0c8 | return_rsci_d_mx0c9 | return_rsci_d_mx0c10)
        ) begin
      return_rsci_d <= MUX1HOT_v_64_11_2(result_rem_12_cmp_1_z, result_rem_12_cmp_2_z,
          result_rem_12_cmp_3_z, result_rem_12_cmp_4_z, result_rem_12_cmp_5_z, result_rem_12_cmp_6_z,
          result_rem_12_cmp_7_z, result_rem_12_cmp_8_z, result_rem_12_cmp_9_z, result_rem_12_cmp_10_z,
          result_rem_12_cmp_z, {return_rsci_d_mx0c0 , return_rsci_d_mx0c1 , return_rsci_d_mx0c2
          , return_rsci_d_mx0c3 , return_rsci_d_mx0c4 , return_rsci_d_mx0c5 , return_rsci_d_mx0c6
          , return_rsci_d_mx0c7 , return_rsci_d_mx0c8 , return_rsci_d_mx0c9 , return_rsci_d_mx0c10});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_11 <= 4'b0000;
    end
    else if ( ccs_ccore_en & main_stage_0_11 & asn_itm_10 ) begin
      result_rem_11cyc_st_11 <= result_rem_11cyc_st_10;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      asn_itm_11 <= 1'b0;
      asn_itm_10 <= 1'b0;
      asn_itm_9 <= 1'b0;
      asn_itm_8 <= 1'b0;
      asn_itm_7 <= 1'b0;
      asn_itm_6 <= 1'b0;
      asn_itm_5 <= 1'b0;
      asn_itm_4 <= 1'b0;
      asn_itm_3 <= 1'b0;
      asn_itm_2 <= 1'b0;
      asn_itm_1 <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      main_stage_0_6 <= 1'b0;
      main_stage_0_7 <= 1'b0;
      main_stage_0_8 <= 1'b0;
      main_stage_0_9 <= 1'b0;
      main_stage_0_10 <= 1'b0;
      main_stage_0_11 <= 1'b0;
      main_stage_0_12 <= 1'b0;
    end
    else if ( ccs_ccore_en ) begin
      asn_itm_11 <= asn_itm_10;
      asn_itm_10 <= asn_itm_9;
      asn_itm_9 <= asn_itm_8;
      asn_itm_8 <= asn_itm_7;
      asn_itm_7 <= asn_itm_6;
      asn_itm_6 <= asn_itm_5;
      asn_itm_5 <= asn_itm_4;
      asn_itm_4 <= asn_itm_3;
      asn_itm_3 <= asn_itm_2;
      asn_itm_2 <= asn_itm_1;
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      main_stage_0_6 <= main_stage_0_5;
      main_stage_0_7 <= main_stage_0_6;
      main_stage_0_8 <= main_stage_0_7;
      main_stage_0_9 <= main_stage_0_8;
      main_stage_0_10 <= main_stage_0_9;
      main_stage_0_11 <= main_stage_0_10;
      main_stage_0_12 <= main_stage_0_11;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_1_cse ) begin
      result_rem_12_cmp_1_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_1_2,
          m_buf_sva_mut_1_3, m_buf_sva_mut_1_4, m_buf_sva_mut_1_5, m_buf_sva_mut_1_6,
          m_buf_sva_mut_1_7, m_buf_sva_mut_1_8, m_buf_sva_mut_1_9, m_buf_sva_mut_1_10,
          {and_dcpl_263 , and_dcpl_269 , and_dcpl_275 , and_dcpl_281 , and_dcpl_287
          , and_dcpl_293 , and_dcpl_299 , and_dcpl_305 , and_dcpl_311 , mux_tmp_37});
      result_rem_12_cmp_1_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_1_2,
          base_buf_sva_mut_1_3, base_buf_sva_mut_1_4, base_buf_sva_mut_1_5, base_buf_sva_mut_1_6,
          base_buf_sva_mut_1_7, base_buf_sva_mut_1_8, base_buf_sva_mut_1_9, base_buf_sva_mut_1_10,
          {and_dcpl_263 , and_dcpl_269 , and_dcpl_275 , and_dcpl_281 , and_dcpl_287
          , and_dcpl_293 , and_dcpl_299 , and_dcpl_305 , and_dcpl_311 , mux_tmp_37});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_3_cse ) begin
      result_rem_12_cmp_2_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2_2,
          m_buf_sva_mut_2_3, m_buf_sva_mut_2_4, m_buf_sva_mut_2_5, m_buf_sva_mut_2_6,
          m_buf_sva_mut_2_7, m_buf_sva_mut_2_8, m_buf_sva_mut_2_9, m_buf_sva_mut_2_10,
          {and_dcpl_319 , and_dcpl_322 , and_dcpl_325 , and_dcpl_329 , and_dcpl_333
          , and_dcpl_337 , and_dcpl_341 , and_dcpl_344 , and_dcpl_347 , mux_tmp_75});
      result_rem_12_cmp_2_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2_2,
          base_buf_sva_mut_2_3, base_buf_sva_mut_2_4, base_buf_sva_mut_2_5, base_buf_sva_mut_2_6,
          base_buf_sva_mut_2_7, base_buf_sva_mut_2_8, base_buf_sva_mut_2_9, base_buf_sva_mut_2_10,
          {and_dcpl_319 , and_dcpl_322 , and_dcpl_325 , and_dcpl_329 , and_dcpl_333
          , and_dcpl_337 , and_dcpl_341 , and_dcpl_344 , and_dcpl_347 , mux_tmp_75});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_5_cse ) begin
      result_rem_12_cmp_3_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_3_2,
          m_buf_sva_mut_3_3, m_buf_sva_mut_3_4, m_buf_sva_mut_3_5, m_buf_sva_mut_3_6,
          m_buf_sva_mut_3_7, m_buf_sva_mut_3_8, m_buf_sva_mut_3_9, m_buf_sva_mut_3_10,
          {and_dcpl_353 , and_dcpl_357 , and_dcpl_361 , and_dcpl_364 , and_dcpl_367
          , and_dcpl_370 , and_dcpl_373 , and_dcpl_377 , and_dcpl_381 , mux_tmp_113});
      result_rem_12_cmp_3_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_3_2,
          base_buf_sva_mut_3_3, base_buf_sva_mut_3_4, base_buf_sva_mut_3_5, base_buf_sva_mut_3_6,
          base_buf_sva_mut_3_7, base_buf_sva_mut_3_8, base_buf_sva_mut_3_9, base_buf_sva_mut_3_10,
          {and_dcpl_353 , and_dcpl_357 , and_dcpl_361 , and_dcpl_364 , and_dcpl_367
          , and_dcpl_370 , and_dcpl_373 , and_dcpl_377 , and_dcpl_381 , mux_tmp_113});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_7_cse ) begin
      result_rem_12_cmp_4_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_4_2,
          m_buf_sva_mut_4_3, m_buf_sva_mut_4_4, m_buf_sva_mut_4_5, m_buf_sva_mut_4_6,
          m_buf_sva_mut_4_7, m_buf_sva_mut_4_8, m_buf_sva_mut_4_9, m_buf_sva_mut_4_10,
          {and_dcpl_387 , and_dcpl_390 , and_dcpl_393 , and_dcpl_396 , and_dcpl_399
          , and_dcpl_402 , and_dcpl_405 , and_dcpl_408 , and_dcpl_411 , mux_tmp_151});
      result_rem_12_cmp_4_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_4_2,
          base_buf_sva_mut_4_3, base_buf_sva_mut_4_4, base_buf_sva_mut_4_5, base_buf_sva_mut_4_6,
          base_buf_sva_mut_4_7, base_buf_sva_mut_4_8, base_buf_sva_mut_4_9, base_buf_sva_mut_4_10,
          {and_dcpl_387 , and_dcpl_390 , and_dcpl_393 , and_dcpl_396 , and_dcpl_399
          , and_dcpl_402 , and_dcpl_405 , and_dcpl_408 , and_dcpl_411 , mux_tmp_151});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_9_cse ) begin
      result_rem_12_cmp_5_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_5_2,
          m_buf_sva_mut_5_3, m_buf_sva_mut_5_4, m_buf_sva_mut_5_5, m_buf_sva_mut_5_6,
          m_buf_sva_mut_5_7, m_buf_sva_mut_5_8, m_buf_sva_mut_5_9, m_buf_sva_mut_5_10,
          {and_dcpl_418 , and_dcpl_422 , and_dcpl_426 , and_dcpl_430 , and_dcpl_433
          , and_dcpl_437 , and_dcpl_441 , and_dcpl_444 , and_dcpl_447 , mux_tmp_189});
      result_rem_12_cmp_5_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_5_2,
          base_buf_sva_mut_5_3, base_buf_sva_mut_5_4, base_buf_sva_mut_5_5, base_buf_sva_mut_5_6,
          base_buf_sva_mut_5_7, base_buf_sva_mut_5_8, base_buf_sva_mut_5_9, base_buf_sva_mut_5_10,
          {and_dcpl_418 , and_dcpl_422 , and_dcpl_426 , and_dcpl_430 , and_dcpl_433
          , and_dcpl_437 , and_dcpl_441 , and_dcpl_444 , and_dcpl_447 , mux_tmp_189});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_11_cse ) begin
      result_rem_12_cmp_6_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_6_2,
          m_buf_sva_mut_6_3, m_buf_sva_mut_6_4, m_buf_sva_mut_6_5, m_buf_sva_mut_6_6,
          m_buf_sva_mut_6_7, m_buf_sva_mut_6_8, m_buf_sva_mut_6_9, m_buf_sva_mut_6_10,
          {and_dcpl_452 , and_dcpl_455 , and_dcpl_458 , and_dcpl_462 , and_dcpl_464
          , and_dcpl_468 , and_dcpl_472 , and_dcpl_474 , and_dcpl_476 , mux_tmp_227});
      result_rem_12_cmp_6_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_6_2,
          base_buf_sva_mut_6_3, base_buf_sva_mut_6_4, base_buf_sva_mut_6_5, base_buf_sva_mut_6_6,
          base_buf_sva_mut_6_7, base_buf_sva_mut_6_8, base_buf_sva_mut_6_9, base_buf_sva_mut_6_10,
          {and_dcpl_452 , and_dcpl_455 , and_dcpl_458 , and_dcpl_462 , and_dcpl_464
          , and_dcpl_468 , and_dcpl_472 , and_dcpl_474 , and_dcpl_476 , mux_tmp_227});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_13_cse ) begin
      result_rem_12_cmp_7_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_7_2,
          m_buf_sva_mut_7_3, m_buf_sva_mut_7_4, m_buf_sva_mut_7_5, m_buf_sva_mut_7_6,
          m_buf_sva_mut_7_7, m_buf_sva_mut_7_8, m_buf_sva_mut_7_9, m_buf_sva_mut_7_10,
          {and_dcpl_480 , and_dcpl_484 , and_dcpl_488 , and_dcpl_491 , and_dcpl_493
          , and_dcpl_496 , and_dcpl_499 , and_dcpl_501 , and_dcpl_503 , mux_tmp_265});
      result_rem_12_cmp_7_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_7_2,
          base_buf_sva_mut_7_3, base_buf_sva_mut_7_4, base_buf_sva_mut_7_5, base_buf_sva_mut_7_6,
          base_buf_sva_mut_7_7, base_buf_sva_mut_7_8, base_buf_sva_mut_7_9, base_buf_sva_mut_7_10,
          {and_dcpl_480 , and_dcpl_484 , and_dcpl_488 , and_dcpl_491 , and_dcpl_493
          , and_dcpl_496 , and_dcpl_499 , and_dcpl_501 , and_dcpl_503 , mux_tmp_265});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_15_cse ) begin
      result_rem_12_cmp_8_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_8_2,
          m_buf_sva_mut_8_3, m_buf_sva_mut_8_4, m_buf_sva_mut_8_5, m_buf_sva_mut_8_6,
          m_buf_sva_mut_8_7, m_buf_sva_mut_8_8, m_buf_sva_mut_8_9, m_buf_sva_mut_8_10,
          {and_dcpl_507 , and_dcpl_510 , and_dcpl_513 , and_dcpl_516 , and_dcpl_518
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_526 , and_dcpl_528 , mux_tmp_303});
      result_rem_12_cmp_8_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_8_2,
          base_buf_sva_mut_8_3, base_buf_sva_mut_8_4, base_buf_sva_mut_8_5, base_buf_sva_mut_8_6,
          base_buf_sva_mut_8_7, base_buf_sva_mut_8_8, base_buf_sva_mut_8_9, base_buf_sva_mut_8_10,
          {and_dcpl_507 , and_dcpl_510 , and_dcpl_513 , and_dcpl_516 , and_dcpl_518
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_526 , and_dcpl_528 , mux_tmp_303});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_17_cse ) begin
      result_rem_12_cmp_9_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_9_2,
          m_buf_sva_mut_9_3, m_buf_sva_mut_9_4, m_buf_sva_mut_9_5, m_buf_sva_mut_9_6,
          m_buf_sva_mut_9_7, m_buf_sva_mut_9_8, m_buf_sva_mut_9_9, m_buf_sva_mut_9_10,
          {and_dcpl_533 , and_dcpl_536 , and_dcpl_539 , and_dcpl_542 , and_dcpl_546
          , and_dcpl_549 , and_dcpl_552 , and_dcpl_556 , and_dcpl_560 , mux_tmp_348});
      result_rem_12_cmp_9_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_9_2,
          base_buf_sva_mut_9_3, base_buf_sva_mut_9_4, base_buf_sva_mut_9_5, base_buf_sva_mut_9_6,
          base_buf_sva_mut_9_7, base_buf_sva_mut_9_8, base_buf_sva_mut_9_9, base_buf_sva_mut_9_10,
          {and_dcpl_533 , and_dcpl_536 , and_dcpl_539 , and_dcpl_542 , and_dcpl_546
          , and_dcpl_549 , and_dcpl_552 , and_dcpl_556 , and_dcpl_560 , mux_tmp_348});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_19_cse ) begin
      result_rem_12_cmp_10_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_10_2,
          m_buf_sva_mut_10_3, m_buf_sva_mut_10_4, m_buf_sva_mut_10_5, m_buf_sva_mut_10_6,
          m_buf_sva_mut_10_7, m_buf_sva_mut_10_8, m_buf_sva_mut_10_9, m_buf_sva_mut_10_10,
          {and_dcpl_566 , and_dcpl_568 , and_dcpl_570 , and_dcpl_572 , and_dcpl_576
          , and_dcpl_578 , and_dcpl_580 , and_dcpl_583 , and_dcpl_586 , mux_tmp_393});
      result_rem_12_cmp_10_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_10_2,
          base_buf_sva_mut_10_3, base_buf_sva_mut_10_4, base_buf_sva_mut_10_5, base_buf_sva_mut_10_6,
          base_buf_sva_mut_10_7, base_buf_sva_mut_10_8, base_buf_sva_mut_10_9, base_buf_sva_mut_10_10,
          {and_dcpl_566 , and_dcpl_568 , and_dcpl_570 , and_dcpl_572 , and_dcpl_576
          , and_dcpl_578 , and_dcpl_580 , and_dcpl_583 , and_dcpl_586 , mux_tmp_393});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( result_and_21_cse ) begin
      result_rem_12_cmp_b <= MUX1HOT_v_64_10_2(m_rsci_idat, m_buf_sva_mut_2, m_buf_sva_mut_3,
          m_buf_sva_mut_4, m_buf_sva_mut_5, m_buf_sva_mut_6, m_buf_sva_mut_7, m_buf_sva_mut_8,
          m_buf_sva_mut_9, m_buf_sva_mut_10, {and_dcpl_590 , and_dcpl_592 , and_dcpl_594
          , and_dcpl_596 , and_dcpl_599 , and_dcpl_601 , and_dcpl_603 , and_dcpl_607
          , and_dcpl_611 , mux_tmp_438});
      result_rem_12_cmp_a <= MUX1HOT_v_64_10_2(base_rsci_idat, base_buf_sva_mut_2,
          base_buf_sva_mut_3, base_buf_sva_mut_4, base_buf_sva_mut_5, base_buf_sva_mut_6,
          base_buf_sva_mut_7, base_buf_sva_mut_8, base_buf_sva_mut_9, base_buf_sva_mut_10,
          {and_dcpl_590 , and_dcpl_592 , and_dcpl_594 , and_dcpl_596 , and_dcpl_599
          , and_dcpl_601 , and_dcpl_603 , and_dcpl_607 , and_dcpl_611 , mux_tmp_438});
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_cse ) begin
      m_buf_sva_mut_1_10 <= m_buf_sva_mut_1_9;
      base_buf_sva_mut_1_10 <= base_buf_sva_mut_1_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_1_cse ) begin
      m_buf_sva_mut_2_10 <= m_buf_sva_mut_2_9;
      base_buf_sva_mut_2_10 <= base_buf_sva_mut_2_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_2_cse ) begin
      m_buf_sva_mut_3_10 <= m_buf_sva_mut_3_9;
      base_buf_sva_mut_3_10 <= base_buf_sva_mut_3_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_3_cse ) begin
      m_buf_sva_mut_4_10 <= m_buf_sva_mut_4_9;
      base_buf_sva_mut_4_10 <= base_buf_sva_mut_4_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_4_cse ) begin
      m_buf_sva_mut_5_10 <= m_buf_sva_mut_5_9;
      base_buf_sva_mut_5_10 <= base_buf_sva_mut_5_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_5_cse ) begin
      m_buf_sva_mut_6_10 <= m_buf_sva_mut_6_9;
      base_buf_sva_mut_6_10 <= base_buf_sva_mut_6_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_6_cse ) begin
      m_buf_sva_mut_7_10 <= m_buf_sva_mut_7_9;
      base_buf_sva_mut_7_10 <= base_buf_sva_mut_7_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_7_cse ) begin
      m_buf_sva_mut_8_10 <= m_buf_sva_mut_8_9;
      base_buf_sva_mut_8_10 <= base_buf_sva_mut_8_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_8_cse ) begin
      m_buf_sva_mut_9_10 <= m_buf_sva_mut_9_9;
      base_buf_sva_mut_9_10 <= base_buf_sva_mut_9_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_9_cse ) begin
      m_buf_sva_mut_10_10 <= m_buf_sva_mut_10_9;
      base_buf_sva_mut_10_10 <= base_buf_sva_mut_10_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_10_cse ) begin
      m_buf_sva_mut_10 <= m_buf_sva_mut_9;
      base_buf_sva_mut_10 <= base_buf_sva_mut_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_10 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_3 ) begin
      result_rem_11cyc_st_10 <= result_rem_11cyc_st_9;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_11_cse ) begin
      m_buf_sva_mut_1_9 <= m_buf_sva_mut_1_8;
      base_buf_sva_mut_1_9 <= base_buf_sva_mut_1_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_12_cse ) begin
      m_buf_sva_mut_2_9 <= m_buf_sva_mut_2_8;
      base_buf_sva_mut_2_9 <= base_buf_sva_mut_2_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_13_cse ) begin
      m_buf_sva_mut_3_9 <= m_buf_sva_mut_3_8;
      base_buf_sva_mut_3_9 <= base_buf_sva_mut_3_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_14_cse ) begin
      m_buf_sva_mut_4_9 <= m_buf_sva_mut_4_8;
      base_buf_sva_mut_4_9 <= base_buf_sva_mut_4_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_15_cse ) begin
      m_buf_sva_mut_5_9 <= m_buf_sva_mut_5_8;
      base_buf_sva_mut_5_9 <= base_buf_sva_mut_5_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_16_cse ) begin
      m_buf_sva_mut_6_9 <= m_buf_sva_mut_6_8;
      base_buf_sva_mut_6_9 <= base_buf_sva_mut_6_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_17_cse ) begin
      m_buf_sva_mut_7_9 <= m_buf_sva_mut_7_8;
      base_buf_sva_mut_7_9 <= base_buf_sva_mut_7_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_18_cse ) begin
      m_buf_sva_mut_8_9 <= m_buf_sva_mut_8_8;
      base_buf_sva_mut_8_9 <= base_buf_sva_mut_8_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_19_cse ) begin
      m_buf_sva_mut_9_9 <= m_buf_sva_mut_9_8;
      base_buf_sva_mut_9_9 <= base_buf_sva_mut_9_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_20_cse ) begin
      m_buf_sva_mut_10_9 <= m_buf_sva_mut_10_8;
      base_buf_sva_mut_10_9 <= base_buf_sva_mut_10_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_21_cse ) begin
      m_buf_sva_mut_9 <= m_buf_sva_mut_8;
      base_buf_sva_mut_9 <= base_buf_sva_mut_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_9 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_28 ) begin
      result_rem_11cyc_st_9 <= result_rem_11cyc_st_8;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_22_cse ) begin
      m_buf_sva_mut_1_8 <= m_buf_sva_mut_1_7;
      base_buf_sva_mut_1_8 <= base_buf_sva_mut_1_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_23_cse ) begin
      m_buf_sva_mut_2_8 <= m_buf_sva_mut_2_7;
      base_buf_sva_mut_2_8 <= base_buf_sva_mut_2_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_24_cse ) begin
      m_buf_sva_mut_3_8 <= m_buf_sva_mut_3_7;
      base_buf_sva_mut_3_8 <= base_buf_sva_mut_3_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_25_cse ) begin
      m_buf_sva_mut_4_8 <= m_buf_sva_mut_4_7;
      base_buf_sva_mut_4_8 <= base_buf_sva_mut_4_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_26_cse ) begin
      m_buf_sva_mut_5_8 <= m_buf_sva_mut_5_7;
      base_buf_sva_mut_5_8 <= base_buf_sva_mut_5_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_27_cse ) begin
      m_buf_sva_mut_6_8 <= m_buf_sva_mut_6_7;
      base_buf_sva_mut_6_8 <= base_buf_sva_mut_6_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_28_cse ) begin
      m_buf_sva_mut_7_8 <= m_buf_sva_mut_7_7;
      base_buf_sva_mut_7_8 <= base_buf_sva_mut_7_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_29_cse ) begin
      m_buf_sva_mut_8_8 <= m_buf_sva_mut_8_7;
      base_buf_sva_mut_8_8 <= base_buf_sva_mut_8_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_30_cse ) begin
      m_buf_sva_mut_9_8 <= m_buf_sva_mut_9_7;
      base_buf_sva_mut_9_8 <= base_buf_sva_mut_9_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_31_cse ) begin
      m_buf_sva_mut_10_8 <= m_buf_sva_mut_10_7;
      base_buf_sva_mut_10_8 <= base_buf_sva_mut_10_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_32_cse ) begin
      m_buf_sva_mut_8 <= m_buf_sva_mut_7;
      base_buf_sva_mut_8 <= base_buf_sva_mut_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_8 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_53 ) begin
      result_rem_11cyc_st_8 <= result_rem_11cyc_st_7;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_33_cse ) begin
      m_buf_sva_mut_1_7 <= m_buf_sva_mut_1_6;
      base_buf_sva_mut_1_7 <= base_buf_sva_mut_1_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_34_cse ) begin
      m_buf_sva_mut_2_7 <= m_buf_sva_mut_2_6;
      base_buf_sva_mut_2_7 <= base_buf_sva_mut_2_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_35_cse ) begin
      m_buf_sva_mut_3_7 <= m_buf_sva_mut_3_6;
      base_buf_sva_mut_3_7 <= base_buf_sva_mut_3_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_36_cse ) begin
      m_buf_sva_mut_4_7 <= m_buf_sva_mut_4_6;
      base_buf_sva_mut_4_7 <= base_buf_sva_mut_4_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_37_cse ) begin
      m_buf_sva_mut_5_7 <= m_buf_sva_mut_5_6;
      base_buf_sva_mut_5_7 <= base_buf_sva_mut_5_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_38_cse ) begin
      m_buf_sva_mut_6_7 <= m_buf_sva_mut_6_6;
      base_buf_sva_mut_6_7 <= base_buf_sva_mut_6_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_39_cse ) begin
      m_buf_sva_mut_7_7 <= m_buf_sva_mut_7_6;
      base_buf_sva_mut_7_7 <= base_buf_sva_mut_7_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_40_cse ) begin
      m_buf_sva_mut_8_7 <= m_buf_sva_mut_8_6;
      base_buf_sva_mut_8_7 <= base_buf_sva_mut_8_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_41_cse ) begin
      m_buf_sva_mut_9_7 <= m_buf_sva_mut_9_6;
      base_buf_sva_mut_9_7 <= base_buf_sva_mut_9_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_42_cse ) begin
      m_buf_sva_mut_10_7 <= m_buf_sva_mut_10_6;
      base_buf_sva_mut_10_7 <= base_buf_sva_mut_10_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_43_cse ) begin
      m_buf_sva_mut_7 <= m_buf_sva_mut_6;
      base_buf_sva_mut_7 <= base_buf_sva_mut_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_7 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_79 ) begin
      result_rem_11cyc_st_7 <= result_rem_11cyc_st_6;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_44_cse ) begin
      m_buf_sva_mut_1_6 <= m_buf_sva_mut_1_5;
      base_buf_sva_mut_1_6 <= base_buf_sva_mut_1_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_45_cse ) begin
      m_buf_sva_mut_2_6 <= m_buf_sva_mut_2_5;
      base_buf_sva_mut_2_6 <= base_buf_sva_mut_2_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_46_cse ) begin
      m_buf_sva_mut_3_6 <= m_buf_sva_mut_3_5;
      base_buf_sva_mut_3_6 <= base_buf_sva_mut_3_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_47_cse ) begin
      m_buf_sva_mut_4_6 <= m_buf_sva_mut_4_5;
      base_buf_sva_mut_4_6 <= base_buf_sva_mut_4_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_48_cse ) begin
      m_buf_sva_mut_5_6 <= m_buf_sva_mut_5_5;
      base_buf_sva_mut_5_6 <= base_buf_sva_mut_5_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_49_cse ) begin
      m_buf_sva_mut_6_6 <= m_buf_sva_mut_6_5;
      base_buf_sva_mut_6_6 <= base_buf_sva_mut_6_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_50_cse ) begin
      m_buf_sva_mut_7_6 <= m_buf_sva_mut_7_5;
      base_buf_sva_mut_7_6 <= base_buf_sva_mut_7_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_51_cse ) begin
      m_buf_sva_mut_8_6 <= m_buf_sva_mut_8_5;
      base_buf_sva_mut_8_6 <= base_buf_sva_mut_8_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_52_cse ) begin
      m_buf_sva_mut_9_6 <= m_buf_sva_mut_9_5;
      base_buf_sva_mut_9_6 <= base_buf_sva_mut_9_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_53_cse ) begin
      m_buf_sva_mut_10_6 <= m_buf_sva_mut_10_5;
      base_buf_sva_mut_10_6 <= base_buf_sva_mut_10_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_54_cse ) begin
      m_buf_sva_mut_6 <= m_buf_sva_mut_5;
      base_buf_sva_mut_6 <= base_buf_sva_mut_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_6 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_105 ) begin
      result_rem_11cyc_st_6 <= result_rem_11cyc_st_5;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_55_cse ) begin
      m_buf_sva_mut_1_5 <= m_buf_sva_mut_1_4;
      base_buf_sva_mut_1_5 <= base_buf_sva_mut_1_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_56_cse ) begin
      m_buf_sva_mut_2_5 <= m_buf_sva_mut_2_4;
      base_buf_sva_mut_2_5 <= base_buf_sva_mut_2_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_57_cse ) begin
      m_buf_sva_mut_3_5 <= m_buf_sva_mut_3_4;
      base_buf_sva_mut_3_5 <= base_buf_sva_mut_3_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_58_cse ) begin
      m_buf_sva_mut_4_5 <= m_buf_sva_mut_4_4;
      base_buf_sva_mut_4_5 <= base_buf_sva_mut_4_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_59_cse ) begin
      m_buf_sva_mut_5_5 <= m_buf_sva_mut_5_4;
      base_buf_sva_mut_5_5 <= base_buf_sva_mut_5_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_60_cse ) begin
      m_buf_sva_mut_6_5 <= m_buf_sva_mut_6_4;
      base_buf_sva_mut_6_5 <= base_buf_sva_mut_6_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_61_cse ) begin
      m_buf_sva_mut_7_5 <= m_buf_sva_mut_7_4;
      base_buf_sva_mut_7_5 <= base_buf_sva_mut_7_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_62_cse ) begin
      m_buf_sva_mut_8_5 <= m_buf_sva_mut_8_4;
      base_buf_sva_mut_8_5 <= base_buf_sva_mut_8_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_63_cse ) begin
      m_buf_sva_mut_9_5 <= m_buf_sva_mut_9_4;
      base_buf_sva_mut_9_5 <= base_buf_sva_mut_9_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_64_cse ) begin
      m_buf_sva_mut_10_5 <= m_buf_sva_mut_10_4;
      base_buf_sva_mut_10_5 <= base_buf_sva_mut_10_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_65_cse ) begin
      m_buf_sva_mut_5 <= m_buf_sva_mut_4;
      base_buf_sva_mut_5 <= base_buf_sva_mut_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_5 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_130 ) begin
      result_rem_11cyc_st_5 <= result_rem_11cyc_st_4;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_66_cse ) begin
      m_buf_sva_mut_1_4 <= m_buf_sva_mut_1_3;
      base_buf_sva_mut_1_4 <= base_buf_sva_mut_1_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_67_cse ) begin
      m_buf_sva_mut_2_4 <= m_buf_sva_mut_2_3;
      base_buf_sva_mut_2_4 <= base_buf_sva_mut_2_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_68_cse ) begin
      m_buf_sva_mut_3_4 <= m_buf_sva_mut_3_3;
      base_buf_sva_mut_3_4 <= base_buf_sva_mut_3_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_69_cse ) begin
      m_buf_sva_mut_4_4 <= m_buf_sva_mut_4_3;
      base_buf_sva_mut_4_4 <= base_buf_sva_mut_4_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_70_cse ) begin
      m_buf_sva_mut_5_4 <= m_buf_sva_mut_5_3;
      base_buf_sva_mut_5_4 <= base_buf_sva_mut_5_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_71_cse ) begin
      m_buf_sva_mut_6_4 <= m_buf_sva_mut_6_3;
      base_buf_sva_mut_6_4 <= base_buf_sva_mut_6_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_72_cse ) begin
      m_buf_sva_mut_7_4 <= m_buf_sva_mut_7_3;
      base_buf_sva_mut_7_4 <= base_buf_sva_mut_7_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_73_cse ) begin
      m_buf_sva_mut_8_4 <= m_buf_sva_mut_8_3;
      base_buf_sva_mut_8_4 <= base_buf_sva_mut_8_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_74_cse ) begin
      m_buf_sva_mut_9_4 <= m_buf_sva_mut_9_3;
      base_buf_sva_mut_9_4 <= base_buf_sva_mut_9_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_75_cse ) begin
      m_buf_sva_mut_10_4 <= m_buf_sva_mut_10_3;
      base_buf_sva_mut_10_4 <= base_buf_sva_mut_10_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_76_cse ) begin
      m_buf_sva_mut_4 <= m_buf_sva_mut_3;
      base_buf_sva_mut_4 <= base_buf_sva_mut_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_4 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_156 ) begin
      result_rem_11cyc_st_4 <= result_rem_11cyc_st_3;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_77_cse ) begin
      m_buf_sva_mut_1_3 <= m_buf_sva_mut_1_2;
      base_buf_sva_mut_1_3 <= base_buf_sva_mut_1_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_78_cse ) begin
      m_buf_sva_mut_2_3 <= m_buf_sva_mut_2_2;
      base_buf_sva_mut_2_3 <= base_buf_sva_mut_2_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_79_cse ) begin
      m_buf_sva_mut_3_3 <= m_buf_sva_mut_3_2;
      base_buf_sva_mut_3_3 <= base_buf_sva_mut_3_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_80_cse ) begin
      m_buf_sva_mut_4_3 <= m_buf_sva_mut_4_2;
      base_buf_sva_mut_4_3 <= base_buf_sva_mut_4_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_81_cse ) begin
      m_buf_sva_mut_5_3 <= m_buf_sva_mut_5_2;
      base_buf_sva_mut_5_3 <= base_buf_sva_mut_5_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_82_cse ) begin
      m_buf_sva_mut_6_3 <= m_buf_sva_mut_6_2;
      base_buf_sva_mut_6_3 <= base_buf_sva_mut_6_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_83_cse ) begin
      m_buf_sva_mut_7_3 <= m_buf_sva_mut_7_2;
      base_buf_sva_mut_7_3 <= base_buf_sva_mut_7_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_84_cse ) begin
      m_buf_sva_mut_8_3 <= m_buf_sva_mut_8_2;
      base_buf_sva_mut_8_3 <= base_buf_sva_mut_8_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_85_cse ) begin
      m_buf_sva_mut_9_3 <= m_buf_sva_mut_9_2;
      base_buf_sva_mut_9_3 <= base_buf_sva_mut_9_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_86_cse ) begin
      m_buf_sva_mut_10_3 <= m_buf_sva_mut_10_2;
      base_buf_sva_mut_10_3 <= base_buf_sva_mut_10_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_87_cse ) begin
      m_buf_sva_mut_3 <= m_buf_sva_mut_2;
      base_buf_sva_mut_3 <= base_buf_sva_mut_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_3 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_182 ) begin
      result_rem_11cyc_st_3 <= result_rem_11cyc_st_2;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_88_cse ) begin
      m_buf_sva_mut_1_2 <= result_rem_12_cmp_1_b;
      base_buf_sva_mut_1_2 <= result_rem_12_cmp_1_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_89_cse ) begin
      m_buf_sva_mut_2_2 <= result_rem_12_cmp_2_b;
      base_buf_sva_mut_2_2 <= result_rem_12_cmp_2_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_90_cse ) begin
      m_buf_sva_mut_3_2 <= result_rem_12_cmp_3_b;
      base_buf_sva_mut_3_2 <= result_rem_12_cmp_3_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_91_cse ) begin
      m_buf_sva_mut_4_2 <= result_rem_12_cmp_4_b;
      base_buf_sva_mut_4_2 <= result_rem_12_cmp_4_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_92_cse ) begin
      m_buf_sva_mut_5_2 <= result_rem_12_cmp_5_b;
      base_buf_sva_mut_5_2 <= result_rem_12_cmp_5_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_93_cse ) begin
      m_buf_sva_mut_6_2 <= result_rem_12_cmp_6_b;
      base_buf_sva_mut_6_2 <= result_rem_12_cmp_6_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_94_cse ) begin
      m_buf_sva_mut_7_2 <= result_rem_12_cmp_7_b;
      base_buf_sva_mut_7_2 <= result_rem_12_cmp_7_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_95_cse ) begin
      m_buf_sva_mut_8_2 <= result_rem_12_cmp_8_b;
      base_buf_sva_mut_8_2 <= result_rem_12_cmp_8_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_96_cse ) begin
      m_buf_sva_mut_9_2 <= result_rem_12_cmp_9_b;
      base_buf_sva_mut_9_2 <= result_rem_12_cmp_9_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_97_cse ) begin
      m_buf_sva_mut_10_2 <= result_rem_12_cmp_10_b;
      base_buf_sva_mut_10_2 <= result_rem_12_cmp_10_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( m_and_98_cse ) begin
      m_buf_sva_mut_2 <= result_rem_12_cmp_b;
      base_buf_sva_mut_2 <= result_rem_12_cmp_a;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc_st_2 <= 4'b0000;
    end
    else if ( ccs_ccore_en & and_dcpl_208 ) begin
      result_rem_11cyc_st_2 <= result_rem_11cyc;
    end
  end
  always @(posedge ccs_ccore_clk) begin
    if ( ccs_ccore_srst ) begin
      result_rem_11cyc <= 4'b0000;
    end
    else if ( ccs_ccore_en & ccs_ccore_start_rsci_idat ) begin
      result_rem_11cyc <= result_result_acc_tmp;
    end
  end

  function automatic [63:0] MUX1HOT_v_64_10_2;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [9:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    MUX1HOT_v_64_10_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_11_2;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [10:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    MUX1HOT_v_64_11_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] conv_s2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_s2s_3_4 = {vector[2], vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    modulo_dev
// ------------------------------------------------------------------


module modulo_dev (
  base_rsc_dat, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_clk,
      ccs_ccore_srst, ccs_ccore_en
);
  input [63:0] base_rsc_dat;
  input [63:0] m_rsc_dat;
  output [63:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_ccore_clk;
  input ccs_ccore_srst;
  input ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  modulo_dev_core modulo_dev_core_inst (
      .base_rsc_dat(base_rsc_dat),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_clk(ccs_ccore_clk),
      .ccs_ccore_srst(ccs_ccore_srst),
      .ccs_ccore_en(ccs_ccore_en)
    );
endmodule




//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Fri Aug 27 10:20:37 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen (
  q, radr, q_d, radr_d, readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output [63:0] q_d;
  input [3:0] radr_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen (
  q, radr, we, d, wadr, d_d, q_d, radr_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d,
      readA_r_ram_ir_internal_RMASK_B_d
);
  input [63:0] q;
  output [3:0] radr;
  output we;
  output [63:0] d;
  output [3:0] wadr;
  input [63:0] d_d;
  output [63:0] q_d;
  input [3:0] radr_d;
  input [3:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign q_d = q;
  assign radr = (radr_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_core_fsm (
  clk, rst, fsm_output, COMP_LOOP_C_28_tr0, COMP_LOOP_C_56_tr0, COMP_LOOP_C_84_tr0,
      COMP_LOOP_C_112_tr0, COMP_LOOP_C_140_tr0, COMP_LOOP_C_168_tr0, COMP_LOOP_C_196_tr0,
      COMP_LOOP_C_224_tr0, VEC_LOOP_C_0_tr0, STAGE_LOOP_C_1_tr0
);
  input clk;
  input rst;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;
  input COMP_LOOP_C_28_tr0;
  input COMP_LOOP_C_56_tr0;
  input COMP_LOOP_C_84_tr0;
  input COMP_LOOP_C_112_tr0;
  input COMP_LOOP_C_140_tr0;
  input COMP_LOOP_C_168_tr0;
  input COMP_LOOP_C_196_tr0;
  input COMP_LOOP_C_224_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_1_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIF_core_core_fsm_1
  parameter
    main_C_0 = 8'd0,
    STAGE_LOOP_C_0 = 8'd1,
    COMP_LOOP_C_0 = 8'd2,
    COMP_LOOP_C_1 = 8'd3,
    COMP_LOOP_C_2 = 8'd4,
    COMP_LOOP_C_3 = 8'd5,
    COMP_LOOP_C_4 = 8'd6,
    COMP_LOOP_C_5 = 8'd7,
    COMP_LOOP_C_6 = 8'd8,
    COMP_LOOP_C_7 = 8'd9,
    COMP_LOOP_C_8 = 8'd10,
    COMP_LOOP_C_9 = 8'd11,
    COMP_LOOP_C_10 = 8'd12,
    COMP_LOOP_C_11 = 8'd13,
    COMP_LOOP_C_12 = 8'd14,
    COMP_LOOP_C_13 = 8'd15,
    COMP_LOOP_C_14 = 8'd16,
    COMP_LOOP_C_15 = 8'd17,
    COMP_LOOP_C_16 = 8'd18,
    COMP_LOOP_C_17 = 8'd19,
    COMP_LOOP_C_18 = 8'd20,
    COMP_LOOP_C_19 = 8'd21,
    COMP_LOOP_C_20 = 8'd22,
    COMP_LOOP_C_21 = 8'd23,
    COMP_LOOP_C_22 = 8'd24,
    COMP_LOOP_C_23 = 8'd25,
    COMP_LOOP_C_24 = 8'd26,
    COMP_LOOP_C_25 = 8'd27,
    COMP_LOOP_C_26 = 8'd28,
    COMP_LOOP_C_27 = 8'd29,
    COMP_LOOP_C_28 = 8'd30,
    COMP_LOOP_C_29 = 8'd31,
    COMP_LOOP_C_30 = 8'd32,
    COMP_LOOP_C_31 = 8'd33,
    COMP_LOOP_C_32 = 8'd34,
    COMP_LOOP_C_33 = 8'd35,
    COMP_LOOP_C_34 = 8'd36,
    COMP_LOOP_C_35 = 8'd37,
    COMP_LOOP_C_36 = 8'd38,
    COMP_LOOP_C_37 = 8'd39,
    COMP_LOOP_C_38 = 8'd40,
    COMP_LOOP_C_39 = 8'd41,
    COMP_LOOP_C_40 = 8'd42,
    COMP_LOOP_C_41 = 8'd43,
    COMP_LOOP_C_42 = 8'd44,
    COMP_LOOP_C_43 = 8'd45,
    COMP_LOOP_C_44 = 8'd46,
    COMP_LOOP_C_45 = 8'd47,
    COMP_LOOP_C_46 = 8'd48,
    COMP_LOOP_C_47 = 8'd49,
    COMP_LOOP_C_48 = 8'd50,
    COMP_LOOP_C_49 = 8'd51,
    COMP_LOOP_C_50 = 8'd52,
    COMP_LOOP_C_51 = 8'd53,
    COMP_LOOP_C_52 = 8'd54,
    COMP_LOOP_C_53 = 8'd55,
    COMP_LOOP_C_54 = 8'd56,
    COMP_LOOP_C_55 = 8'd57,
    COMP_LOOP_C_56 = 8'd58,
    COMP_LOOP_C_57 = 8'd59,
    COMP_LOOP_C_58 = 8'd60,
    COMP_LOOP_C_59 = 8'd61,
    COMP_LOOP_C_60 = 8'd62,
    COMP_LOOP_C_61 = 8'd63,
    COMP_LOOP_C_62 = 8'd64,
    COMP_LOOP_C_63 = 8'd65,
    COMP_LOOP_C_64 = 8'd66,
    COMP_LOOP_C_65 = 8'd67,
    COMP_LOOP_C_66 = 8'd68,
    COMP_LOOP_C_67 = 8'd69,
    COMP_LOOP_C_68 = 8'd70,
    COMP_LOOP_C_69 = 8'd71,
    COMP_LOOP_C_70 = 8'd72,
    COMP_LOOP_C_71 = 8'd73,
    COMP_LOOP_C_72 = 8'd74,
    COMP_LOOP_C_73 = 8'd75,
    COMP_LOOP_C_74 = 8'd76,
    COMP_LOOP_C_75 = 8'd77,
    COMP_LOOP_C_76 = 8'd78,
    COMP_LOOP_C_77 = 8'd79,
    COMP_LOOP_C_78 = 8'd80,
    COMP_LOOP_C_79 = 8'd81,
    COMP_LOOP_C_80 = 8'd82,
    COMP_LOOP_C_81 = 8'd83,
    COMP_LOOP_C_82 = 8'd84,
    COMP_LOOP_C_83 = 8'd85,
    COMP_LOOP_C_84 = 8'd86,
    COMP_LOOP_C_85 = 8'd87,
    COMP_LOOP_C_86 = 8'd88,
    COMP_LOOP_C_87 = 8'd89,
    COMP_LOOP_C_88 = 8'd90,
    COMP_LOOP_C_89 = 8'd91,
    COMP_LOOP_C_90 = 8'd92,
    COMP_LOOP_C_91 = 8'd93,
    COMP_LOOP_C_92 = 8'd94,
    COMP_LOOP_C_93 = 8'd95,
    COMP_LOOP_C_94 = 8'd96,
    COMP_LOOP_C_95 = 8'd97,
    COMP_LOOP_C_96 = 8'd98,
    COMP_LOOP_C_97 = 8'd99,
    COMP_LOOP_C_98 = 8'd100,
    COMP_LOOP_C_99 = 8'd101,
    COMP_LOOP_C_100 = 8'd102,
    COMP_LOOP_C_101 = 8'd103,
    COMP_LOOP_C_102 = 8'd104,
    COMP_LOOP_C_103 = 8'd105,
    COMP_LOOP_C_104 = 8'd106,
    COMP_LOOP_C_105 = 8'd107,
    COMP_LOOP_C_106 = 8'd108,
    COMP_LOOP_C_107 = 8'd109,
    COMP_LOOP_C_108 = 8'd110,
    COMP_LOOP_C_109 = 8'd111,
    COMP_LOOP_C_110 = 8'd112,
    COMP_LOOP_C_111 = 8'd113,
    COMP_LOOP_C_112 = 8'd114,
    COMP_LOOP_C_113 = 8'd115,
    COMP_LOOP_C_114 = 8'd116,
    COMP_LOOP_C_115 = 8'd117,
    COMP_LOOP_C_116 = 8'd118,
    COMP_LOOP_C_117 = 8'd119,
    COMP_LOOP_C_118 = 8'd120,
    COMP_LOOP_C_119 = 8'd121,
    COMP_LOOP_C_120 = 8'd122,
    COMP_LOOP_C_121 = 8'd123,
    COMP_LOOP_C_122 = 8'd124,
    COMP_LOOP_C_123 = 8'd125,
    COMP_LOOP_C_124 = 8'd126,
    COMP_LOOP_C_125 = 8'd127,
    COMP_LOOP_C_126 = 8'd128,
    COMP_LOOP_C_127 = 8'd129,
    COMP_LOOP_C_128 = 8'd130,
    COMP_LOOP_C_129 = 8'd131,
    COMP_LOOP_C_130 = 8'd132,
    COMP_LOOP_C_131 = 8'd133,
    COMP_LOOP_C_132 = 8'd134,
    COMP_LOOP_C_133 = 8'd135,
    COMP_LOOP_C_134 = 8'd136,
    COMP_LOOP_C_135 = 8'd137,
    COMP_LOOP_C_136 = 8'd138,
    COMP_LOOP_C_137 = 8'd139,
    COMP_LOOP_C_138 = 8'd140,
    COMP_LOOP_C_139 = 8'd141,
    COMP_LOOP_C_140 = 8'd142,
    COMP_LOOP_C_141 = 8'd143,
    COMP_LOOP_C_142 = 8'd144,
    COMP_LOOP_C_143 = 8'd145,
    COMP_LOOP_C_144 = 8'd146,
    COMP_LOOP_C_145 = 8'd147,
    COMP_LOOP_C_146 = 8'd148,
    COMP_LOOP_C_147 = 8'd149,
    COMP_LOOP_C_148 = 8'd150,
    COMP_LOOP_C_149 = 8'd151,
    COMP_LOOP_C_150 = 8'd152,
    COMP_LOOP_C_151 = 8'd153,
    COMP_LOOP_C_152 = 8'd154,
    COMP_LOOP_C_153 = 8'd155,
    COMP_LOOP_C_154 = 8'd156,
    COMP_LOOP_C_155 = 8'd157,
    COMP_LOOP_C_156 = 8'd158,
    COMP_LOOP_C_157 = 8'd159,
    COMP_LOOP_C_158 = 8'd160,
    COMP_LOOP_C_159 = 8'd161,
    COMP_LOOP_C_160 = 8'd162,
    COMP_LOOP_C_161 = 8'd163,
    COMP_LOOP_C_162 = 8'd164,
    COMP_LOOP_C_163 = 8'd165,
    COMP_LOOP_C_164 = 8'd166,
    COMP_LOOP_C_165 = 8'd167,
    COMP_LOOP_C_166 = 8'd168,
    COMP_LOOP_C_167 = 8'd169,
    COMP_LOOP_C_168 = 8'd170,
    COMP_LOOP_C_169 = 8'd171,
    COMP_LOOP_C_170 = 8'd172,
    COMP_LOOP_C_171 = 8'd173,
    COMP_LOOP_C_172 = 8'd174,
    COMP_LOOP_C_173 = 8'd175,
    COMP_LOOP_C_174 = 8'd176,
    COMP_LOOP_C_175 = 8'd177,
    COMP_LOOP_C_176 = 8'd178,
    COMP_LOOP_C_177 = 8'd179,
    COMP_LOOP_C_178 = 8'd180,
    COMP_LOOP_C_179 = 8'd181,
    COMP_LOOP_C_180 = 8'd182,
    COMP_LOOP_C_181 = 8'd183,
    COMP_LOOP_C_182 = 8'd184,
    COMP_LOOP_C_183 = 8'd185,
    COMP_LOOP_C_184 = 8'd186,
    COMP_LOOP_C_185 = 8'd187,
    COMP_LOOP_C_186 = 8'd188,
    COMP_LOOP_C_187 = 8'd189,
    COMP_LOOP_C_188 = 8'd190,
    COMP_LOOP_C_189 = 8'd191,
    COMP_LOOP_C_190 = 8'd192,
    COMP_LOOP_C_191 = 8'd193,
    COMP_LOOP_C_192 = 8'd194,
    COMP_LOOP_C_193 = 8'd195,
    COMP_LOOP_C_194 = 8'd196,
    COMP_LOOP_C_195 = 8'd197,
    COMP_LOOP_C_196 = 8'd198,
    COMP_LOOP_C_197 = 8'd199,
    COMP_LOOP_C_198 = 8'd200,
    COMP_LOOP_C_199 = 8'd201,
    COMP_LOOP_C_200 = 8'd202,
    COMP_LOOP_C_201 = 8'd203,
    COMP_LOOP_C_202 = 8'd204,
    COMP_LOOP_C_203 = 8'd205,
    COMP_LOOP_C_204 = 8'd206,
    COMP_LOOP_C_205 = 8'd207,
    COMP_LOOP_C_206 = 8'd208,
    COMP_LOOP_C_207 = 8'd209,
    COMP_LOOP_C_208 = 8'd210,
    COMP_LOOP_C_209 = 8'd211,
    COMP_LOOP_C_210 = 8'd212,
    COMP_LOOP_C_211 = 8'd213,
    COMP_LOOP_C_212 = 8'd214,
    COMP_LOOP_C_213 = 8'd215,
    COMP_LOOP_C_214 = 8'd216,
    COMP_LOOP_C_215 = 8'd217,
    COMP_LOOP_C_216 = 8'd218,
    COMP_LOOP_C_217 = 8'd219,
    COMP_LOOP_C_218 = 8'd220,
    COMP_LOOP_C_219 = 8'd221,
    COMP_LOOP_C_220 = 8'd222,
    COMP_LOOP_C_221 = 8'd223,
    COMP_LOOP_C_222 = 8'd224,
    COMP_LOOP_C_223 = 8'd225,
    COMP_LOOP_C_224 = 8'd226,
    VEC_LOOP_C_0 = 8'd227,
    STAGE_LOOP_C_1 = 8'd228,
    main_C_1 = 8'd229;

  reg [7:0] state_var;
  reg [7:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIF_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 8'b00000001;
        state_var_NS = COMP_LOOP_C_0;
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 8'b00000010;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 8'b00000011;
        state_var_NS = COMP_LOOP_C_2;
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 8'b00000100;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 8'b00000101;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 8'b00000110;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 8'b00000111;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 8'b00001000;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 8'b00001001;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 8'b00001010;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 8'b00001011;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 8'b00001100;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 8'b00001101;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 8'b00001110;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 8'b00001111;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 8'b00010000;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 8'b00010001;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 8'b00010010;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 8'b00010011;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 8'b00010100;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 8'b00010101;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 8'b00010110;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 8'b00010111;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 8'b00011000;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 8'b00011001;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 8'b00011010;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 8'b00011011;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 8'b00011100;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 8'b00011101;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 8'b00011110;
        if ( COMP_LOOP_C_28_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_29;
        end
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 8'b00011111;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 8'b00100000;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 8'b00100001;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 8'b00100010;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 8'b00100011;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 8'b00100100;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 8'b00100101;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 8'b00100110;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 8'b00100111;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 8'b00101000;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 8'b00101001;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 8'b00101010;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 8'b00101011;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 8'b00101100;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 8'b00101101;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 8'b00101110;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 8'b00101111;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 8'b00110000;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 8'b00110001;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 8'b00110010;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 8'b00110011;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 8'b00110100;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 8'b00110101;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 8'b00110110;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 8'b00110111;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 8'b00111000;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 8'b00111001;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 8'b00111010;
        if ( COMP_LOOP_C_56_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_57;
        end
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 8'b00111011;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 8'b00111100;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 8'b00111101;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 8'b00111110;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 8'b00111111;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 8'b01000000;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 8'b01000001;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 8'b01000010;
        state_var_NS = COMP_LOOP_C_65;
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 8'b01000011;
        state_var_NS = COMP_LOOP_C_66;
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 8'b01000100;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 8'b01000101;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 8'b01000110;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 8'b01000111;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 8'b01001000;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 8'b01001001;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 8'b01001010;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 8'b01001011;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 8'b01001100;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 8'b01001101;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 8'b01001110;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 8'b01001111;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 8'b01010000;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 8'b01010001;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 8'b01010010;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 8'b01010011;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 8'b01010100;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 8'b01010101;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 8'b01010110;
        if ( COMP_LOOP_C_84_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_85;
        end
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 8'b01010111;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 8'b01011000;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 8'b01011001;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 8'b01011010;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 8'b01011011;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 8'b01011100;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 8'b01011101;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 8'b01011110;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 8'b01011111;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 8'b01100000;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 8'b01100001;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 8'b01100010;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 8'b01100011;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 8'b01100100;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 8'b01100101;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 8'b01100110;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 8'b01100111;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 8'b01101000;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 8'b01101001;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 8'b01101010;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 8'b01101011;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 8'b01101100;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 8'b01101101;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 8'b01101110;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 8'b01101111;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 8'b01110000;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 8'b01110001;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 8'b01110010;
        if ( COMP_LOOP_C_112_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_113;
        end
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 8'b01110011;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 8'b01110100;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 8'b01110101;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 8'b01110110;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 8'b01110111;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 8'b01111000;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 8'b01111001;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 8'b01111010;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 8'b01111011;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 8'b01111100;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 8'b01111101;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 8'b01111110;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 8'b01111111;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 8'b10000000;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 8'b10000001;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 8'b10000010;
        state_var_NS = COMP_LOOP_C_129;
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 8'b10000011;
        state_var_NS = COMP_LOOP_C_130;
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 8'b10000100;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 8'b10000101;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 8'b10000110;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 8'b10000111;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 8'b10001000;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 8'b10001001;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 8'b10001010;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 8'b10001011;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 8'b10001100;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 8'b10001101;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 8'b10001110;
        if ( COMP_LOOP_C_140_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_141;
        end
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 8'b10001111;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 8'b10010000;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 8'b10010001;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 8'b10010010;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 8'b10010011;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 8'b10010100;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 8'b10010101;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 8'b10010110;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 8'b10010111;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 8'b10011000;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 8'b10011001;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 8'b10011010;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 8'b10011011;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 8'b10011100;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 8'b10011101;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 8'b10011110;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 8'b10011111;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 8'b10100000;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 8'b10100001;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 8'b10100010;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 8'b10100011;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 8'b10100100;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 8'b10100101;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 8'b10100110;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 8'b10100111;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 8'b10101000;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 8'b10101001;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 8'b10101010;
        if ( COMP_LOOP_C_168_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_169;
        end
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 8'b10101011;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 8'b10101100;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 8'b10101101;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 8'b10101110;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 8'b10101111;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 8'b10110000;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 8'b10110001;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 8'b10110010;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 8'b10110011;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 8'b10110100;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 8'b10110101;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 8'b10110110;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 8'b10110111;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 8'b10111000;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 8'b10111001;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 8'b10111010;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 8'b10111011;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 8'b10111100;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 8'b10111101;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 8'b10111110;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 8'b10111111;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 8'b11000000;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 8'b11000001;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 8'b11000010;
        state_var_NS = COMP_LOOP_C_193;
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 8'b11000011;
        state_var_NS = COMP_LOOP_C_194;
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 8'b11000100;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 8'b11000101;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 8'b11000110;
        if ( COMP_LOOP_C_196_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_197;
        end
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 8'b11000111;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 8'b11001000;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 8'b11001001;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 8'b11001010;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 8'b11001011;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 8'b11001100;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 8'b11001101;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 8'b11001110;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 8'b11001111;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 8'b11010000;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 8'b11010001;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 8'b11010010;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 8'b11010011;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 8'b11010100;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 8'b11010101;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 8'b11010110;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 8'b11010111;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 8'b11011000;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 8'b11011001;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 8'b11011010;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 8'b11011011;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 8'b11011100;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 8'b11011101;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 8'b11011110;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 8'b11011111;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 8'b11100000;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 8'b11100001;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 8'b11100010;
        if ( COMP_LOOP_C_224_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 8'b11100011;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 8'b11100100;
        if ( STAGE_LOOP_C_1_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 8'b11100101;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 8'b00000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core_wait_dp
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core_wait_dp (
  ensig_cgo_iro, ensig_cgo, COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en
);
  input ensig_cgo_iro;
  input ensig_cgo;
  output COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en;



  // Interconnect Declarations for Component Instantiations 
  assign COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en = ensig_cgo | ensig_cgo_iro;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF_core
// ------------------------------------------------------------------


module inPlaceNTT_DIF_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, vec_rsc_triosy_0_16_lz, vec_rsc_triosy_0_17_lz, vec_rsc_triosy_0_18_lz,
      vec_rsc_triosy_0_19_lz, vec_rsc_triosy_0_20_lz, vec_rsc_triosy_0_21_lz, vec_rsc_triosy_0_22_lz,
      vec_rsc_triosy_0_23_lz, vec_rsc_triosy_0_24_lz, vec_rsc_triosy_0_25_lz, vec_rsc_triosy_0_26_lz,
      vec_rsc_triosy_0_27_lz, vec_rsc_triosy_0_28_lz, vec_rsc_triosy_0_29_lz, vec_rsc_triosy_0_30_lz,
      vec_rsc_triosy_0_31_lz, vec_rsc_triosy_0_32_lz, vec_rsc_triosy_0_33_lz, vec_rsc_triosy_0_34_lz,
      vec_rsc_triosy_0_35_lz, vec_rsc_triosy_0_36_lz, vec_rsc_triosy_0_37_lz, vec_rsc_triosy_0_38_lz,
      vec_rsc_triosy_0_39_lz, vec_rsc_triosy_0_40_lz, vec_rsc_triosy_0_41_lz, vec_rsc_triosy_0_42_lz,
      vec_rsc_triosy_0_43_lz, vec_rsc_triosy_0_44_lz, vec_rsc_triosy_0_45_lz, vec_rsc_triosy_0_46_lz,
      vec_rsc_triosy_0_47_lz, vec_rsc_triosy_0_48_lz, vec_rsc_triosy_0_49_lz, vec_rsc_triosy_0_50_lz,
      vec_rsc_triosy_0_51_lz, vec_rsc_triosy_0_52_lz, vec_rsc_triosy_0_53_lz, vec_rsc_triosy_0_54_lz,
      vec_rsc_triosy_0_55_lz, vec_rsc_triosy_0_56_lz, vec_rsc_triosy_0_57_lz, vec_rsc_triosy_0_58_lz,
      vec_rsc_triosy_0_59_lz, vec_rsc_triosy_0_60_lz, vec_rsc_triosy_0_61_lz, vec_rsc_triosy_0_62_lz,
      vec_rsc_triosy_0_63_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_triosy_0_2_lz, twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_triosy_0_4_lz, twiddle_rsc_triosy_0_5_lz, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_triosy_0_7_lz, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_triosy_0_10_lz, twiddle_rsc_triosy_0_11_lz, twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_triosy_0_13_lz, twiddle_rsc_triosy_0_14_lz, twiddle_rsc_triosy_0_15_lz,
      twiddle_rsc_triosy_0_16_lz, twiddle_rsc_triosy_0_17_lz, twiddle_rsc_triosy_0_18_lz,
      twiddle_rsc_triosy_0_19_lz, twiddle_rsc_triosy_0_20_lz, twiddle_rsc_triosy_0_21_lz,
      twiddle_rsc_triosy_0_22_lz, twiddle_rsc_triosy_0_23_lz, twiddle_rsc_triosy_0_24_lz,
      twiddle_rsc_triosy_0_25_lz, twiddle_rsc_triosy_0_26_lz, twiddle_rsc_triosy_0_27_lz,
      twiddle_rsc_triosy_0_28_lz, twiddle_rsc_triosy_0_29_lz, twiddle_rsc_triosy_0_30_lz,
      twiddle_rsc_triosy_0_31_lz, twiddle_rsc_triosy_0_32_lz, twiddle_rsc_triosy_0_33_lz,
      twiddle_rsc_triosy_0_34_lz, twiddle_rsc_triosy_0_35_lz, twiddle_rsc_triosy_0_36_lz,
      twiddle_rsc_triosy_0_37_lz, twiddle_rsc_triosy_0_38_lz, twiddle_rsc_triosy_0_39_lz,
      twiddle_rsc_triosy_0_40_lz, twiddle_rsc_triosy_0_41_lz, twiddle_rsc_triosy_0_42_lz,
      twiddle_rsc_triosy_0_43_lz, twiddle_rsc_triosy_0_44_lz, twiddle_rsc_triosy_0_45_lz,
      twiddle_rsc_triosy_0_46_lz, twiddle_rsc_triosy_0_47_lz, twiddle_rsc_triosy_0_48_lz,
      twiddle_rsc_triosy_0_49_lz, twiddle_rsc_triosy_0_50_lz, twiddle_rsc_triosy_0_51_lz,
      twiddle_rsc_triosy_0_52_lz, twiddle_rsc_triosy_0_53_lz, twiddle_rsc_triosy_0_54_lz,
      twiddle_rsc_triosy_0_55_lz, twiddle_rsc_triosy_0_56_lz, twiddle_rsc_triosy_0_57_lz,
      twiddle_rsc_triosy_0_58_lz, twiddle_rsc_triosy_0_59_lz, twiddle_rsc_triosy_0_60_lz,
      twiddle_rsc_triosy_0_61_lz, twiddle_rsc_triosy_0_62_lz, twiddle_rsc_triosy_0_63_lz,
      vec_rsc_0_0_i_q_d, vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_q_d,
      vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_q_d, vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_q_d,
      vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_q_d, vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_q_d, vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_q_d,
      vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_q_d, vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_q_d, vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_q_d, vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_q_d, vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_13_i_q_d,
      vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_q_d, vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_16_i_q_d,
      vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_17_i_q_d, vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_18_i_q_d, vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_19_i_q_d,
      vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_20_i_q_d, vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_21_i_q_d, vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_22_i_q_d,
      vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_23_i_q_d, vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_24_i_q_d, vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_25_i_q_d,
      vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_26_i_q_d, vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_27_i_q_d, vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_28_i_q_d,
      vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_29_i_q_d, vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_30_i_q_d, vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_31_i_q_d,
      vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_32_i_q_d, vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_33_i_q_d, vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_34_i_q_d,
      vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_35_i_q_d, vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_36_i_q_d, vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_37_i_q_d,
      vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_38_i_q_d, vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_39_i_q_d, vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_40_i_q_d,
      vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_41_i_q_d, vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_42_i_q_d, vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_43_i_q_d,
      vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_44_i_q_d, vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_45_i_q_d, vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_46_i_q_d,
      vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_47_i_q_d, vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_48_i_q_d, vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_49_i_q_d,
      vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_50_i_q_d, vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_51_i_q_d, vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_52_i_q_d,
      vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_53_i_q_d, vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_54_i_q_d, vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_55_i_q_d,
      vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_56_i_q_d, vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_57_i_q_d, vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_58_i_q_d,
      vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_59_i_q_d, vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_60_i_q_d, vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_61_i_q_d,
      vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_62_i_q_d, vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_63_i_q_d, vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_0_i_q_d,
      twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_1_i_q_d,
      twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_2_i_q_d,
      twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_3_i_q_d,
      twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_4_i_q_d,
      twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_5_i_q_d,
      twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_6_i_q_d,
      twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_7_i_q_d,
      twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_8_i_q_d,
      twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_9_i_q_d,
      twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_10_i_q_d,
      twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_11_i_q_d,
      twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_12_i_q_d,
      twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_13_i_q_d,
      twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_14_i_q_d,
      twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_15_i_q_d,
      twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_16_i_q_d,
      twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_17_i_q_d,
      twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_18_i_q_d,
      twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_19_i_q_d,
      twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_20_i_q_d,
      twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_21_i_q_d,
      twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_22_i_q_d,
      twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_23_i_q_d,
      twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_24_i_q_d,
      twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_25_i_q_d,
      twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_26_i_q_d,
      twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_27_i_q_d,
      twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_28_i_q_d,
      twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_29_i_q_d,
      twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_30_i_q_d,
      twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_31_i_q_d,
      twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_32_i_q_d,
      twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_33_i_q_d,
      twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_34_i_q_d,
      twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_35_i_q_d,
      twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_36_i_q_d,
      twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_37_i_q_d,
      twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_38_i_q_d,
      twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_39_i_q_d,
      twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_40_i_q_d,
      twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_41_i_q_d,
      twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_42_i_q_d,
      twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_43_i_q_d,
      twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_44_i_q_d,
      twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_45_i_q_d,
      twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_46_i_q_d,
      twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_47_i_q_d,
      twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_48_i_q_d,
      twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_49_i_q_d,
      twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_50_i_q_d,
      twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_51_i_q_d,
      twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_52_i_q_d,
      twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_53_i_q_d,
      twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_54_i_q_d,
      twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_55_i_q_d,
      twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_56_i_q_d,
      twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_57_i_q_d,
      twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_58_i_q_d,
      twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_59_i_q_d,
      twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_60_i_q_d,
      twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_61_i_q_d,
      twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_62_i_q_d,
      twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d, twiddle_rsc_0_63_i_q_d,
      twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_d_d_pff,
      vec_rsc_0_0_i_radr_d_pff, vec_rsc_0_0_i_wadr_d_pff, vec_rsc_0_0_i_we_d_pff,
      vec_rsc_0_1_i_we_d_pff, vec_rsc_0_2_i_we_d_pff, vec_rsc_0_3_i_we_d_pff, vec_rsc_0_4_i_we_d_pff,
      vec_rsc_0_5_i_we_d_pff, vec_rsc_0_6_i_we_d_pff, vec_rsc_0_7_i_we_d_pff, vec_rsc_0_8_i_we_d_pff,
      vec_rsc_0_9_i_we_d_pff, vec_rsc_0_10_i_we_d_pff, vec_rsc_0_11_i_we_d_pff, vec_rsc_0_12_i_we_d_pff,
      vec_rsc_0_13_i_we_d_pff, vec_rsc_0_14_i_we_d_pff, vec_rsc_0_15_i_we_d_pff,
      vec_rsc_0_16_i_we_d_pff, vec_rsc_0_17_i_we_d_pff, vec_rsc_0_18_i_we_d_pff,
      vec_rsc_0_19_i_we_d_pff, vec_rsc_0_20_i_we_d_pff, vec_rsc_0_21_i_we_d_pff,
      vec_rsc_0_22_i_we_d_pff, vec_rsc_0_23_i_we_d_pff, vec_rsc_0_24_i_we_d_pff,
      vec_rsc_0_25_i_we_d_pff, vec_rsc_0_26_i_we_d_pff, vec_rsc_0_27_i_we_d_pff,
      vec_rsc_0_28_i_we_d_pff, vec_rsc_0_29_i_we_d_pff, vec_rsc_0_30_i_we_d_pff,
      vec_rsc_0_31_i_we_d_pff, vec_rsc_0_32_i_we_d_pff, vec_rsc_0_33_i_we_d_pff,
      vec_rsc_0_34_i_we_d_pff, vec_rsc_0_35_i_we_d_pff, vec_rsc_0_36_i_we_d_pff,
      vec_rsc_0_37_i_we_d_pff, vec_rsc_0_38_i_we_d_pff, vec_rsc_0_39_i_we_d_pff,
      vec_rsc_0_40_i_we_d_pff, vec_rsc_0_41_i_we_d_pff, vec_rsc_0_42_i_we_d_pff,
      vec_rsc_0_43_i_we_d_pff, vec_rsc_0_44_i_we_d_pff, vec_rsc_0_45_i_we_d_pff,
      vec_rsc_0_46_i_we_d_pff, vec_rsc_0_47_i_we_d_pff, vec_rsc_0_48_i_we_d_pff,
      vec_rsc_0_49_i_we_d_pff, vec_rsc_0_50_i_we_d_pff, vec_rsc_0_51_i_we_d_pff,
      vec_rsc_0_52_i_we_d_pff, vec_rsc_0_53_i_we_d_pff, vec_rsc_0_54_i_we_d_pff,
      vec_rsc_0_55_i_we_d_pff, vec_rsc_0_56_i_we_d_pff, vec_rsc_0_57_i_we_d_pff,
      vec_rsc_0_58_i_we_d_pff, vec_rsc_0_59_i_we_d_pff, vec_rsc_0_60_i_we_d_pff,
      vec_rsc_0_61_i_we_d_pff, vec_rsc_0_62_i_we_d_pff, vec_rsc_0_63_i_we_d_pff,
      twiddle_rsc_0_0_i_radr_d_pff, twiddle_rsc_0_1_i_radr_d_pff, twiddle_rsc_0_2_i_radr_d_pff,
      twiddle_rsc_0_4_i_radr_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  output vec_rsc_triosy_0_16_lz;
  output vec_rsc_triosy_0_17_lz;
  output vec_rsc_triosy_0_18_lz;
  output vec_rsc_triosy_0_19_lz;
  output vec_rsc_triosy_0_20_lz;
  output vec_rsc_triosy_0_21_lz;
  output vec_rsc_triosy_0_22_lz;
  output vec_rsc_triosy_0_23_lz;
  output vec_rsc_triosy_0_24_lz;
  output vec_rsc_triosy_0_25_lz;
  output vec_rsc_triosy_0_26_lz;
  output vec_rsc_triosy_0_27_lz;
  output vec_rsc_triosy_0_28_lz;
  output vec_rsc_triosy_0_29_lz;
  output vec_rsc_triosy_0_30_lz;
  output vec_rsc_triosy_0_31_lz;
  output vec_rsc_triosy_0_32_lz;
  output vec_rsc_triosy_0_33_lz;
  output vec_rsc_triosy_0_34_lz;
  output vec_rsc_triosy_0_35_lz;
  output vec_rsc_triosy_0_36_lz;
  output vec_rsc_triosy_0_37_lz;
  output vec_rsc_triosy_0_38_lz;
  output vec_rsc_triosy_0_39_lz;
  output vec_rsc_triosy_0_40_lz;
  output vec_rsc_triosy_0_41_lz;
  output vec_rsc_triosy_0_42_lz;
  output vec_rsc_triosy_0_43_lz;
  output vec_rsc_triosy_0_44_lz;
  output vec_rsc_triosy_0_45_lz;
  output vec_rsc_triosy_0_46_lz;
  output vec_rsc_triosy_0_47_lz;
  output vec_rsc_triosy_0_48_lz;
  output vec_rsc_triosy_0_49_lz;
  output vec_rsc_triosy_0_50_lz;
  output vec_rsc_triosy_0_51_lz;
  output vec_rsc_triosy_0_52_lz;
  output vec_rsc_triosy_0_53_lz;
  output vec_rsc_triosy_0_54_lz;
  output vec_rsc_triosy_0_55_lz;
  output vec_rsc_triosy_0_56_lz;
  output vec_rsc_triosy_0_57_lz;
  output vec_rsc_triosy_0_58_lz;
  output vec_rsc_triosy_0_59_lz;
  output vec_rsc_triosy_0_60_lz;
  output vec_rsc_triosy_0_61_lz;
  output vec_rsc_triosy_0_62_lz;
  output vec_rsc_triosy_0_63_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_0_0_lz;
  output twiddle_rsc_triosy_0_1_lz;
  output twiddle_rsc_triosy_0_2_lz;
  output twiddle_rsc_triosy_0_3_lz;
  output twiddle_rsc_triosy_0_4_lz;
  output twiddle_rsc_triosy_0_5_lz;
  output twiddle_rsc_triosy_0_6_lz;
  output twiddle_rsc_triosy_0_7_lz;
  output twiddle_rsc_triosy_0_8_lz;
  output twiddle_rsc_triosy_0_9_lz;
  output twiddle_rsc_triosy_0_10_lz;
  output twiddle_rsc_triosy_0_11_lz;
  output twiddle_rsc_triosy_0_12_lz;
  output twiddle_rsc_triosy_0_13_lz;
  output twiddle_rsc_triosy_0_14_lz;
  output twiddle_rsc_triosy_0_15_lz;
  output twiddle_rsc_triosy_0_16_lz;
  output twiddle_rsc_triosy_0_17_lz;
  output twiddle_rsc_triosy_0_18_lz;
  output twiddle_rsc_triosy_0_19_lz;
  output twiddle_rsc_triosy_0_20_lz;
  output twiddle_rsc_triosy_0_21_lz;
  output twiddle_rsc_triosy_0_22_lz;
  output twiddle_rsc_triosy_0_23_lz;
  output twiddle_rsc_triosy_0_24_lz;
  output twiddle_rsc_triosy_0_25_lz;
  output twiddle_rsc_triosy_0_26_lz;
  output twiddle_rsc_triosy_0_27_lz;
  output twiddle_rsc_triosy_0_28_lz;
  output twiddle_rsc_triosy_0_29_lz;
  output twiddle_rsc_triosy_0_30_lz;
  output twiddle_rsc_triosy_0_31_lz;
  output twiddle_rsc_triosy_0_32_lz;
  output twiddle_rsc_triosy_0_33_lz;
  output twiddle_rsc_triosy_0_34_lz;
  output twiddle_rsc_triosy_0_35_lz;
  output twiddle_rsc_triosy_0_36_lz;
  output twiddle_rsc_triosy_0_37_lz;
  output twiddle_rsc_triosy_0_38_lz;
  output twiddle_rsc_triosy_0_39_lz;
  output twiddle_rsc_triosy_0_40_lz;
  output twiddle_rsc_triosy_0_41_lz;
  output twiddle_rsc_triosy_0_42_lz;
  output twiddle_rsc_triosy_0_43_lz;
  output twiddle_rsc_triosy_0_44_lz;
  output twiddle_rsc_triosy_0_45_lz;
  output twiddle_rsc_triosy_0_46_lz;
  output twiddle_rsc_triosy_0_47_lz;
  output twiddle_rsc_triosy_0_48_lz;
  output twiddle_rsc_triosy_0_49_lz;
  output twiddle_rsc_triosy_0_50_lz;
  output twiddle_rsc_triosy_0_51_lz;
  output twiddle_rsc_triosy_0_52_lz;
  output twiddle_rsc_triosy_0_53_lz;
  output twiddle_rsc_triosy_0_54_lz;
  output twiddle_rsc_triosy_0_55_lz;
  output twiddle_rsc_triosy_0_56_lz;
  output twiddle_rsc_triosy_0_57_lz;
  output twiddle_rsc_triosy_0_58_lz;
  output twiddle_rsc_triosy_0_59_lz;
  output twiddle_rsc_triosy_0_60_lz;
  output twiddle_rsc_triosy_0_61_lz;
  output twiddle_rsc_triosy_0_62_lz;
  output twiddle_rsc_triosy_0_63_lz;
  input [63:0] vec_rsc_0_0_i_q_d;
  output vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_q_d;
  output vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_q_d;
  output vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_q_d;
  output vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_q_d;
  output vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_q_d;
  output vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_q_d;
  output vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_q_d;
  output vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_q_d;
  output vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_q_d;
  output vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_q_d;
  output vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_q_d;
  output vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_q_d;
  output vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_q_d;
  output vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_q_d;
  output vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_q_d;
  output vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_16_i_q_d;
  output vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_17_i_q_d;
  output vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_18_i_q_d;
  output vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_19_i_q_d;
  output vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_20_i_q_d;
  output vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_21_i_q_d;
  output vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_22_i_q_d;
  output vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_23_i_q_d;
  output vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_24_i_q_d;
  output vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_25_i_q_d;
  output vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_26_i_q_d;
  output vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_27_i_q_d;
  output vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_28_i_q_d;
  output vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_29_i_q_d;
  output vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_30_i_q_d;
  output vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_31_i_q_d;
  output vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_32_i_q_d;
  output vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_33_i_q_d;
  output vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_34_i_q_d;
  output vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_35_i_q_d;
  output vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_36_i_q_d;
  output vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_37_i_q_d;
  output vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_38_i_q_d;
  output vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_39_i_q_d;
  output vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_40_i_q_d;
  output vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_41_i_q_d;
  output vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_42_i_q_d;
  output vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_43_i_q_d;
  output vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_44_i_q_d;
  output vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_45_i_q_d;
  output vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_46_i_q_d;
  output vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_47_i_q_d;
  output vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_48_i_q_d;
  output vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_49_i_q_d;
  output vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_50_i_q_d;
  output vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_51_i_q_d;
  output vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_52_i_q_d;
  output vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_53_i_q_d;
  output vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_54_i_q_d;
  output vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_55_i_q_d;
  output vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_56_i_q_d;
  output vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_57_i_q_d;
  output vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_58_i_q_d;
  output vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_59_i_q_d;
  output vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_60_i_q_d;
  output vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_61_i_q_d;
  output vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_62_i_q_d;
  output vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_63_i_q_d;
  output vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_0_i_q_d;
  output twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_1_i_q_d;
  output twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_2_i_q_d;
  output twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_3_i_q_d;
  output twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_4_i_q_d;
  output twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_5_i_q_d;
  output twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_6_i_q_d;
  output twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_7_i_q_d;
  output twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_8_i_q_d;
  output twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_9_i_q_d;
  output twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_10_i_q_d;
  output twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_11_i_q_d;
  output twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_12_i_q_d;
  output twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_13_i_q_d;
  output twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_14_i_q_d;
  output twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_15_i_q_d;
  output twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_16_i_q_d;
  output twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_17_i_q_d;
  output twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_18_i_q_d;
  output twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_19_i_q_d;
  output twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_20_i_q_d;
  output twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_21_i_q_d;
  output twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_22_i_q_d;
  output twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_23_i_q_d;
  output twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_24_i_q_d;
  output twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_25_i_q_d;
  output twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_26_i_q_d;
  output twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_27_i_q_d;
  output twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_28_i_q_d;
  output twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_29_i_q_d;
  output twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_30_i_q_d;
  output twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_31_i_q_d;
  output twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_32_i_q_d;
  output twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_33_i_q_d;
  output twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_34_i_q_d;
  output twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_35_i_q_d;
  output twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_36_i_q_d;
  output twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_37_i_q_d;
  output twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_38_i_q_d;
  output twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_39_i_q_d;
  output twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_40_i_q_d;
  output twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_41_i_q_d;
  output twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_42_i_q_d;
  output twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_43_i_q_d;
  output twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_44_i_q_d;
  output twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_45_i_q_d;
  output twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_46_i_q_d;
  output twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_47_i_q_d;
  output twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_48_i_q_d;
  output twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_49_i_q_d;
  output twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_50_i_q_d;
  output twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_51_i_q_d;
  output twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_52_i_q_d;
  output twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_53_i_q_d;
  output twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_54_i_q_d;
  output twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_55_i_q_d;
  output twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_56_i_q_d;
  output twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_57_i_q_d;
  output twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_58_i_q_d;
  output twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_59_i_q_d;
  output twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_60_i_q_d;
  output twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_61_i_q_d;
  output twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_62_i_q_d;
  output twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d;
  input [63:0] twiddle_rsc_0_63_i_q_d;
  output twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d;
  output [63:0] vec_rsc_0_0_i_d_d_pff;
  output [3:0] vec_rsc_0_0_i_radr_d_pff;
  output [3:0] vec_rsc_0_0_i_wadr_d_pff;
  output vec_rsc_0_0_i_we_d_pff;
  output vec_rsc_0_1_i_we_d_pff;
  output vec_rsc_0_2_i_we_d_pff;
  output vec_rsc_0_3_i_we_d_pff;
  output vec_rsc_0_4_i_we_d_pff;
  output vec_rsc_0_5_i_we_d_pff;
  output vec_rsc_0_6_i_we_d_pff;
  output vec_rsc_0_7_i_we_d_pff;
  output vec_rsc_0_8_i_we_d_pff;
  output vec_rsc_0_9_i_we_d_pff;
  output vec_rsc_0_10_i_we_d_pff;
  output vec_rsc_0_11_i_we_d_pff;
  output vec_rsc_0_12_i_we_d_pff;
  output vec_rsc_0_13_i_we_d_pff;
  output vec_rsc_0_14_i_we_d_pff;
  output vec_rsc_0_15_i_we_d_pff;
  output vec_rsc_0_16_i_we_d_pff;
  output vec_rsc_0_17_i_we_d_pff;
  output vec_rsc_0_18_i_we_d_pff;
  output vec_rsc_0_19_i_we_d_pff;
  output vec_rsc_0_20_i_we_d_pff;
  output vec_rsc_0_21_i_we_d_pff;
  output vec_rsc_0_22_i_we_d_pff;
  output vec_rsc_0_23_i_we_d_pff;
  output vec_rsc_0_24_i_we_d_pff;
  output vec_rsc_0_25_i_we_d_pff;
  output vec_rsc_0_26_i_we_d_pff;
  output vec_rsc_0_27_i_we_d_pff;
  output vec_rsc_0_28_i_we_d_pff;
  output vec_rsc_0_29_i_we_d_pff;
  output vec_rsc_0_30_i_we_d_pff;
  output vec_rsc_0_31_i_we_d_pff;
  output vec_rsc_0_32_i_we_d_pff;
  output vec_rsc_0_33_i_we_d_pff;
  output vec_rsc_0_34_i_we_d_pff;
  output vec_rsc_0_35_i_we_d_pff;
  output vec_rsc_0_36_i_we_d_pff;
  output vec_rsc_0_37_i_we_d_pff;
  output vec_rsc_0_38_i_we_d_pff;
  output vec_rsc_0_39_i_we_d_pff;
  output vec_rsc_0_40_i_we_d_pff;
  output vec_rsc_0_41_i_we_d_pff;
  output vec_rsc_0_42_i_we_d_pff;
  output vec_rsc_0_43_i_we_d_pff;
  output vec_rsc_0_44_i_we_d_pff;
  output vec_rsc_0_45_i_we_d_pff;
  output vec_rsc_0_46_i_we_d_pff;
  output vec_rsc_0_47_i_we_d_pff;
  output vec_rsc_0_48_i_we_d_pff;
  output vec_rsc_0_49_i_we_d_pff;
  output vec_rsc_0_50_i_we_d_pff;
  output vec_rsc_0_51_i_we_d_pff;
  output vec_rsc_0_52_i_we_d_pff;
  output vec_rsc_0_53_i_we_d_pff;
  output vec_rsc_0_54_i_we_d_pff;
  output vec_rsc_0_55_i_we_d_pff;
  output vec_rsc_0_56_i_we_d_pff;
  output vec_rsc_0_57_i_we_d_pff;
  output vec_rsc_0_58_i_we_d_pff;
  output vec_rsc_0_59_i_we_d_pff;
  output vec_rsc_0_60_i_we_d_pff;
  output vec_rsc_0_61_i_we_d_pff;
  output vec_rsc_0_62_i_we_d_pff;
  output vec_rsc_0_63_i_we_d_pff;
  output [3:0] twiddle_rsc_0_0_i_radr_d_pff;
  output [3:0] twiddle_rsc_0_1_i_radr_d_pff;
  output [3:0] twiddle_rsc_0_2_i_radr_d_pff;
  output [3:0] twiddle_rsc_0_4_i_radr_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] COMP_LOOP_1_modulo_dev_cmp_return_rsc_z;
  wire COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en;
  wire [7:0] fsm_output;
  wire nor_tmp_1;
  wire mux_tmp_6;
  wire and_dcpl_8;
  wire and_tmp_10;
  wire or_tmp_105;
  wire or_tmp_118;
  wire or_tmp_119;
  wire not_tmp_88;
  wire nor_tmp_99;
  wire mux_tmp_206;
  wire mux_tmp_293;
  wire mux_tmp_444;
  wire or_tmp_404;
  wire mux_tmp_656;
  wire and_dcpl_55;
  wire and_dcpl_57;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_62;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_tmp_29;
  wire mux_tmp_720;
  wire and_dcpl_72;
  wire and_dcpl_73;
  wire and_dcpl_74;
  wire and_dcpl_75;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_78;
  wire and_dcpl_79;
  wire and_dcpl_80;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_87;
  wire and_dcpl_88;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_94;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire and_dcpl_97;
  wire and_dcpl_99;
  wire and_dcpl_101;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire and_dcpl_106;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_110;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire or_tmp_491;
  wire or_tmp_495;
  wire or_tmp_497;
  wire or_tmp_501;
  wire or_tmp_535;
  wire or_tmp_539;
  wire or_tmp_541;
  wire or_tmp_545;
  wire not_tmp_321;
  wire or_tmp_579;
  wire or_tmp_583;
  wire or_tmp_585;
  wire or_tmp_589;
  wire or_tmp_623;
  wire or_tmp_627;
  wire or_tmp_629;
  wire or_tmp_633;
  wire not_tmp_330;
  wire or_tmp_667;
  wire or_tmp_671;
  wire or_tmp_673;
  wire or_tmp_677;
  wire or_tmp_711;
  wire or_tmp_715;
  wire or_tmp_717;
  wire or_tmp_721;
  wire or_tmp_755;
  wire or_tmp_759;
  wire or_tmp_761;
  wire or_tmp_765;
  wire or_tmp_799;
  wire or_tmp_803;
  wire or_tmp_805;
  wire or_tmp_809;
  wire not_tmp_347;
  wire or_tmp_843;
  wire or_tmp_847;
  wire or_tmp_849;
  wire or_tmp_853;
  wire or_tmp_887;
  wire or_tmp_891;
  wire or_tmp_893;
  wire or_tmp_897;
  wire or_tmp_931;
  wire or_tmp_935;
  wire or_tmp_937;
  wire or_tmp_941;
  wire or_tmp_975;
  wire or_tmp_979;
  wire or_tmp_981;
  wire or_tmp_985;
  wire or_tmp_1019;
  wire or_tmp_1023;
  wire or_tmp_1025;
  wire or_tmp_1029;
  wire or_tmp_1063;
  wire or_tmp_1067;
  wire or_tmp_1069;
  wire or_tmp_1073;
  wire or_tmp_1107;
  wire or_tmp_1111;
  wire or_tmp_1113;
  wire or_tmp_1117;
  wire or_tmp_1151;
  wire or_tmp_1155;
  wire or_tmp_1157;
  wire or_tmp_1161;
  wire or_tmp_1195;
  wire or_tmp_1199;
  wire or_tmp_1201;
  wire or_tmp_1205;
  wire not_tmp_384;
  wire not_tmp_388;
  wire or_tmp_1239;
  wire or_tmp_1243;
  wire or_tmp_1245;
  wire or_tmp_1249;
  wire or_tmp_1283;
  wire or_tmp_1287;
  wire or_tmp_1289;
  wire or_tmp_1293;
  wire or_tmp_1327;
  wire or_tmp_1331;
  wire or_tmp_1333;
  wire or_tmp_1337;
  wire or_tmp_1371;
  wire or_tmp_1375;
  wire or_tmp_1377;
  wire or_tmp_1381;
  wire or_tmp_1415;
  wire or_tmp_1419;
  wire or_tmp_1421;
  wire or_tmp_1425;
  wire or_tmp_1459;
  wire or_tmp_1463;
  wire or_tmp_1465;
  wire or_tmp_1469;
  wire or_tmp_1503;
  wire or_tmp_1507;
  wire or_tmp_1509;
  wire or_tmp_1513;
  wire not_tmp_414;
  wire or_tmp_1547;
  wire or_tmp_1551;
  wire or_tmp_1553;
  wire or_tmp_1557;
  wire or_tmp_1591;
  wire or_tmp_1595;
  wire or_tmp_1597;
  wire or_tmp_1601;
  wire or_tmp_1635;
  wire or_tmp_1639;
  wire or_tmp_1641;
  wire or_tmp_1645;
  wire or_tmp_1679;
  wire or_tmp_1683;
  wire or_tmp_1685;
  wire or_tmp_1689;
  wire or_tmp_1723;
  wire or_tmp_1727;
  wire or_tmp_1729;
  wire or_tmp_1733;
  wire or_tmp_1767;
  wire or_tmp_1771;
  wire or_tmp_1773;
  wire or_tmp_1777;
  wire or_tmp_1811;
  wire or_tmp_1815;
  wire or_tmp_1817;
  wire or_tmp_1821;
  wire or_tmp_1855;
  wire or_tmp_1859;
  wire or_tmp_1861;
  wire or_tmp_1865;
  wire or_tmp_1898;
  wire or_tmp_1902;
  wire or_tmp_1904;
  wire not_tmp_452;
  wire not_tmp_453;
  wire or_tmp_1908;
  wire or_tmp_1942;
  wire or_tmp_1946;
  wire or_tmp_1948;
  wire not_tmp_458;
  wire or_tmp_1952;
  wire or_tmp_1986;
  wire or_tmp_1990;
  wire or_tmp_1992;
  wire or_tmp_1996;
  wire or_tmp_2030;
  wire or_tmp_2034;
  wire or_tmp_2036;
  wire not_tmp_467;
  wire or_tmp_2040;
  wire or_tmp_2074;
  wire or_tmp_2078;
  wire or_tmp_2080;
  wire or_tmp_2084;
  wire or_tmp_2118;
  wire or_tmp_2122;
  wire or_tmp_2124;
  wire or_tmp_2128;
  wire or_tmp_2162;
  wire or_tmp_2166;
  wire or_tmp_2168;
  wire or_tmp_2172;
  wire or_tmp_2206;
  wire or_tmp_2210;
  wire or_tmp_2212;
  wire not_tmp_484;
  wire or_tmp_2216;
  wire or_tmp_2250;
  wire or_tmp_2254;
  wire or_tmp_2256;
  wire or_tmp_2260;
  wire or_tmp_2294;
  wire or_tmp_2298;
  wire or_tmp_2300;
  wire or_tmp_2304;
  wire or_tmp_2338;
  wire or_tmp_2342;
  wire or_tmp_2344;
  wire or_tmp_2348;
  wire or_tmp_2382;
  wire or_tmp_2386;
  wire or_tmp_2388;
  wire or_tmp_2392;
  wire or_tmp_2426;
  wire or_tmp_2430;
  wire or_tmp_2432;
  wire or_tmp_2436;
  wire or_tmp_2470;
  wire or_tmp_2474;
  wire or_tmp_2476;
  wire or_tmp_2480;
  wire or_tmp_2514;
  wire or_tmp_2518;
  wire or_tmp_2520;
  wire or_tmp_2524;
  wire or_tmp_2558;
  wire or_tmp_2562;
  wire or_tmp_2564;
  wire or_tmp_2567;
  wire or_tmp_2601;
  wire or_tmp_2605;
  wire or_tmp_2607;
  wire not_tmp_522;
  wire or_tmp_2611;
  wire not_tmp_523;
  wire not_tmp_527;
  wire or_tmp_2645;
  wire or_tmp_2649;
  wire or_tmp_2651;
  wire or_tmp_2655;
  wire or_tmp_2689;
  wire or_tmp_2693;
  wire or_tmp_2695;
  wire or_tmp_2699;
  wire or_tmp_2733;
  wire or_tmp_2737;
  wire or_tmp_2739;
  wire or_tmp_2743;
  wire or_tmp_2777;
  wire or_tmp_2781;
  wire or_tmp_2783;
  wire or_tmp_2787;
  wire not_tmp_544;
  wire or_tmp_2821;
  wire or_tmp_2825;
  wire or_tmp_2827;
  wire or_tmp_2831;
  wire not_tmp_549;
  wire or_tmp_2865;
  wire or_tmp_2869;
  wire or_tmp_2871;
  wire or_tmp_2875;
  wire or_tmp_2909;
  wire or_tmp_2913;
  wire or_tmp_2915;
  wire or_tmp_2919;
  wire or_tmp_2953;
  wire or_tmp_2957;
  wire or_tmp_2959;
  wire not_tmp_559;
  wire or_tmp_2963;
  wire not_tmp_560;
  wire or_tmp_2997;
  wire or_tmp_3001;
  wire or_tmp_3003;
  wire not_tmp_565;
  wire or_tmp_3007;
  wire or_tmp_3041;
  wire or_tmp_3045;
  wire or_tmp_3047;
  wire or_tmp_3051;
  wire not_tmp_570;
  wire or_tmp_3085;
  wire or_tmp_3089;
  wire or_tmp_3091;
  wire not_tmp_575;
  wire or_tmp_3094;
  wire or_tmp_3128;
  wire or_tmp_3132;
  wire or_tmp_3134;
  wire or_tmp_3138;
  wire or_tmp_3172;
  wire or_tmp_3176;
  wire or_tmp_3178;
  wire or_tmp_3182;
  wire or_tmp_3215;
  wire or_tmp_3219;
  wire or_tmp_3221;
  wire or_tmp_3225;
  wire or_tmp_3258;
  wire or_tmp_3262;
  wire or_tmp_3264;
  wire nor_tmp_306;
  wire nor_tmp_307;
  wire and_dcpl_258;
  wire and_dcpl_259;
  wire and_dcpl_260;
  wire and_dcpl_261;
  wire and_dcpl_262;
  wire and_dcpl_263;
  wire and_dcpl_264;
  wire and_dcpl_265;
  wire and_dcpl_268;
  wire mux_tmp_2924;
  wire or_tmp_3717;
  wire mux_tmp_2927;
  wire or_tmp_3718;
  wire and_dcpl_340;
  wire or_tmp_3721;
  wire and_dcpl_343;
  wire and_dcpl_344;
  wire and_dcpl_346;
  wire and_dcpl_347;
  wire and_dcpl_349;
  wire and_dcpl_351;
  wire and_dcpl_353;
  wire and_dcpl_354;
  wire and_dcpl_355;
  wire and_dcpl_357;
  wire and_dcpl_359;
  wire nand_tmp_142;
  wire mux_tmp_2939;
  wire or_tmp_3734;
  wire and_dcpl_365;
  wire or_dcpl_122;
  wire or_dcpl_125;
  wire mux_tmp_2953;
  wire mux_tmp_2955;
  wire mux_tmp_2956;
  wire mux_tmp_2959;
  wire mux_tmp_2960;
  wire mux_tmp_2961;
  wire mux_tmp_2965;
  wire mux_tmp_2966;
  wire mux_tmp_2968;
  wire and_dcpl_370;
  wire mux_tmp_2971;
  wire or_tmp_3744;
  wire mux_tmp_2975;
  wire or_tmp_3746;
  wire mux_tmp_2976;
  wire and_dcpl_375;
  wire or_tmp_3747;
  wire and_dcpl_377;
  wire and_dcpl_382;
  wire and_dcpl_384;
  wire mux_tmp_2993;
  wire mux_tmp_2994;
  wire or_tmp_3757;
  wire or_tmp_3760;
  wire mux_tmp_3001;
  wire mux_tmp_3003;
  wire mux_tmp_3009;
  wire mux_tmp_3012;
  wire mux_tmp_3013;
  wire mux_tmp_3016;
  wire and_dcpl_387;
  wire or_tmp_3773;
  wire and_dcpl_388;
  wire mux_tmp_3042;
  wire and_tmp_31;
  wire mux_tmp_3049;
  wire and_dcpl_390;
  wire and_dcpl_392;
  wire and_dcpl_396;
  wire and_dcpl_399;
  wire and_dcpl_402;
  wire mux_tmp_3069;
  wire mux_tmp_3070;
  wire mux_tmp_3078;
  wire and_dcpl_403;
  wire and_dcpl_404;
  wire and_dcpl_406;
  wire and_dcpl_407;
  wire mux_tmp_3098;
  wire mux_tmp_3100;
  wire mux_tmp_3101;
  wire mux_tmp_3102;
  wire and_dcpl_410;
  wire and_dcpl_411;
  wire mux_tmp_3119;
  wire not_tmp_811;
  wire mux_tmp_3133;
  wire or_tmp_3801;
  wire and_tmp_33;
  wire and_dcpl_421;
  wire mux_tmp_3169;
  wire mux_tmp_3193;
  wire mux_tmp_3196;
  wire and_tmp_35;
  wire mux_tmp_3210;
  wire and_tmp_36;
  wire mux_tmp_3213;
  wire mux_tmp_3214;
  wire mux_tmp_3218;
  wire or_dcpl_134;
  wire and_dcpl_432;
  wire or_tmp_3833;
  wire nor_tmp_391;
  wire mux_tmp_3280;
  wire not_tmp_868;
  wire or_dcpl_150;
  wire mux_tmp_3288;
  reg COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  wire [8:0] COMP_LOOP_acc_14_psp_sva_1;
  wire [9:0] nl_COMP_LOOP_acc_14_psp_sva_1;
  reg [9:0] VEC_LOOP_j_10_0_sva_9_0;
  reg [6:0] COMP_LOOP_k_10_3_sva_6_0;
  reg COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_nor_315_itm;
  reg COMP_LOOP_nor_289_itm;
  reg COMP_LOOP_nor_313_itm;
  reg COMP_LOOP_nor_326_itm;
  reg COMP_LOOP_nor_319_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  reg COMP_LOOP_nor_521_itm;
  reg COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_nor_767_itm;
  reg COMP_LOOP_nor_760_itm;
  reg COMP_LOOP_nor_734_itm;
  reg COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_nor_970_itm;
  reg COMP_LOOP_nor_969_itm;
  reg COMP_LOOP_nor_984_itm;
  reg COMP_LOOP_nor_964_itm;
  reg COMP_LOOP_nor_961_itm;
  reg COMP_LOOP_nor_955_itm;
  reg COMP_LOOP_nor_962_itm;
  reg COMP_LOOP_nor_957_itm;
  reg COMP_LOOP_nor_976_itm;
  reg COMP_LOOP_nor_958_itm;
  reg COMP_LOOP_nor_998_itm;
  reg COMP_LOOP_nor_972_itm;
  reg COMP_LOOP_nor_987_itm;
  reg COMP_LOOP_nor_985_itm;
  reg COMP_LOOP_nor_991_itm;
  reg COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_nor_1185_itm;
  reg COMP_LOOP_nor_1211_itm;
  reg COMP_LOOP_nor_1209_itm;
  reg COMP_LOOP_nor_1196_itm;
  reg COMP_LOOP_nor_1208_itm;
  reg COMP_LOOP_nor_1186_itm;
  reg COMP_LOOP_nor_1182_itm;
  reg COMP_LOOP_nor_1222_itm;
  reg COMP_LOOP_nor_1188_itm;
  reg COMP_LOOP_nor_1215_itm;
  reg COMP_LOOP_nor_1194_itm;
  reg COMP_LOOP_nor_1193_itm;
  reg COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  reg COMP_LOOP_nor_1435_itm;
  reg COMP_LOOP_nor_1446_itm;
  reg COMP_LOOP_nor_1439_itm;
  reg COMP_LOOP_nor_1420_itm;
  reg COMP_LOOP_nor_1432_itm;
  reg COMP_LOOP_nor_1424_itm;
  reg COMP_LOOP_nor_1410_itm;
  reg COMP_LOOP_nor_1403_itm;
  reg COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  reg COMP_LOOP_nor_1663_itm;
  reg COMP_LOOP_nor_1659_itm;
  reg COMP_LOOP_nor_1633_itm;
  reg COMP_LOOP_nor_1642_itm;
  reg COMP_LOOP_nor_1648_itm;
  reg COMP_LOOP_nor_1630_itm;
  reg COMP_LOOP_nor_1670_itm;
  reg COMP_LOOP_nor_1629_itm;
  reg [9:0] COMP_LOOP_2_tmp_mul_idiv_sva;
  reg [9:0] COMP_LOOP_2_tmp_lshift_ncse_sva;
  reg COMP_LOOP_tmp_nor_10_itm;
  reg [8:0] COMP_LOOP_3_tmp_lshift_ncse_sva;
  reg COMP_LOOP_tmp_nor_206_itm;
  reg COMP_LOOP_tmp_nor_151_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm;
  reg COMP_LOOP_COMP_LOOP_and_119_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm;
  reg COMP_LOOP_COMP_LOOP_and_109_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm;
  reg COMP_LOOP_COMP_LOOP_and_1106_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm;
  reg COMP_LOOP_COMP_LOOP_and_102_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm;
  reg COMP_LOOP_COMP_LOOP_and_117_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm;
  reg COMP_LOOP_COMP_LOOP_and_1370_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm;
  reg COMP_LOOP_COMP_LOOP_and_122_itm;
  reg [9:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_4_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_2_sva;
  reg [9:0] COMP_LOOP_acc_1_cse_6_sva;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_6_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_6_sva;
  reg [8:0] COMP_LOOP_acc_11_psp_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_3_sva;
  reg [8:0] COMP_LOOP_acc_14_psp_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_7_sva;
  reg [6:0] COMP_LOOP_acc_psp_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_1_sva;
  reg [7:0] COMP_LOOP_acc_13_psp_sva;
  wire [8:0] nl_COMP_LOOP_acc_13_psp_sva;
  reg [9:0] COMP_LOOP_acc_10_cse_10_1_5_sva;
  reg [7:0] COMP_LOOP_5_tmp_mul_idiv_sva;
  reg [10:0] STAGE_LOOP_lshift_psp_sva;
  wire [9:0] COMP_LOOP_acc_1_cse_4_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_4_sva_1;
  wire [9:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [10:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire [6:0] COMP_LOOP_acc_psp_sva_mx0w0;
  wire [7:0] nl_COMP_LOOP_acc_psp_sva_mx0w0;
  wire [8:0] COMP_LOOP_acc_11_psp_sva_1;
  wire [9:0] nl_COMP_LOOP_acc_11_psp_sva_1;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt;
  wire mux_3360_tmp;
  wire and_478_m1c;
  wire nor_tmp_396;
  wire and_476_tmp;
  wire nor_1579_tmp;
  wire and_474_tmp;
  reg [6:0] reg_COMP_LOOP_k_10_3_ftd;
  wire nand_191_cse;
  wire nand_190_cse;
  wire nand_188_cse;
  wire nand_174_cse;
  wire nand_175_cse;
  wire nand_184_cse;
  reg reg_vec_rsc_triosy_0_63_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire or_595_cse;
  wire and_507_cse;
  wire or_341_cse;
  wire or_359_cse;
  wire mux_297_cse;
  wire or_4057_cse;
  wire and_677_cse;
  wire nor_358_cse;
  wire nor_412_cse;
  wire and_493_cse;
  wire and_640_cse;
  wire or_564_cse;
  wire COMP_LOOP_tmp_or_cse;
  wire COMP_LOOP_tmp_or_5_cse;
  wire COMP_LOOP_tmp_or_36_cse;
  wire COMP_LOOP_tmp_or_43_cse;
  wire nor_399_cse;
  wire or_4007_cse;
  wire or_80_cse;
  wire and_705_cse;
  wire nor_1683_cse;
  wire and_673_cse;
  wire and_639_cse;
  wire and_735_cse;
  wire or_364_cse;
  wire and_763_cse;
  wire or_477_cse;
  wire nor_1674_cse;
  wire and_808_cse;
  wire or_150_cse;
  wire nor_398_cse;
  wire mux_742_cse;
  wire and_779_cse;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm;
  wire and_655_cse;
  wire or_4050_cse;
  wire and_78_cse;
  wire mux_180_cse;
  wire mux_221_cse;
  wire and_736_cse;
  wire mux_3095_cse;
  wire mux_2997_rmff;
  reg [63:0] COMP_LOOP_1_acc_8_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_1_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_2_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_3_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_4_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_5_itm;
  reg [63:0] COMP_LOOP_tmp_mux1h_6_itm;
  reg [63:0] tmp_21_sva_1;
  reg [63:0] p_sva;
  wire mux_3025_itm;
  wire mux_3058_itm;
  wire mux_3114_itm;
  wire mux_3175_itm;
  wire mux_3185_itm;
  wire mux_3187_itm;
  wire mux_3201_itm;
  wire mux_3305_itm;
  wire [10:0] z_out;
  wire [9:0] z_out_1;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  wire and_dcpl_477;
  wire and_dcpl_488;
  wire [10:0] z_out_3;
  wire and_dcpl_501;
  wire [3:0] z_out_4;
  wire [4:0] nl_z_out_4;
  wire and_dcpl_503;
  wire and_dcpl_509;
  wire and_dcpl_513;
  wire and_dcpl_514;
  wire and_dcpl_519;
  wire and_dcpl_526;
  wire and_dcpl_570;
  wire and_dcpl_573;
  wire and_dcpl_574;
  wire and_dcpl_576;
  wire and_dcpl_577;
  wire and_dcpl_579;
  wire and_dcpl_580;
  wire and_dcpl_582;
  wire and_dcpl_583;
  wire and_dcpl_588;
  wire and_dcpl_589;
  wire and_dcpl_590;
  wire [9:0] z_out_7;
  wire [19:0] nl_z_out_7;
  wire and_dcpl_599;
  wire and_dcpl_602;
  wire and_dcpl_605;
  wire and_dcpl_608;
  wire and_dcpl_611;
  wire and_dcpl_612;
  wire and_dcpl_614;
  wire and_dcpl_615;
  wire and_dcpl_617;
  wire and_dcpl_618;
  wire and_dcpl_619;
  wire and_dcpl_620;
  wire and_dcpl_623;
  wire and_dcpl_625;
  wire [63:0] z_out_8;
  wire [127:0] nl_z_out_8;
  wire and_dcpl_632;
  wire and_dcpl_636;
  wire [63:0] z_out_9;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [3:0] COMP_LOOP_1_tmp_acc_cse_sva;
  reg [63:0] tmp_21_sva_2;
  reg [63:0] tmp_21_sva_3;
  reg [63:0] tmp_21_sva_5;
  reg [63:0] tmp_21_sva_6;
  reg [63:0] tmp_21_sva_7;
  reg [63:0] tmp_21_sva_9;
  reg [63:0] tmp_21_sva_11;
  reg [63:0] tmp_21_sva_13;
  reg [63:0] tmp_21_sva_14;
  reg [63:0] tmp_21_sva_15;
  reg [63:0] tmp_21_sva_17;
  reg [63:0] tmp_21_sva_18;
  reg [63:0] tmp_21_sva_19;
  reg [63:0] tmp_21_sva_21;
  reg [63:0] tmp_21_sva_22;
  reg [63:0] tmp_21_sva_23;
  reg [63:0] tmp_21_sva_25;
  reg [63:0] tmp_21_sva_26;
  reg [63:0] tmp_21_sva_27;
  reg [63:0] tmp_21_sva_29;
  reg [63:0] tmp_21_sva_30;
  reg [63:0] tmp_21_sva_31;
  reg [63:0] tmp_21_sva_33;
  reg [63:0] tmp_21_sva_34;
  reg [63:0] tmp_21_sva_35;
  reg [63:0] tmp_21_sva_37;
  reg [63:0] tmp_21_sva_38;
  reg [63:0] tmp_21_sva_39;
  reg [63:0] tmp_21_sva_41;
  reg [63:0] tmp_21_sva_42;
  reg [63:0] tmp_21_sva_43;
  reg [63:0] tmp_21_sva_45;
  reg [63:0] tmp_21_sva_46;
  reg [63:0] tmp_21_sva_47;
  reg [63:0] tmp_21_sva_49;
  reg [63:0] tmp_21_sva_50;
  reg [63:0] tmp_21_sva_51;
  reg [63:0] tmp_21_sva_53;
  reg [63:0] tmp_21_sva_54;
  reg [63:0] tmp_21_sva_55;
  reg [63:0] tmp_21_sva_57;
  reg [63:0] tmp_21_sva_58;
  reg [63:0] tmp_21_sva_59;
  reg [63:0] tmp_21_sva_61;
  reg [63:0] tmp_21_sva_62;
  reg [63:0] tmp_21_sva_63;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg COMP_LOOP_COMP_LOOP_and_18_itm;
  reg COMP_LOOP_COMP_LOOP_and_20_itm;
  reg COMP_LOOP_COMP_LOOP_and_21_itm;
  reg COMP_LOOP_COMP_LOOP_and_22_itm;
  reg COMP_LOOP_COMP_LOOP_and_23_itm;
  reg COMP_LOOP_COMP_LOOP_and_24_itm;
  reg COMP_LOOP_COMP_LOOP_and_25_itm;
  reg COMP_LOOP_COMP_LOOP_and_26_itm;
  reg COMP_LOOP_COMP_LOOP_and_27_itm;
  reg COMP_LOOP_COMP_LOOP_and_28_itm;
  reg COMP_LOOP_COMP_LOOP_and_29_itm;
  reg COMP_LOOP_COMP_LOOP_and_30_itm;
  reg COMP_LOOP_COMP_LOOP_and_34_itm;
  reg COMP_LOOP_COMP_LOOP_and_36_itm;
  reg COMP_LOOP_COMP_LOOP_and_37_itm;
  reg COMP_LOOP_COMP_LOOP_and_38_itm;
  reg COMP_LOOP_COMP_LOOP_and_39_itm;
  reg COMP_LOOP_COMP_LOOP_and_40_itm;
  reg COMP_LOOP_COMP_LOOP_and_41_itm;
  reg COMP_LOOP_COMP_LOOP_and_42_itm;
  reg COMP_LOOP_COMP_LOOP_and_43_itm;
  reg COMP_LOOP_COMP_LOOP_and_44_itm;
  reg COMP_LOOP_COMP_LOOP_and_45_itm;
  reg COMP_LOOP_COMP_LOOP_and_46_itm;
  reg COMP_LOOP_COMP_LOOP_and_47_itm;
  reg COMP_LOOP_COMP_LOOP_and_48_itm;
  reg COMP_LOOP_COMP_LOOP_and_49_itm;
  reg COMP_LOOP_COMP_LOOP_and_50_itm;
  reg COMP_LOOP_COMP_LOOP_and_51_itm;
  reg COMP_LOOP_COMP_LOOP_and_52_itm;
  reg COMP_LOOP_COMP_LOOP_and_53_itm;
  reg COMP_LOOP_COMP_LOOP_and_54_itm;
  reg COMP_LOOP_COMP_LOOP_and_55_itm;
  reg COMP_LOOP_COMP_LOOP_and_56_itm;
  reg COMP_LOOP_COMP_LOOP_and_57_itm;
  reg COMP_LOOP_COMP_LOOP_and_58_itm;
  reg COMP_LOOP_COMP_LOOP_and_59_itm;
  reg COMP_LOOP_COMP_LOOP_and_60_itm;
  reg COMP_LOOP_COMP_LOOP_and_61_itm;
  reg COMP_LOOP_COMP_LOOP_and_62_itm;
  reg COMP_LOOP_COMP_LOOP_and_73_itm;
  reg COMP_LOOP_COMP_LOOP_and_74_itm;
  reg COMP_LOOP_COMP_LOOP_and_75_itm;
  reg COMP_LOOP_COMP_LOOP_and_100_itm;
  reg COMP_LOOP_COMP_LOOP_and_101_itm;
  reg COMP_LOOP_COMP_LOOP_and_103_itm;
  reg COMP_LOOP_COMP_LOOP_and_104_itm;
  reg COMP_LOOP_COMP_LOOP_and_105_itm;
  reg COMP_LOOP_COMP_LOOP_and_106_itm;
  reg COMP_LOOP_COMP_LOOP_and_107_itm;
  reg COMP_LOOP_COMP_LOOP_and_108_itm;
  reg COMP_LOOP_COMP_LOOP_and_110_itm;
  reg COMP_LOOP_COMP_LOOP_and_115_itm;
  reg COMP_LOOP_COMP_LOOP_and_116_itm;
  reg COMP_LOOP_COMP_LOOP_and_118_itm;
  reg COMP_LOOP_COMP_LOOP_and_120_itm;
  reg COMP_LOOP_COMP_LOOP_and_121_itm;
  reg COMP_LOOP_COMP_LOOP_and_123_itm;
  reg COMP_LOOP_COMP_LOOP_and_124_itm;
  reg COMP_LOOP_COMP_LOOP_and_125_itm;
  reg COMP_LOOP_COMP_LOOP_and_258_itm;
  reg COMP_LOOP_COMP_LOOP_and_260_itm;
  reg COMP_LOOP_COMP_LOOP_and_261_itm;
  reg COMP_LOOP_COMP_LOOP_and_262_itm;
  reg COMP_LOOP_COMP_LOOP_and_264_itm;
  reg COMP_LOOP_COMP_LOOP_and_268_itm;
  reg COMP_LOOP_COMP_LOOP_and_270_itm;
  reg COMP_LOOP_COMP_LOOP_and_272_itm;
  reg COMP_LOOP_COMP_LOOP_and_284_itm;
  reg COMP_LOOP_COMP_LOOP_and_285_itm;
  reg COMP_LOOP_COMP_LOOP_and_286_itm;
  reg COMP_LOOP_COMP_LOOP_and_288_itm;
  reg COMP_LOOP_COMP_LOOP_nor_5_itm;
  reg COMP_LOOP_nor_281_itm;
  reg COMP_LOOP_nor_282_itm;
  reg COMP_LOOP_nor_284_itm;
  reg COMP_LOOP_nor_288_itm;
  reg COMP_LOOP_nor_296_itm;
  reg COMP_LOOP_COMP_LOOP_and_333_itm;
  reg COMP_LOOP_COMP_LOOP_and_334_itm;
  reg COMP_LOOP_COMP_LOOP_and_335_itm;
  reg COMP_LOOP_COMP_LOOP_and_336_itm;
  reg COMP_LOOP_COMP_LOOP_and_337_itm;
  reg COMP_LOOP_COMP_LOOP_and_338_itm;
  reg COMP_LOOP_COMP_LOOP_and_339_itm;
  reg COMP_LOOP_COMP_LOOP_and_340_itm;
  reg COMP_LOOP_COMP_LOOP_and_341_itm;
  reg COMP_LOOP_COMP_LOOP_and_342_itm;
  reg COMP_LOOP_COMP_LOOP_and_343_itm;
  reg COMP_LOOP_COMP_LOOP_and_344_itm;
  reg COMP_LOOP_COMP_LOOP_and_345_itm;
  reg COMP_LOOP_nor_311_itm;
  reg COMP_LOOP_COMP_LOOP_and_347_itm;
  reg COMP_LOOP_COMP_LOOP_and_349_itm;
  reg COMP_LOOP_COMP_LOOP_and_351_itm;
  reg COMP_LOOP_COMP_LOOP_and_352_itm;
  reg COMP_LOOP_COMP_LOOP_and_353_itm;
  reg COMP_LOOP_COMP_LOOP_and_355_itm;
  reg COMP_LOOP_COMP_LOOP_and_356_itm;
  reg COMP_LOOP_COMP_LOOP_and_357_itm;
  reg COMP_LOOP_COMP_LOOP_and_358_itm;
  reg COMP_LOOP_COMP_LOOP_and_359_itm;
  reg COMP_LOOP_COMP_LOOP_and_360_itm;
  reg COMP_LOOP_COMP_LOOP_and_361_itm;
  reg COMP_LOOP_COMP_LOOP_and_363_itm;
  reg COMP_LOOP_COMP_LOOP_and_364_itm;
  reg COMP_LOOP_COMP_LOOP_and_365_itm;
  reg COMP_LOOP_COMP_LOOP_and_366_itm;
  reg COMP_LOOP_COMP_LOOP_and_367_itm;
  reg COMP_LOOP_COMP_LOOP_and_368_itm;
  reg COMP_LOOP_COMP_LOOP_and_369_itm;
  reg COMP_LOOP_COMP_LOOP_and_370_itm;
  reg COMP_LOOP_COMP_LOOP_and_371_itm;
  reg COMP_LOOP_COMP_LOOP_and_372_itm;
  reg COMP_LOOP_COMP_LOOP_and_373_itm;
  reg COMP_LOOP_COMP_LOOP_and_374_itm;
  reg COMP_LOOP_COMP_LOOP_and_375_itm;
  reg COMP_LOOP_COMP_LOOP_and_376_itm;
  reg COMP_LOOP_COMP_LOOP_and_377_itm;
  reg COMP_LOOP_COMP_LOOP_and_509_itm;
  reg COMP_LOOP_COMP_LOOP_and_510_itm;
  reg COMP_LOOP_COMP_LOOP_and_522_itm;
  reg COMP_LOOP_COMP_LOOP_nor_9_itm;
  reg COMP_LOOP_nor_505_itm;
  reg COMP_LOOP_nor_506_itm;
  reg COMP_LOOP_COMP_LOOP_and_569_itm;
  reg COMP_LOOP_nor_508_itm;
  reg COMP_LOOP_COMP_LOOP_and_571_itm;
  reg COMP_LOOP_COMP_LOOP_and_572_itm;
  reg COMP_LOOP_COMP_LOOP_and_573_itm;
  reg COMP_LOOP_nor_512_itm;
  reg COMP_LOOP_COMP_LOOP_and_575_itm;
  reg COMP_LOOP_COMP_LOOP_and_576_itm;
  reg COMP_LOOP_COMP_LOOP_and_577_itm;
  reg COMP_LOOP_COMP_LOOP_and_578_itm;
  reg COMP_LOOP_COMP_LOOP_and_579_itm;
  reg COMP_LOOP_COMP_LOOP_and_580_itm;
  reg COMP_LOOP_COMP_LOOP_and_581_itm;
  reg COMP_LOOP_nor_520_itm;
  reg COMP_LOOP_COMP_LOOP_and_583_itm;
  reg COMP_LOOP_COMP_LOOP_and_584_itm;
  reg COMP_LOOP_COMP_LOOP_and_585_itm;
  reg COMP_LOOP_COMP_LOOP_and_586_itm;
  reg COMP_LOOP_COMP_LOOP_and_587_itm;
  reg COMP_LOOP_COMP_LOOP_and_588_itm;
  reg COMP_LOOP_COMP_LOOP_and_589_itm;
  reg COMP_LOOP_COMP_LOOP_and_590_itm;
  reg COMP_LOOP_COMP_LOOP_and_591_itm;
  reg COMP_LOOP_COMP_LOOP_and_592_itm;
  reg COMP_LOOP_COMP_LOOP_and_593_itm;
  reg COMP_LOOP_COMP_LOOP_and_594_itm;
  reg COMP_LOOP_COMP_LOOP_and_595_itm;
  reg COMP_LOOP_COMP_LOOP_and_596_itm;
  reg COMP_LOOP_COMP_LOOP_and_597_itm;
  reg COMP_LOOP_nor_535_itm;
  reg COMP_LOOP_COMP_LOOP_and_599_itm;
  reg COMP_LOOP_COMP_LOOP_and_600_itm;
  reg COMP_LOOP_COMP_LOOP_and_601_itm;
  reg COMP_LOOP_COMP_LOOP_and_602_itm;
  reg COMP_LOOP_COMP_LOOP_and_603_itm;
  reg COMP_LOOP_COMP_LOOP_and_604_itm;
  reg COMP_LOOP_COMP_LOOP_and_605_itm;
  reg COMP_LOOP_COMP_LOOP_and_606_itm;
  reg COMP_LOOP_COMP_LOOP_and_607_itm;
  reg COMP_LOOP_COMP_LOOP_and_608_itm;
  reg COMP_LOOP_COMP_LOOP_and_609_itm;
  reg COMP_LOOP_COMP_LOOP_and_610_itm;
  reg COMP_LOOP_COMP_LOOP_and_611_itm;
  reg COMP_LOOP_COMP_LOOP_and_612_itm;
  reg COMP_LOOP_COMP_LOOP_and_613_itm;
  reg COMP_LOOP_COMP_LOOP_and_614_itm;
  reg COMP_LOOP_COMP_LOOP_and_615_itm;
  reg COMP_LOOP_COMP_LOOP_and_616_itm;
  reg COMP_LOOP_COMP_LOOP_and_617_itm;
  reg COMP_LOOP_COMP_LOOP_and_618_itm;
  reg COMP_LOOP_COMP_LOOP_and_619_itm;
  reg COMP_LOOP_COMP_LOOP_and_620_itm;
  reg COMP_LOOP_COMP_LOOP_and_621_itm;
  reg COMP_LOOP_COMP_LOOP_and_622_itm;
  reg COMP_LOOP_COMP_LOOP_and_623_itm;
  reg COMP_LOOP_COMP_LOOP_and_624_itm;
  reg COMP_LOOP_COMP_LOOP_and_625_itm;
  reg COMP_LOOP_COMP_LOOP_and_626_itm;
  reg COMP_LOOP_COMP_LOOP_and_627_itm;
  reg COMP_LOOP_COMP_LOOP_and_628_itm;
  reg COMP_LOOP_COMP_LOOP_and_629_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm;
  reg COMP_LOOP_COMP_LOOP_and_760_itm;
  reg COMP_LOOP_COMP_LOOP_and_761_itm;
  reg COMP_LOOP_COMP_LOOP_nor_13_itm;
  reg COMP_LOOP_nor_729_itm;
  reg COMP_LOOP_nor_730_itm;
  reg COMP_LOOP_COMP_LOOP_and_821_itm;
  reg COMP_LOOP_nor_732_itm;
  reg COMP_LOOP_COMP_LOOP_and_823_itm;
  reg COMP_LOOP_COMP_LOOP_and_825_itm;
  reg COMP_LOOP_nor_736_itm;
  reg COMP_LOOP_COMP_LOOP_and_827_itm;
  reg COMP_LOOP_COMP_LOOP_and_828_itm;
  reg COMP_LOOP_COMP_LOOP_and_829_itm;
  reg COMP_LOOP_COMP_LOOP_and_830_itm;
  reg COMP_LOOP_COMP_LOOP_and_831_itm;
  reg COMP_LOOP_COMP_LOOP_and_832_itm;
  reg COMP_LOOP_COMP_LOOP_and_833_itm;
  reg COMP_LOOP_nor_744_itm;
  reg COMP_LOOP_COMP_LOOP_and_835_itm;
  reg COMP_LOOP_COMP_LOOP_and_836_itm;
  reg COMP_LOOP_COMP_LOOP_and_837_itm;
  reg COMP_LOOP_COMP_LOOP_and_838_itm;
  reg COMP_LOOP_COMP_LOOP_and_839_itm;
  reg COMP_LOOP_COMP_LOOP_and_840_itm;
  reg COMP_LOOP_COMP_LOOP_and_841_itm;
  reg COMP_LOOP_COMP_LOOP_and_842_itm;
  reg COMP_LOOP_COMP_LOOP_and_843_itm;
  reg COMP_LOOP_COMP_LOOP_and_844_itm;
  reg COMP_LOOP_COMP_LOOP_and_845_itm;
  reg COMP_LOOP_COMP_LOOP_and_846_itm;
  reg COMP_LOOP_COMP_LOOP_and_847_itm;
  reg COMP_LOOP_COMP_LOOP_and_848_itm;
  reg COMP_LOOP_COMP_LOOP_and_849_itm;
  reg COMP_LOOP_nor_759_itm;
  reg COMP_LOOP_COMP_LOOP_and_852_itm;
  reg COMP_LOOP_COMP_LOOP_and_853_itm;
  reg COMP_LOOP_COMP_LOOP_and_854_itm;
  reg COMP_LOOP_COMP_LOOP_and_855_itm;
  reg COMP_LOOP_COMP_LOOP_and_856_itm;
  reg COMP_LOOP_COMP_LOOP_and_857_itm;
  reg COMP_LOOP_COMP_LOOP_and_859_itm;
  reg COMP_LOOP_COMP_LOOP_and_860_itm;
  reg COMP_LOOP_COMP_LOOP_and_861_itm;
  reg COMP_LOOP_COMP_LOOP_and_862_itm;
  reg COMP_LOOP_COMP_LOOP_and_863_itm;
  reg COMP_LOOP_COMP_LOOP_and_864_itm;
  reg COMP_LOOP_COMP_LOOP_and_865_itm;
  reg COMP_LOOP_COMP_LOOP_and_866_itm;
  reg COMP_LOOP_COMP_LOOP_and_867_itm;
  reg COMP_LOOP_COMP_LOOP_and_868_itm;
  reg COMP_LOOP_COMP_LOOP_and_869_itm;
  reg COMP_LOOP_COMP_LOOP_and_870_itm;
  reg COMP_LOOP_COMP_LOOP_and_871_itm;
  reg COMP_LOOP_COMP_LOOP_and_872_itm;
  reg COMP_LOOP_COMP_LOOP_and_873_itm;
  reg COMP_LOOP_COMP_LOOP_and_874_itm;
  reg COMP_LOOP_COMP_LOOP_and_875_itm;
  reg COMP_LOOP_COMP_LOOP_and_876_itm;
  reg COMP_LOOP_COMP_LOOP_and_877_itm;
  reg COMP_LOOP_COMP_LOOP_and_878_itm;
  reg COMP_LOOP_COMP_LOOP_and_879_itm;
  reg COMP_LOOP_COMP_LOOP_and_880_itm;
  reg COMP_LOOP_COMP_LOOP_and_881_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm;
  reg COMP_LOOP_COMP_LOOP_nor_17_itm;
  reg COMP_LOOP_nor_953_itm;
  reg COMP_LOOP_nor_954_itm;
  reg COMP_LOOP_nor_956_itm;
  reg COMP_LOOP_COMP_LOOP_and_1077_itm;
  reg COMP_LOOP_nor_960_itm;
  reg COMP_LOOP_COMP_LOOP_and_1081_itm;
  reg COMP_LOOP_COMP_LOOP_and_1083_itm;
  reg COMP_LOOP_COMP_LOOP_and_1084_itm;
  reg COMP_LOOP_COMP_LOOP_and_1085_itm;
  reg COMP_LOOP_nor_968_itm;
  reg COMP_LOOP_COMP_LOOP_and_1089_itm;
  reg COMP_LOOP_COMP_LOOP_and_1091_itm;
  reg COMP_LOOP_COMP_LOOP_and_1092_itm;
  reg COMP_LOOP_COMP_LOOP_and_1093_itm;
  reg COMP_LOOP_COMP_LOOP_and_1095_itm;
  reg COMP_LOOP_COMP_LOOP_and_1096_itm;
  reg COMP_LOOP_COMP_LOOP_and_1097_itm;
  reg COMP_LOOP_COMP_LOOP_and_1098_itm;
  reg COMP_LOOP_COMP_LOOP_and_1099_itm;
  reg COMP_LOOP_COMP_LOOP_and_1100_itm;
  reg COMP_LOOP_COMP_LOOP_and_1101_itm;
  reg COMP_LOOP_nor_983_itm;
  reg COMP_LOOP_COMP_LOOP_and_1104_itm;
  reg COMP_LOOP_COMP_LOOP_and_1105_itm;
  reg COMP_LOOP_COMP_LOOP_and_1107_itm;
  reg COMP_LOOP_COMP_LOOP_and_1108_itm;
  reg COMP_LOOP_COMP_LOOP_and_1109_itm;
  reg COMP_LOOP_COMP_LOOP_and_1110_itm;
  reg COMP_LOOP_COMP_LOOP_and_1111_itm;
  reg COMP_LOOP_COMP_LOOP_and_1112_itm;
  reg COMP_LOOP_COMP_LOOP_and_1113_itm;
  reg COMP_LOOP_COMP_LOOP_and_1114_itm;
  reg COMP_LOOP_COMP_LOOP_and_1115_itm;
  reg COMP_LOOP_COMP_LOOP_and_1116_itm;
  reg COMP_LOOP_COMP_LOOP_and_1117_itm;
  reg COMP_LOOP_COMP_LOOP_and_1118_itm;
  reg COMP_LOOP_COMP_LOOP_and_1119_itm;
  reg COMP_LOOP_COMP_LOOP_and_1120_itm;
  reg COMP_LOOP_COMP_LOOP_and_1121_itm;
  reg COMP_LOOP_COMP_LOOP_and_1122_itm;
  reg COMP_LOOP_COMP_LOOP_and_1123_itm;
  reg COMP_LOOP_COMP_LOOP_and_1124_itm;
  reg COMP_LOOP_COMP_LOOP_and_1125_itm;
  reg COMP_LOOP_COMP_LOOP_and_1126_itm;
  reg COMP_LOOP_COMP_LOOP_and_1127_itm;
  reg COMP_LOOP_COMP_LOOP_and_1128_itm;
  reg COMP_LOOP_COMP_LOOP_and_1129_itm;
  reg COMP_LOOP_COMP_LOOP_and_1130_itm;
  reg COMP_LOOP_COMP_LOOP_and_1131_itm;
  reg COMP_LOOP_COMP_LOOP_and_1132_itm;
  reg COMP_LOOP_COMP_LOOP_and_1133_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm;
  reg COMP_LOOP_tmp_nor_140_itm;
  reg COMP_LOOP_tmp_nor_141_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm;
  reg COMP_LOOP_tmp_nor_143_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm;
  reg COMP_LOOP_tmp_nor_146_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm;
  reg COMP_LOOP_COMP_LOOP_nor_21_itm;
  reg COMP_LOOP_nor_1177_itm;
  reg COMP_LOOP_nor_1178_itm;
  reg COMP_LOOP_COMP_LOOP_and_1325_itm;
  reg COMP_LOOP_nor_1180_itm;
  reg COMP_LOOP_COMP_LOOP_and_1327_itm;
  reg COMP_LOOP_COMP_LOOP_and_1329_itm;
  reg COMP_LOOP_nor_1184_itm;
  reg COMP_LOOP_COMP_LOOP_and_1333_itm;
  reg COMP_LOOP_COMP_LOOP_and_1335_itm;
  reg COMP_LOOP_COMP_LOOP_and_1336_itm;
  reg COMP_LOOP_COMP_LOOP_and_1337_itm;
  reg COMP_LOOP_nor_1192_itm;
  reg COMP_LOOP_COMP_LOOP_and_1341_itm;
  reg COMP_LOOP_COMP_LOOP_and_1343_itm;
  reg COMP_LOOP_COMP_LOOP_and_1344_itm;
  reg COMP_LOOP_COMP_LOOP_and_1345_itm;
  reg COMP_LOOP_COMP_LOOP_and_1346_itm;
  reg COMP_LOOP_COMP_LOOP_and_1347_itm;
  reg COMP_LOOP_COMP_LOOP_and_1348_itm;
  reg COMP_LOOP_COMP_LOOP_and_1349_itm;
  reg COMP_LOOP_COMP_LOOP_and_1350_itm;
  reg COMP_LOOP_COMP_LOOP_and_1351_itm;
  reg COMP_LOOP_COMP_LOOP_and_1352_itm;
  reg COMP_LOOP_COMP_LOOP_and_1353_itm;
  reg COMP_LOOP_nor_1207_itm;
  reg COMP_LOOP_COMP_LOOP_and_1357_itm;
  reg COMP_LOOP_COMP_LOOP_and_1359_itm;
  reg COMP_LOOP_COMP_LOOP_and_1360_itm;
  reg COMP_LOOP_COMP_LOOP_and_1361_itm;
  reg COMP_LOOP_COMP_LOOP_and_1363_itm;
  reg COMP_LOOP_COMP_LOOP_and_1364_itm;
  reg COMP_LOOP_COMP_LOOP_and_1365_itm;
  reg COMP_LOOP_COMP_LOOP_and_1366_itm;
  reg COMP_LOOP_COMP_LOOP_and_1367_itm;
  reg COMP_LOOP_COMP_LOOP_and_1368_itm;
  reg COMP_LOOP_COMP_LOOP_and_1369_itm;
  reg COMP_LOOP_COMP_LOOP_and_1371_itm;
  reg COMP_LOOP_COMP_LOOP_and_1372_itm;
  reg COMP_LOOP_COMP_LOOP_and_1373_itm;
  reg COMP_LOOP_COMP_LOOP_and_1374_itm;
  reg COMP_LOOP_COMP_LOOP_and_1375_itm;
  reg COMP_LOOP_COMP_LOOP_and_1376_itm;
  reg COMP_LOOP_COMP_LOOP_and_1377_itm;
  reg COMP_LOOP_COMP_LOOP_and_1378_itm;
  reg COMP_LOOP_COMP_LOOP_and_1379_itm;
  reg COMP_LOOP_COMP_LOOP_and_1380_itm;
  reg COMP_LOOP_COMP_LOOP_and_1381_itm;
  reg COMP_LOOP_COMP_LOOP_and_1382_itm;
  reg COMP_LOOP_COMP_LOOP_and_1383_itm;
  reg COMP_LOOP_COMP_LOOP_and_1384_itm;
  reg COMP_LOOP_COMP_LOOP_and_1385_itm;
  reg COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm;
  reg COMP_LOOP_tmp_nor_153_itm;
  reg COMP_LOOP_tmp_nor_157_itm;
  reg COMP_LOOP_tmp_nor_165_itm;
  reg COMP_LOOP_tmp_nor_180_itm;
  reg COMP_LOOP_COMP_LOOP_and_1518_itm;
  reg COMP_LOOP_COMP_LOOP_nor_25_itm;
  reg COMP_LOOP_nor_1401_itm;
  reg COMP_LOOP_nor_1402_itm;
  reg COMP_LOOP_COMP_LOOP_and_1577_itm;
  reg COMP_LOOP_nor_1404_itm;
  reg COMP_LOOP_COMP_LOOP_and_1579_itm;
  reg COMP_LOOP_COMP_LOOP_and_1580_itm;
  reg COMP_LOOP_COMP_LOOP_and_1581_itm;
  reg COMP_LOOP_nor_1408_itm;
  reg COMP_LOOP_COMP_LOOP_and_1583_itm;
  reg COMP_LOOP_COMP_LOOP_and_1584_itm;
  reg COMP_LOOP_COMP_LOOP_and_1585_itm;
  reg COMP_LOOP_COMP_LOOP_and_1586_itm;
  reg COMP_LOOP_COMP_LOOP_and_1587_itm;
  reg COMP_LOOP_COMP_LOOP_and_1588_itm;
  reg COMP_LOOP_COMP_LOOP_and_1589_itm;
  reg COMP_LOOP_nor_1416_itm;
  reg COMP_LOOP_COMP_LOOP_and_1591_itm;
  reg COMP_LOOP_COMP_LOOP_and_1592_itm;
  reg COMP_LOOP_COMP_LOOP_and_1593_itm;
  reg COMP_LOOP_COMP_LOOP_and_1594_itm;
  reg COMP_LOOP_COMP_LOOP_and_1595_itm;
  reg COMP_LOOP_COMP_LOOP_and_1596_itm;
  reg COMP_LOOP_COMP_LOOP_and_1597_itm;
  reg COMP_LOOP_COMP_LOOP_and_1598_itm;
  reg COMP_LOOP_COMP_LOOP_and_1599_itm;
  reg COMP_LOOP_COMP_LOOP_and_1600_itm;
  reg COMP_LOOP_COMP_LOOP_and_1601_itm;
  reg COMP_LOOP_COMP_LOOP_and_1602_itm;
  reg COMP_LOOP_COMP_LOOP_and_1603_itm;
  reg COMP_LOOP_COMP_LOOP_and_1604_itm;
  reg COMP_LOOP_COMP_LOOP_and_1605_itm;
  reg COMP_LOOP_nor_1431_itm;
  reg COMP_LOOP_COMP_LOOP_and_1607_itm;
  reg COMP_LOOP_COMP_LOOP_and_1608_itm;
  reg COMP_LOOP_COMP_LOOP_and_1609_itm;
  reg COMP_LOOP_COMP_LOOP_and_1610_itm;
  reg COMP_LOOP_COMP_LOOP_and_1611_itm;
  reg COMP_LOOP_COMP_LOOP_and_1612_itm;
  reg COMP_LOOP_COMP_LOOP_and_1613_itm;
  reg COMP_LOOP_COMP_LOOP_and_1614_itm;
  reg COMP_LOOP_COMP_LOOP_and_1615_itm;
  reg COMP_LOOP_COMP_LOOP_and_1616_itm;
  reg COMP_LOOP_COMP_LOOP_and_1617_itm;
  reg COMP_LOOP_COMP_LOOP_and_1618_itm;
  reg COMP_LOOP_COMP_LOOP_and_1619_itm;
  reg COMP_LOOP_COMP_LOOP_and_1620_itm;
  reg COMP_LOOP_COMP_LOOP_and_1621_itm;
  reg COMP_LOOP_COMP_LOOP_and_1622_itm;
  reg COMP_LOOP_COMP_LOOP_and_1623_itm;
  reg COMP_LOOP_COMP_LOOP_and_1624_itm;
  reg COMP_LOOP_COMP_LOOP_and_1625_itm;
  reg COMP_LOOP_COMP_LOOP_and_1626_itm;
  reg COMP_LOOP_COMP_LOOP_and_1627_itm;
  reg COMP_LOOP_COMP_LOOP_and_1628_itm;
  reg COMP_LOOP_COMP_LOOP_and_1629_itm;
  reg COMP_LOOP_COMP_LOOP_and_1630_itm;
  reg COMP_LOOP_COMP_LOOP_and_1631_itm;
  reg COMP_LOOP_COMP_LOOP_and_1632_itm;
  reg COMP_LOOP_COMP_LOOP_and_1633_itm;
  reg COMP_LOOP_COMP_LOOP_and_1634_itm;
  reg COMP_LOOP_COMP_LOOP_and_1635_itm;
  reg COMP_LOOP_COMP_LOOP_and_1636_itm;
  reg COMP_LOOP_COMP_LOOP_and_1637_itm;
  reg COMP_LOOP_tmp_nor_207_itm;
  reg COMP_LOOP_tmp_nor_209_itm;
  reg COMP_LOOP_tmp_nor_213_itm;
  reg COMP_LOOP_tmp_nor_220_itm;
  reg COMP_LOOP_COMP_LOOP_nor_29_itm;
  reg COMP_LOOP_nor_1625_itm;
  reg COMP_LOOP_nor_1626_itm;
  reg COMP_LOOP_COMP_LOOP_and_1829_itm;
  reg COMP_LOOP_nor_1628_itm;
  reg COMP_LOOP_COMP_LOOP_and_1831_itm;
  reg COMP_LOOP_COMP_LOOP_and_1832_itm;
  reg COMP_LOOP_COMP_LOOP_and_1833_itm;
  reg COMP_LOOP_nor_1632_itm;
  reg COMP_LOOP_COMP_LOOP_and_1835_itm;
  reg COMP_LOOP_COMP_LOOP_and_1836_itm;
  reg COMP_LOOP_COMP_LOOP_and_1837_itm;
  reg COMP_LOOP_COMP_LOOP_and_1838_itm;
  reg COMP_LOOP_COMP_LOOP_and_1839_itm;
  reg COMP_LOOP_COMP_LOOP_and_1840_itm;
  reg COMP_LOOP_COMP_LOOP_and_1841_itm;
  reg COMP_LOOP_nor_1640_itm;
  reg COMP_LOOP_COMP_LOOP_and_1843_itm;
  reg COMP_LOOP_COMP_LOOP_and_1844_itm;
  reg COMP_LOOP_COMP_LOOP_and_1845_itm;
  reg COMP_LOOP_COMP_LOOP_and_1846_itm;
  reg COMP_LOOP_COMP_LOOP_and_1847_itm;
  reg COMP_LOOP_COMP_LOOP_and_1848_itm;
  reg COMP_LOOP_COMP_LOOP_and_1849_itm;
  reg COMP_LOOP_COMP_LOOP_and_1850_itm;
  reg COMP_LOOP_COMP_LOOP_and_1851_itm;
  reg COMP_LOOP_COMP_LOOP_and_1852_itm;
  reg COMP_LOOP_COMP_LOOP_and_1853_itm;
  reg COMP_LOOP_COMP_LOOP_and_1854_itm;
  reg COMP_LOOP_COMP_LOOP_and_1855_itm;
  reg COMP_LOOP_COMP_LOOP_and_1856_itm;
  reg COMP_LOOP_COMP_LOOP_and_1857_itm;
  reg COMP_LOOP_nor_1655_itm;
  reg COMP_LOOP_COMP_LOOP_and_1859_itm;
  reg COMP_LOOP_COMP_LOOP_and_1860_itm;
  reg COMP_LOOP_COMP_LOOP_and_1861_itm;
  reg COMP_LOOP_COMP_LOOP_and_1862_itm;
  reg COMP_LOOP_COMP_LOOP_and_1863_itm;
  reg COMP_LOOP_COMP_LOOP_and_1864_itm;
  reg COMP_LOOP_COMP_LOOP_and_1865_itm;
  reg COMP_LOOP_COMP_LOOP_and_1866_itm;
  reg COMP_LOOP_COMP_LOOP_and_1867_itm;
  reg COMP_LOOP_COMP_LOOP_and_1868_itm;
  reg COMP_LOOP_COMP_LOOP_and_1869_itm;
  reg COMP_LOOP_COMP_LOOP_and_1870_itm;
  reg COMP_LOOP_COMP_LOOP_and_1871_itm;
  reg COMP_LOOP_COMP_LOOP_and_1872_itm;
  reg COMP_LOOP_COMP_LOOP_and_1873_itm;
  reg COMP_LOOP_COMP_LOOP_and_1874_itm;
  reg COMP_LOOP_COMP_LOOP_and_1875_itm;
  reg COMP_LOOP_COMP_LOOP_and_1876_itm;
  reg COMP_LOOP_COMP_LOOP_and_1877_itm;
  reg COMP_LOOP_COMP_LOOP_and_1878_itm;
  reg COMP_LOOP_COMP_LOOP_and_1879_itm;
  reg COMP_LOOP_COMP_LOOP_and_1880_itm;
  reg COMP_LOOP_COMP_LOOP_and_1881_itm;
  reg COMP_LOOP_COMP_LOOP_and_1882_itm;
  reg COMP_LOOP_COMP_LOOP_and_1883_itm;
  reg COMP_LOOP_COMP_LOOP_and_1884_itm;
  reg COMP_LOOP_COMP_LOOP_and_1885_itm;
  reg COMP_LOOP_COMP_LOOP_and_1886_itm;
  reg COMP_LOOP_COMP_LOOP_and_1887_itm;
  reg COMP_LOOP_COMP_LOOP_and_1888_itm;
  reg COMP_LOOP_COMP_LOOP_and_1889_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  wire COMP_LOOP_1_acc_8_itm_mx0c4;
  reg [2:0] COMP_LOOP_1_tmp_mul_idiv_sva_2_0;
  reg [4:0] COMP_LOOP_3_tmp_mul_idiv_sva_4_0;
  wire COMP_LOOP_or_120_rgt;
  wire COMP_LOOP_or_110_rgt;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse;
  wire COMP_LOOP_tmp_nor_76_cse;
  wire COMP_LOOP_tmp_nor_77_cse;
  wire COMP_LOOP_tmp_nor_78_cse;
  wire COMP_LOOP_tmp_nor_79_cse;
  wire COMP_LOOP_tmp_nor_80_cse;
  wire COMP_LOOP_tmp_nor_81_cse;
  wire COMP_LOOP_tmp_nor_82_cse;
  wire COMP_LOOP_tmp_nor_83_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse;
  wire COMP_LOOP_tmp_nor_140_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse;
  wire COMP_LOOP_tmp_nor_141_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse;
  wire COMP_LOOP_tmp_nor_208_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse;
  wire COMP_LOOP_tmp_nor_63_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse;
  wire COMP_LOOP_tmp_nor_64_cse;
  wire COMP_LOOP_tmp_nor_65_cse;
  wire COMP_LOOP_tmp_nor_67_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse;
  wire COMP_LOOP_tmp_nor_68_cse;
  wire COMP_LOOP_tmp_nor_69_cse;
  wire COMP_LOOP_tmp_nor_70_cse;
  wire COMP_LOOP_tmp_nor_71_cse;
  wire COMP_LOOP_tmp_nor_72_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse;
  wire COMP_LOOP_tmp_nor_150_cse;
  wire COMP_LOOP_or_74_cse;
  wire COMP_LOOP_tmp_nor_151_cse;
  wire COMP_LOOP_tmp_nor_153_cse;
  wire COMP_LOOP_tmp_nor_10_cse;
  wire COMP_LOOP_tmp_nor_18_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse;
  wire COMP_LOOP_tmp_nor_34_cse;
  wire COMP_LOOP_tmp_nor_35_cse;
  wire COMP_LOOP_tmp_nor_37_cse;
  wire COMP_LOOP_tmp_nor_41_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse;
  wire nor_746_cse;
  wire nor_740_cse;
  wire nor_735_cse;
  wire nor_734_cse;
  wire nor_730_cse;
  wire nor_719_cse;
  wire nor_714_cse;
  wire nor_713_cse;
  wire nor_709_cse;
  wire nor_703_cse;
  wire nor_697_cse;
  wire nor_692_cse;
  wire nor_691_cse;
  wire nor_687_cse;
  wire nor_676_cse;
  wire nor_671_cse;
  wire nor_670_cse;
  wire nor_666_cse;
  wire nor_660_cse;
  wire nor_654_cse;
  wire nor_649_cse;
  wire nor_648_cse;
  wire nor_644_cse;
  wire nor_633_cse;
  wire nor_628_cse;
  wire nor_627_cse;
  wire nor_623_cse;
  wire nor_617_cse;
  wire nor_611_cse;
  wire nor_606_cse;
  wire nor_605_cse;
  wire nor_601_cse;
  wire nor_590_cse;
  wire nor_585_cse;
  wire nor_584_cse;
  wire and_533_cse;
  wire nor_576_cse;
  wire nor_570_cse;
  wire nor_565_cse;
  wire nor_564_cse;
  wire nor_560_cse;
  wire nor_549_cse;
  wire nor_544_cse;
  wire nor_543_cse;
  wire nor_539_cse;
  wire nor_533_cse;
  wire nor_527_cse;
  wire nor_522_cse;
  wire nor_521_cse;
  wire nor_517_cse;
  wire nor_506_cse;
  wire nor_501_cse;
  wire nor_500_cse;
  wire and_531_cse;
  wire nor_492_cse;
  wire nor_486_cse;
  wire nor_481_cse;
  wire nor_480_cse;
  wire nor_476_cse;
  wire nor_465_cse;
  wire nor_460_cse;
  wire nor_459_cse;
  wire and_529_cse;
  wire nor_451_cse;
  wire nor_446_cse;
  wire nor_441_cse;
  wire nor_440_cse;
  wire and_526_cse;
  wire and_523_cse;
  wire and_519_cse;
  wire and_518_cse;
  wire and_515_cse;
  wire nor_1716_cse;
  wire nor_1715_cse;
  wire COMP_LOOP_or_121_cse;
  wire COMP_LOOP_or_126_cse;
  wire COMP_LOOP_or_135_cse;
  wire COMP_LOOP_or_151_cse;
  wire COMP_LOOP_or_153_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse;
  wire COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse;
  wire and_907_cse;
  wire and_918_cse;
  wire and_903_cse;
  wire and_910_cse;
  wire and_914_cse;
  wire and_920_cse;
  wire nor_1744_cse;
  wire and_1046_cse;
  wire COMP_LOOP_or_68_itm;
  wire COMP_LOOP_or_65_itm;
  wire COMP_LOOP_tmp_or_83_itm;
  wire [9:0] COMP_LOOP_1_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_2_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_3_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_4_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_5_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_6_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_7_acc_10_itm_10_1_1;
  wire [9:0] COMP_LOOP_8_acc_10_itm_10_1_1;
  wire COMP_LOOP_tmp_or_54_ssc;
  wire [63:0] COMP_LOOP_mux_724_cse;
  wire COMP_LOOP_tmp_nor_300_cse;

  wire[0:0] nor_1423_nl;
  wire[0:0] mux_789_nl;
  wire[0:0] mux_788_nl;
  wire[0:0] mux_2996_nl;
  wire[0:0] mux_2995_nl;
  wire[0:0] mux_2993_nl;
  wire[0:0] mux_2992_nl;
  wire[0:0] nor_425_nl;
  wire[0:0] VEC_LOOP_j_not_1_nl;
  wire[0:0] nor_422_nl;
  wire[0:0] nand_480_nl;
  wire[0:0] mux_781_nl;
  wire[0:0] nor_1426_nl;
  wire[0:0] and_637_nl;
  wire[0:0] or_4159_nl;
  wire[0:0] nand_493_nl;
  wire[0:0] mux_3365_nl;
  wire[0:0] mux_nl;
  wire[0:0] nor_1745_nl;
  wire[0:0] or_4154_nl;
  wire[0:0] mux_3031_nl;
  wire[0:0] mux_3030_nl;
  wire[0:0] mux_3029_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_73_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_824_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_74_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_851_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_75_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_858_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_100_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_323_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1073_nl;
  wire[0:0] mux_3037_nl;
  wire[0:0] mux_3036_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_101_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_348_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1075_nl;
  wire[0:0] and_403_nl;
  wire[0:0] mux_3039_nl;
  wire[0:0] nor_420_nl;
  wire[0:0] mux_3045_nl;
  wire[0:0] mux_3044_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_102_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1076_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_103_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_350_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1079_nl;
  wire[0:0] mux_3046_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_104_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_354_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1080_nl;
  wire[0:0] and_409_nl;
  wire[0:0] mux_3047_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_105_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_362_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1082_nl;
  wire[0:0] mux_3048_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_106_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1087_nl;
  wire[0:0] and_411_nl;
  wire[0:0] mux_3053_nl;
  wire[0:0] mux_3052_nl;
  wire[0:0] mux_3051_nl;
  wire[0:0] or_3878_nl;
  wire[0:0] or_3877_nl;
  wire[0:0] mux_3050_nl;
  wire[0:0] mux_3049_nl;
  wire[0:0] nor_418_nl;
  wire[0:0] or_3874_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_107_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1088_nl;
  wire[0:0] mux_3059_nl;
  wire[0:0] mux_3056_nl;
  wire[0:0] mux_3055_nl;
  wire[0:0] mux_3054_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_108_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1090_nl;
  wire[0:0] mux_3063_nl;
  wire[0:0] mux_3062_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_109_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1094_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_110_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1103_nl;
  wire[0:0] mux_3064_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_115_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1328_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_116_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1331_nl;
  wire[0:0] mux_3073_nl;
  wire[0:0] or_3889_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_117_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1332_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_118_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1334_nl;
  wire[0:0] mux_3081_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_119_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1339_nl;
  wire[0:0] mux_3085_nl;
  wire[0:0] mux_3084_nl;
  wire[0:0] nor_414_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_120_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1340_nl;
  wire[0:0] mux_3092_nl;
  wire[0:0] mux_3091_nl;
  wire[0:0] mux_3090_nl;
  wire[0:0] mux_3089_nl;
  wire[0:0] mux_3087_nl;
  wire[0:0] mux_3094_nl;
  wire[0:0] or_3900_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_121_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1342_nl;
  wire[0:0] mux_3097_nl;
  wire[0:0] mux_3096_nl;
  wire[0:0] and_503_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_122_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1355_nl;
  wire[0:0] or_560_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_123_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1356_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_124_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1358_nl;
  wire[0:0] mux_3102_nl;
  wire[0:0] or_3904_nl;
  wire[0:0] nand_145_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_125_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1362_nl;
  wire[0:0] mux_3107_nl;
  wire[0:0] mux_3106_nl;
  wire[0:0] mux_3105_nl;
  wire[0:0] mux_3104_nl;
  wire[0:0] mux_3111_nl;
  wire[0:0] mux_3110_nl;
  wire[0:0] mux_3115_nl;
  wire[0:0] mux_3113_nl;
  wire[0:0] mux_3123_nl;
  wire[10:0] COMP_LOOP_3_acc_nl;
  wire[11:0] nl_COMP_LOOP_3_acc_nl;
  wire[0:0] mux_3124_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] mux_3126_nl;
  wire[0:0] mux_3125_nl;
  wire[8:0] COMP_LOOP_acc_12_nl;
  wire[9:0] nl_COMP_LOOP_acc_12_nl;
  wire[0:0] mux_3128_nl;
  wire[0:0] mux_3127_nl;
  wire[0:0] mux_3130_nl;
  wire[10:0] COMP_LOOP_5_acc_nl;
  wire[11:0] nl_COMP_LOOP_5_acc_nl;
  wire[0:0] mux_3132_nl;
  wire[0:0] mux_3131_nl;
  wire[0:0] mux_3140_nl;
  wire[0:0] mux_3139_nl;
  wire[0:0] mux_3138_nl;
  wire[0:0] and_497_nl;
  wire[0:0] mux_3143_nl;
  wire[0:0] mux_3142_nl;
  wire[10:0] COMP_LOOP_6_acc_nl;
  wire[11:0] nl_COMP_LOOP_6_acc_nl;
  wire[0:0] mux_3146_nl;
  wire[0:0] mux_3152_nl;
  wire[0:0] mux_212_nl;
  wire[0:0] mux_3160_nl;
  wire[0:0] mux_219_nl;
  wire[0:0] or_154_nl;
  wire[0:0] mux_3163_nl;
  wire[0:0] mux_3162_nl;
  wire[0:0] mux_3161_nl;
  wire[0:0] nor_410_nl;
  wire[0:0] and_491_nl;
  wire[0:0] and_492_nl;
  wire[10:0] COMP_LOOP_7_acc_nl;
  wire[11:0] nl_COMP_LOOP_7_acc_nl;
  wire[0:0] mux_3171_nl;
  wire[0:0] mux_3182_nl;
  wire[0:0] mux_3181_nl;
  wire[7:0] COMP_LOOP_acc_15_nl;
  wire[8:0] nl_COMP_LOOP_acc_15_nl;
  wire[0:0] mux_3188_nl;
  wire[0:0] nand_148_nl;
  wire[0:0] mux_3192_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] mux_3193_nl;
  wire[10:0] COMP_LOOP_1_acc_nl;
  wire[11:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] mux_3197_nl;
  wire[0:0] mux_3205_nl;
  wire[0:0] mux_3204_nl;
  wire[0:0] mux_3203_nl;
  wire[0:0] and_489_nl;
  wire[0:0] mux_3202_nl;
  wire[0:0] mux_3210_nl;
  wire[0:0] mux_3209_nl;
  wire[0:0] mux_3208_nl;
  wire[0:0] and_449_nl;
  wire[0:0] mux_3207_nl;
  wire[0:0] mux_3206_nl;
  wire[0:0] mux_3216_nl;
  wire[0:0] mux_3215_nl;
  wire[0:0] mux_3214_nl;
  wire[0:0] mux_3213_nl;
  wire[0:0] mux_3212_nl;
  wire[0:0] mux_3211_nl;
  wire[0:0] mux_3219_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_111_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1104_nl;
  wire[0:0] mux_3223_nl;
  wire[0:0] mux_3222_nl;
  wire[0:0] mux_3221_nl;
  wire[0:0] or_3932_nl;
  wire[0:0] mux_3220_nl;
  wire[0:0] or_3929_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_112_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1106_nl;
  wire[0:0] mux_3226_nl;
  wire[0:0] mux_3225_nl;
  wire[0:0] mux_3224_nl;
  wire[0:0] or_3934_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_113_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1110_nl;
  wire[0:0] mux_3227_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_114_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1118_nl;
  wire[0:0] mux_3229_nl;
  wire[0:0] mux_3228_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_65_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1370_nl;
  wire[0:0] mux_3231_nl;
  wire[0:0] mux_3230_nl;
  wire[0:0] mux_3234_nl;
  wire[0:0] mux_3233_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_67_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1577_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_68_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1584_nl;
  wire[0:0] mux_3238_nl;
  wire[0:0] mux_3237_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_317_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1594_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_319_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1598_nl;
  wire[0:0] mux_3243_nl;
  wire[0:0] mux_3242_nl;
  wire[0:0] mux_3241_nl;
  wire[0:0] nor_403_nl;
  wire[0:0] nor_405_nl;
  wire[0:0] mux_3240_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_320_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1607_nl;
  wire[0:0] and_458_nl;
  wire[0:0] mux_3246_nl;
  wire[0:0] mux_3245_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_321_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1610_nl;
  wire[0:0] mux_3253_nl;
  wire[0:0] mux_3252_nl;
  wire[0:0] mux_3251_nl;
  wire[0:0] or_3946_nl;
  wire[0:0] mux_582_nl;
  wire[0:0] mux_3249_nl;
  wire[0:0] mux_3248_nl;
  wire[0:0] or_3943_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_324_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1614_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_325_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1622_nl;
  wire[0:0] and_459_nl;
  wire[0:0] mux_3256_nl;
  wire[0:0] mux_3255_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_69_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1831_nl;
  wire[0:0] mux_3264_nl;
  wire[0:0] mux_3261_nl;
  wire[0:0] mux_3259_nl;
  wire[0:0] mux_3258_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_326_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1832_nl;
  wire[0:0] and_461_nl;
  wire[0:0] mux_3274_nl;
  wire[0:0] mux_3273_nl;
  wire[0:0] mux_3272_nl;
  wire[0:0] mux_3271_nl;
  wire[0:0] mux_3270_nl;
  wire[0:0] mux_3269_nl;
  wire[0:0] mux_3268_nl;
  wire[0:0] nor_386_nl;
  wire[0:0] mux_3267_nl;
  wire[0:0] nor_384_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_327_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1835_nl;
  wire[0:0] and_463_nl;
  wire[0:0] mux_3283_nl;
  wire[0:0] mux_3282_nl;
  wire[0:0] mux_3279_nl;
  wire[0:0] mux_3278_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_328_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1844_nl;
  wire[0:0] mux_3286_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_329_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1850_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_331_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1862_nl;
  wire[0:0] and_465_nl;
  wire[0:0] mux_3292_nl;
  wire[0:0] mux_3291_nl;
  wire[0:0] and_464_nl;
  wire[0:0] mux_3290_nl;
  wire[0:0] mux_3289_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_332_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1866_nl;
  wire[0:0] and_468_nl;
  wire[0:0] mux_3298_nl;
  wire[0:0] mux_3297_nl;
  wire[0:0] mux_3296_nl;
  wire[0:0] and_73_nl;
  wire[0:0] mux_3295_nl;
  wire[0:0] mux_3294_nl;
  wire[0:0] and_466_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_71_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1874_nl;
  wire[0:0] mux_3302_nl;
  wire[0:0] mux_3301_nl;
  wire[0:0] mux_3300_nl;
  wire[0:0] nor_397_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_72_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_583_nl;
  wire[0:0] mux_3306_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_nor_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_76_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_79_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_80_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_81_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_82_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_83_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_86_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_87_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_88_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_89_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_90_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_91_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_92_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_93_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_95_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_96_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_97_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_98_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nor_1_nl;
  wire[0:0] COMP_LOOP_nor_57_nl;
  wire[0:0] COMP_LOOP_nor_58_nl;
  wire[0:0] COMP_LOOP_nor_60_nl;
  wire[0:0] COMP_LOOP_nor_64_nl;
  wire[0:0] COMP_LOOP_nor_72_nl;
  wire[0:0] COMP_LOOP_nor_87_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl;
  wire[63:0] COMP_LOOP_acc_17_nl;
  wire[64:0] nl_COMP_LOOP_acc_17_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_mux_21_nl;
  wire[0:0] COMP_LOOP_or_nl;
  wire[0:0] COMP_LOOP_or_1_nl;
  wire[0:0] COMP_LOOP_or_2_nl;
  wire[0:0] COMP_LOOP_or_3_nl;
  wire[0:0] COMP_LOOP_or_4_nl;
  wire[0:0] COMP_LOOP_or_5_nl;
  wire[0:0] COMP_LOOP_or_6_nl;
  wire[0:0] COMP_LOOP_or_7_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_or_23_nl;
  wire[0:0] COMP_LOOP_or_24_nl;
  wire[0:0] COMP_LOOP_or_25_nl;
  wire[0:0] COMP_LOOP_or_26_nl;
  wire[0:0] COMP_LOOP_or_27_nl;
  wire[0:0] COMP_LOOP_or_28_nl;
  wire[0:0] COMP_LOOP_or_29_nl;
  wire[0:0] COMP_LOOP_or_30_nl;
  wire[0:0] COMP_LOOP_or_31_nl;
  wire[0:0] COMP_LOOP_or_32_nl;
  wire[0:0] COMP_LOOP_or_33_nl;
  wire[0:0] COMP_LOOP_or_34_nl;
  wire[0:0] COMP_LOOP_or_35_nl;
  wire[0:0] COMP_LOOP_or_36_nl;
  wire[0:0] COMP_LOOP_or_37_nl;
  wire[0:0] COMP_LOOP_or_38_nl;
  wire[0:0] COMP_LOOP_or_39_nl;
  wire[0:0] COMP_LOOP_or_40_nl;
  wire[0:0] COMP_LOOP_or_41_nl;
  wire[0:0] COMP_LOOP_or_42_nl;
  wire[0:0] COMP_LOOP_or_43_nl;
  wire[0:0] COMP_LOOP_or_44_nl;
  wire[0:0] COMP_LOOP_or_45_nl;
  wire[0:0] COMP_LOOP_or_46_nl;
  wire[0:0] COMP_LOOP_or_47_nl;
  wire[0:0] COMP_LOOP_or_48_nl;
  wire[0:0] COMP_LOOP_or_49_nl;
  wire[0:0] COMP_LOOP_or_50_nl;
  wire[0:0] COMP_LOOP_or_51_nl;
  wire[0:0] COMP_LOOP_or_52_nl;
  wire[0:0] COMP_LOOP_or_53_nl;
  wire[0:0] COMP_LOOP_or_54_nl;
  wire[0:0] COMP_LOOP_or_55_nl;
  wire[0:0] COMP_LOOP_or_56_nl;
  wire[0:0] COMP_LOOP_or_57_nl;
  wire[0:0] COMP_LOOP_or_58_nl;
  wire[0:0] COMP_LOOP_or_59_nl;
  wire[0:0] COMP_LOOP_or_60_nl;
  wire[0:0] COMP_LOOP_or_61_nl;
  wire[0:0] COMP_LOOP_or_62_nl;
  wire[0:0] COMP_LOOP_or_63_nl;
  wire[0:0] COMP_LOOP_tmp_and_249_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_nl;
  wire[0:0] COMP_LOOP_tmp_and_250_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_nl;
  wire[0:0] COMP_LOOP_tmp_and_251_nl;
  wire[0:0] COMP_LOOP_tmp_and_252_nl;
  wire[0:0] COMP_LOOP_tmp_and_253_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_nl;
  wire[0:0] COMP_LOOP_tmp_and_254_nl;
  wire[0:0] COMP_LOOP_tmp_and_255_nl;
  wire[0:0] COMP_LOOP_tmp_and_256_nl;
  wire[0:0] COMP_LOOP_tmp_and_257_nl;
  wire[0:0] COMP_LOOP_tmp_and_258_nl;
  wire[0:0] COMP_LOOP_tmp_and_259_nl;
  wire[0:0] COMP_LOOP_tmp_and_260_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_22_nl;
  wire[0:0] COMP_LOOP_tmp_and_261_nl;
  wire[0:0] COMP_LOOP_tmp_and_262_nl;
  wire[0:0] COMP_LOOP_tmp_and_263_nl;
  wire[0:0] COMP_LOOP_tmp_and_264_nl;
  wire[0:0] COMP_LOOP_tmp_and_265_nl;
  wire[0:0] COMP_LOOP_tmp_and_266_nl;
  wire[0:0] COMP_LOOP_tmp_and_267_nl;
  wire[0:0] COMP_LOOP_tmp_and_268_nl;
  wire[0:0] COMP_LOOP_tmp_and_269_nl;
  wire[0:0] COMP_LOOP_tmp_and_270_nl;
  wire[0:0] COMP_LOOP_tmp_and_271_nl;
  wire[0:0] COMP_LOOP_tmp_and_272_nl;
  wire[0:0] COMP_LOOP_tmp_and_273_nl;
  wire[0:0] COMP_LOOP_tmp_and_274_nl;
  wire[0:0] COMP_LOOP_tmp_and_275_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_nl;
  wire[0:0] COMP_LOOP_tmp_and_276_nl;
  wire[0:0] COMP_LOOP_tmp_and_277_nl;
  wire[0:0] COMP_LOOP_tmp_and_278_nl;
  wire[0:0] COMP_LOOP_tmp_and_279_nl;
  wire[0:0] COMP_LOOP_tmp_and_280_nl;
  wire[0:0] COMP_LOOP_tmp_and_281_nl;
  wire[0:0] COMP_LOOP_tmp_and_282_nl;
  wire[0:0] COMP_LOOP_tmp_and_283_nl;
  wire[0:0] COMP_LOOP_tmp_and_284_nl;
  wire[0:0] COMP_LOOP_tmp_and_285_nl;
  wire[0:0] COMP_LOOP_tmp_and_286_nl;
  wire[0:0] COMP_LOOP_tmp_and_287_nl;
  wire[0:0] COMP_LOOP_tmp_and_288_nl;
  wire[0:0] COMP_LOOP_tmp_and_289_nl;
  wire[0:0] COMP_LOOP_tmp_and_290_nl;
  wire[0:0] COMP_LOOP_tmp_and_291_nl;
  wire[0:0] COMP_LOOP_tmp_and_292_nl;
  wire[0:0] COMP_LOOP_tmp_and_293_nl;
  wire[0:0] COMP_LOOP_tmp_and_294_nl;
  wire[0:0] COMP_LOOP_tmp_and_295_nl;
  wire[0:0] COMP_LOOP_tmp_and_296_nl;
  wire[0:0] COMP_LOOP_tmp_and_297_nl;
  wire[0:0] COMP_LOOP_tmp_and_298_nl;
  wire[0:0] COMP_LOOP_tmp_and_299_nl;
  wire[0:0] COMP_LOOP_tmp_and_300_nl;
  wire[0:0] COMP_LOOP_tmp_and_301_nl;
  wire[0:0] COMP_LOOP_tmp_and_302_nl;
  wire[0:0] COMP_LOOP_tmp_and_303_nl;
  wire[0:0] COMP_LOOP_tmp_and_304_nl;
  wire[0:0] COMP_LOOP_tmp_and_305_nl;
  wire[0:0] COMP_LOOP_tmp_and_306_nl;
  wire[0:0] COMP_LOOP_tmp_and_222_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_70_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_71_nl;
  wire[0:0] COMP_LOOP_tmp_and_223_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_73_nl;
  wire[0:0] COMP_LOOP_tmp_and_224_nl;
  wire[0:0] COMP_LOOP_tmp_and_225_nl;
  wire[0:0] COMP_LOOP_tmp_and_226_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_77_nl;
  wire[0:0] COMP_LOOP_tmp_and_227_nl;
  wire[0:0] COMP_LOOP_tmp_and_228_nl;
  wire[0:0] COMP_LOOP_tmp_and_229_nl;
  wire[0:0] COMP_LOOP_tmp_and_230_nl;
  wire[0:0] COMP_LOOP_tmp_and_231_nl;
  wire[0:0] COMP_LOOP_tmp_and_232_nl;
  wire[0:0] COMP_LOOP_tmp_and_233_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_nl;
  wire[0:0] COMP_LOOP_tmp_and_234_nl;
  wire[0:0] COMP_LOOP_tmp_and_235_nl;
  wire[0:0] COMP_LOOP_tmp_and_236_nl;
  wire[0:0] COMP_LOOP_tmp_and_237_nl;
  wire[0:0] COMP_LOOP_tmp_and_238_nl;
  wire[0:0] COMP_LOOP_tmp_and_239_nl;
  wire[0:0] COMP_LOOP_tmp_and_240_nl;
  wire[0:0] COMP_LOOP_tmp_and_241_nl;
  wire[0:0] COMP_LOOP_tmp_and_242_nl;
  wire[0:0] COMP_LOOP_tmp_and_243_nl;
  wire[0:0] COMP_LOOP_tmp_and_244_nl;
  wire[0:0] COMP_LOOP_tmp_and_245_nl;
  wire[0:0] COMP_LOOP_tmp_and_246_nl;
  wire[0:0] COMP_LOOP_tmp_and_247_nl;
  wire[0:0] COMP_LOOP_tmp_and_248_nl;
  wire[0:0] COMP_LOOP_tmp_and_164_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_102_nl;
  wire[0:0] COMP_LOOP_tmp_and_165_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_nl;
  wire[0:0] COMP_LOOP_tmp_and_166_nl;
  wire[0:0] COMP_LOOP_tmp_and_167_nl;
  wire[0:0] COMP_LOOP_tmp_and_168_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_nl;
  wire[0:0] COMP_LOOP_tmp_and_169_nl;
  wire[0:0] COMP_LOOP_tmp_and_170_nl;
  wire[0:0] COMP_LOOP_tmp_and_171_nl;
  wire[0:0] COMP_LOOP_tmp_and_172_nl;
  wire[0:0] COMP_LOOP_tmp_and_173_nl;
  wire[0:0] COMP_LOOP_tmp_and_174_nl;
  wire[0:0] COMP_LOOP_tmp_and_175_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_nl;
  wire[0:0] COMP_LOOP_tmp_and_176_nl;
  wire[0:0] COMP_LOOP_tmp_and_177_nl;
  wire[0:0] COMP_LOOP_tmp_and_178_nl;
  wire[0:0] COMP_LOOP_tmp_and_179_nl;
  wire[0:0] COMP_LOOP_tmp_and_180_nl;
  wire[0:0] COMP_LOOP_tmp_and_181_nl;
  wire[0:0] COMP_LOOP_tmp_and_182_nl;
  wire[0:0] COMP_LOOP_tmp_and_183_nl;
  wire[0:0] COMP_LOOP_tmp_and_184_nl;
  wire[0:0] COMP_LOOP_tmp_and_185_nl;
  wire[0:0] COMP_LOOP_tmp_and_186_nl;
  wire[0:0] COMP_LOOP_tmp_and_187_nl;
  wire[0:0] COMP_LOOP_tmp_and_188_nl;
  wire[0:0] COMP_LOOP_tmp_and_189_nl;
  wire[0:0] COMP_LOOP_tmp_and_190_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_nl;
  wire[0:0] COMP_LOOP_tmp_and_191_nl;
  wire[0:0] COMP_LOOP_tmp_and_192_nl;
  wire[0:0] COMP_LOOP_tmp_and_193_nl;
  wire[0:0] COMP_LOOP_tmp_and_194_nl;
  wire[0:0] COMP_LOOP_tmp_and_195_nl;
  wire[0:0] COMP_LOOP_tmp_and_196_nl;
  wire[0:0] COMP_LOOP_tmp_and_197_nl;
  wire[0:0] COMP_LOOP_tmp_and_198_nl;
  wire[0:0] COMP_LOOP_tmp_and_199_nl;
  wire[0:0] COMP_LOOP_tmp_and_200_nl;
  wire[0:0] COMP_LOOP_tmp_and_201_nl;
  wire[0:0] COMP_LOOP_tmp_and_202_nl;
  wire[0:0] COMP_LOOP_tmp_and_203_nl;
  wire[0:0] COMP_LOOP_tmp_and_204_nl;
  wire[0:0] COMP_LOOP_tmp_and_205_nl;
  wire[0:0] COMP_LOOP_tmp_and_206_nl;
  wire[0:0] COMP_LOOP_tmp_and_207_nl;
  wire[0:0] COMP_LOOP_tmp_and_208_nl;
  wire[0:0] COMP_LOOP_tmp_and_209_nl;
  wire[0:0] COMP_LOOP_tmp_and_210_nl;
  wire[0:0] COMP_LOOP_tmp_and_211_nl;
  wire[0:0] COMP_LOOP_tmp_and_212_nl;
  wire[0:0] COMP_LOOP_tmp_and_213_nl;
  wire[0:0] COMP_LOOP_tmp_and_214_nl;
  wire[0:0] COMP_LOOP_tmp_and_215_nl;
  wire[0:0] COMP_LOOP_tmp_and_216_nl;
  wire[0:0] COMP_LOOP_tmp_and_217_nl;
  wire[0:0] COMP_LOOP_tmp_and_218_nl;
  wire[0:0] COMP_LOOP_tmp_and_219_nl;
  wire[0:0] COMP_LOOP_tmp_and_220_nl;
  wire[0:0] COMP_LOOP_tmp_and_221_nl;
  wire[0:0] COMP_LOOP_tmp_and_152_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_164_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_165_nl;
  wire[0:0] COMP_LOOP_tmp_and_153_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_167_nl;
  wire[0:0] COMP_LOOP_tmp_and_154_nl;
  wire[0:0] COMP_LOOP_tmp_and_155_nl;
  wire[0:0] COMP_LOOP_tmp_and_156_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_171_nl;
  wire[0:0] COMP_LOOP_tmp_and_157_nl;
  wire[0:0] COMP_LOOP_tmp_and_158_nl;
  wire[0:0] COMP_LOOP_tmp_and_159_nl;
  wire[0:0] COMP_LOOP_tmp_and_160_nl;
  wire[0:0] COMP_LOOP_tmp_and_161_nl;
  wire[0:0] COMP_LOOP_tmp_and_162_nl;
  wire[0:0] COMP_LOOP_tmp_and_163_nl;
  wire[0:0] COMP_LOOP_tmp_and_89_nl;
  wire[0:0] COMP_LOOP_tmp_and_90_nl;
  wire[0:0] COMP_LOOP_tmp_and_91_nl;
  wire[0:0] COMP_LOOP_tmp_and_92_nl;
  wire[0:0] COMP_LOOP_tmp_and_93_nl;
  wire[0:0] COMP_LOOP_tmp_and_94_nl;
  wire[0:0] COMP_LOOP_tmp_and_95_nl;
  wire[0:0] COMP_LOOP_tmp_and_96_nl;
  wire[0:0] COMP_LOOP_tmp_and_97_nl;
  wire[0:0] COMP_LOOP_tmp_and_98_nl;
  wire[0:0] COMP_LOOP_tmp_and_99_nl;
  wire[0:0] COMP_LOOP_tmp_and_100_nl;
  wire[0:0] COMP_LOOP_tmp_and_101_nl;
  wire[0:0] COMP_LOOP_tmp_and_102_nl;
  wire[0:0] COMP_LOOP_tmp_and_103_nl;
  wire[0:0] COMP_LOOP_tmp_and_104_nl;
  wire[0:0] COMP_LOOP_tmp_and_105_nl;
  wire[0:0] COMP_LOOP_tmp_and_106_nl;
  wire[0:0] COMP_LOOP_tmp_and_107_nl;
  wire[0:0] COMP_LOOP_tmp_and_108_nl;
  wire[0:0] COMP_LOOP_tmp_and_109_nl;
  wire[0:0] COMP_LOOP_tmp_and_110_nl;
  wire[0:0] COMP_LOOP_tmp_and_111_nl;
  wire[0:0] COMP_LOOP_tmp_and_112_nl;
  wire[0:0] COMP_LOOP_tmp_and_113_nl;
  wire[0:0] COMP_LOOP_tmp_and_114_nl;
  wire[0:0] COMP_LOOP_tmp_and_115_nl;
  wire[0:0] COMP_LOOP_tmp_and_116_nl;
  wire[0:0] COMP_LOOP_tmp_and_117_nl;
  wire[0:0] COMP_LOOP_tmp_and_118_nl;
  wire[0:0] COMP_LOOP_tmp_and_119_nl;
  wire[0:0] COMP_LOOP_tmp_and_120_nl;
  wire[0:0] COMP_LOOP_tmp_and_121_nl;
  wire[0:0] COMP_LOOP_tmp_and_122_nl;
  wire[0:0] COMP_LOOP_tmp_and_123_nl;
  wire[0:0] COMP_LOOP_tmp_and_124_nl;
  wire[0:0] COMP_LOOP_tmp_and_125_nl;
  wire[0:0] COMP_LOOP_tmp_and_126_nl;
  wire[0:0] COMP_LOOP_tmp_and_127_nl;
  wire[0:0] COMP_LOOP_tmp_and_128_nl;
  wire[0:0] COMP_LOOP_tmp_and_129_nl;
  wire[0:0] COMP_LOOP_tmp_and_130_nl;
  wire[0:0] COMP_LOOP_tmp_and_131_nl;
  wire[0:0] COMP_LOOP_tmp_and_132_nl;
  wire[0:0] COMP_LOOP_tmp_and_133_nl;
  wire[0:0] COMP_LOOP_tmp_and_134_nl;
  wire[0:0] COMP_LOOP_tmp_and_135_nl;
  wire[0:0] COMP_LOOP_tmp_and_136_nl;
  wire[0:0] COMP_LOOP_tmp_and_137_nl;
  wire[0:0] COMP_LOOP_tmp_and_138_nl;
  wire[0:0] COMP_LOOP_tmp_and_139_nl;
  wire[0:0] COMP_LOOP_tmp_and_140_nl;
  wire[0:0] COMP_LOOP_tmp_and_141_nl;
  wire[0:0] COMP_LOOP_tmp_and_142_nl;
  wire[0:0] COMP_LOOP_tmp_and_143_nl;
  wire[0:0] COMP_LOOP_tmp_and_144_nl;
  wire[0:0] COMP_LOOP_tmp_and_145_nl;
  wire[0:0] COMP_LOOP_tmp_and_146_nl;
  wire[0:0] COMP_LOOP_tmp_and_147_nl;
  wire[0:0] COMP_LOOP_tmp_and_148_nl;
  wire[0:0] COMP_LOOP_tmp_and_149_nl;
  wire[0:0] COMP_LOOP_tmp_and_150_nl;
  wire[0:0] COMP_LOOP_tmp_and_151_nl;
  wire[0:0] mux_3353_nl;
  wire[0:0] mux_3352_nl;
  wire[0:0] mux_3351_nl;
  wire[0:0] mux_3350_nl;
  wire[0:0] mux_3349_nl;
  wire[0:0] mux_3348_nl;
  wire[0:0] mux_3359_nl;
  wire[0:0] mux_3358_nl;
  wire[0:0] mux_3357_nl;
  wire[0:0] mux_3356_nl;
  wire[0:0] COMP_LOOP_tmp_and_31_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_179_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_180_nl;
  wire[0:0] COMP_LOOP_tmp_and_32_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_182_nl;
  wire[0:0] COMP_LOOP_tmp_and_33_nl;
  wire[0:0] COMP_LOOP_tmp_and_34_nl;
  wire[0:0] COMP_LOOP_tmp_and_35_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_186_nl;
  wire[0:0] COMP_LOOP_tmp_and_36_nl;
  wire[0:0] COMP_LOOP_tmp_and_37_nl;
  wire[0:0] COMP_LOOP_tmp_and_38_nl;
  wire[0:0] COMP_LOOP_tmp_and_39_nl;
  wire[0:0] COMP_LOOP_tmp_and_40_nl;
  wire[0:0] COMP_LOOP_tmp_and_41_nl;
  wire[0:0] COMP_LOOP_tmp_and_42_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_194_nl;
  wire[0:0] COMP_LOOP_tmp_and_43_nl;
  wire[0:0] COMP_LOOP_tmp_and_44_nl;
  wire[0:0] COMP_LOOP_tmp_and_45_nl;
  wire[0:0] COMP_LOOP_tmp_and_46_nl;
  wire[0:0] COMP_LOOP_tmp_and_47_nl;
  wire[0:0] COMP_LOOP_tmp_and_48_nl;
  wire[0:0] COMP_LOOP_tmp_and_49_nl;
  wire[0:0] COMP_LOOP_tmp_and_50_nl;
  wire[0:0] COMP_LOOP_tmp_and_51_nl;
  wire[0:0] COMP_LOOP_tmp_and_52_nl;
  wire[0:0] COMP_LOOP_tmp_and_53_nl;
  wire[0:0] COMP_LOOP_tmp_and_54_nl;
  wire[0:0] COMP_LOOP_tmp_and_55_nl;
  wire[0:0] COMP_LOOP_tmp_and_56_nl;
  wire[0:0] COMP_LOOP_tmp_and_57_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_210_nl;
  wire[0:0] COMP_LOOP_tmp_and_58_nl;
  wire[0:0] COMP_LOOP_tmp_and_59_nl;
  wire[0:0] COMP_LOOP_tmp_and_60_nl;
  wire[0:0] COMP_LOOP_tmp_and_61_nl;
  wire[0:0] COMP_LOOP_tmp_and_62_nl;
  wire[0:0] COMP_LOOP_tmp_and_63_nl;
  wire[0:0] COMP_LOOP_tmp_and_64_nl;
  wire[0:0] COMP_LOOP_tmp_and_65_nl;
  wire[0:0] COMP_LOOP_tmp_and_66_nl;
  wire[0:0] COMP_LOOP_tmp_and_67_nl;
  wire[0:0] COMP_LOOP_tmp_and_68_nl;
  wire[0:0] COMP_LOOP_tmp_and_69_nl;
  wire[0:0] COMP_LOOP_tmp_and_70_nl;
  wire[0:0] COMP_LOOP_tmp_and_71_nl;
  wire[0:0] COMP_LOOP_tmp_and_72_nl;
  wire[0:0] COMP_LOOP_tmp_and_73_nl;
  wire[0:0] COMP_LOOP_tmp_and_74_nl;
  wire[0:0] COMP_LOOP_tmp_and_75_nl;
  wire[0:0] COMP_LOOP_tmp_and_76_nl;
  wire[0:0] COMP_LOOP_tmp_and_77_nl;
  wire[0:0] COMP_LOOP_tmp_and_78_nl;
  wire[0:0] COMP_LOOP_tmp_and_79_nl;
  wire[0:0] COMP_LOOP_tmp_and_80_nl;
  wire[0:0] COMP_LOOP_tmp_and_81_nl;
  wire[0:0] COMP_LOOP_tmp_and_82_nl;
  wire[0:0] COMP_LOOP_tmp_and_83_nl;
  wire[0:0] COMP_LOOP_tmp_and_84_nl;
  wire[0:0] COMP_LOOP_tmp_and_85_nl;
  wire[0:0] COMP_LOOP_tmp_and_86_nl;
  wire[0:0] COMP_LOOP_tmp_and_87_nl;
  wire[0:0] COMP_LOOP_tmp_and_88_nl;
  wire[0:0] COMP_LOOP_tmp_and_nl;
  wire[0:0] COMP_LOOP_tmp_and_1_nl;
  wire[0:0] COMP_LOOP_tmp_and_2_nl;
  wire[0:0] COMP_LOOP_tmp_and_3_nl;
  wire[0:0] COMP_LOOP_tmp_and_4_nl;
  wire[0:0] COMP_LOOP_tmp_and_5_nl;
  wire[0:0] COMP_LOOP_tmp_and_6_nl;
  wire[0:0] COMP_LOOP_tmp_and_7_nl;
  wire[0:0] COMP_LOOP_tmp_and_8_nl;
  wire[0:0] COMP_LOOP_tmp_and_9_nl;
  wire[0:0] COMP_LOOP_tmp_and_10_nl;
  wire[0:0] COMP_LOOP_tmp_and_11_nl;
  wire[0:0] COMP_LOOP_tmp_and_12_nl;
  wire[0:0] COMP_LOOP_tmp_and_13_nl;
  wire[0:0] COMP_LOOP_tmp_and_14_nl;
  wire[0:0] COMP_LOOP_tmp_and_15_nl;
  wire[0:0] COMP_LOOP_tmp_and_16_nl;
  wire[0:0] COMP_LOOP_tmp_and_17_nl;
  wire[0:0] COMP_LOOP_tmp_and_18_nl;
  wire[0:0] COMP_LOOP_tmp_and_19_nl;
  wire[0:0] COMP_LOOP_tmp_and_20_nl;
  wire[0:0] COMP_LOOP_tmp_and_21_nl;
  wire[0:0] COMP_LOOP_tmp_and_22_nl;
  wire[0:0] COMP_LOOP_tmp_and_23_nl;
  wire[0:0] COMP_LOOP_tmp_and_24_nl;
  wire[0:0] COMP_LOOP_tmp_and_25_nl;
  wire[0:0] COMP_LOOP_tmp_and_26_nl;
  wire[0:0] COMP_LOOP_tmp_and_27_nl;
  wire[0:0] COMP_LOOP_tmp_and_28_nl;
  wire[0:0] COMP_LOOP_tmp_and_29_nl;
  wire[0:0] COMP_LOOP_tmp_and_30_nl;
  wire[0:0] mux_3364_nl;
  wire[0:0] mux_3363_nl;
  wire[0:0] mux_3362_nl;
  wire[0:0] mux_3361_nl;
  wire[10:0] COMP_LOOP_1_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_1_acc_10_nl;
  wire[10:0] COMP_LOOP_2_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_2_acc_10_nl;
  wire[10:0] COMP_LOOP_3_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_3_acc_10_nl;
  wire[10:0] COMP_LOOP_4_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_4_acc_10_nl;
  wire[10:0] COMP_LOOP_5_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_5_acc_10_nl;
  wire[10:0] COMP_LOOP_6_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_6_acc_10_nl;
  wire[10:0] COMP_LOOP_7_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_7_acc_10_nl;
  wire[10:0] COMP_LOOP_8_acc_10_nl;
  wire[12:0] nl_COMP_LOOP_8_acc_10_nl;
  wire[0:0] mux_510_nl;
  wire[0:0] or_201_nl;
  wire[0:0] mux_3004_nl;
  wire[0:0] mux_522_nl;
  wire[0:0] or_3843_nl;
  wire[0:0] mux_3024_nl;
  wire[0:0] mux_3021_nl;
  wire[0:0] mux_3034_nl;
  wire[0:0] mux_3041_nl;
  wire[0:0] mux_3057_nl;
  wire[0:0] or_3880_nl;
  wire[0:0] or_3887_nl;
  wire[0:0] mux_3069_nl;
  wire[0:0] mux_3067_nl;
  wire[0:0] mux_3065_nl;
  wire[0:0] or_3884_nl;
  wire[0:0] mux_3075_nl;
  wire[0:0] or_3906_nl;
  wire[0:0] mux_3119_nl;
  wire[0:0] mux_3118_nl;
  wire[0:0] mux_3117_nl;
  wire[0:0] mux_3122_nl;
  wire[0:0] mux_67_nl;
  wire[0:0] mux_3129_nl;
  wire[0:0] mux_3135_nl;
  wire[0:0] mux_3134_nl;
  wire[0:0] mux_3133_nl;
  wire[0:0] nor_1425_nl;
  wire[0:0] mux_3148_nl;
  wire[0:0] mux_3150_nl;
  wire[0:0] mux_210_nl;
  wire[0:0] mux_3156_nl;
  wire[0:0] mux_215_nl;
  wire[0:0] mux_214_nl;
  wire[0:0] mux_3158_nl;
  wire[0:0] mux_217_nl;
  wire[0:0] mux_3166_nl;
  wire[0:0] mux_3174_nl;
  wire[0:0] mux_3173_nl;
  wire[0:0] mux_3178_nl;
  wire[0:0] mux_3177_nl;
  wire[0:0] mux_3176_nl;
  wire[0:0] mux_3180_nl;
  wire[0:0] mux_3179_nl;
  wire[0:0] mux_3184_nl;
  wire[0:0] nor_1524_nl;
  wire[0:0] nor_409_nl;
  wire[0:0] mux_3199_nl;
  wire[0:0] mux_3262_nl;
  wire[0:0] nor_400_nl;
  wire[0:0] nor_1474_nl;
  wire[0:0] mux_75_nl;
  wire[0:0] mux_3314_nl;
  wire[0:0] nor_1709_nl;
  wire[0:0] nor_1710_nl;
  wire[0:0] mux_3354_nl;
  wire[0:0] mux_3320_nl;
  wire[0:0] mux_3319_nl;
  wire[0:0] mux_3318_nl;
  wire[0:0] mux_3317_nl;
  wire[0:0] mux_3316_nl;
  wire[0:0] or_3973_nl;
  wire[0:0] mux_3315_nl;
  wire[0:0] mux_3340_nl;
  wire[0:0] mux_3343_nl;
  wire[0:0] mux_3342_nl;
  wire[0:0] mux_104_nl;
  wire[0:0] mux_3346_nl;
  wire[0:0] mux_3345_nl;
  wire[0:0] mux_3344_nl;
  wire[0:0] and_102_nl;
  wire[0:0] and_114_nl;
  wire[0:0] and_120_nl;
  wire[0:0] and_124_nl;
  wire[0:0] and_129_nl;
  wire[0:0] and_133_nl;
  wire[0:0] and_136_nl;
  wire[0:0] and_138_nl;
  wire[0:0] and_142_nl;
  wire[0:0] and_145_nl;
  wire[0:0] and_148_nl;
  wire[0:0] and_151_nl;
  wire[0:0] and_152_nl;
  wire[0:0] and_153_nl;
  wire[0:0] and_154_nl;
  wire[0:0] and_155_nl;
  wire[0:0] and_156_nl;
  wire[0:0] and_157_nl;
  wire[0:0] and_158_nl;
  wire[0:0] and_159_nl;
  wire[0:0] and_160_nl;
  wire[0:0] mux_805_nl;
  wire[0:0] nand_469_nl;
  wire[0:0] mux_804_nl;
  wire[0:0] mux_803_nl;
  wire[0:0] mux_802_nl;
  wire[0:0] nor_1414_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] mux_801_nl;
  wire[0:0] nor_1416_nl;
  wire[0:0] nor_1417_nl;
  wire[0:0] mux_800_nl;
  wire[0:0] mux_799_nl;
  wire[0:0] nor_1418_nl;
  wire[0:0] nor_1419_nl;
  wire[0:0] mux_798_nl;
  wire[0:0] nor_1420_nl;
  wire[0:0] nor_1421_nl;
  wire[0:0] or_4142_nl;
  wire[0:0] mux_797_nl;
  wire[0:0] mux_796_nl;
  wire[0:0] mux_795_nl;
  wire[0:0] or_615_nl;
  wire[0:0] mux_794_nl;
  wire[0:0] or_612_nl;
  wire[0:0] mux_793_nl;
  wire[0:0] mux_792_nl;
  wire[0:0] or_609_nl;
  wire[0:0] mux_791_nl;
  wire[0:0] or_606_nl;
  wire[0:0] mux_820_nl;
  wire[0:0] mux_819_nl;
  wire[0:0] or_649_nl;
  wire[0:0] mux_818_nl;
  wire[0:0] or_648_nl;
  wire[0:0] or_647_nl;
  wire[0:0] mux_817_nl;
  wire[0:0] mux_816_nl;
  wire[0:0] mux_815_nl;
  wire[0:0] or_645_nl;
  wire[0:0] mux_814_nl;
  wire[0:0] or_643_nl;
  wire[0:0] mux_813_nl;
  wire[0:0] mux_812_nl;
  wire[0:0] or_642_nl;
  wire[0:0] mux_811_nl;
  wire[0:0] or_640_nl;
  wire[0:0] or_639_nl;
  wire[0:0] mux_810_nl;
  wire[0:0] mux_809_nl;
  wire[0:0] mux_808_nl;
  wire[0:0] or_638_nl;
  wire[0:0] or_636_nl;
  wire[0:0] mux_807_nl;
  wire[0:0] or_634_nl;
  wire[0:0] or_633_nl;
  wire[0:0] nand_15_nl;
  wire[0:0] mux_806_nl;
  wire[0:0] nor_1412_nl;
  wire[0:0] nor_1413_nl;
  wire[0:0] mux_835_nl;
  wire[0:0] nand_468_nl;
  wire[0:0] mux_834_nl;
  wire[0:0] mux_833_nl;
  wire[0:0] mux_832_nl;
  wire[0:0] nor_1403_nl;
  wire[0:0] nor_1404_nl;
  wire[0:0] mux_831_nl;
  wire[0:0] nor_1405_nl;
  wire[0:0] nor_1406_nl;
  wire[0:0] mux_830_nl;
  wire[0:0] mux_829_nl;
  wire[0:0] nor_1407_nl;
  wire[0:0] nor_1408_nl;
  wire[0:0] mux_828_nl;
  wire[0:0] nor_1409_nl;
  wire[0:0] nor_1410_nl;
  wire[0:0] or_4141_nl;
  wire[0:0] mux_827_nl;
  wire[0:0] mux_826_nl;
  wire[0:0] mux_825_nl;
  wire[0:0] or_659_nl;
  wire[0:0] mux_824_nl;
  wire[0:0] or_656_nl;
  wire[0:0] mux_823_nl;
  wire[0:0] mux_822_nl;
  wire[0:0] or_653_nl;
  wire[0:0] mux_821_nl;
  wire[0:0] or_650_nl;
  wire[0:0] mux_850_nl;
  wire[0:0] mux_849_nl;
  wire[0:0] or_693_nl;
  wire[0:0] mux_848_nl;
  wire[0:0] or_692_nl;
  wire[0:0] or_691_nl;
  wire[0:0] mux_847_nl;
  wire[0:0] mux_846_nl;
  wire[0:0] mux_845_nl;
  wire[0:0] or_689_nl;
  wire[0:0] mux_844_nl;
  wire[0:0] or_687_nl;
  wire[0:0] mux_843_nl;
  wire[0:0] mux_842_nl;
  wire[0:0] or_686_nl;
  wire[0:0] mux_841_nl;
  wire[0:0] or_684_nl;
  wire[0:0] or_683_nl;
  wire[0:0] mux_840_nl;
  wire[0:0] mux_839_nl;
  wire[0:0] mux_838_nl;
  wire[0:0] or_682_nl;
  wire[0:0] or_680_nl;
  wire[0:0] mux_837_nl;
  wire[0:0] or_678_nl;
  wire[0:0] or_677_nl;
  wire[0:0] nand_17_nl;
  wire[0:0] mux_836_nl;
  wire[0:0] nor_1401_nl;
  wire[0:0] nor_1402_nl;
  wire[0:0] mux_865_nl;
  wire[0:0] nand_467_nl;
  wire[0:0] mux_864_nl;
  wire[0:0] mux_863_nl;
  wire[0:0] mux_862_nl;
  wire[0:0] nor_1392_nl;
  wire[0:0] nor_1393_nl;
  wire[0:0] mux_861_nl;
  wire[0:0] nor_1394_nl;
  wire[0:0] nor_1395_nl;
  wire[0:0] mux_860_nl;
  wire[0:0] mux_859_nl;
  wire[0:0] nor_1396_nl;
  wire[0:0] nor_1397_nl;
  wire[0:0] mux_858_nl;
  wire[0:0] nor_1398_nl;
  wire[0:0] nor_1399_nl;
  wire[0:0] or_4140_nl;
  wire[0:0] mux_857_nl;
  wire[0:0] mux_856_nl;
  wire[0:0] mux_855_nl;
  wire[0:0] or_703_nl;
  wire[0:0] mux_854_nl;
  wire[0:0] or_700_nl;
  wire[0:0] mux_853_nl;
  wire[0:0] mux_852_nl;
  wire[0:0] or_697_nl;
  wire[0:0] mux_851_nl;
  wire[0:0] or_694_nl;
  wire[0:0] mux_880_nl;
  wire[0:0] mux_879_nl;
  wire[0:0] or_737_nl;
  wire[0:0] mux_878_nl;
  wire[0:0] or_736_nl;
  wire[0:0] or_735_nl;
  wire[0:0] mux_877_nl;
  wire[0:0] mux_876_nl;
  wire[0:0] mux_875_nl;
  wire[0:0] or_733_nl;
  wire[0:0] mux_874_nl;
  wire[0:0] or_731_nl;
  wire[0:0] mux_873_nl;
  wire[0:0] mux_872_nl;
  wire[0:0] or_730_nl;
  wire[0:0] mux_871_nl;
  wire[0:0] or_728_nl;
  wire[0:0] or_727_nl;
  wire[0:0] mux_870_nl;
  wire[0:0] mux_869_nl;
  wire[0:0] mux_868_nl;
  wire[0:0] or_726_nl;
  wire[0:0] or_724_nl;
  wire[0:0] mux_867_nl;
  wire[0:0] or_722_nl;
  wire[0:0] or_721_nl;
  wire[0:0] nand_19_nl;
  wire[0:0] mux_866_nl;
  wire[0:0] nor_1390_nl;
  wire[0:0] nor_1391_nl;
  wire[0:0] mux_895_nl;
  wire[0:0] nand_466_nl;
  wire[0:0] mux_894_nl;
  wire[0:0] mux_893_nl;
  wire[0:0] mux_892_nl;
  wire[0:0] nor_1381_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] mux_891_nl;
  wire[0:0] nor_1383_nl;
  wire[0:0] nor_1384_nl;
  wire[0:0] mux_890_nl;
  wire[0:0] mux_889_nl;
  wire[0:0] nor_1385_nl;
  wire[0:0] nor_1386_nl;
  wire[0:0] mux_888_nl;
  wire[0:0] nor_1387_nl;
  wire[0:0] nor_1388_nl;
  wire[0:0] or_4139_nl;
  wire[0:0] mux_887_nl;
  wire[0:0] mux_886_nl;
  wire[0:0] mux_885_nl;
  wire[0:0] or_747_nl;
  wire[0:0] mux_884_nl;
  wire[0:0] or_744_nl;
  wire[0:0] mux_883_nl;
  wire[0:0] mux_882_nl;
  wire[0:0] or_741_nl;
  wire[0:0] mux_881_nl;
  wire[0:0] or_738_nl;
  wire[0:0] mux_910_nl;
  wire[0:0] mux_909_nl;
  wire[0:0] or_781_nl;
  wire[0:0] mux_908_nl;
  wire[0:0] or_780_nl;
  wire[0:0] or_779_nl;
  wire[0:0] mux_907_nl;
  wire[0:0] mux_906_nl;
  wire[0:0] mux_905_nl;
  wire[0:0] or_777_nl;
  wire[0:0] mux_904_nl;
  wire[0:0] or_775_nl;
  wire[0:0] mux_903_nl;
  wire[0:0] mux_902_nl;
  wire[0:0] or_774_nl;
  wire[0:0] mux_901_nl;
  wire[0:0] or_772_nl;
  wire[0:0] or_771_nl;
  wire[0:0] mux_900_nl;
  wire[0:0] mux_899_nl;
  wire[0:0] mux_898_nl;
  wire[0:0] or_770_nl;
  wire[0:0] or_768_nl;
  wire[0:0] mux_897_nl;
  wire[0:0] or_766_nl;
  wire[0:0] or_765_nl;
  wire[0:0] nand_21_nl;
  wire[0:0] mux_896_nl;
  wire[0:0] nor_1379_nl;
  wire[0:0] nor_1380_nl;
  wire[0:0] mux_925_nl;
  wire[0:0] nand_465_nl;
  wire[0:0] mux_924_nl;
  wire[0:0] mux_923_nl;
  wire[0:0] mux_922_nl;
  wire[0:0] nor_1370_nl;
  wire[0:0] nor_1371_nl;
  wire[0:0] mux_921_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] mux_920_nl;
  wire[0:0] mux_919_nl;
  wire[0:0] nor_1374_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] mux_918_nl;
  wire[0:0] nor_1376_nl;
  wire[0:0] nor_1377_nl;
  wire[0:0] or_4138_nl;
  wire[0:0] mux_917_nl;
  wire[0:0] mux_916_nl;
  wire[0:0] mux_915_nl;
  wire[0:0] or_791_nl;
  wire[0:0] mux_914_nl;
  wire[0:0] or_788_nl;
  wire[0:0] mux_913_nl;
  wire[0:0] mux_912_nl;
  wire[0:0] or_785_nl;
  wire[0:0] mux_911_nl;
  wire[0:0] or_782_nl;
  wire[0:0] mux_940_nl;
  wire[0:0] mux_939_nl;
  wire[0:0] or_825_nl;
  wire[0:0] mux_938_nl;
  wire[0:0] or_824_nl;
  wire[0:0] or_823_nl;
  wire[0:0] mux_937_nl;
  wire[0:0] mux_936_nl;
  wire[0:0] mux_935_nl;
  wire[0:0] or_821_nl;
  wire[0:0] mux_934_nl;
  wire[0:0] or_819_nl;
  wire[0:0] mux_933_nl;
  wire[0:0] mux_932_nl;
  wire[0:0] or_818_nl;
  wire[0:0] mux_931_nl;
  wire[0:0] or_816_nl;
  wire[0:0] or_815_nl;
  wire[0:0] mux_930_nl;
  wire[0:0] mux_929_nl;
  wire[0:0] mux_928_nl;
  wire[0:0] or_814_nl;
  wire[0:0] or_812_nl;
  wire[0:0] mux_927_nl;
  wire[0:0] or_810_nl;
  wire[0:0] or_809_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] mux_926_nl;
  wire[0:0] nor_1368_nl;
  wire[0:0] nor_1369_nl;
  wire[0:0] mux_955_nl;
  wire[0:0] nand_464_nl;
  wire[0:0] mux_954_nl;
  wire[0:0] mux_953_nl;
  wire[0:0] mux_952_nl;
  wire[0:0] nor_1359_nl;
  wire[0:0] nor_1360_nl;
  wire[0:0] mux_951_nl;
  wire[0:0] nor_1361_nl;
  wire[0:0] nor_1362_nl;
  wire[0:0] mux_950_nl;
  wire[0:0] mux_949_nl;
  wire[0:0] nor_1363_nl;
  wire[0:0] nor_1364_nl;
  wire[0:0] mux_948_nl;
  wire[0:0] nor_1365_nl;
  wire[0:0] nor_1366_nl;
  wire[0:0] or_4137_nl;
  wire[0:0] mux_947_nl;
  wire[0:0] mux_946_nl;
  wire[0:0] mux_945_nl;
  wire[0:0] or_835_nl;
  wire[0:0] mux_944_nl;
  wire[0:0] or_832_nl;
  wire[0:0] mux_943_nl;
  wire[0:0] mux_942_nl;
  wire[0:0] or_829_nl;
  wire[0:0] mux_941_nl;
  wire[0:0] or_826_nl;
  wire[0:0] mux_970_nl;
  wire[0:0] mux_969_nl;
  wire[0:0] or_869_nl;
  wire[0:0] mux_968_nl;
  wire[0:0] or_868_nl;
  wire[0:0] or_867_nl;
  wire[0:0] mux_967_nl;
  wire[0:0] mux_966_nl;
  wire[0:0] mux_965_nl;
  wire[0:0] or_865_nl;
  wire[0:0] mux_964_nl;
  wire[0:0] or_863_nl;
  wire[0:0] mux_963_nl;
  wire[0:0] mux_962_nl;
  wire[0:0] or_862_nl;
  wire[0:0] mux_961_nl;
  wire[0:0] or_860_nl;
  wire[0:0] or_859_nl;
  wire[0:0] mux_960_nl;
  wire[0:0] mux_959_nl;
  wire[0:0] mux_958_nl;
  wire[0:0] or_858_nl;
  wire[0:0] or_856_nl;
  wire[0:0] mux_957_nl;
  wire[0:0] or_854_nl;
  wire[0:0] or_853_nl;
  wire[0:0] nand_25_nl;
  wire[0:0] mux_956_nl;
  wire[0:0] nor_1357_nl;
  wire[0:0] nor_1358_nl;
  wire[0:0] mux_985_nl;
  wire[0:0] nand_463_nl;
  wire[0:0] mux_984_nl;
  wire[0:0] mux_983_nl;
  wire[0:0] mux_982_nl;
  wire[0:0] nor_1348_nl;
  wire[0:0] nor_1349_nl;
  wire[0:0] mux_981_nl;
  wire[0:0] nor_1350_nl;
  wire[0:0] nor_1351_nl;
  wire[0:0] mux_980_nl;
  wire[0:0] mux_979_nl;
  wire[0:0] nor_1352_nl;
  wire[0:0] nor_1353_nl;
  wire[0:0] mux_978_nl;
  wire[0:0] nor_1354_nl;
  wire[0:0] nor_1355_nl;
  wire[0:0] or_4136_nl;
  wire[0:0] mux_977_nl;
  wire[0:0] mux_976_nl;
  wire[0:0] mux_975_nl;
  wire[0:0] or_879_nl;
  wire[0:0] mux_974_nl;
  wire[0:0] or_876_nl;
  wire[0:0] mux_973_nl;
  wire[0:0] mux_972_nl;
  wire[0:0] or_873_nl;
  wire[0:0] mux_971_nl;
  wire[0:0] or_870_nl;
  wire[0:0] mux_1000_nl;
  wire[0:0] mux_999_nl;
  wire[0:0] or_913_nl;
  wire[0:0] mux_998_nl;
  wire[0:0] or_912_nl;
  wire[0:0] or_911_nl;
  wire[0:0] mux_997_nl;
  wire[0:0] mux_996_nl;
  wire[0:0] mux_995_nl;
  wire[0:0] or_909_nl;
  wire[0:0] mux_994_nl;
  wire[0:0] or_907_nl;
  wire[0:0] mux_993_nl;
  wire[0:0] mux_992_nl;
  wire[0:0] or_906_nl;
  wire[0:0] mux_991_nl;
  wire[0:0] or_904_nl;
  wire[0:0] or_903_nl;
  wire[0:0] mux_990_nl;
  wire[0:0] mux_989_nl;
  wire[0:0] mux_988_nl;
  wire[0:0] or_902_nl;
  wire[0:0] or_900_nl;
  wire[0:0] mux_987_nl;
  wire[0:0] or_898_nl;
  wire[0:0] or_897_nl;
  wire[0:0] nand_27_nl;
  wire[0:0] mux_986_nl;
  wire[0:0] nor_1346_nl;
  wire[0:0] nor_1347_nl;
  wire[0:0] mux_1015_nl;
  wire[0:0] nand_462_nl;
  wire[0:0] mux_1014_nl;
  wire[0:0] mux_1013_nl;
  wire[0:0] mux_1012_nl;
  wire[0:0] nor_1337_nl;
  wire[0:0] nor_1338_nl;
  wire[0:0] mux_1011_nl;
  wire[0:0] nor_1339_nl;
  wire[0:0] nor_1340_nl;
  wire[0:0] mux_1010_nl;
  wire[0:0] mux_1009_nl;
  wire[0:0] nor_1341_nl;
  wire[0:0] nor_1342_nl;
  wire[0:0] mux_1008_nl;
  wire[0:0] nor_1343_nl;
  wire[0:0] nor_1344_nl;
  wire[0:0] or_4135_nl;
  wire[0:0] mux_1007_nl;
  wire[0:0] mux_1006_nl;
  wire[0:0] mux_1005_nl;
  wire[0:0] or_923_nl;
  wire[0:0] mux_1004_nl;
  wire[0:0] or_920_nl;
  wire[0:0] mux_1003_nl;
  wire[0:0] mux_1002_nl;
  wire[0:0] or_917_nl;
  wire[0:0] mux_1001_nl;
  wire[0:0] or_914_nl;
  wire[0:0] mux_1030_nl;
  wire[0:0] mux_1029_nl;
  wire[0:0] or_957_nl;
  wire[0:0] mux_1028_nl;
  wire[0:0] or_956_nl;
  wire[0:0] or_955_nl;
  wire[0:0] mux_1027_nl;
  wire[0:0] mux_1026_nl;
  wire[0:0] mux_1025_nl;
  wire[0:0] or_953_nl;
  wire[0:0] mux_1024_nl;
  wire[0:0] or_951_nl;
  wire[0:0] mux_1023_nl;
  wire[0:0] mux_1022_nl;
  wire[0:0] or_950_nl;
  wire[0:0] mux_1021_nl;
  wire[0:0] or_948_nl;
  wire[0:0] or_947_nl;
  wire[0:0] mux_1020_nl;
  wire[0:0] mux_1019_nl;
  wire[0:0] mux_1018_nl;
  wire[0:0] or_946_nl;
  wire[0:0] or_944_nl;
  wire[0:0] mux_1017_nl;
  wire[0:0] or_942_nl;
  wire[0:0] or_941_nl;
  wire[0:0] nand_29_nl;
  wire[0:0] mux_1016_nl;
  wire[0:0] nor_1335_nl;
  wire[0:0] nor_1336_nl;
  wire[0:0] mux_1045_nl;
  wire[0:0] nand_461_nl;
  wire[0:0] mux_1044_nl;
  wire[0:0] mux_1043_nl;
  wire[0:0] mux_1042_nl;
  wire[0:0] nor_1326_nl;
  wire[0:0] nor_1327_nl;
  wire[0:0] mux_1041_nl;
  wire[0:0] nor_1328_nl;
  wire[0:0] nor_1329_nl;
  wire[0:0] mux_1040_nl;
  wire[0:0] mux_1039_nl;
  wire[0:0] nor_1330_nl;
  wire[0:0] nor_1331_nl;
  wire[0:0] mux_1038_nl;
  wire[0:0] nor_1332_nl;
  wire[0:0] nor_1333_nl;
  wire[0:0] or_4134_nl;
  wire[0:0] mux_1037_nl;
  wire[0:0] mux_1036_nl;
  wire[0:0] mux_1035_nl;
  wire[0:0] or_967_nl;
  wire[0:0] mux_1034_nl;
  wire[0:0] or_964_nl;
  wire[0:0] mux_1033_nl;
  wire[0:0] mux_1032_nl;
  wire[0:0] or_961_nl;
  wire[0:0] mux_1031_nl;
  wire[0:0] or_958_nl;
  wire[0:0] mux_1060_nl;
  wire[0:0] mux_1059_nl;
  wire[0:0] or_1001_nl;
  wire[0:0] mux_1058_nl;
  wire[0:0] or_1000_nl;
  wire[0:0] or_999_nl;
  wire[0:0] mux_1057_nl;
  wire[0:0] mux_1056_nl;
  wire[0:0] mux_1055_nl;
  wire[0:0] or_997_nl;
  wire[0:0] mux_1054_nl;
  wire[0:0] or_995_nl;
  wire[0:0] mux_1053_nl;
  wire[0:0] mux_1052_nl;
  wire[0:0] or_994_nl;
  wire[0:0] mux_1051_nl;
  wire[0:0] or_992_nl;
  wire[0:0] or_991_nl;
  wire[0:0] mux_1050_nl;
  wire[0:0] mux_1049_nl;
  wire[0:0] mux_1048_nl;
  wire[0:0] or_990_nl;
  wire[0:0] or_988_nl;
  wire[0:0] mux_1047_nl;
  wire[0:0] or_986_nl;
  wire[0:0] or_985_nl;
  wire[0:0] nand_31_nl;
  wire[0:0] mux_1046_nl;
  wire[0:0] nor_1324_nl;
  wire[0:0] nor_1325_nl;
  wire[0:0] mux_1075_nl;
  wire[0:0] nand_460_nl;
  wire[0:0] mux_1074_nl;
  wire[0:0] mux_1073_nl;
  wire[0:0] mux_1072_nl;
  wire[0:0] nor_1315_nl;
  wire[0:0] nor_1316_nl;
  wire[0:0] mux_1071_nl;
  wire[0:0] nor_1317_nl;
  wire[0:0] nor_1318_nl;
  wire[0:0] mux_1070_nl;
  wire[0:0] mux_1069_nl;
  wire[0:0] nor_1319_nl;
  wire[0:0] nor_1320_nl;
  wire[0:0] mux_1068_nl;
  wire[0:0] nor_1321_nl;
  wire[0:0] nor_1322_nl;
  wire[0:0] or_4133_nl;
  wire[0:0] mux_1067_nl;
  wire[0:0] mux_1066_nl;
  wire[0:0] mux_1065_nl;
  wire[0:0] or_1011_nl;
  wire[0:0] mux_1064_nl;
  wire[0:0] or_1008_nl;
  wire[0:0] mux_1063_nl;
  wire[0:0] mux_1062_nl;
  wire[0:0] or_1005_nl;
  wire[0:0] mux_1061_nl;
  wire[0:0] or_1002_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] or_1045_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] or_1043_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] or_1041_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] or_1039_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] mux_1082_nl;
  wire[0:0] or_1038_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] or_1036_nl;
  wire[0:0] or_1035_nl;
  wire[0:0] mux_1080_nl;
  wire[0:0] mux_1079_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] or_1034_nl;
  wire[0:0] or_1032_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] or_1030_nl;
  wire[0:0] or_1029_nl;
  wire[0:0] nand_33_nl;
  wire[0:0] mux_1076_nl;
  wire[0:0] nor_1313_nl;
  wire[0:0] nor_1314_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] nand_459_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] nor_1304_nl;
  wire[0:0] nor_1305_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] nor_1306_nl;
  wire[0:0] nor_1307_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] nor_1308_nl;
  wire[0:0] nor_1309_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] nor_1310_nl;
  wire[0:0] nor_1311_nl;
  wire[0:0] or_4132_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] or_1055_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] or_1052_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] or_1049_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] or_1046_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_1089_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] or_1088_nl;
  wire[0:0] or_1087_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] mux_1116_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] or_1085_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] or_1083_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] or_1082_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] or_1080_nl;
  wire[0:0] or_1079_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] or_1078_nl;
  wire[0:0] or_1076_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] or_1074_nl;
  wire[0:0] or_1073_nl;
  wire[0:0] nand_35_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] nor_1302_nl;
  wire[0:0] nor_1303_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] nand_458_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_1293_nl;
  wire[0:0] nor_1294_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] nor_1295_nl;
  wire[0:0] nor_1296_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] nor_1297_nl;
  wire[0:0] nor_1298_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] nor_1299_nl;
  wire[0:0] nor_1300_nl;
  wire[0:0] or_4131_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] or_1099_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] or_1096_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] or_1093_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] or_1090_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] mux_1149_nl;
  wire[0:0] or_1133_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] or_1132_nl;
  wire[0:0] or_1131_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] or_1127_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] or_1126_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] or_1124_nl;
  wire[0:0] or_1123_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] mux_1139_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] or_1122_nl;
  wire[0:0] or_1120_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] or_1118_nl;
  wire[0:0] or_1117_nl;
  wire[0:0] nand_37_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] nor_1291_nl;
  wire[0:0] nor_1292_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] nand_457_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] nor_1282_nl;
  wire[0:0] nor_1283_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] nor_1284_nl;
  wire[0:0] nor_1285_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] nor_1286_nl;
  wire[0:0] nor_1287_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] nor_1288_nl;
  wire[0:0] nor_1289_nl;
  wire[0:0] or_4130_nl;
  wire[0:0] mux_1157_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] or_1143_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] or_1140_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] or_1137_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] or_1134_nl;
  wire[0:0] mux_1180_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] or_1177_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] or_1176_nl;
  wire[0:0] or_1175_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] or_1173_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] or_1171_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] mux_1172_nl;
  wire[0:0] or_1170_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] or_1168_nl;
  wire[0:0] or_1167_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] or_1166_nl;
  wire[0:0] or_1164_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] or_1162_nl;
  wire[0:0] or_1161_nl;
  wire[0:0] nand_39_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] nor_1281_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] nand_456_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] nor_1271_nl;
  wire[0:0] nor_1272_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] nor_1273_nl;
  wire[0:0] nor_1274_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] nor_1275_nl;
  wire[0:0] nor_1276_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] nor_1277_nl;
  wire[0:0] nor_1278_nl;
  wire[0:0] or_4129_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] or_1187_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] or_1184_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] or_1181_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] or_1178_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] or_1221_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] or_1220_nl;
  wire[0:0] or_1219_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] or_1217_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] or_1215_nl;
  wire[0:0] mux_1203_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] or_1214_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] or_1212_nl;
  wire[0:0] or_1211_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] or_1210_nl;
  wire[0:0] or_1208_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] or_1206_nl;
  wire[0:0] or_1205_nl;
  wire[0:0] nand_41_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] nor_1269_nl;
  wire[0:0] nor_1270_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] nand_455_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] nor_1260_nl;
  wire[0:0] nor_1261_nl;
  wire[0:0] mux_1221_nl;
  wire[0:0] nor_1262_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] nor_1264_nl;
  wire[0:0] nor_1265_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] nor_1267_nl;
  wire[0:0] or_4128_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] or_1231_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] or_1228_nl;
  wire[0:0] mux_1213_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] or_1225_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] or_1222_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] or_1265_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] or_1264_nl;
  wire[0:0] or_1263_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] mux_1236_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] or_1261_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] or_1259_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] or_1258_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] or_1256_nl;
  wire[0:0] or_1255_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] or_1254_nl;
  wire[0:0] or_1252_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] or_1250_nl;
  wire[0:0] or_1249_nl;
  wire[0:0] nand_43_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] nor_1258_nl;
  wire[0:0] nor_1259_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] nand_454_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] and_618_nl;
  wire[0:0] nor_1250_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] nor_1251_nl;
  wire[0:0] nor_1252_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] nor_1255_nl;
  wire[0:0] nor_1256_nl;
  wire[0:0] or_4127_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] nand_332_nl;
  wire[0:0] mux_1244_nl;
  wire[0:0] or_1272_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] or_1269_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] or_1266_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] or_1309_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] or_1308_nl;
  wire[0:0] or_1307_nl;
  wire[0:0] mux_1267_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] nand_330_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] or_1303_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] or_1302_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] or_1300_nl;
  wire[0:0] or_1299_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] or_1298_nl;
  wire[0:0] nand_331_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] or_1294_nl;
  wire[0:0] or_1293_nl;
  wire[0:0] nand_45_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] nor_1249_nl;
  wire[0:0] mux_1285_nl;
  wire[0:0] nand_453_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] nor_1239_nl;
  wire[0:0] nor_1240_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] nor_1242_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] nor_1243_nl;
  wire[0:0] nor_1244_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] nor_1245_nl;
  wire[0:0] nor_1246_nl;
  wire[0:0] or_4126_nl;
  wire[0:0] mux_1277_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] or_1319_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] or_1316_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] or_1313_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] or_1310_nl;
  wire[0:0] mux_1300_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] or_1353_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] or_1352_nl;
  wire[0:0] or_1351_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] or_1349_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] or_1347_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] or_1346_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] or_1344_nl;
  wire[0:0] or_1343_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] or_1342_nl;
  wire[0:0] or_1340_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] or_1338_nl;
  wire[0:0] or_1337_nl;
  wire[0:0] nand_47_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] nor_1237_nl;
  wire[0:0] nor_1238_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] nand_452_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] nor_1228_nl;
  wire[0:0] nor_1229_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] nor_1230_nl;
  wire[0:0] nor_1231_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] nor_1232_nl;
  wire[0:0] nor_1233_nl;
  wire[0:0] mux_1308_nl;
  wire[0:0] nor_1234_nl;
  wire[0:0] nor_1235_nl;
  wire[0:0] or_4125_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] or_1363_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] or_1360_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] or_1357_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] or_1354_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] or_1397_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] or_1396_nl;
  wire[0:0] or_1395_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] or_1393_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] or_1391_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] or_1390_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] or_1388_nl;
  wire[0:0] or_1387_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] or_1386_nl;
  wire[0:0] or_1384_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] or_1382_nl;
  wire[0:0] or_1381_nl;
  wire[0:0] nand_49_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] nor_1226_nl;
  wire[0:0] nor_1227_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] nand_451_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] nor_1217_nl;
  wire[0:0] nor_1218_nl;
  wire[0:0] mux_1341_nl;
  wire[0:0] nor_1219_nl;
  wire[0:0] nor_1220_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] nor_1221_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] nor_1223_nl;
  wire[0:0] nor_1224_nl;
  wire[0:0] or_4124_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] or_1407_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] or_1404_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] or_1401_nl;
  wire[0:0] mux_1331_nl;
  wire[0:0] or_1398_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] or_1441_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] or_1440_nl;
  wire[0:0] or_1439_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] or_1437_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] or_1435_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] or_1434_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] or_1432_nl;
  wire[0:0] or_1431_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] mux_1349_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] or_1430_nl;
  wire[0:0] or_1428_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] or_1426_nl;
  wire[0:0] or_1425_nl;
  wire[0:0] nand_51_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] nor_1215_nl;
  wire[0:0] nor_1216_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] nand_450_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] mux_1372_nl;
  wire[0:0] nor_1206_nl;
  wire[0:0] nor_1207_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] nor_1208_nl;
  wire[0:0] nor_1209_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] nor_1210_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] nor_1212_nl;
  wire[0:0] nor_1213_nl;
  wire[0:0] or_4123_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] or_1451_nl;
  wire[0:0] mux_1364_nl;
  wire[0:0] or_1448_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] or_1445_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] or_1442_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] or_1485_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] or_1484_nl;
  wire[0:0] or_1483_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] or_1481_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] or_1479_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] or_1478_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] or_1476_nl;
  wire[0:0] or_1475_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] or_1474_nl;
  wire[0:0] or_1472_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] or_1470_nl;
  wire[0:0] or_1469_nl;
  wire[0:0] nand_53_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] nor_1204_nl;
  wire[0:0] nor_1205_nl;
  wire[0:0] mux_1405_nl;
  wire[0:0] nand_449_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] nor_1195_nl;
  wire[0:0] nor_1196_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] nor_1200_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] nor_1202_nl;
  wire[0:0] or_4122_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] mux_1395_nl;
  wire[0:0] or_1495_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] or_1492_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] or_1489_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] or_1486_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] or_1529_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] or_1528_nl;
  wire[0:0] or_1527_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] or_1525_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] or_1523_nl;
  wire[0:0] mux_1413_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] or_1522_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] or_1520_nl;
  wire[0:0] or_1519_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] or_1518_nl;
  wire[0:0] or_1516_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] or_1514_nl;
  wire[0:0] or_1513_nl;
  wire[0:0] nand_55_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] nor_1193_nl;
  wire[0:0] nor_1194_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] nand_448_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] nor_1184_nl;
  wire[0:0] nor_1185_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] nor_1186_nl;
  wire[0:0] nor_1187_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] nor_1188_nl;
  wire[0:0] nor_1189_nl;
  wire[0:0] mux_1428_nl;
  wire[0:0] nor_1190_nl;
  wire[0:0] nor_1191_nl;
  wire[0:0] or_4121_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] or_1539_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] or_1536_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] or_1533_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] or_1530_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] or_1573_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] or_1572_nl;
  wire[0:0] or_1571_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] or_1569_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] or_1567_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] or_1566_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] or_1564_nl;
  wire[0:0] or_1563_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] or_1562_nl;
  wire[0:0] or_1560_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] or_1558_nl;
  wire[0:0] or_1557_nl;
  wire[0:0] nand_57_nl;
  wire[0:0] mux_1436_nl;
  wire[0:0] nor_1182_nl;
  wire[0:0] nor_1183_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] nand_447_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] nor_1173_nl;
  wire[0:0] nor_1174_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] nor_1175_nl;
  wire[0:0] nor_1176_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] mux_1459_nl;
  wire[0:0] nor_1177_nl;
  wire[0:0] nor_1178_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] nor_1180_nl;
  wire[0:0] or_4120_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] or_1583_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] or_1580_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] or_1577_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] or_1574_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] or_1617_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] or_1616_nl;
  wire[0:0] or_1615_nl;
  wire[0:0] mux_1477_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] or_1613_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] or_1611_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] or_1610_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] or_1608_nl;
  wire[0:0] or_1607_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] mux_1469_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] or_1606_nl;
  wire[0:0] or_1604_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] or_1602_nl;
  wire[0:0] or_1601_nl;
  wire[0:0] nand_59_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] nor_1171_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] nand_446_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] mux_1492_nl;
  wire[0:0] nor_1162_nl;
  wire[0:0] nor_1163_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] nor_1164_nl;
  wire[0:0] nor_1165_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] nor_1166_nl;
  wire[0:0] nor_1167_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] nor_1168_nl;
  wire[0:0] nor_1169_nl;
  wire[0:0] or_4119_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] nand_326_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] or_1624_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] or_1621_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] or_1618_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] or_1661_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] or_1660_nl;
  wire[0:0] or_1659_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] nand_325_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] or_1655_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] or_1654_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] or_1652_nl;
  wire[0:0] or_1651_nl;
  wire[0:0] mux_1500_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] or_1650_nl;
  wire[0:0] or_1648_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] or_1646_nl;
  wire[0:0] or_1645_nl;
  wire[0:0] nand_61_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] nor_1161_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] nand_445_nl;
  wire[0:0] mux_1524_nl;
  wire[0:0] mux_1523_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] nor_1151_nl;
  wire[0:0] nor_1152_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] nor_1154_nl;
  wire[0:0] mux_1520_nl;
  wire[0:0] mux_1519_nl;
  wire[0:0] nor_1155_nl;
  wire[0:0] nor_1156_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] nor_1158_nl;
  wire[0:0] or_4118_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] or_1671_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] or_1668_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] or_1665_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] or_1662_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] or_1705_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] or_1704_nl;
  wire[0:0] or_1703_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] or_1701_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] or_1699_nl;
  wire[0:0] mux_1533_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] or_1698_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] or_1696_nl;
  wire[0:0] or_1695_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] or_1694_nl;
  wire[0:0] or_1692_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] or_1690_nl;
  wire[0:0] or_1689_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] nor_1149_nl;
  wire[0:0] nor_1150_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] nand_444_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] nor_1140_nl;
  wire[0:0] nor_1141_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] nor_1142_nl;
  wire[0:0] nor_1143_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] nor_1144_nl;
  wire[0:0] nor_1145_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] nor_1146_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] or_4117_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] or_1715_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] or_1712_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] or_1709_nl;
  wire[0:0] mux_1541_nl;
  wire[0:0] or_1706_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] or_1749_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] or_1748_nl;
  wire[0:0] or_1747_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] mux_1566_nl;
  wire[0:0] mux_1565_nl;
  wire[0:0] or_1745_nl;
  wire[0:0] mux_1564_nl;
  wire[0:0] or_1743_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] or_1742_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] or_1740_nl;
  wire[0:0] or_1739_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] or_1738_nl;
  wire[0:0] or_1736_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] or_1734_nl;
  wire[0:0] or_1733_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_1556_nl;
  wire[0:0] nor_1138_nl;
  wire[0:0] nor_1139_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] nand_443_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] nor_1130_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] nor_1131_nl;
  wire[0:0] nor_1132_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] nor_1134_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] nor_1135_nl;
  wire[0:0] nor_1136_nl;
  wire[0:0] or_4116_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] or_1759_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] or_1756_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] or_1753_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] or_1750_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] or_1793_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] or_1792_nl;
  wire[0:0] or_1791_nl;
  wire[0:0] mux_1597_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] or_1789_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] or_1787_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] or_1786_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] or_1784_nl;
  wire[0:0] or_1783_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] or_1782_nl;
  wire[0:0] or_1780_nl;
  wire[0:0] mux_1587_nl;
  wire[0:0] or_1778_nl;
  wire[0:0] or_1777_nl;
  wire[0:0] nand_67_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] nor_1127_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] nand_442_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] nor_1118_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] nor_1120_nl;
  wire[0:0] nor_1121_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] nor_1123_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] nor_1124_nl;
  wire[0:0] nor_1125_nl;
  wire[0:0] or_4115_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] mux_1605_nl;
  wire[0:0] nand_324_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] or_1800_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] or_1797_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] or_1794_nl;
  wire[0:0] mux_1630_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] or_1837_nl;
  wire[0:0] mux_1628_nl;
  wire[0:0] or_1836_nl;
  wire[0:0] or_1835_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] nand_323_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] or_1831_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] or_1828_nl;
  wire[0:0] or_1827_nl;
  wire[0:0] mux_1620_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] or_1826_nl;
  wire[0:0] or_1824_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] or_1822_nl;
  wire[0:0] or_1821_nl;
  wire[0:0] nand_69_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] nor_1116_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] nand_441_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] nor_1107_nl;
  wire[0:0] nor_1108_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] nor_1109_nl;
  wire[0:0] nor_1110_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] nor_1111_nl;
  wire[0:0] nor_1112_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] nor_1113_nl;
  wire[0:0] nor_1114_nl;
  wire[0:0] or_4114_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] or_1847_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] or_1844_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] or_1841_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] or_1838_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] mux_1659_nl;
  wire[0:0] or_1881_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] or_1880_nl;
  wire[0:0] or_1879_nl;
  wire[0:0] mux_1657_nl;
  wire[0:0] mux_1656_nl;
  wire[0:0] mux_1655_nl;
  wire[0:0] or_1877_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] or_1875_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] or_1874_nl;
  wire[0:0] mux_1651_nl;
  wire[0:0] or_1872_nl;
  wire[0:0] or_1871_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] or_1870_nl;
  wire[0:0] or_1868_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] or_1866_nl;
  wire[0:0] or_1865_nl;
  wire[0:0] nand_71_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] nor_1105_nl;
  wire[0:0] nor_1106_nl;
  wire[0:0] mux_1675_nl;
  wire[0:0] nand_440_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] mux_1672_nl;
  wire[0:0] nor_1096_nl;
  wire[0:0] nor_1097_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] nor_1098_nl;
  wire[0:0] nor_1099_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] mux_1669_nl;
  wire[0:0] nor_1100_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] mux_1668_nl;
  wire[0:0] nor_1102_nl;
  wire[0:0] nor_1103_nl;
  wire[0:0] or_4113_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] mux_1666_nl;
  wire[0:0] mux_1665_nl;
  wire[0:0] nand_322_nl;
  wire[0:0] mux_1664_nl;
  wire[0:0] or_1888_nl;
  wire[0:0] mux_1663_nl;
  wire[0:0] mux_1662_nl;
  wire[0:0] or_1885_nl;
  wire[0:0] mux_1661_nl;
  wire[0:0] or_1882_nl;
  wire[0:0] mux_1690_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] or_1925_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] or_1924_nl;
  wire[0:0] or_1923_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] nand_321_nl;
  wire[0:0] mux_1684_nl;
  wire[0:0] or_1919_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] mux_1682_nl;
  wire[0:0] or_1918_nl;
  wire[0:0] mux_1681_nl;
  wire[0:0] or_1916_nl;
  wire[0:0] or_1915_nl;
  wire[0:0] mux_1680_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] mux_1678_nl;
  wire[0:0] or_1914_nl;
  wire[0:0] or_1912_nl;
  wire[0:0] mux_1677_nl;
  wire[0:0] or_1910_nl;
  wire[0:0] or_1909_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] mux_1676_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] nor_1095_nl;
  wire[0:0] mux_1705_nl;
  wire[0:0] nand_439_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] mux_1702_nl;
  wire[0:0] nor_1086_nl;
  wire[0:0] and_602_nl;
  wire[0:0] mux_1701_nl;
  wire[0:0] nor_1087_nl;
  wire[0:0] nor_1088_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] nor_1089_nl;
  wire[0:0] nor_1090_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] nor_1091_nl;
  wire[0:0] nor_1092_nl;
  wire[0:0] or_4112_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] nand_320_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] or_1932_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] mux_1692_nl;
  wire[0:0] or_1929_nl;
  wire[0:0] mux_1691_nl;
  wire[0:0] or_1926_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] or_1969_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] or_1968_nl;
  wire[0:0] or_1967_nl;
  wire[0:0] mux_1717_nl;
  wire[0:0] mux_1716_nl;
  wire[0:0] mux_1715_nl;
  wire[0:0] nand_318_nl;
  wire[0:0] mux_1714_nl;
  wire[0:0] or_1963_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] mux_1712_nl;
  wire[0:0] or_1962_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] or_1960_nl;
  wire[0:0] or_1959_nl;
  wire[0:0] mux_1710_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] nand_319_nl;
  wire[0:0] or_1956_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] or_1954_nl;
  wire[0:0] or_1953_nl;
  wire[0:0] nand_75_nl;
  wire[0:0] mux_1706_nl;
  wire[0:0] nor_1084_nl;
  wire[0:0] nor_1085_nl;
  wire[0:0] mux_1735_nl;
  wire[0:0] nand_438_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] mux_1733_nl;
  wire[0:0] mux_1732_nl;
  wire[0:0] nor_1077_nl;
  wire[0:0] nor_1078_nl;
  wire[0:0] mux_1731_nl;
  wire[0:0] and_599_nl;
  wire[0:0] and_600_nl;
  wire[0:0] mux_1730_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] and_811_nl;
  wire[0:0] and_818_nl;
  wire[0:0] mux_1728_nl;
  wire[0:0] nor_1081_nl;
  wire[0:0] nor_1082_nl;
  wire[0:0] or_4111_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] mux_1726_nl;
  wire[0:0] mux_1725_nl;
  wire[0:0] nand_313_nl;
  wire[0:0] mux_1724_nl;
  wire[0:0] nand_314_nl;
  wire[0:0] mux_1723_nl;
  wire[0:0] mux_1722_nl;
  wire[0:0] nand_478_nl;
  wire[0:0] mux_1721_nl;
  wire[0:0] or_1970_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] or_2012_nl;
  wire[0:0] mux_1748_nl;
  wire[0:0] or_2011_nl;
  wire[0:0] or_2010_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] mux_1745_nl;
  wire[0:0] nand_302_nl;
  wire[0:0] mux_1744_nl;
  wire[0:0] nand_303_nl;
  wire[0:0] mux_1743_nl;
  wire[0:0] mux_1742_nl;
  wire[0:0] nand_404_nl;
  wire[0:0] mux_1741_nl;
  wire[0:0] or_2003_nl;
  wire[0:0] or_2002_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] mux_1739_nl;
  wire[0:0] mux_1738_nl;
  wire[0:0] or_2001_nl;
  wire[0:0] or_1999_nl;
  wire[0:0] mux_1737_nl;
  wire[0:0] nand_307_nl;
  wire[0:0] nand_308_nl;
  wire[0:0] nand_77_nl;
  wire[0:0] mux_1736_nl;
  wire[0:0] nor_1075_nl;
  wire[0:0] nor_1076_nl;
  wire[0:0] mux_1765_nl;
  wire[0:0] nand_437_nl;
  wire[0:0] mux_1764_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] nor_1066_nl;
  wire[0:0] nor_1067_nl;
  wire[0:0] mux_1761_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] nor_1069_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] mux_1759_nl;
  wire[0:0] nor_1070_nl;
  wire[0:0] nor_1071_nl;
  wire[0:0] mux_1758_nl;
  wire[0:0] nor_1072_nl;
  wire[0:0] nor_1073_nl;
  wire[0:0] or_4110_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] mux_1756_nl;
  wire[0:0] mux_1755_nl;
  wire[0:0] or_2022_nl;
  wire[0:0] mux_1754_nl;
  wire[0:0] or_2019_nl;
  wire[0:0] mux_1753_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] or_2016_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] or_2013_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] mux_1779_nl;
  wire[0:0] or_2056_nl;
  wire[0:0] mux_1778_nl;
  wire[0:0] or_2055_nl;
  wire[0:0] or_2054_nl;
  wire[0:0] mux_1777_nl;
  wire[0:0] mux_1776_nl;
  wire[0:0] mux_1775_nl;
  wire[0:0] or_2052_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] or_2050_nl;
  wire[0:0] mux_1773_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] or_2049_nl;
  wire[0:0] mux_1771_nl;
  wire[0:0] or_2047_nl;
  wire[0:0] or_2046_nl;
  wire[0:0] mux_1770_nl;
  wire[0:0] mux_1769_nl;
  wire[0:0] mux_1768_nl;
  wire[0:0] or_2045_nl;
  wire[0:0] or_2043_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] or_2041_nl;
  wire[0:0] or_2040_nl;
  wire[0:0] nand_79_nl;
  wire[0:0] mux_1766_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] nor_1065_nl;
  wire[0:0] mux_1795_nl;
  wire[0:0] nand_436_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] mux_1793_nl;
  wire[0:0] mux_1792_nl;
  wire[0:0] nor_1055_nl;
  wire[0:0] nor_1056_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] nor_1057_nl;
  wire[0:0] nor_1058_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] mux_1789_nl;
  wire[0:0] nor_1059_nl;
  wire[0:0] nor_1060_nl;
  wire[0:0] mux_1788_nl;
  wire[0:0] nor_1061_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] or_4109_nl;
  wire[0:0] mux_1787_nl;
  wire[0:0] mux_1786_nl;
  wire[0:0] mux_1785_nl;
  wire[0:0] or_2066_nl;
  wire[0:0] mux_1784_nl;
  wire[0:0] or_2063_nl;
  wire[0:0] mux_1783_nl;
  wire[0:0] mux_1782_nl;
  wire[0:0] or_2060_nl;
  wire[0:0] mux_1781_nl;
  wire[0:0] or_2057_nl;
  wire[0:0] mux_1810_nl;
  wire[0:0] mux_1809_nl;
  wire[0:0] or_2100_nl;
  wire[0:0] mux_1808_nl;
  wire[0:0] or_2099_nl;
  wire[0:0] or_2098_nl;
  wire[0:0] mux_1807_nl;
  wire[0:0] mux_1806_nl;
  wire[0:0] mux_1805_nl;
  wire[0:0] or_2096_nl;
  wire[0:0] mux_1804_nl;
  wire[0:0] or_2094_nl;
  wire[0:0] mux_1803_nl;
  wire[0:0] mux_1802_nl;
  wire[0:0] or_2093_nl;
  wire[0:0] mux_1801_nl;
  wire[0:0] or_2091_nl;
  wire[0:0] or_2090_nl;
  wire[0:0] mux_1800_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] or_2089_nl;
  wire[0:0] or_2087_nl;
  wire[0:0] mux_1797_nl;
  wire[0:0] or_2085_nl;
  wire[0:0] or_2084_nl;
  wire[0:0] nand_81_nl;
  wire[0:0] mux_1796_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] nor_1054_nl;
  wire[0:0] mux_1825_nl;
  wire[0:0] nand_435_nl;
  wire[0:0] mux_1824_nl;
  wire[0:0] mux_1823_nl;
  wire[0:0] mux_1822_nl;
  wire[0:0] nor_1044_nl;
  wire[0:0] nor_1045_nl;
  wire[0:0] mux_1821_nl;
  wire[0:0] nor_1046_nl;
  wire[0:0] nor_1047_nl;
  wire[0:0] mux_1820_nl;
  wire[0:0] mux_1819_nl;
  wire[0:0] nor_1048_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] mux_1818_nl;
  wire[0:0] nor_1050_nl;
  wire[0:0] nor_1051_nl;
  wire[0:0] or_4108_nl;
  wire[0:0] mux_1817_nl;
  wire[0:0] mux_1816_nl;
  wire[0:0] mux_1815_nl;
  wire[0:0] or_2110_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] or_2107_nl;
  wire[0:0] mux_1813_nl;
  wire[0:0] mux_1812_nl;
  wire[0:0] or_2104_nl;
  wire[0:0] mux_1811_nl;
  wire[0:0] or_2101_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] mux_1839_nl;
  wire[0:0] or_2144_nl;
  wire[0:0] mux_1838_nl;
  wire[0:0] or_2143_nl;
  wire[0:0] or_2142_nl;
  wire[0:0] mux_1837_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] or_2140_nl;
  wire[0:0] mux_1834_nl;
  wire[0:0] or_2138_nl;
  wire[0:0] mux_1833_nl;
  wire[0:0] mux_1832_nl;
  wire[0:0] or_2137_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] or_2135_nl;
  wire[0:0] or_2134_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] or_2133_nl;
  wire[0:0] or_2131_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] or_2129_nl;
  wire[0:0] or_2128_nl;
  wire[0:0] nand_83_nl;
  wire[0:0] mux_1826_nl;
  wire[0:0] nor_1042_nl;
  wire[0:0] nor_1043_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] nand_434_nl;
  wire[0:0] mux_1854_nl;
  wire[0:0] mux_1853_nl;
  wire[0:0] mux_1852_nl;
  wire[0:0] nor_1033_nl;
  wire[0:0] nor_1034_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] nor_1036_nl;
  wire[0:0] mux_1850_nl;
  wire[0:0] mux_1849_nl;
  wire[0:0] nor_1037_nl;
  wire[0:0] nor_1038_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] nor_1039_nl;
  wire[0:0] nor_1040_nl;
  wire[0:0] or_4107_nl;
  wire[0:0] mux_1847_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] or_2154_nl;
  wire[0:0] mux_1844_nl;
  wire[0:0] or_2151_nl;
  wire[0:0] mux_1843_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] or_2148_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] or_2145_nl;
  wire[0:0] mux_1870_nl;
  wire[0:0] mux_1869_nl;
  wire[0:0] or_2188_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] or_2187_nl;
  wire[0:0] or_2186_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] mux_1866_nl;
  wire[0:0] mux_1865_nl;
  wire[0:0] or_2184_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] or_2182_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] or_2181_nl;
  wire[0:0] mux_1861_nl;
  wire[0:0] or_2179_nl;
  wire[0:0] or_2178_nl;
  wire[0:0] mux_1860_nl;
  wire[0:0] mux_1859_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] or_2177_nl;
  wire[0:0] or_2175_nl;
  wire[0:0] mux_1857_nl;
  wire[0:0] or_2173_nl;
  wire[0:0] or_2172_nl;
  wire[0:0] nand_85_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] nor_1032_nl;
  wire[0:0] mux_1885_nl;
  wire[0:0] nand_433_nl;
  wire[0:0] mux_1884_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] mux_1882_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] nor_1023_nl;
  wire[0:0] mux_1881_nl;
  wire[0:0] nor_1024_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] mux_1879_nl;
  wire[0:0] nor_1026_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] mux_1878_nl;
  wire[0:0] nor_1028_nl;
  wire[0:0] nor_1029_nl;
  wire[0:0] or_4106_nl;
  wire[0:0] mux_1877_nl;
  wire[0:0] mux_1876_nl;
  wire[0:0] mux_1875_nl;
  wire[0:0] or_2198_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] or_2195_nl;
  wire[0:0] mux_1873_nl;
  wire[0:0] mux_1872_nl;
  wire[0:0] or_2192_nl;
  wire[0:0] mux_1871_nl;
  wire[0:0] or_2189_nl;
  wire[0:0] mux_1900_nl;
  wire[0:0] mux_1899_nl;
  wire[0:0] or_2232_nl;
  wire[0:0] mux_1898_nl;
  wire[0:0] or_2231_nl;
  wire[0:0] or_2230_nl;
  wire[0:0] mux_1897_nl;
  wire[0:0] mux_1896_nl;
  wire[0:0] mux_1895_nl;
  wire[0:0] or_2228_nl;
  wire[0:0] mux_1894_nl;
  wire[0:0] or_2226_nl;
  wire[0:0] mux_1893_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] or_2225_nl;
  wire[0:0] mux_1891_nl;
  wire[0:0] or_2223_nl;
  wire[0:0] or_2222_nl;
  wire[0:0] mux_1890_nl;
  wire[0:0] mux_1889_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] or_2221_nl;
  wire[0:0] or_2219_nl;
  wire[0:0] mux_1887_nl;
  wire[0:0] or_2217_nl;
  wire[0:0] or_2216_nl;
  wire[0:0] nand_87_nl;
  wire[0:0] mux_1886_nl;
  wire[0:0] nor_1020_nl;
  wire[0:0] nor_1021_nl;
  wire[0:0] mux_1915_nl;
  wire[0:0] nand_432_nl;
  wire[0:0] mux_1914_nl;
  wire[0:0] mux_1913_nl;
  wire[0:0] mux_1912_nl;
  wire[0:0] nor_1011_nl;
  wire[0:0] nor_1012_nl;
  wire[0:0] mux_1911_nl;
  wire[0:0] nor_1013_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] mux_1910_nl;
  wire[0:0] mux_1909_nl;
  wire[0:0] nor_1015_nl;
  wire[0:0] nor_1016_nl;
  wire[0:0] mux_1908_nl;
  wire[0:0] nor_1017_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] or_4105_nl;
  wire[0:0] mux_1907_nl;
  wire[0:0] mux_1906_nl;
  wire[0:0] mux_1905_nl;
  wire[0:0] or_2242_nl;
  wire[0:0] mux_1904_nl;
  wire[0:0] or_2239_nl;
  wire[0:0] mux_1903_nl;
  wire[0:0] mux_1902_nl;
  wire[0:0] or_2236_nl;
  wire[0:0] mux_1901_nl;
  wire[0:0] or_2233_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] or_2276_nl;
  wire[0:0] mux_1928_nl;
  wire[0:0] or_2275_nl;
  wire[0:0] or_2274_nl;
  wire[0:0] mux_1927_nl;
  wire[0:0] mux_1926_nl;
  wire[0:0] mux_1925_nl;
  wire[0:0] or_2272_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] or_2270_nl;
  wire[0:0] mux_1923_nl;
  wire[0:0] mux_1922_nl;
  wire[0:0] or_2269_nl;
  wire[0:0] mux_1921_nl;
  wire[0:0] or_2267_nl;
  wire[0:0] or_2266_nl;
  wire[0:0] mux_1920_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] mux_1918_nl;
  wire[0:0] or_2265_nl;
  wire[0:0] or_2263_nl;
  wire[0:0] mux_1917_nl;
  wire[0:0] or_2261_nl;
  wire[0:0] or_2260_nl;
  wire[0:0] nand_89_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] nor_1009_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] mux_1945_nl;
  wire[0:0] nand_431_nl;
  wire[0:0] mux_1944_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] mux_1942_nl;
  wire[0:0] nor_1000_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] mux_1941_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] nor_1003_nl;
  wire[0:0] mux_1940_nl;
  wire[0:0] mux_1939_nl;
  wire[0:0] nor_1004_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] mux_1938_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] or_4104_nl;
  wire[0:0] mux_1937_nl;
  wire[0:0] mux_1936_nl;
  wire[0:0] mux_1935_nl;
  wire[0:0] or_2286_nl;
  wire[0:0] mux_1934_nl;
  wire[0:0] or_2283_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] mux_1932_nl;
  wire[0:0] or_2280_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] or_2277_nl;
  wire[0:0] mux_1960_nl;
  wire[0:0] mux_1959_nl;
  wire[0:0] or_2320_nl;
  wire[0:0] mux_1958_nl;
  wire[0:0] or_2319_nl;
  wire[0:0] or_2318_nl;
  wire[0:0] mux_1957_nl;
  wire[0:0] mux_1956_nl;
  wire[0:0] mux_1955_nl;
  wire[0:0] or_2316_nl;
  wire[0:0] mux_1954_nl;
  wire[0:0] or_2314_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] or_2313_nl;
  wire[0:0] mux_1951_nl;
  wire[0:0] or_2311_nl;
  wire[0:0] or_2310_nl;
  wire[0:0] mux_1950_nl;
  wire[0:0] mux_1949_nl;
  wire[0:0] mux_1948_nl;
  wire[0:0] or_2309_nl;
  wire[0:0] or_2307_nl;
  wire[0:0] mux_1947_nl;
  wire[0:0] or_2305_nl;
  wire[0:0] or_2304_nl;
  wire[0:0] nand_91_nl;
  wire[0:0] mux_1946_nl;
  wire[0:0] nor_998_nl;
  wire[0:0] nor_999_nl;
  wire[0:0] mux_1975_nl;
  wire[0:0] nand_430_nl;
  wire[0:0] mux_1974_nl;
  wire[0:0] mux_1973_nl;
  wire[0:0] mux_1972_nl;
  wire[0:0] and_590_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_1971_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] mux_1970_nl;
  wire[0:0] mux_1969_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] mux_1968_nl;
  wire[0:0] nor_995_nl;
  wire[0:0] nor_996_nl;
  wire[0:0] or_4103_nl;
  wire[0:0] mux_1967_nl;
  wire[0:0] mux_1966_nl;
  wire[0:0] mux_1965_nl;
  wire[0:0] or_2330_nl;
  wire[0:0] mux_1964_nl;
  wire[0:0] or_2327_nl;
  wire[0:0] mux_1963_nl;
  wire[0:0] mux_1962_nl;
  wire[0:0] or_2324_nl;
  wire[0:0] mux_1961_nl;
  wire[0:0] or_2321_nl;
  wire[0:0] mux_1990_nl;
  wire[0:0] mux_1989_nl;
  wire[0:0] or_2364_nl;
  wire[0:0] mux_1988_nl;
  wire[0:0] or_2363_nl;
  wire[0:0] or_2362_nl;
  wire[0:0] mux_1987_nl;
  wire[0:0] mux_1986_nl;
  wire[0:0] mux_1985_nl;
  wire[0:0] or_2360_nl;
  wire[0:0] mux_1984_nl;
  wire[0:0] or_2358_nl;
  wire[0:0] mux_1983_nl;
  wire[0:0] mux_1982_nl;
  wire[0:0] or_2357_nl;
  wire[0:0] mux_1981_nl;
  wire[0:0] or_2355_nl;
  wire[0:0] or_2354_nl;
  wire[0:0] mux_1980_nl;
  wire[0:0] mux_1979_nl;
  wire[0:0] mux_1978_nl;
  wire[0:0] or_2353_nl;
  wire[0:0] nand_296_nl;
  wire[0:0] mux_1977_nl;
  wire[0:0] or_2349_nl;
  wire[0:0] or_2348_nl;
  wire[0:0] nand_93_nl;
  wire[0:0] mux_1976_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] mux_2005_nl;
  wire[0:0] nand_429_nl;
  wire[0:0] mux_2004_nl;
  wire[0:0] mux_2003_nl;
  wire[0:0] mux_2002_nl;
  wire[0:0] nor_979_nl;
  wire[0:0] nor_980_nl;
  wire[0:0] mux_2001_nl;
  wire[0:0] nor_981_nl;
  wire[0:0] nor_982_nl;
  wire[0:0] mux_2000_nl;
  wire[0:0] mux_1999_nl;
  wire[0:0] nor_983_nl;
  wire[0:0] nor_984_nl;
  wire[0:0] mux_1998_nl;
  wire[0:0] nor_985_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] or_4102_nl;
  wire[0:0] mux_1997_nl;
  wire[0:0] mux_1996_nl;
  wire[0:0] mux_1995_nl;
  wire[0:0] or_2374_nl;
  wire[0:0] mux_1994_nl;
  wire[0:0] or_2371_nl;
  wire[0:0] mux_1993_nl;
  wire[0:0] mux_1992_nl;
  wire[0:0] or_2368_nl;
  wire[0:0] mux_1991_nl;
  wire[0:0] or_2365_nl;
  wire[0:0] mux_2020_nl;
  wire[0:0] mux_2019_nl;
  wire[0:0] or_2408_nl;
  wire[0:0] mux_2018_nl;
  wire[0:0] or_2407_nl;
  wire[0:0] or_2406_nl;
  wire[0:0] mux_2017_nl;
  wire[0:0] mux_2016_nl;
  wire[0:0] mux_2015_nl;
  wire[0:0] or_2404_nl;
  wire[0:0] mux_2014_nl;
  wire[0:0] or_2402_nl;
  wire[0:0] mux_2013_nl;
  wire[0:0] mux_2012_nl;
  wire[0:0] or_2401_nl;
  wire[0:0] mux_2011_nl;
  wire[0:0] or_2399_nl;
  wire[0:0] or_2398_nl;
  wire[0:0] mux_2010_nl;
  wire[0:0] mux_2009_nl;
  wire[0:0] mux_2008_nl;
  wire[0:0] or_2397_nl;
  wire[0:0] or_2395_nl;
  wire[0:0] mux_2007_nl;
  wire[0:0] or_2393_nl;
  wire[0:0] or_2392_nl;
  wire[0:0] nand_95_nl;
  wire[0:0] mux_2006_nl;
  wire[0:0] nor_977_nl;
  wire[0:0] nor_978_nl;
  wire[0:0] mux_2035_nl;
  wire[0:0] nand_428_nl;
  wire[0:0] mux_2034_nl;
  wire[0:0] mux_2033_nl;
  wire[0:0] mux_2032_nl;
  wire[0:0] nor_968_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] mux_2031_nl;
  wire[0:0] nor_970_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] mux_2030_nl;
  wire[0:0] mux_2029_nl;
  wire[0:0] nor_972_nl;
  wire[0:0] nor_973_nl;
  wire[0:0] mux_2028_nl;
  wire[0:0] nor_974_nl;
  wire[0:0] nor_975_nl;
  wire[0:0] or_4101_nl;
  wire[0:0] mux_2027_nl;
  wire[0:0] mux_2026_nl;
  wire[0:0] mux_2025_nl;
  wire[0:0] or_2418_nl;
  wire[0:0] mux_2024_nl;
  wire[0:0] or_2415_nl;
  wire[0:0] mux_2023_nl;
  wire[0:0] mux_2022_nl;
  wire[0:0] or_2412_nl;
  wire[0:0] mux_2021_nl;
  wire[0:0] or_2409_nl;
  wire[0:0] mux_2050_nl;
  wire[0:0] mux_2049_nl;
  wire[0:0] or_2452_nl;
  wire[0:0] mux_2048_nl;
  wire[0:0] or_2451_nl;
  wire[0:0] or_2450_nl;
  wire[0:0] mux_2047_nl;
  wire[0:0] mux_2046_nl;
  wire[0:0] mux_2045_nl;
  wire[0:0] or_2448_nl;
  wire[0:0] mux_2044_nl;
  wire[0:0] or_2446_nl;
  wire[0:0] mux_2043_nl;
  wire[0:0] mux_2042_nl;
  wire[0:0] or_2445_nl;
  wire[0:0] mux_2041_nl;
  wire[0:0] or_2443_nl;
  wire[0:0] or_2442_nl;
  wire[0:0] mux_2040_nl;
  wire[0:0] mux_2039_nl;
  wire[0:0] mux_2038_nl;
  wire[0:0] or_2441_nl;
  wire[0:0] or_2439_nl;
  wire[0:0] mux_2037_nl;
  wire[0:0] or_2437_nl;
  wire[0:0] or_2436_nl;
  wire[0:0] nand_97_nl;
  wire[0:0] mux_2036_nl;
  wire[0:0] nor_966_nl;
  wire[0:0] nor_967_nl;
  wire[0:0] mux_2065_nl;
  wire[0:0] nand_427_nl;
  wire[0:0] mux_2064_nl;
  wire[0:0] mux_2063_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] nor_957_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] mux_2061_nl;
  wire[0:0] nor_959_nl;
  wire[0:0] nor_960_nl;
  wire[0:0] mux_2060_nl;
  wire[0:0] mux_2059_nl;
  wire[0:0] nor_961_nl;
  wire[0:0] nor_962_nl;
  wire[0:0] mux_2058_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] or_4100_nl;
  wire[0:0] mux_2057_nl;
  wire[0:0] mux_2056_nl;
  wire[0:0] mux_2055_nl;
  wire[0:0] or_2462_nl;
  wire[0:0] mux_2054_nl;
  wire[0:0] or_2459_nl;
  wire[0:0] mux_2053_nl;
  wire[0:0] mux_2052_nl;
  wire[0:0] or_2456_nl;
  wire[0:0] mux_2051_nl;
  wire[0:0] or_2453_nl;
  wire[0:0] mux_2080_nl;
  wire[0:0] mux_2079_nl;
  wire[0:0] or_2496_nl;
  wire[0:0] mux_2078_nl;
  wire[0:0] or_2495_nl;
  wire[0:0] or_2494_nl;
  wire[0:0] mux_2077_nl;
  wire[0:0] mux_2076_nl;
  wire[0:0] mux_2075_nl;
  wire[0:0] or_2492_nl;
  wire[0:0] mux_2074_nl;
  wire[0:0] or_2490_nl;
  wire[0:0] mux_2073_nl;
  wire[0:0] mux_2072_nl;
  wire[0:0] or_2489_nl;
  wire[0:0] mux_2071_nl;
  wire[0:0] or_2487_nl;
  wire[0:0] or_2486_nl;
  wire[0:0] mux_2070_nl;
  wire[0:0] mux_2069_nl;
  wire[0:0] mux_2068_nl;
  wire[0:0] or_2485_nl;
  wire[0:0] or_2483_nl;
  wire[0:0] mux_2067_nl;
  wire[0:0] or_2481_nl;
  wire[0:0] or_2480_nl;
  wire[0:0] nand_99_nl;
  wire[0:0] mux_2066_nl;
  wire[0:0] nor_955_nl;
  wire[0:0] nor_956_nl;
  wire[0:0] mux_2095_nl;
  wire[0:0] nand_426_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] mux_2093_nl;
  wire[0:0] mux_2092_nl;
  wire[0:0] and_585_nl;
  wire[0:0] nor_947_nl;
  wire[0:0] mux_2091_nl;
  wire[0:0] nor_948_nl;
  wire[0:0] nor_949_nl;
  wire[0:0] mux_2090_nl;
  wire[0:0] mux_2089_nl;
  wire[0:0] nor_950_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] mux_2088_nl;
  wire[0:0] nor_952_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] or_4099_nl;
  wire[0:0] mux_2087_nl;
  wire[0:0] mux_2086_nl;
  wire[0:0] mux_2085_nl;
  wire[0:0] or_2506_nl;
  wire[0:0] mux_2084_nl;
  wire[0:0] or_2503_nl;
  wire[0:0] mux_2083_nl;
  wire[0:0] mux_2082_nl;
  wire[0:0] or_2500_nl;
  wire[0:0] mux_2081_nl;
  wire[0:0] or_2497_nl;
  wire[0:0] mux_2110_nl;
  wire[0:0] mux_2109_nl;
  wire[0:0] or_2540_nl;
  wire[0:0] mux_2108_nl;
  wire[0:0] or_2539_nl;
  wire[0:0] or_2538_nl;
  wire[0:0] mux_2107_nl;
  wire[0:0] mux_2106_nl;
  wire[0:0] mux_2105_nl;
  wire[0:0] or_2536_nl;
  wire[0:0] mux_2104_nl;
  wire[0:0] or_2534_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] or_2533_nl;
  wire[0:0] mux_2101_nl;
  wire[0:0] or_2531_nl;
  wire[0:0] or_2530_nl;
  wire[0:0] mux_2100_nl;
  wire[0:0] mux_2099_nl;
  wire[0:0] mux_2098_nl;
  wire[0:0] or_2529_nl;
  wire[0:0] nand_295_nl;
  wire[0:0] mux_2097_nl;
  wire[0:0] or_2525_nl;
  wire[0:0] or_2524_nl;
  wire[0:0] nand_101_nl;
  wire[0:0] mux_2096_nl;
  wire[0:0] nor_945_nl;
  wire[0:0] nor_946_nl;
  wire[0:0] mux_2125_nl;
  wire[0:0] nand_425_nl;
  wire[0:0] mux_2124_nl;
  wire[0:0] mux_2123_nl;
  wire[0:0] mux_2122_nl;
  wire[0:0] nor_936_nl;
  wire[0:0] nor_937_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] nor_938_nl;
  wire[0:0] nor_939_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] mux_2119_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] nor_941_nl;
  wire[0:0] mux_2118_nl;
  wire[0:0] nor_942_nl;
  wire[0:0] nor_943_nl;
  wire[0:0] or_4098_nl;
  wire[0:0] mux_2117_nl;
  wire[0:0] mux_2116_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] or_2550_nl;
  wire[0:0] mux_2114_nl;
  wire[0:0] or_2547_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] or_2544_nl;
  wire[0:0] mux_2111_nl;
  wire[0:0] or_2541_nl;
  wire[0:0] mux_2140_nl;
  wire[0:0] mux_2139_nl;
  wire[0:0] or_2584_nl;
  wire[0:0] mux_2138_nl;
  wire[0:0] or_2583_nl;
  wire[0:0] or_2582_nl;
  wire[0:0] mux_2137_nl;
  wire[0:0] mux_2136_nl;
  wire[0:0] mux_2135_nl;
  wire[0:0] or_2580_nl;
  wire[0:0] mux_2134_nl;
  wire[0:0] or_2578_nl;
  wire[0:0] mux_2133_nl;
  wire[0:0] mux_2132_nl;
  wire[0:0] or_2577_nl;
  wire[0:0] mux_2131_nl;
  wire[0:0] or_2575_nl;
  wire[0:0] or_2574_nl;
  wire[0:0] mux_2130_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] mux_2128_nl;
  wire[0:0] or_2573_nl;
  wire[0:0] or_2571_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] or_2569_nl;
  wire[0:0] or_2568_nl;
  wire[0:0] nand_103_nl;
  wire[0:0] mux_2126_nl;
  wire[0:0] nor_934_nl;
  wire[0:0] nor_935_nl;
  wire[0:0] mux_2155_nl;
  wire[0:0] nand_424_nl;
  wire[0:0] mux_2154_nl;
  wire[0:0] mux_2153_nl;
  wire[0:0] mux_2152_nl;
  wire[0:0] and_582_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] mux_2151_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] nor_928_nl;
  wire[0:0] mux_2150_nl;
  wire[0:0] mux_2149_nl;
  wire[0:0] nor_929_nl;
  wire[0:0] nor_930_nl;
  wire[0:0] mux_2148_nl;
  wire[0:0] nor_931_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] or_4097_nl;
  wire[0:0] mux_2147_nl;
  wire[0:0] mux_2146_nl;
  wire[0:0] mux_2145_nl;
  wire[0:0] or_2594_nl;
  wire[0:0] mux_2144_nl;
  wire[0:0] or_2591_nl;
  wire[0:0] mux_2143_nl;
  wire[0:0] mux_2142_nl;
  wire[0:0] or_2588_nl;
  wire[0:0] mux_2141_nl;
  wire[0:0] or_2585_nl;
  wire[0:0] mux_2170_nl;
  wire[0:0] mux_2169_nl;
  wire[0:0] or_2628_nl;
  wire[0:0] mux_2168_nl;
  wire[0:0] or_2627_nl;
  wire[0:0] or_2626_nl;
  wire[0:0] mux_2167_nl;
  wire[0:0] mux_2166_nl;
  wire[0:0] mux_2165_nl;
  wire[0:0] or_2624_nl;
  wire[0:0] mux_2164_nl;
  wire[0:0] or_2622_nl;
  wire[0:0] mux_2163_nl;
  wire[0:0] mux_2162_nl;
  wire[0:0] or_2621_nl;
  wire[0:0] mux_2161_nl;
  wire[0:0] or_2619_nl;
  wire[0:0] or_2618_nl;
  wire[0:0] mux_2160_nl;
  wire[0:0] mux_2159_nl;
  wire[0:0] mux_2158_nl;
  wire[0:0] or_2617_nl;
  wire[0:0] nand_294_nl;
  wire[0:0] mux_2157_nl;
  wire[0:0] or_2613_nl;
  wire[0:0] or_2612_nl;
  wire[0:0] nand_105_nl;
  wire[0:0] mux_2156_nl;
  wire[0:0] nor_924_nl;
  wire[0:0] nor_925_nl;
  wire[0:0] mux_2185_nl;
  wire[0:0] nand_423_nl;
  wire[0:0] mux_2184_nl;
  wire[0:0] mux_2183_nl;
  wire[0:0] mux_2182_nl;
  wire[0:0] and_579_nl;
  wire[0:0] and_580_nl;
  wire[0:0] mux_2181_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] mux_2180_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] mux_2178_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] nor_922_nl;
  wire[0:0] or_4096_nl;
  wire[0:0] mux_2177_nl;
  wire[0:0] mux_2176_nl;
  wire[0:0] mux_2175_nl;
  wire[0:0] or_2638_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] or_2635_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] mux_2172_nl;
  wire[0:0] or_2632_nl;
  wire[0:0] mux_2171_nl;
  wire[0:0] or_2629_nl;
  wire[0:0] mux_2200_nl;
  wire[0:0] mux_2199_nl;
  wire[0:0] or_2672_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] or_2671_nl;
  wire[0:0] or_2670_nl;
  wire[0:0] mux_2197_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] or_2668_nl;
  wire[0:0] mux_2194_nl;
  wire[0:0] or_2666_nl;
  wire[0:0] mux_2193_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] or_2665_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] or_2663_nl;
  wire[0:0] or_2662_nl;
  wire[0:0] mux_2190_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] mux_2188_nl;
  wire[0:0] nand_292_nl;
  wire[0:0] nand_293_nl;
  wire[0:0] mux_2187_nl;
  wire[0:0] or_2657_nl;
  wire[0:0] or_2656_nl;
  wire[0:0] nand_107_nl;
  wire[0:0] mux_2186_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] nand_422_nl;
  wire[0:0] mux_2214_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] and_575_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] and_576_nl;
  wire[0:0] and_577_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] mux_2209_nl;
  wire[0:0] and_812_nl;
  wire[0:0] and_819_nl;
  wire[0:0] mux_2208_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] or_4095_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] mux_2206_nl;
  wire[0:0] mux_2205_nl;
  wire[0:0] or_2682_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] nand_287_nl;
  wire[0:0] mux_2203_nl;
  wire[0:0] mux_2202_nl;
  wire[0:0] nand_477_nl;
  wire[0:0] mux_2201_nl;
  wire[0:0] or_2673_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2229_nl;
  wire[0:0] or_2715_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] or_2714_nl;
  wire[0:0] or_2713_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] mux_2226_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] or_2711_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] nand_278_nl;
  wire[0:0] mux_2223_nl;
  wire[0:0] mux_2222_nl;
  wire[0:0] nand_402_nl;
  wire[0:0] mux_2221_nl;
  wire[0:0] or_2706_nl;
  wire[0:0] or_2705_nl;
  wire[0:0] mux_2220_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] or_2704_nl;
  wire[0:0] nand_281_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] nand_282_nl;
  wire[0:0] nand_283_nl;
  wire[0:0] nand_109_nl;
  wire[0:0] mux_2216_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] mux_2245_nl;
  wire[0:0] nand_421_nl;
  wire[0:0] mux_2244_nl;
  wire[0:0] mux_2243_nl;
  wire[0:0] mux_2242_nl;
  wire[0:0] nor_898_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] mux_2241_nl;
  wire[0:0] nor_900_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] mux_2240_nl;
  wire[0:0] mux_2239_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] nor_903_nl;
  wire[0:0] mux_2238_nl;
  wire[0:0] nor_904_nl;
  wire[0:0] nor_905_nl;
  wire[0:0] or_4094_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] mux_2235_nl;
  wire[0:0] or_2725_nl;
  wire[0:0] mux_2234_nl;
  wire[0:0] or_2722_nl;
  wire[0:0] mux_2233_nl;
  wire[0:0] mux_2232_nl;
  wire[0:0] or_2719_nl;
  wire[0:0] mux_2231_nl;
  wire[0:0] or_2716_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] or_2759_nl;
  wire[0:0] mux_2258_nl;
  wire[0:0] or_2758_nl;
  wire[0:0] or_2757_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] mux_2256_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] or_2755_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] or_2753_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] mux_2252_nl;
  wire[0:0] or_2752_nl;
  wire[0:0] mux_2251_nl;
  wire[0:0] or_2750_nl;
  wire[0:0] or_2749_nl;
  wire[0:0] mux_2250_nl;
  wire[0:0] mux_2249_nl;
  wire[0:0] mux_2248_nl;
  wire[0:0] or_2748_nl;
  wire[0:0] or_2746_nl;
  wire[0:0] mux_2247_nl;
  wire[0:0] or_2744_nl;
  wire[0:0] or_2743_nl;
  wire[0:0] nand_111_nl;
  wire[0:0] mux_2246_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] nor_897_nl;
  wire[0:0] mux_2275_nl;
  wire[0:0] nand_420_nl;
  wire[0:0] mux_2274_nl;
  wire[0:0] mux_2273_nl;
  wire[0:0] mux_2272_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_2271_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] mux_2270_nl;
  wire[0:0] mux_2269_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] mux_2268_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] nor_894_nl;
  wire[0:0] or_4093_nl;
  wire[0:0] mux_2267_nl;
  wire[0:0] mux_2266_nl;
  wire[0:0] mux_2265_nl;
  wire[0:0] or_2769_nl;
  wire[0:0] mux_2264_nl;
  wire[0:0] or_2766_nl;
  wire[0:0] mux_2263_nl;
  wire[0:0] mux_2262_nl;
  wire[0:0] or_2763_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] or_2760_nl;
  wire[0:0] mux_2290_nl;
  wire[0:0] mux_2289_nl;
  wire[0:0] or_2803_nl;
  wire[0:0] mux_2288_nl;
  wire[0:0] or_2802_nl;
  wire[0:0] or_2801_nl;
  wire[0:0] mux_2287_nl;
  wire[0:0] mux_2286_nl;
  wire[0:0] mux_2285_nl;
  wire[0:0] or_2799_nl;
  wire[0:0] mux_2284_nl;
  wire[0:0] or_2797_nl;
  wire[0:0] mux_2283_nl;
  wire[0:0] mux_2282_nl;
  wire[0:0] or_2796_nl;
  wire[0:0] mux_2281_nl;
  wire[0:0] or_2794_nl;
  wire[0:0] or_2793_nl;
  wire[0:0] mux_2280_nl;
  wire[0:0] mux_2279_nl;
  wire[0:0] mux_2278_nl;
  wire[0:0] or_2792_nl;
  wire[0:0] or_2790_nl;
  wire[0:0] mux_2277_nl;
  wire[0:0] or_2788_nl;
  wire[0:0] or_2787_nl;
  wire[0:0] nand_113_nl;
  wire[0:0] mux_2276_nl;
  wire[0:0] nor_885_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] mux_2305_nl;
  wire[0:0] nand_419_nl;
  wire[0:0] mux_2304_nl;
  wire[0:0] mux_2303_nl;
  wire[0:0] mux_2302_nl;
  wire[0:0] nor_876_nl;
  wire[0:0] nor_877_nl;
  wire[0:0] mux_2301_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] mux_2300_nl;
  wire[0:0] mux_2299_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] mux_2298_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] or_4092_nl;
  wire[0:0] mux_2297_nl;
  wire[0:0] mux_2296_nl;
  wire[0:0] mux_2295_nl;
  wire[0:0] or_2813_nl;
  wire[0:0] mux_2294_nl;
  wire[0:0] or_2810_nl;
  wire[0:0] mux_2293_nl;
  wire[0:0] mux_2292_nl;
  wire[0:0] or_2807_nl;
  wire[0:0] mux_2291_nl;
  wire[0:0] or_2804_nl;
  wire[0:0] mux_2320_nl;
  wire[0:0] mux_2319_nl;
  wire[0:0] or_2847_nl;
  wire[0:0] mux_2318_nl;
  wire[0:0] or_2846_nl;
  wire[0:0] or_2845_nl;
  wire[0:0] mux_2317_nl;
  wire[0:0] mux_2316_nl;
  wire[0:0] mux_2315_nl;
  wire[0:0] or_2843_nl;
  wire[0:0] mux_2314_nl;
  wire[0:0] or_2841_nl;
  wire[0:0] mux_2313_nl;
  wire[0:0] mux_2312_nl;
  wire[0:0] or_2840_nl;
  wire[0:0] mux_2311_nl;
  wire[0:0] or_2838_nl;
  wire[0:0] or_2837_nl;
  wire[0:0] mux_2310_nl;
  wire[0:0] mux_2309_nl;
  wire[0:0] mux_2308_nl;
  wire[0:0] or_2836_nl;
  wire[0:0] or_2834_nl;
  wire[0:0] mux_2307_nl;
  wire[0:0] or_2832_nl;
  wire[0:0] or_2831_nl;
  wire[0:0] nand_115_nl;
  wire[0:0] mux_2306_nl;
  wire[0:0] nor_874_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] mux_2335_nl;
  wire[0:0] nand_418_nl;
  wire[0:0] mux_2334_nl;
  wire[0:0] mux_2333_nl;
  wire[0:0] mux_2332_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] nor_866_nl;
  wire[0:0] mux_2331_nl;
  wire[0:0] nor_867_nl;
  wire[0:0] nor_868_nl;
  wire[0:0] mux_2330_nl;
  wire[0:0] mux_2329_nl;
  wire[0:0] nor_869_nl;
  wire[0:0] nor_870_nl;
  wire[0:0] mux_2328_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] nor_872_nl;
  wire[0:0] or_4091_nl;
  wire[0:0] mux_2327_nl;
  wire[0:0] mux_2326_nl;
  wire[0:0] mux_2325_nl;
  wire[0:0] or_2857_nl;
  wire[0:0] mux_2324_nl;
  wire[0:0] or_2854_nl;
  wire[0:0] mux_2323_nl;
  wire[0:0] mux_2322_nl;
  wire[0:0] or_2851_nl;
  wire[0:0] mux_2321_nl;
  wire[0:0] or_2848_nl;
  wire[0:0] mux_2350_nl;
  wire[0:0] mux_2349_nl;
  wire[0:0] or_2891_nl;
  wire[0:0] mux_2348_nl;
  wire[0:0] or_2890_nl;
  wire[0:0] or_2889_nl;
  wire[0:0] mux_2347_nl;
  wire[0:0] mux_2346_nl;
  wire[0:0] mux_2345_nl;
  wire[0:0] or_2887_nl;
  wire[0:0] mux_2344_nl;
  wire[0:0] or_2885_nl;
  wire[0:0] mux_2343_nl;
  wire[0:0] mux_2342_nl;
  wire[0:0] or_2884_nl;
  wire[0:0] mux_2341_nl;
  wire[0:0] or_2882_nl;
  wire[0:0] or_2881_nl;
  wire[0:0] mux_2340_nl;
  wire[0:0] mux_2339_nl;
  wire[0:0] mux_2338_nl;
  wire[0:0] or_2880_nl;
  wire[0:0] or_2878_nl;
  wire[0:0] mux_2337_nl;
  wire[0:0] or_2876_nl;
  wire[0:0] or_2875_nl;
  wire[0:0] nand_117_nl;
  wire[0:0] mux_2336_nl;
  wire[0:0] nor_863_nl;
  wire[0:0] nor_864_nl;
  wire[0:0] mux_2365_nl;
  wire[0:0] nand_417_nl;
  wire[0:0] mux_2364_nl;
  wire[0:0] mux_2363_nl;
  wire[0:0] mux_2362_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] nor_855_nl;
  wire[0:0] mux_2361_nl;
  wire[0:0] nor_856_nl;
  wire[0:0] nor_857_nl;
  wire[0:0] mux_2360_nl;
  wire[0:0] mux_2359_nl;
  wire[0:0] nor_858_nl;
  wire[0:0] nor_859_nl;
  wire[0:0] mux_2358_nl;
  wire[0:0] nor_860_nl;
  wire[0:0] nor_861_nl;
  wire[0:0] or_4090_nl;
  wire[0:0] mux_2357_nl;
  wire[0:0] mux_2356_nl;
  wire[0:0] mux_2355_nl;
  wire[0:0] or_2901_nl;
  wire[0:0] mux_2354_nl;
  wire[0:0] or_2898_nl;
  wire[0:0] mux_2353_nl;
  wire[0:0] mux_2352_nl;
  wire[0:0] or_2895_nl;
  wire[0:0] mux_2351_nl;
  wire[0:0] or_2892_nl;
  wire[0:0] mux_2380_nl;
  wire[0:0] mux_2379_nl;
  wire[0:0] or_2935_nl;
  wire[0:0] mux_2378_nl;
  wire[0:0] or_2934_nl;
  wire[0:0] or_2933_nl;
  wire[0:0] mux_2377_nl;
  wire[0:0] mux_2376_nl;
  wire[0:0] mux_2375_nl;
  wire[0:0] or_2931_nl;
  wire[0:0] mux_2374_nl;
  wire[0:0] or_2929_nl;
  wire[0:0] mux_2373_nl;
  wire[0:0] mux_2372_nl;
  wire[0:0] or_2928_nl;
  wire[0:0] mux_2371_nl;
  wire[0:0] or_2926_nl;
  wire[0:0] or_2925_nl;
  wire[0:0] mux_2370_nl;
  wire[0:0] mux_2369_nl;
  wire[0:0] mux_2368_nl;
  wire[0:0] or_2924_nl;
  wire[0:0] or_2922_nl;
  wire[0:0] mux_2367_nl;
  wire[0:0] or_2920_nl;
  wire[0:0] or_2919_nl;
  wire[0:0] nand_119_nl;
  wire[0:0] mux_2366_nl;
  wire[0:0] nor_852_nl;
  wire[0:0] nor_853_nl;
  wire[0:0] mux_2395_nl;
  wire[0:0] nand_416_nl;
  wire[0:0] mux_2394_nl;
  wire[0:0] mux_2393_nl;
  wire[0:0] mux_2392_nl;
  wire[0:0] nor_843_nl;
  wire[0:0] nor_844_nl;
  wire[0:0] mux_2391_nl;
  wire[0:0] nor_845_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] mux_2390_nl;
  wire[0:0] mux_2389_nl;
  wire[0:0] nor_847_nl;
  wire[0:0] nor_848_nl;
  wire[0:0] mux_2388_nl;
  wire[0:0] nor_849_nl;
  wire[0:0] nor_850_nl;
  wire[0:0] or_4089_nl;
  wire[0:0] mux_2387_nl;
  wire[0:0] mux_2386_nl;
  wire[0:0] mux_2385_nl;
  wire[0:0] or_2945_nl;
  wire[0:0] mux_2384_nl;
  wire[0:0] or_2942_nl;
  wire[0:0] mux_2383_nl;
  wire[0:0] mux_2382_nl;
  wire[0:0] or_2939_nl;
  wire[0:0] mux_2381_nl;
  wire[0:0] or_2936_nl;
  wire[0:0] mux_2410_nl;
  wire[0:0] mux_2409_nl;
  wire[0:0] or_2979_nl;
  wire[0:0] mux_2408_nl;
  wire[0:0] or_2978_nl;
  wire[0:0] or_2977_nl;
  wire[0:0] mux_2407_nl;
  wire[0:0] mux_2406_nl;
  wire[0:0] mux_2405_nl;
  wire[0:0] or_2975_nl;
  wire[0:0] mux_2404_nl;
  wire[0:0] or_2973_nl;
  wire[0:0] mux_2403_nl;
  wire[0:0] mux_2402_nl;
  wire[0:0] or_2972_nl;
  wire[0:0] mux_2401_nl;
  wire[0:0] or_2970_nl;
  wire[0:0] or_2969_nl;
  wire[0:0] mux_2400_nl;
  wire[0:0] mux_2399_nl;
  wire[0:0] mux_2398_nl;
  wire[0:0] or_2968_nl;
  wire[0:0] or_2966_nl;
  wire[0:0] mux_2397_nl;
  wire[0:0] or_2964_nl;
  wire[0:0] or_2963_nl;
  wire[0:0] nand_121_nl;
  wire[0:0] mux_2396_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] nor_842_nl;
  wire[0:0] mux_2425_nl;
  wire[0:0] nand_415_nl;
  wire[0:0] mux_2424_nl;
  wire[0:0] mux_2423_nl;
  wire[0:0] mux_2422_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] and_567_nl;
  wire[0:0] mux_2421_nl;
  wire[0:0] nor_834_nl;
  wire[0:0] nor_835_nl;
  wire[0:0] mux_2420_nl;
  wire[0:0] mux_2419_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] nor_837_nl;
  wire[0:0] mux_2418_nl;
  wire[0:0] nor_838_nl;
  wire[0:0] nor_839_nl;
  wire[0:0] or_4088_nl;
  wire[0:0] mux_2417_nl;
  wire[0:0] mux_2416_nl;
  wire[0:0] mux_2415_nl;
  wire[0:0] or_2989_nl;
  wire[0:0] mux_2414_nl;
  wire[0:0] or_2986_nl;
  wire[0:0] mux_2413_nl;
  wire[0:0] mux_2412_nl;
  wire[0:0] or_2983_nl;
  wire[0:0] mux_2411_nl;
  wire[0:0] or_2980_nl;
  wire[0:0] mux_2440_nl;
  wire[0:0] mux_2439_nl;
  wire[0:0] or_3023_nl;
  wire[0:0] mux_2438_nl;
  wire[0:0] or_3022_nl;
  wire[0:0] or_3021_nl;
  wire[0:0] mux_2437_nl;
  wire[0:0] mux_2436_nl;
  wire[0:0] mux_2435_nl;
  wire[0:0] or_3019_nl;
  wire[0:0] mux_2434_nl;
  wire[0:0] or_3017_nl;
  wire[0:0] mux_2433_nl;
  wire[0:0] mux_2432_nl;
  wire[0:0] or_3016_nl;
  wire[0:0] mux_2431_nl;
  wire[0:0] or_3014_nl;
  wire[0:0] or_3013_nl;
  wire[0:0] mux_2430_nl;
  wire[0:0] mux_2429_nl;
  wire[0:0] mux_2428_nl;
  wire[0:0] nand_271_nl;
  wire[0:0] or_3010_nl;
  wire[0:0] mux_2427_nl;
  wire[0:0] or_3008_nl;
  wire[0:0] or_3007_nl;
  wire[0:0] nand_123_nl;
  wire[0:0] mux_2426_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] nor_832_nl;
  wire[0:0] mux_2455_nl;
  wire[0:0] nand_414_nl;
  wire[0:0] mux_2454_nl;
  wire[0:0] mux_2453_nl;
  wire[0:0] mux_2452_nl;
  wire[0:0] nor_824_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] mux_2451_nl;
  wire[0:0] and_564_nl;
  wire[0:0] and_565_nl;
  wire[0:0] mux_2450_nl;
  wire[0:0] mux_2449_nl;
  wire[0:0] and_813_nl;
  wire[0:0] and_820_nl;
  wire[0:0] mux_2448_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] nor_829_nl;
  wire[0:0] or_4087_nl;
  wire[0:0] mux_2447_nl;
  wire[0:0] mux_2446_nl;
  wire[0:0] mux_2445_nl;
  wire[0:0] or_3033_nl;
  wire[0:0] mux_2444_nl;
  wire[0:0] nand_267_nl;
  wire[0:0] mux_2443_nl;
  wire[0:0] mux_2442_nl;
  wire[0:0] nand_476_nl;
  wire[0:0] mux_2441_nl;
  wire[0:0] or_3024_nl;
  wire[0:0] mux_2470_nl;
  wire[0:0] mux_2469_nl;
  wire[0:0] or_3067_nl;
  wire[0:0] mux_2468_nl;
  wire[0:0] or_3066_nl;
  wire[0:0] or_3065_nl;
  wire[0:0] mux_2467_nl;
  wire[0:0] mux_2466_nl;
  wire[0:0] mux_2465_nl;
  wire[0:0] or_3063_nl;
  wire[0:0] mux_2464_nl;
  wire[0:0] nand_258_nl;
  wire[0:0] mux_2463_nl;
  wire[0:0] mux_2462_nl;
  wire[0:0] nand_400_nl;
  wire[0:0] mux_2461_nl;
  wire[0:0] or_3058_nl;
  wire[0:0] or_3057_nl;
  wire[0:0] mux_2460_nl;
  wire[0:0] mux_2459_nl;
  wire[0:0] mux_2458_nl;
  wire[0:0] or_3056_nl;
  wire[0:0] or_3054_nl;
  wire[0:0] mux_2457_nl;
  wire[0:0] nand_261_nl;
  wire[0:0] nand_262_nl;
  wire[0:0] nand_125_nl;
  wire[0:0] mux_2456_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] nor_823_nl;
  wire[0:0] mux_2485_nl;
  wire[0:0] nand_413_nl;
  wire[0:0] mux_2484_nl;
  wire[0:0] mux_2483_nl;
  wire[0:0] mux_2482_nl;
  wire[0:0] nor_813_nl;
  wire[0:0] nor_814_nl;
  wire[0:0] mux_2481_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] nor_816_nl;
  wire[0:0] mux_2480_nl;
  wire[0:0] mux_2479_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] nor_818_nl;
  wire[0:0] mux_2478_nl;
  wire[0:0] nor_819_nl;
  wire[0:0] nor_820_nl;
  wire[0:0] or_4086_nl;
  wire[0:0] mux_2477_nl;
  wire[0:0] mux_2476_nl;
  wire[0:0] mux_2475_nl;
  wire[0:0] or_3077_nl;
  wire[0:0] mux_2474_nl;
  wire[0:0] or_3074_nl;
  wire[0:0] mux_2473_nl;
  wire[0:0] mux_2472_nl;
  wire[0:0] or_3071_nl;
  wire[0:0] mux_2471_nl;
  wire[0:0] or_3068_nl;
  wire[0:0] mux_2500_nl;
  wire[0:0] mux_2499_nl;
  wire[0:0] or_3111_nl;
  wire[0:0] mux_2498_nl;
  wire[0:0] or_3110_nl;
  wire[0:0] or_3109_nl;
  wire[0:0] mux_2497_nl;
  wire[0:0] mux_2496_nl;
  wire[0:0] mux_2495_nl;
  wire[0:0] or_3107_nl;
  wire[0:0] mux_2494_nl;
  wire[0:0] or_3105_nl;
  wire[0:0] mux_2493_nl;
  wire[0:0] mux_2492_nl;
  wire[0:0] or_3104_nl;
  wire[0:0] mux_2491_nl;
  wire[0:0] or_3102_nl;
  wire[0:0] or_3101_nl;
  wire[0:0] mux_2490_nl;
  wire[0:0] mux_2489_nl;
  wire[0:0] mux_2488_nl;
  wire[0:0] or_3100_nl;
  wire[0:0] or_3098_nl;
  wire[0:0] mux_2487_nl;
  wire[0:0] or_3096_nl;
  wire[0:0] or_3095_nl;
  wire[0:0] nand_127_nl;
  wire[0:0] mux_2486_nl;
  wire[0:0] nor_811_nl;
  wire[0:0] nor_812_nl;
  wire[0:0] mux_2515_nl;
  wire[0:0] nand_412_nl;
  wire[0:0] mux_2514_nl;
  wire[0:0] mux_2513_nl;
  wire[0:0] mux_2512_nl;
  wire[0:0] nor_802_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] mux_2511_nl;
  wire[0:0] nor_804_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] mux_2510_nl;
  wire[0:0] mux_2509_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] nor_807_nl;
  wire[0:0] mux_2508_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] nor_809_nl;
  wire[0:0] or_4085_nl;
  wire[0:0] mux_2507_nl;
  wire[0:0] mux_2506_nl;
  wire[0:0] mux_2505_nl;
  wire[0:0] or_3121_nl;
  wire[0:0] mux_2504_nl;
  wire[0:0] or_3118_nl;
  wire[0:0] mux_2503_nl;
  wire[0:0] mux_2502_nl;
  wire[0:0] or_3115_nl;
  wire[0:0] mux_2501_nl;
  wire[0:0] or_3112_nl;
  wire[0:0] mux_2530_nl;
  wire[0:0] mux_2529_nl;
  wire[0:0] or_3155_nl;
  wire[0:0] mux_2528_nl;
  wire[0:0] or_3154_nl;
  wire[0:0] or_3153_nl;
  wire[0:0] mux_2527_nl;
  wire[0:0] mux_2526_nl;
  wire[0:0] mux_2525_nl;
  wire[0:0] or_3151_nl;
  wire[0:0] mux_2524_nl;
  wire[0:0] or_3149_nl;
  wire[0:0] mux_2523_nl;
  wire[0:0] mux_2522_nl;
  wire[0:0] or_3148_nl;
  wire[0:0] mux_2521_nl;
  wire[0:0] or_3146_nl;
  wire[0:0] or_3145_nl;
  wire[0:0] mux_2520_nl;
  wire[0:0] mux_2519_nl;
  wire[0:0] mux_2518_nl;
  wire[0:0] or_3144_nl;
  wire[0:0] or_3142_nl;
  wire[0:0] mux_2517_nl;
  wire[0:0] or_3140_nl;
  wire[0:0] or_3139_nl;
  wire[0:0] nand_129_nl;
  wire[0:0] mux_2516_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] nor_801_nl;
  wire[0:0] mux_2545_nl;
  wire[0:0] nand_411_nl;
  wire[0:0] mux_2544_nl;
  wire[0:0] mux_2543_nl;
  wire[0:0] mux_2542_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] and_560_nl;
  wire[0:0] mux_2541_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] nor_794_nl;
  wire[0:0] mux_2540_nl;
  wire[0:0] mux_2539_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] mux_2538_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] or_4084_nl;
  wire[0:0] mux_2537_nl;
  wire[0:0] mux_2536_nl;
  wire[0:0] mux_2535_nl;
  wire[0:0] or_3165_nl;
  wire[0:0] mux_2534_nl;
  wire[0:0] or_3162_nl;
  wire[0:0] mux_2533_nl;
  wire[0:0] mux_2532_nl;
  wire[0:0] or_3159_nl;
  wire[0:0] mux_2531_nl;
  wire[0:0] or_3156_nl;
  wire[0:0] mux_2560_nl;
  wire[0:0] mux_2559_nl;
  wire[0:0] or_3199_nl;
  wire[0:0] mux_2558_nl;
  wire[0:0] or_3198_nl;
  wire[0:0] or_3197_nl;
  wire[0:0] mux_2557_nl;
  wire[0:0] mux_2556_nl;
  wire[0:0] mux_2555_nl;
  wire[0:0] or_3195_nl;
  wire[0:0] mux_2554_nl;
  wire[0:0] or_3193_nl;
  wire[0:0] mux_2553_nl;
  wire[0:0] mux_2552_nl;
  wire[0:0] or_3192_nl;
  wire[0:0] mux_2551_nl;
  wire[0:0] or_3190_nl;
  wire[0:0] or_3189_nl;
  wire[0:0] mux_2550_nl;
  wire[0:0] mux_2549_nl;
  wire[0:0] mux_2548_nl;
  wire[0:0] nand_252_nl;
  wire[0:0] or_3186_nl;
  wire[0:0] mux_2547_nl;
  wire[0:0] or_3184_nl;
  wire[0:0] or_3183_nl;
  wire[0:0] nand_131_nl;
  wire[0:0] mux_2546_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] mux_2575_nl;
  wire[0:0] nand_410_nl;
  wire[0:0] mux_2574_nl;
  wire[0:0] mux_2573_nl;
  wire[0:0] mux_2572_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] nor_784_nl;
  wire[0:0] mux_2571_nl;
  wire[0:0] and_557_nl;
  wire[0:0] and_558_nl;
  wire[0:0] mux_2570_nl;
  wire[0:0] mux_2569_nl;
  wire[0:0] and_814_nl;
  wire[0:0] and_821_nl;
  wire[0:0] mux_2568_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] or_4083_nl;
  wire[0:0] mux_2567_nl;
  wire[0:0] mux_2566_nl;
  wire[0:0] mux_2565_nl;
  wire[0:0] or_3208_nl;
  wire[0:0] mux_2564_nl;
  wire[0:0] nand_247_nl;
  wire[0:0] mux_2563_nl;
  wire[0:0] mux_2562_nl;
  wire[0:0] nand_475_nl;
  wire[0:0] mux_2561_nl;
  wire[0:0] or_3200_nl;
  wire[0:0] mux_2590_nl;
  wire[0:0] mux_2589_nl;
  wire[0:0] or_3242_nl;
  wire[0:0] mux_2588_nl;
  wire[0:0] or_3241_nl;
  wire[0:0] or_3240_nl;
  wire[0:0] mux_2587_nl;
  wire[0:0] mux_2586_nl;
  wire[0:0] mux_2585_nl;
  wire[0:0] or_3238_nl;
  wire[0:0] mux_2584_nl;
  wire[0:0] nand_238_nl;
  wire[0:0] mux_2583_nl;
  wire[0:0] mux_2582_nl;
  wire[0:0] nand_398_nl;
  wire[0:0] mux_2581_nl;
  wire[0:0] or_3233_nl;
  wire[0:0] or_3232_nl;
  wire[0:0] mux_2580_nl;
  wire[0:0] mux_2579_nl;
  wire[0:0] mux_2578_nl;
  wire[0:0] or_3231_nl;
  wire[0:0] or_3229_nl;
  wire[0:0] mux_2577_nl;
  wire[0:0] nand_242_nl;
  wire[0:0] nand_243_nl;
  wire[0:0] nand_133_nl;
  wire[0:0] mux_2576_nl;
  wire[0:0] nor_781_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] mux_2605_nl;
  wire[0:0] nand_409_nl;
  wire[0:0] mux_2604_nl;
  wire[0:0] mux_2603_nl;
  wire[0:0] mux_2602_nl;
  wire[0:0] nor_773_nl;
  wire[0:0] and_555_nl;
  wire[0:0] mux_2601_nl;
  wire[0:0] nor_774_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] mux_2600_nl;
  wire[0:0] mux_2599_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] nor_777_nl;
  wire[0:0] mux_2598_nl;
  wire[0:0] nor_778_nl;
  wire[0:0] nor_779_nl;
  wire[0:0] or_4082_nl;
  wire[0:0] mux_2597_nl;
  wire[0:0] mux_2596_nl;
  wire[0:0] mux_2595_nl;
  wire[0:0] or_3252_nl;
  wire[0:0] mux_2594_nl;
  wire[0:0] or_3249_nl;
  wire[0:0] mux_2593_nl;
  wire[0:0] mux_2592_nl;
  wire[0:0] or_3246_nl;
  wire[0:0] mux_2591_nl;
  wire[0:0] or_3243_nl;
  wire[0:0] mux_2620_nl;
  wire[0:0] mux_2619_nl;
  wire[0:0] or_3286_nl;
  wire[0:0] mux_2618_nl;
  wire[0:0] or_3285_nl;
  wire[0:0] or_3284_nl;
  wire[0:0] mux_2617_nl;
  wire[0:0] mux_2616_nl;
  wire[0:0] mux_2615_nl;
  wire[0:0] or_3282_nl;
  wire[0:0] mux_2614_nl;
  wire[0:0] or_3280_nl;
  wire[0:0] mux_2613_nl;
  wire[0:0] mux_2612_nl;
  wire[0:0] or_3279_nl;
  wire[0:0] mux_2611_nl;
  wire[0:0] or_3277_nl;
  wire[0:0] or_3276_nl;
  wire[0:0] mux_2610_nl;
  wire[0:0] mux_2609_nl;
  wire[0:0] mux_2608_nl;
  wire[0:0] nand_237_nl;
  wire[0:0] or_3273_nl;
  wire[0:0] mux_2607_nl;
  wire[0:0] or_3271_nl;
  wire[0:0] or_3270_nl;
  wire[0:0] nand_135_nl;
  wire[0:0] mux_2606_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] mux_2635_nl;
  wire[0:0] nand_408_nl;
  wire[0:0] mux_2634_nl;
  wire[0:0] mux_2633_nl;
  wire[0:0] mux_2632_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] mux_2631_nl;
  wire[0:0] and_552_nl;
  wire[0:0] and_553_nl;
  wire[0:0] mux_2630_nl;
  wire[0:0] mux_2629_nl;
  wire[0:0] and_815_nl;
  wire[0:0] and_822_nl;
  wire[0:0] mux_2628_nl;
  wire[0:0] nor_768_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] or_4081_nl;
  wire[0:0] mux_2627_nl;
  wire[0:0] mux_2626_nl;
  wire[0:0] mux_2625_nl;
  wire[0:0] or_3296_nl;
  wire[0:0] mux_2624_nl;
  wire[0:0] nand_232_nl;
  wire[0:0] mux_2623_nl;
  wire[0:0] mux_2622_nl;
  wire[0:0] nand_474_nl;
  wire[0:0] mux_2621_nl;
  wire[0:0] or_3287_nl;
  wire[0:0] mux_2650_nl;
  wire[0:0] mux_2649_nl;
  wire[0:0] or_3329_nl;
  wire[0:0] mux_2648_nl;
  wire[0:0] or_3328_nl;
  wire[0:0] or_3327_nl;
  wire[0:0] mux_2647_nl;
  wire[0:0] mux_2646_nl;
  wire[0:0] mux_2645_nl;
  wire[0:0] or_3325_nl;
  wire[0:0] mux_2644_nl;
  wire[0:0] nand_223_nl;
  wire[0:0] mux_2643_nl;
  wire[0:0] mux_2642_nl;
  wire[0:0] nand_396_nl;
  wire[0:0] mux_2641_nl;
  wire[0:0] or_3320_nl;
  wire[0:0] or_3319_nl;
  wire[0:0] mux_2640_nl;
  wire[0:0] mux_2639_nl;
  wire[0:0] mux_2638_nl;
  wire[0:0] or_3318_nl;
  wire[0:0] or_3316_nl;
  wire[0:0] mux_2637_nl;
  wire[0:0] nand_227_nl;
  wire[0:0] nand_228_nl;
  wire[0:0] nand_137_nl;
  wire[0:0] mux_2636_nl;
  wire[0:0] nor_762_nl;
  wire[0:0] nor_763_nl;
  wire[0:0] mux_2665_nl;
  wire[0:0] nand_407_nl;
  wire[0:0] mux_2664_nl;
  wire[0:0] mux_2663_nl;
  wire[0:0] mux_2662_nl;
  wire[0:0] nor_756_nl;
  wire[0:0] and_548_nl;
  wire[0:0] mux_2661_nl;
  wire[0:0] and_549_nl;
  wire[0:0] and_550_nl;
  wire[0:0] mux_2660_nl;
  wire[0:0] mux_2659_nl;
  wire[0:0] and_816_nl;
  wire[0:0] and_823_nl;
  wire[0:0] mux_2658_nl;
  wire[0:0] nor_759_nl;
  wire[0:0] nor_760_nl;
  wire[0:0] or_4080_nl;
  wire[0:0] mux_2657_nl;
  wire[0:0] mux_2656_nl;
  wire[0:0] mux_2655_nl;
  wire[0:0] or_3339_nl;
  wire[0:0] mux_2654_nl;
  wire[0:0] nand_218_nl;
  wire[0:0] mux_2653_nl;
  wire[0:0] mux_2652_nl;
  wire[0:0] nand_473_nl;
  wire[0:0] mux_2651_nl;
  wire[0:0] or_3330_nl;
  wire[0:0] mux_2680_nl;
  wire[0:0] mux_2679_nl;
  wire[0:0] or_3372_nl;
  wire[0:0] mux_2678_nl;
  wire[0:0] or_3371_nl;
  wire[0:0] or_3370_nl;
  wire[0:0] mux_2677_nl;
  wire[0:0] mux_2676_nl;
  wire[0:0] mux_2675_nl;
  wire[0:0] or_3368_nl;
  wire[0:0] mux_2674_nl;
  wire[0:0] nand_210_nl;
  wire[0:0] mux_2673_nl;
  wire[0:0] mux_2672_nl;
  wire[0:0] nand_394_nl;
  wire[0:0] mux_2671_nl;
  wire[0:0] or_3363_nl;
  wire[0:0] or_3362_nl;
  wire[0:0] mux_2670_nl;
  wire[0:0] mux_2669_nl;
  wire[0:0] mux_2668_nl;
  wire[0:0] nand_212_nl;
  wire[0:0] or_3359_nl;
  wire[0:0] mux_2667_nl;
  wire[0:0] nand_213_nl;
  wire[0:0] nand_214_nl;
  wire[0:0] nand_139_nl;
  wire[0:0] mux_2666_nl;
  wire[0:0] nor_754_nl;
  wire[0:0] nor_755_nl;
  wire[0:0] mux_2695_nl;
  wire[0:0] nand_406_nl;
  wire[0:0] mux_2694_nl;
  wire[0:0] mux_2693_nl;
  wire[0:0] mux_2692_nl;
  wire[0:0] and_539_nl;
  wire[0:0] and_540_nl;
  wire[0:0] mux_2691_nl;
  wire[0:0] and_541_nl;
  wire[0:0] and_542_nl;
  wire[0:0] mux_2690_nl;
  wire[0:0] mux_2689_nl;
  wire[0:0] and_817_nl;
  wire[0:0] and_824_nl;
  wire[0:0] mux_2688_nl;
  wire[0:0] and_543_nl;
  wire[0:0] and_544_nl;
  wire[0:0] or_4079_nl;
  wire[0:0] mux_2687_nl;
  wire[0:0] mux_2686_nl;
  wire[0:0] mux_2685_nl;
  wire[0:0] mux_2684_nl;
  wire[0:0] nand_203_nl;
  wire[0:0] mux_2683_nl;
  wire[0:0] mux_2682_nl;
  wire[0:0] nand_nl;
  wire[0:0] mux_2681_nl;
  wire[0:0] nand_205_nl;
  wire[0:0] mux_2710_nl;
  wire[0:0] mux_2709_nl;
  wire[0:0] or_3405_nl;
  wire[0:0] mux_2708_nl;
  wire[0:0] nand_192_nl;
  wire[0:0] nand_193_nl;
  wire[0:0] mux_2707_nl;
  wire[0:0] mux_2706_nl;
  wire[0:0] mux_2705_nl;
  wire[0:0] and_535_nl;
  wire[0:0] mux_2704_nl;
  wire[0:0] nand_194_nl;
  wire[0:0] mux_2703_nl;
  wire[0:0] mux_2702_nl;
  wire[0:0] nand_392_nl;
  wire[0:0] mux_2701_nl;
  wire[0:0] nand_196_nl;
  wire[0:0] or_3396_nl;
  wire[0:0] mux_2700_nl;
  wire[0:0] mux_2699_nl;
  wire[0:0] mux_2698_nl;
  wire[0:0] or_4002_nl;
  wire[0:0] nand_198_nl;
  wire[0:0] mux_2697_nl;
  wire[0:0] nand_199_nl;
  wire[0:0] nand_200_nl;
  wire[0:0] nand_141_nl;
  wire[0:0] mux_2696_nl;
  wire[0:0] and_536_nl;
  wire[0:0] and_537_nl;
  wire[0:0] mux_2717_nl;
  wire[0:0] mux_2716_nl;
  wire[0:0] mux_2715_nl;
  wire[0:0] nor_743_nl;
  wire[0:0] nor_744_nl;
  wire[0:0] mux_2714_nl;
  wire[0:0] nor_745_nl;
  wire[0:0] mux_2713_nl;
  wire[0:0] mux_2712_nl;
  wire[0:0] nor_747_nl;
  wire[0:0] mux_2711_nl;
  wire[0:0] nor_749_nl;
  wire[0:0] nor_750_nl;
  wire[0:0] mux_2720_nl;
  wire[0:0] mux_2719_nl;
  wire[0:0] nor_739_nl;
  wire[0:0] mux_2718_nl;
  wire[0:0] nor_742_nl;
  wire[0:0] mux_2725_nl;
  wire[0:0] mux_2724_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] mux_2723_nl;
  wire[0:0] mux_2722_nl;
  wire[0:0] nor_736_nl;
  wire[0:0] mux_2721_nl;
  wire[0:0] mux_2728_nl;
  wire[0:0] mux_2727_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] mux_2726_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] mux_2734_nl;
  wire[0:0] mux_2733_nl;
  wire[0:0] mux_2732_nl;
  wire[0:0] nor_722_nl;
  wire[0:0] nor_723_nl;
  wire[0:0] mux_2731_nl;
  wire[0:0] nor_724_nl;
  wire[0:0] nor_725_nl;
  wire[0:0] mux_2730_nl;
  wire[0:0] nor_726_nl;
  wire[0:0] mux_2729_nl;
  wire[0:0] nor_727_nl;
  wire[0:0] nor_728_nl;
  wire[0:0] mux_2737_nl;
  wire[0:0] mux_2736_nl;
  wire[0:0] nor_718_nl;
  wire[0:0] mux_2735_nl;
  wire[0:0] nor_721_nl;
  wire[0:0] mux_2742_nl;
  wire[0:0] mux_2741_nl;
  wire[0:0] nor_712_nl;
  wire[0:0] mux_2740_nl;
  wire[0:0] mux_2739_nl;
  wire[0:0] nor_715_nl;
  wire[0:0] mux_2738_nl;
  wire[0:0] mux_2745_nl;
  wire[0:0] mux_2744_nl;
  wire[0:0] nor_708_nl;
  wire[0:0] mux_2743_nl;
  wire[0:0] nor_711_nl;
  wire[0:0] mux_2752_nl;
  wire[0:0] mux_2751_nl;
  wire[0:0] mux_2750_nl;
  wire[0:0] nor_700_nl;
  wire[0:0] nor_701_nl;
  wire[0:0] mux_2749_nl;
  wire[0:0] nor_702_nl;
  wire[0:0] mux_2748_nl;
  wire[0:0] mux_2747_nl;
  wire[0:0] nor_704_nl;
  wire[0:0] mux_2746_nl;
  wire[0:0] nor_706_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] mux_2755_nl;
  wire[0:0] mux_2754_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] mux_2753_nl;
  wire[0:0] nor_699_nl;
  wire[0:0] mux_2760_nl;
  wire[0:0] mux_2759_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] mux_2758_nl;
  wire[0:0] mux_2757_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] mux_2756_nl;
  wire[0:0] mux_2763_nl;
  wire[0:0] mux_2762_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] mux_2761_nl;
  wire[0:0] nor_689_nl;
  wire[0:0] mux_2769_nl;
  wire[0:0] mux_2768_nl;
  wire[0:0] mux_2767_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_2766_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] mux_2765_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] mux_2764_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] mux_2772_nl;
  wire[0:0] mux_2771_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] mux_2770_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] mux_2777_nl;
  wire[0:0] mux_2776_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] mux_2775_nl;
  wire[0:0] mux_2774_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] mux_2773_nl;
  wire[0:0] mux_2780_nl;
  wire[0:0] mux_2779_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] mux_2778_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] mux_2787_nl;
  wire[0:0] mux_2786_nl;
  wire[0:0] mux_2785_nl;
  wire[0:0] nor_657_nl;
  wire[0:0] nor_658_nl;
  wire[0:0] mux_2784_nl;
  wire[0:0] nor_659_nl;
  wire[0:0] mux_2783_nl;
  wire[0:0] mux_2782_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] mux_2781_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] mux_2790_nl;
  wire[0:0] mux_2789_nl;
  wire[0:0] nor_653_nl;
  wire[0:0] mux_2788_nl;
  wire[0:0] nor_656_nl;
  wire[0:0] mux_2795_nl;
  wire[0:0] mux_2794_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] mux_2793_nl;
  wire[0:0] mux_2792_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_2791_nl;
  wire[0:0] mux_2798_nl;
  wire[0:0] mux_2797_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] mux_2796_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] mux_2804_nl;
  wire[0:0] mux_2803_nl;
  wire[0:0] mux_2802_nl;
  wire[0:0] nor_636_nl;
  wire[0:0] nor_637_nl;
  wire[0:0] mux_2801_nl;
  wire[0:0] nor_638_nl;
  wire[0:0] nor_639_nl;
  wire[0:0] mux_2800_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] mux_2799_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] mux_2807_nl;
  wire[0:0] mux_2806_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_2805_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] mux_2812_nl;
  wire[0:0] mux_2811_nl;
  wire[0:0] nor_626_nl;
  wire[0:0] mux_2810_nl;
  wire[0:0] mux_2809_nl;
  wire[0:0] nor_629_nl;
  wire[0:0] mux_2808_nl;
  wire[0:0] mux_2815_nl;
  wire[0:0] mux_2814_nl;
  wire[0:0] nor_622_nl;
  wire[0:0] mux_2813_nl;
  wire[0:0] nor_625_nl;
  wire[0:0] mux_2822_nl;
  wire[0:0] mux_2821_nl;
  wire[0:0] mux_2820_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] mux_2819_nl;
  wire[0:0] nor_616_nl;
  wire[0:0] mux_2818_nl;
  wire[0:0] mux_2817_nl;
  wire[0:0] nor_618_nl;
  wire[0:0] mux_2816_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] mux_2825_nl;
  wire[0:0] mux_2824_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] mux_2823_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] mux_2830_nl;
  wire[0:0] mux_2829_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] mux_2828_nl;
  wire[0:0] mux_2827_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] mux_2826_nl;
  wire[0:0] mux_2833_nl;
  wire[0:0] mux_2832_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] mux_2831_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] mux_2839_nl;
  wire[0:0] mux_2838_nl;
  wire[0:0] mux_2837_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] nor_594_nl;
  wire[0:0] mux_2836_nl;
  wire[0:0] nor_595_nl;
  wire[0:0] nor_596_nl;
  wire[0:0] mux_2835_nl;
  wire[0:0] nor_597_nl;
  wire[0:0] mux_2834_nl;
  wire[0:0] nor_598_nl;
  wire[0:0] nor_599_nl;
  wire[0:0] mux_2842_nl;
  wire[0:0] mux_2841_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] mux_2840_nl;
  wire[0:0] nor_592_nl;
  wire[0:0] mux_2847_nl;
  wire[0:0] mux_2846_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] mux_2845_nl;
  wire[0:0] mux_2844_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] mux_2843_nl;
  wire[0:0] mux_2850_nl;
  wire[0:0] mux_2849_nl;
  wire[0:0] nor_581_nl;
  wire[0:0] mux_2848_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] mux_2857_nl;
  wire[0:0] mux_2856_nl;
  wire[0:0] mux_2855_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] mux_2854_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] mux_2853_nl;
  wire[0:0] mux_2852_nl;
  wire[0:0] nor_577_nl;
  wire[0:0] mux_2851_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] mux_2860_nl;
  wire[0:0] mux_2859_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] mux_2858_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] mux_2865_nl;
  wire[0:0] mux_2864_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] mux_2863_nl;
  wire[0:0] mux_2862_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] mux_2861_nl;
  wire[0:0] mux_2868_nl;
  wire[0:0] mux_2867_nl;
  wire[0:0] nor_559_nl;
  wire[0:0] mux_2866_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] mux_2874_nl;
  wire[0:0] mux_2873_nl;
  wire[0:0] mux_2872_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] mux_2871_nl;
  wire[0:0] nor_554_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] mux_2870_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_2869_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] nor_558_nl;
  wire[0:0] mux_2877_nl;
  wire[0:0] mux_2876_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] mux_2875_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] mux_2882_nl;
  wire[0:0] mux_2881_nl;
  wire[0:0] nor_542_nl;
  wire[0:0] mux_2880_nl;
  wire[0:0] mux_2879_nl;
  wire[0:0] nor_545_nl;
  wire[0:0] mux_2878_nl;
  wire[0:0] mux_2885_nl;
  wire[0:0] mux_2884_nl;
  wire[0:0] nor_538_nl;
  wire[0:0] mux_2883_nl;
  wire[0:0] nor_541_nl;
  wire[0:0] mux_2892_nl;
  wire[0:0] mux_2891_nl;
  wire[0:0] mux_2890_nl;
  wire[0:0] nor_530_nl;
  wire[0:0] nor_531_nl;
  wire[0:0] mux_2889_nl;
  wire[0:0] nor_532_nl;
  wire[0:0] mux_2888_nl;
  wire[0:0] mux_2887_nl;
  wire[0:0] nor_534_nl;
  wire[0:0] mux_2886_nl;
  wire[0:0] nor_536_nl;
  wire[0:0] nor_537_nl;
  wire[0:0] mux_2895_nl;
  wire[0:0] mux_2894_nl;
  wire[0:0] nor_526_nl;
  wire[0:0] mux_2893_nl;
  wire[0:0] nor_529_nl;
  wire[0:0] mux_2900_nl;
  wire[0:0] mux_2899_nl;
  wire[0:0] nor_520_nl;
  wire[0:0] mux_2898_nl;
  wire[0:0] mux_2897_nl;
  wire[0:0] nor_523_nl;
  wire[0:0] mux_2896_nl;
  wire[0:0] mux_2903_nl;
  wire[0:0] mux_2902_nl;
  wire[0:0] nor_516_nl;
  wire[0:0] mux_2901_nl;
  wire[0:0] nor_519_nl;
  wire[0:0] mux_2909_nl;
  wire[0:0] mux_2908_nl;
  wire[0:0] mux_2907_nl;
  wire[0:0] nor_509_nl;
  wire[0:0] nor_510_nl;
  wire[0:0] mux_2906_nl;
  wire[0:0] nor_511_nl;
  wire[0:0] nor_512_nl;
  wire[0:0] mux_2905_nl;
  wire[0:0] nor_513_nl;
  wire[0:0] mux_2904_nl;
  wire[0:0] nor_514_nl;
  wire[0:0] nor_515_nl;
  wire[0:0] mux_2912_nl;
  wire[0:0] mux_2911_nl;
  wire[0:0] nor_505_nl;
  wire[0:0] mux_2910_nl;
  wire[0:0] nor_508_nl;
  wire[0:0] mux_2917_nl;
  wire[0:0] mux_2916_nl;
  wire[0:0] nor_499_nl;
  wire[0:0] mux_2915_nl;
  wire[0:0] mux_2914_nl;
  wire[0:0] nor_502_nl;
  wire[0:0] mux_2913_nl;
  wire[0:0] mux_2920_nl;
  wire[0:0] mux_2919_nl;
  wire[0:0] nor_497_nl;
  wire[0:0] mux_2918_nl;
  wire[0:0] nor_498_nl;
  wire[0:0] mux_2927_nl;
  wire[0:0] mux_2926_nl;
  wire[0:0] mux_2925_nl;
  wire[0:0] nor_489_nl;
  wire[0:0] nor_490_nl;
  wire[0:0] mux_2924_nl;
  wire[0:0] nor_491_nl;
  wire[0:0] mux_2923_nl;
  wire[0:0] mux_2922_nl;
  wire[0:0] nor_493_nl;
  wire[0:0] mux_2921_nl;
  wire[0:0] nor_495_nl;
  wire[0:0] nor_496_nl;
  wire[0:0] mux_2930_nl;
  wire[0:0] mux_2929_nl;
  wire[0:0] nor_485_nl;
  wire[0:0] mux_2928_nl;
  wire[0:0] nor_488_nl;
  wire[0:0] mux_2935_nl;
  wire[0:0] mux_2934_nl;
  wire[0:0] nor_479_nl;
  wire[0:0] mux_2933_nl;
  wire[0:0] mux_2932_nl;
  wire[0:0] nor_482_nl;
  wire[0:0] mux_2931_nl;
  wire[0:0] mux_2938_nl;
  wire[0:0] mux_2937_nl;
  wire[0:0] nor_475_nl;
  wire[0:0] mux_2936_nl;
  wire[0:0] nor_478_nl;
  wire[0:0] mux_2944_nl;
  wire[0:0] mux_2943_nl;
  wire[0:0] mux_2942_nl;
  wire[0:0] nor_468_nl;
  wire[0:0] nor_469_nl;
  wire[0:0] mux_2941_nl;
  wire[0:0] nor_470_nl;
  wire[0:0] nor_471_nl;
  wire[0:0] mux_2940_nl;
  wire[0:0] nor_472_nl;
  wire[0:0] mux_2939_nl;
  wire[0:0] nor_473_nl;
  wire[0:0] nor_474_nl;
  wire[0:0] mux_2947_nl;
  wire[0:0] mux_2946_nl;
  wire[0:0] nor_464_nl;
  wire[0:0] mux_2945_nl;
  wire[0:0] nor_467_nl;
  wire[0:0] mux_2952_nl;
  wire[0:0] mux_2951_nl;
  wire[0:0] nor_458_nl;
  wire[0:0] mux_2950_nl;
  wire[0:0] mux_2949_nl;
  wire[0:0] nor_461_nl;
  wire[0:0] mux_2948_nl;
  wire[0:0] mux_2955_nl;
  wire[0:0] mux_2954_nl;
  wire[0:0] nor_456_nl;
  wire[0:0] mux_2953_nl;
  wire[0:0] nor_457_nl;
  wire[0:0] mux_2962_nl;
  wire[0:0] mux_2961_nl;
  wire[0:0] mux_2960_nl;
  wire[0:0] nor_449_nl;
  wire[0:0] nor_450_nl;
  wire[0:0] mux_2959_nl;
  wire[0:0] and_528_nl;
  wire[0:0] mux_2958_nl;
  wire[0:0] mux_2957_nl;
  wire[0:0] nor_452_nl;
  wire[0:0] mux_2956_nl;
  wire[0:0] nor_454_nl;
  wire[0:0] nor_455_nl;
  wire[0:0] mux_2965_nl;
  wire[0:0] mux_2964_nl;
  wire[0:0] nor_445_nl;
  wire[0:0] mux_2963_nl;
  wire[0:0] nor_448_nl;
  wire[0:0] mux_2970_nl;
  wire[0:0] mux_2969_nl;
  wire[0:0] nor_439_nl;
  wire[0:0] mux_2968_nl;
  wire[0:0] mux_2967_nl;
  wire[0:0] nor_442_nl;
  wire[0:0] mux_2966_nl;
  wire[0:0] mux_2973_nl;
  wire[0:0] mux_2972_nl;
  wire[0:0] nor_437_nl;
  wire[0:0] mux_2971_nl;
  wire[0:0] nor_438_nl;
  wire[0:0] mux_2979_nl;
  wire[0:0] mux_2978_nl;
  wire[0:0] mux_2977_nl;
  wire[0:0] and_789_nl;
  wire[0:0] and_810_nl;
  wire[0:0] mux_2976_nl;
  wire[0:0] nor_433_nl;
  wire[0:0] nor_434_nl;
  wire[0:0] mux_2975_nl;
  wire[0:0] nor_435_nl;
  wire[0:0] mux_2974_nl;
  wire[0:0] and_525_nl;
  wire[0:0] nor_436_nl;
  wire[0:0] mux_2982_nl;
  wire[0:0] mux_2981_nl;
  wire[0:0] nor_429_nl;
  wire[0:0] mux_2980_nl;
  wire[0:0] nor_430_nl;
  wire[0:0] mux_2987_nl;
  wire[0:0] mux_2986_nl;
  wire[0:0] and_790_nl;
  wire[0:0] mux_2985_nl;
  wire[0:0] mux_2984_nl;
  wire[0:0] and_520_nl;
  wire[0:0] mux_2983_nl;
  wire[0:0] mux_2990_nl;
  wire[0:0] mux_2989_nl;
  wire[0:0] nor_427_nl;
  wire[0:0] mux_2988_nl;
  wire[0:0] and_517_nl;
  wire[6:0] COMP_LOOP_mux_721_nl;
  wire[0:0] and_1047_nl;
  wire[11:0] acc_1_nl;
  wire[12:0] nl_acc_1_nl;
  wire[10:0] COMP_LOOP_mux_722_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_nand_1_nl;
  wire[9:0] COMP_LOOP_mux_723_nl;
  wire[3:0] STAGE_LOOP_mux_4_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_and_337_nl;
  wire[0:0] COMP_LOOP_tmp_mux_64_nl;
  wire[8:0] COMP_LOOP_tmp_mux1h_146_nl;
  wire[0:0] COMP_LOOP_tmp_or_88_nl;
  wire[0:0] COMP_LOOP_tmp_and_312_nl;
  wire[5:0] COMP_LOOP_tmp_mux1h_147_nl;
  wire[0:0] COMP_LOOP_tmp_or_89_nl;
  wire[0:0] COMP_LOOP_tmp_or_90_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_mux_17_nl;
  wire[0:0] COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl;
  wire[63:0] COMP_LOOP_tmp_mux1h_148_nl;
  wire[0:0] and_1048_nl;
  wire[63:0] COMP_LOOP_tmp_mux_65_nl;
  wire[0:0] COMP_LOOP_tmp_or_91_nl;
  wire[0:0] COMP_LOOP_mux1h_1267_nl;
  wire[0:0] COMP_LOOP_mux1h_1268_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1890_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1891_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1892_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1893_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1894_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1895_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1896_nl;
  wire[0:0] COMP_LOOP_mux1h_1269_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1897_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1898_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1899_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1900_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1901_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1902_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1903_nl;
  wire[0:0] COMP_LOOP_mux1h_1270_nl;
  wire[0:0] COMP_LOOP_mux1h_1271_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1904_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1905_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1906_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1907_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1908_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1909_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1910_nl;
  wire[0:0] COMP_LOOP_mux1h_1272_nl;
  wire[0:0] COMP_LOOP_mux1h_1273_nl;
  wire[0:0] COMP_LOOP_mux1h_1274_nl;
  wire[0:0] COMP_LOOP_mux1h_1275_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1911_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1912_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1913_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1914_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1915_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1916_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1917_nl;
  wire[0:0] COMP_LOOP_mux1h_1276_nl;
  wire[0:0] COMP_LOOP_mux1h_1277_nl;
  wire[0:0] COMP_LOOP_mux1h_1278_nl;
  wire[0:0] COMP_LOOP_mux1h_1279_nl;
  wire[0:0] COMP_LOOP_mux1h_1280_nl;
  wire[0:0] COMP_LOOP_mux1h_1281_nl;
  wire[0:0] COMP_LOOP_mux1h_1282_nl;
  wire[0:0] COMP_LOOP_mux1h_1283_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1918_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1919_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1920_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1921_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1922_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1923_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1924_nl;
  wire[0:0] COMP_LOOP_mux1h_1284_nl;
  wire[0:0] COMP_LOOP_mux1h_1285_nl;
  wire[0:0] COMP_LOOP_mux1h_1286_nl;
  wire[0:0] COMP_LOOP_mux1h_1287_nl;
  wire[0:0] COMP_LOOP_mux1h_1288_nl;
  wire[0:0] COMP_LOOP_mux1h_1289_nl;
  wire[0:0] COMP_LOOP_mux1h_1290_nl;
  wire[0:0] COMP_LOOP_mux1h_1291_nl;
  wire[0:0] COMP_LOOP_mux1h_1292_nl;
  wire[0:0] COMP_LOOP_mux1h_1293_nl;
  wire[0:0] COMP_LOOP_mux1h_1294_nl;
  wire[0:0] COMP_LOOP_mux1h_1295_nl;
  wire[0:0] COMP_LOOP_mux1h_1296_nl;
  wire[0:0] COMP_LOOP_mux1h_1297_nl;
  wire[0:0] COMP_LOOP_mux1h_1298_nl;
  wire[0:0] COMP_LOOP_mux1h_1299_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1925_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1926_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1927_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1928_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1929_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1930_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_1931_nl;
  wire[0:0] COMP_LOOP_mux1h_1300_nl;
  wire[0:0] COMP_LOOP_mux1h_1301_nl;
  wire[0:0] COMP_LOOP_mux1h_1302_nl;
  wire[0:0] COMP_LOOP_mux1h_1303_nl;
  wire[0:0] COMP_LOOP_mux1h_1304_nl;
  wire[0:0] COMP_LOOP_mux1h_1305_nl;
  wire[0:0] COMP_LOOP_mux1h_1306_nl;
  wire[0:0] COMP_LOOP_mux1h_1307_nl;
  wire[0:0] COMP_LOOP_mux1h_1308_nl;
  wire[0:0] COMP_LOOP_mux1h_1309_nl;
  wire[0:0] COMP_LOOP_mux1h_1310_nl;
  wire[0:0] COMP_LOOP_mux1h_1311_nl;
  wire[0:0] COMP_LOOP_mux1h_1312_nl;
  wire[0:0] COMP_LOOP_mux1h_1313_nl;
  wire[0:0] COMP_LOOP_mux1h_1314_nl;
  wire[0:0] COMP_LOOP_mux1h_1315_nl;
  wire[0:0] COMP_LOOP_mux1h_1316_nl;
  wire[0:0] COMP_LOOP_mux1h_1317_nl;
  wire[0:0] COMP_LOOP_mux1h_1318_nl;
  wire[0:0] COMP_LOOP_mux1h_1319_nl;
  wire[0:0] COMP_LOOP_mux1h_1320_nl;
  wire[0:0] COMP_LOOP_mux1h_1321_nl;
  wire[0:0] COMP_LOOP_mux1h_1322_nl;
  wire[0:0] COMP_LOOP_mux1h_1323_nl;
  wire[0:0] COMP_LOOP_mux1h_1324_nl;
  wire[0:0] COMP_LOOP_mux1h_1325_nl;
  wire[0:0] COMP_LOOP_mux1h_1326_nl;
  wire[0:0] COMP_LOOP_mux1h_1327_nl;
  wire[0:0] COMP_LOOP_mux1h_1328_nl;
  wire[0:0] COMP_LOOP_mux1h_1329_nl;
  wire[0:0] COMP_LOOP_mux1h_1330_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[64:0] acc_4_nl;
  wire[65:0] nl_acc_4_nl;
  wire[63:0] COMP_LOOP_COMP_LOOP_mux_22_nl;
  wire[0:0] and_372_nl;
  wire[0:0] mux_3002_nl;
  wire[0:0] mux_3001_nl;
  wire[0:0] mux_3000_nl;
  wire[0:0] mux_2999_nl;
  wire[0:0] mux_2998_nl;
  wire[0:0] or_3835_nl;
  wire[0:0] COMP_LOOP_or_169_nl;
  wire [63:0] nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat;
  assign COMP_LOOP_COMP_LOOP_mux_22_nl = MUX_v_64_2_2((~ COMP_LOOP_1_acc_8_itm),
      (~ z_out_9), COMP_LOOP_or_65_itm);
  assign nl_acc_4_nl = ({COMP_LOOP_mux_724_cse , 1'b1}) + ({COMP_LOOP_COMP_LOOP_mux_22_nl
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[64:0];
  assign mux_3000_nl = MUX_s_1_2_2(or_tmp_3721, mux_tmp_2924, fsm_output[6]);
  assign mux_3001_nl = MUX_s_1_2_2(mux_3000_nl, or_tmp_3718, fsm_output[2]);
  assign or_3835_nl = (~ (fsm_output[4])) | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2998_nl = MUX_s_1_2_2(mux_tmp_2924, or_3835_nl, fsm_output[6]);
  assign mux_2999_nl = MUX_s_1_2_2(or_tmp_3718, mux_2998_nl, fsm_output[2]);
  assign mux_3002_nl = MUX_s_1_2_2(mux_3001_nl, mux_2999_nl, fsm_output[5]);
  assign and_372_nl = (~ mux_3002_nl) & and_dcpl_340;
  assign COMP_LOOP_or_169_nl = (and_dcpl_92 & and_dcpl_57) | (and_dcpl_262 & and_dcpl_344)
      | (and_dcpl_262 & and_dcpl_347) | (and_dcpl_60 & and_dcpl_64) | (and_dcpl_66
      & and_dcpl_57) | (and_dcpl_355 & and_dcpl_110) | (and_dcpl_355 & and_dcpl_113)
      | (and_dcpl_353 & and_dcpl_116);
  assign nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat = MUX1HOT_v_64_3_2((readslicef_65_64_1(acc_4_nl)),
      COMP_LOOP_1_acc_8_itm, z_out_8, {COMP_LOOP_or_68_itm , and_372_nl , COMP_LOOP_or_169_nl});
  wire [63:0] nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat;
  assign nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat = p_sva;
  wire[0:0] mux_3012_nl;
  wire[0:0] mux_3011_nl;
  wire[0:0] mux_3010_nl;
  wire[0:0] or_3846_nl;
  wire[0:0] mux_3009_nl;
  wire[0:0] or_3845_nl;
  wire[0:0] mux_3008_nl;
  wire[0:0] mux_3007_nl;
  wire[0:0] or_3842_nl;
  wire[0:0] mux_3005_nl;
  wire[0:0] or_3840_nl;
  wire [0:0] nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat;
  assign mux_3009_nl = MUX_s_1_2_2(or_364_cse, and_735_cse, fsm_output[0]);
  assign or_3846_nl = (fsm_output[3]) | (~ mux_3009_nl);
  assign mux_3010_nl = MUX_s_1_2_2(or_3846_nl, nand_tmp_142, fsm_output[6]);
  assign or_3845_nl = (fsm_output[6]) | mux_tmp_2939;
  assign mux_3011_nl = MUX_s_1_2_2(mux_3010_nl, or_3845_nl, fsm_output[5]);
  assign or_3842_nl = (fsm_output[3]) | (fsm_output[0]) | (~ and_735_cse);
  assign mux_3007_nl = MUX_s_1_2_2(mux_tmp_2939, or_3842_nl, fsm_output[6]);
  assign or_3840_nl = (fsm_output[3]) | (~((~ (fsm_output[0])) | (fsm_output[4])))
      | (fsm_output[7]);
  assign mux_3005_nl = MUX_s_1_2_2(nand_tmp_142, or_3840_nl, fsm_output[6]);
  assign mux_3008_nl = MUX_s_1_2_2(mux_3007_nl, mux_3005_nl, fsm_output[5]);
  assign mux_3012_nl = MUX_s_1_2_2(mux_3011_nl, mux_3008_nl, fsm_output[2]);
  assign nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat = ~(mux_3012_nl |
      (fsm_output[1]));
  wire[0:0] and_835_nl;
  wire [3:0] nl_COMP_LOOP_5_tmp_lshift_rg_s;
  assign and_835_nl = (fsm_output==8'b00000010);
  assign nl_COMP_LOOP_5_tmp_lshift_rg_s = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, z_out_4,
      and_835_nl);
  wire[0:0] COMP_LOOP_tmp_or_56_nl;
  wire [3:0] nl_COMP_LOOP_1_tmp_lshift_rg_s;
  assign COMP_LOOP_tmp_or_56_nl = ((~ (fsm_output[4])) & (fsm_output[0]) & nor_1715_cse
      & (fsm_output[2:1]==2'b01) & nor_1716_cse) | ((~ (fsm_output[4])) & (~ (fsm_output[0]))
      & nor_1715_cse & (fsm_output[2:1]==2'b10) & nor_1716_cse);
  assign nl_COMP_LOOP_1_tmp_lshift_rg_s = MUX_v_4_2_2(z_out_4, COMP_LOOP_1_tmp_acc_cse_sva,
      COMP_LOOP_tmp_or_56_nl);
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0 = ~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0 = ~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0 = ~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0 = ~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0 = ~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0 = ~ COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm;
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out_3[10];
  wire [0:0] nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0 = ~ (z_out_2[4]);
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_63_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_63_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_62_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_62_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_61_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_61_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_60_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_60_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_59_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_59_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_58_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_58_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_57_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_57_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_56_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_56_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_55_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_55_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_54_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_54_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_53_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_53_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_52_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_52_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_51_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_51_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_50_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_50_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_49_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_49_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_48_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_48_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_47_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_47_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_46_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_46_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_45_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_45_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_44_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_44_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_43_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_43_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_42_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_42_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_41_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_41_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_40_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_40_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_39_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_39_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_38_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_38_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_37_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_37_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_36_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_36_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_35_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_35_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_34_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_34_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_33_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_33_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_32_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_32_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_31_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_30_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_29_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_28_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_27_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_26_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_25_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_24_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_23_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_22_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_21_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_20_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_19_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_18_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_17_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_16_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_63_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_63_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_62_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_62_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_61_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_61_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_60_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_60_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_59_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_59_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_58_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_58_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_57_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_57_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_56_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_56_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_55_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_55_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_54_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_54_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_53_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_53_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_52_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_52_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_51_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_51_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_50_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_50_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_49_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_49_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_48_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_48_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_47_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_47_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_46_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_46_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_45_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_45_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_44_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_44_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_43_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_43_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_42_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_42_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_41_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_41_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_40_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_40_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_39_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_39_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_38_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_38_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_37_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_37_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_36_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_36_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_35_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_35_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_34_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_34_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_33_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_33_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_32_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_32_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_31_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_30_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_29_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_28_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_27_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_26_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_25_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_24_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_23_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_22_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_21_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_20_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_19_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_18_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_17_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_16_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_63_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_0_lz)
    );
  modulo_dev  COMP_LOOP_1_modulo_dev_cmp (
      .base_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_base_rsc_dat[63:0]),
      .m_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_m_rsc_dat[63:0]),
      .return_rsc_z(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z),
      .ccs_ccore_start_rsc_dat(nl_COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_start_rsc_dat[0:0]),
      .ccs_ccore_clk(clk),
      .ccs_ccore_srst(rst),
      .ccs_ccore_en(COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd11)) COMP_LOOP_5_tmp_lshift_rg (
      .a(1'b1),
      .s(nl_COMP_LOOP_5_tmp_lshift_rg_s[3:0]),
      .z(z_out)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) COMP_LOOP_1_tmp_lshift_rg (
      .a(1'b1),
      .s(nl_COMP_LOOP_1_tmp_lshift_rg_s[3:0]),
      .z(z_out_1)
    );
  inPlaceNTT_DIF_core_wait_dp inPlaceNTT_DIF_core_wait_dp_inst (
      .ensig_cgo_iro(mux_2997_rmff),
      .ensig_cgo(reg_ensig_cgo_cse),
      .COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en(COMP_LOOP_1_modulo_dev_cmp_ccs_ccore_en)
    );
  inPlaceNTT_DIF_core_core_fsm inPlaceNTT_DIF_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .COMP_LOOP_C_28_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_28_tr0[0:0]),
      .COMP_LOOP_C_56_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_56_tr0[0:0]),
      .COMP_LOOP_C_84_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_84_tr0[0:0]),
      .COMP_LOOP_C_112_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_112_tr0[0:0]),
      .COMP_LOOP_C_140_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_140_tr0[0:0]),
      .COMP_LOOP_C_168_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_168_tr0[0:0]),
      .COMP_LOOP_C_196_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_196_tr0[0:0]),
      .COMP_LOOP_C_224_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_COMP_LOOP_C_224_tr0[0:0]),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_1_tr0(nl_inPlaceNTT_DIF_core_core_fsm_inst_STAGE_LOOP_C_1_tr0[0:0])
    );
  assign or_595_cse = (fsm_output[4:3]!=2'b00);
  assign nand_191_cse = ~((z_out_7[0]) & (fsm_output[3]));
  assign nand_190_cse = ~((z_out_7[1:0]==2'b11) & (fsm_output[3]));
  assign nand_188_cse = ~((z_out_7[2:0]==3'b111) & (fsm_output[3]));
  assign nand_184_cse = ~((z_out_7[3:0]==4'b1111) & (fsm_output[3]));
  assign nand_174_cse = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4]) & (fsm_output[3]));
  assign nand_175_cse = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5]) & (fsm_output[3]));
  assign mux_2995_nl = MUX_s_1_2_2(mux_tmp_2924, mux_tmp_2927, fsm_output[6]);
  assign mux_2996_nl = MUX_s_1_2_2(or_tmp_3718, mux_2995_nl, fsm_output[2]);
  assign nor_425_nl = ~((~((fsm_output[4:3]!=2'b10))) | (fsm_output[7]));
  assign mux_2992_nl = MUX_s_1_2_2(mux_tmp_2924, nor_425_nl, fsm_output[6]);
  assign mux_2993_nl = MUX_s_1_2_2(mux_2992_nl, (~ and_705_cse), fsm_output[2]);
  assign mux_2997_rmff = MUX_s_1_2_2(mux_2996_nl, mux_2993_nl, fsm_output[5]);
  assign or_4007_cse = (fsm_output[4]) | (fsm_output[0]) | (fsm_output[3]);
  assign and_78_cse = (fsm_output[6]) & or_4007_cse & (fsm_output[7]);
  assign nor_1744_cse = ~((fsm_output[2:1]!=2'b00));
  assign and_1046_cse = (fsm_output[1:0]==2'b11);
  assign mux_3029_nl = MUX_s_1_2_2(mux_tmp_2959, mux_tmp_2961, fsm_output[2]);
  assign mux_3030_nl = MUX_s_1_2_2(mux_3029_nl, mux_tmp_2960, fsm_output[1]);
  assign mux_3031_nl = MUX_s_1_2_2(mux_3030_nl, (fsm_output[6]), fsm_output[5]);
  assign COMP_LOOP_or_121_cse = mux_3031_nl | (fsm_output[7]);
  assign and_507_cse = (fsm_output[2:1]==2'b11);
  assign nor_1674_cse = ~((fsm_output[2]) | (fsm_output[6]));
  assign COMP_LOOP_or_120_rgt = and_dcpl_259 | and_dcpl_260 | and_dcpl_263;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse = (z_out_7[5:0]==6'b001011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse = (z_out_7[5:0]==6'b001010);
  assign COMP_LOOP_tmp_nor_67_cse = ~((z_out_7[4]) | (z_out_7[2]) | (z_out_7[1]));
  assign mux_3044_nl = MUX_s_1_2_2(mux_tmp_2976, mux_tmp_2975, fsm_output[1]);
  assign mux_3045_nl = MUX_s_1_2_2(mux_3044_nl, (~ mux_180_cse), fsm_output[5]);
  assign COMP_LOOP_or_126_cse = ~(mux_3045_nl & (~ (fsm_output[7])));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse = (z_out_7[3]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_67_cse;
  assign nor_358_cse = ~((fsm_output[5]) | (~ (fsm_output[0])));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse = (z_out_7[5:0]==6'b001100);
  assign COMP_LOOP_tmp_nor_68_cse = ~((z_out_7[4]) | (z_out_7[2]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse = (z_out_7[3]) & (z_out_7[1]) & COMP_LOOP_tmp_nor_68_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse = (z_out_7[5:0]==6'b001101);
  assign COMP_LOOP_tmp_nor_69_cse = ~((z_out_7[4]) | (z_out_7[2]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse = (z_out_7[3]) & (z_out_7[1]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_69_cse;
  assign or_341_cse = (fsm_output[4]) | (fsm_output[6]);
  assign and_677_cse = (fsm_output[3]) & (fsm_output[4]) & (fsm_output[6]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse = (z_out_7[5:0]==6'b001110);
  assign COMP_LOOP_tmp_nor_70_cse = ~((z_out_7[4]) | (z_out_7[1]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse = (z_out_7[3:2]==2'b11) & COMP_LOOP_tmp_nor_70_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse = (z_out_7[5:0]==6'b001111);
  assign COMP_LOOP_tmp_nor_71_cse = ~((z_out_7[4]) | (z_out_7[1]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse = (z_out_7[3]) & (z_out_7[2]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_71_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse = (z_out_7[5:0]==6'b010001);
  assign COMP_LOOP_tmp_nor_72_cse = ~((z_out_7[4]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse = (z_out_7[3:1]==3'b111) & COMP_LOOP_tmp_nor_72_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse = (z_out_7[5:0]==6'b010101);
  assign COMP_LOOP_tmp_nor_76_cse = ~((z_out_7[3:2]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse = (z_out_7[5:0]==6'b010100);
  assign COMP_LOOP_or_135_cse = MUX_s_1_2_2(mux_tmp_3003, (fsm_output[7]), fsm_output[5]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse = (z_out_7[4]) & (z_out_7[1]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_76_cse;
  assign and_640_cse = (fsm_output[4:3]==2'b11);
  assign and_639_cse = (fsm_output[3]) & (fsm_output[0]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse = (z_out_7[5:0]==6'b010110);
  assign COMP_LOOP_tmp_nor_77_cse = ~((z_out_7[3]) | (z_out_7[1]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse = (z_out_7[4]) & (z_out_7[2]) & COMP_LOOP_tmp_nor_77_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse = (z_out_7[5:0]==6'b010111);
  assign COMP_LOOP_tmp_nor_78_cse = ~((z_out_7[3]) | (z_out_7[1]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse = (z_out_7[4]) & (z_out_7[2]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_78_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse = (z_out_7[5:0]==6'b011000);
  assign COMP_LOOP_tmp_nor_79_cse = ~((z_out_7[3]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse = (z_out_7[4]) & (z_out_7[2]) & (z_out_7[1])
      & COMP_LOOP_tmp_nor_79_cse;
  assign or_359_cse = (fsm_output[2:1]!=2'b00);
  assign and_673_cse = (fsm_output[6]) & (fsm_output[4]);
  assign or_364_cse = (fsm_output[4]) | (fsm_output[7]);
  assign COMP_LOOP_or_110_rgt = and_dcpl_77 | and_dcpl_259;
  assign COMP_LOOP_tmp_nor_208_cse = ~((z_out_7[4:2]!=3'b000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse = (z_out_7[1:0]==2'b11) & COMP_LOOP_tmp_nor_208_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse = ~((z_out_7[5:0]!=6'b000000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse = (z_out_7[5:0]==6'b011001);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse = (z_out_7[4:0]==5'b10111);
  assign nor_412_cse = ~((~ (fsm_output[5])) | (fsm_output[7]));
  assign or_3900_nl = and_507_cse | (fsm_output[7]);
  assign mux_3094_nl = MUX_s_1_2_2(or_3900_nl, or_tmp_3773, fsm_output[3]);
  assign mux_3095_cse = MUX_s_1_2_2((fsm_output[7]), mux_3094_nl, fsm_output[0]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse = (z_out_7[5:0]==6'b011010);
  assign COMP_LOOP_tmp_nor_80_cse = ~((z_out_7[2:0]!=3'b000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse = (z_out_7[4:3]==2'b11) & COMP_LOOP_tmp_nor_80_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse = (z_out_7[5:0]==6'b011011);
  assign COMP_LOOP_tmp_nor_81_cse = ~((z_out_7[2:1]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse = (z_out_7[4]) & (z_out_7[3]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_81_cse;
  assign or_560_nl = (~ (fsm_output[4])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_742_cse = MUX_s_1_2_2(or_560_nl, (fsm_output[7]), fsm_output[6]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse = (z_out_7[5:0]==6'b011100);
  assign COMP_LOOP_tmp_nor_82_cse = ~((z_out_7[2]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse = (z_out_7[4]) & (z_out_7[3]) & (z_out_7[1])
      & COMP_LOOP_tmp_nor_82_cse;
  assign or_564_cse = (~ (fsm_output[5])) | (fsm_output[7]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse = (z_out_7[5:0]==6'b011101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse = (z_out_7[4:0]==5'b11011);
  assign COMP_LOOP_tmp_nor_83_cse = ~((z_out_7[1:0]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse = (z_out_7[5:0]==6'b011110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse = (z_out_7[4:2]==3'b111) & COMP_LOOP_tmp_nor_83_cse;
  assign mux_297_cse = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign and_808_cse = (fsm_output[2]) & (fsm_output[6]);
  assign and_763_cse = (fsm_output[3]) & (fsm_output[7]);
  assign or_154_nl = (fsm_output[2]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[3]);
  assign mux_221_cse = MUX_s_1_2_2(or_80_cse, or_154_nl, fsm_output[1]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse = ~((z_out_7[3:0]!=4'b0000));
  assign COMP_LOOP_tmp_nor_140_cse = ~((z_out_7[3:1]!=3'b000));
  assign COMP_LOOP_tmp_nor_141_cse = ~((z_out_7[3]) | (z_out_7[2]) | (z_out_7[0]));
  assign and_493_cse = (fsm_output[5]) & (fsm_output[7]);
  assign or_4057_cse = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[3]);
  assign and_736_cse = or_4057_cse & (fsm_output[7]);
  assign and_705_cse = (fsm_output[7:6]==2'b11);
  assign mux_180_cse = MUX_s_1_2_2(and_677_cse, and_673_cse, fsm_output[2]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse = (z_out_7[5:0]==6'b010010);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse = (z_out_7[4:0]==5'b01111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse = (z_out_7[5:0]==6'b010011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse = (z_out_7[4]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_140_cse;
  assign nor_1683_cse = ~((fsm_output[6:5]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse = (z_out_7[4]) & (z_out_7[1]) & COMP_LOOP_tmp_nor_141_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse = (z_out_7[5:0]==6'b011111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse = (z_out_7[4:0]==5'b11101);
  assign mux_3233_nl = MUX_s_1_2_2(mux_tmp_3100, mux_tmp_3098, fsm_output[2]);
  assign mux_3234_nl = MUX_s_1_2_2(mux_3233_nl, mux_tmp_3101, fsm_output[1]);
  assign COMP_LOOP_or_151_cse = MUX_s_1_2_2(mux_3234_nl, mux_tmp_3119, fsm_output[5]);
  assign mux_3237_nl = MUX_s_1_2_2(mux_tmp_3169, (fsm_output[7]), fsm_output[6]);
  assign mux_3238_nl = MUX_s_1_2_2(mux_tmp_656, mux_3237_nl, fsm_output[2]);
  assign COMP_LOOP_or_153_cse = MUX_s_1_2_2(mux_tmp_3102, mux_3238_nl, fsm_output[5]);
  assign COMP_LOOP_tmp_nor_34_cse = ~((z_out_7[4:1]!=4'b0000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse = (z_out_7[5]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_34_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse = (z_out_7[4:0]==5'b11110);
  assign nor_399_cse = ~((fsm_output[7:6]!=2'b00));
  assign or_477_cse = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]);
  assign and_655_cse = or_595_cse & (fsm_output[7]);
  assign nor_398_cse = ~((fsm_output[4]) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign COMP_LOOP_tmp_nor_35_cse = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[2])
      | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse = (z_out_7[5]) & (z_out_7[1]) & COMP_LOOP_tmp_nor_35_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse = ~((z_out_7[4:0]!=5'b00000));
  assign COMP_LOOP_tmp_or_cse = and_dcpl_74 | and_dcpl_77 | and_dcpl_258 | and_dcpl_259
      | and_dcpl_260 | and_dcpl_263;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse = (z_out_7[5:0]==6'b000101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse = (z_out_7[5:0]==6'b000011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse = (z_out_7[4:0]==5'b11111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse = (z_out_7[5:0]==6'b000110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse = (z_out_7[5:0]==6'b000111);
  assign COMP_LOOP_tmp_nor_63_cse = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[1]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse = (z_out_7[2]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_63_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse = (z_out_7[5:0]==6'b001001);
  assign COMP_LOOP_tmp_nor_64_cse = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse = (z_out_7[2:1]==2'b11) & COMP_LOOP_tmp_nor_64_cse;
  assign COMP_LOOP_tmp_nor_65_cse = ~((z_out_7[4:3]!=2'b00));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse = (z_out_7[2:0]==3'b111) & COMP_LOOP_tmp_nor_65_cse;
  assign COMP_LOOP_tmp_or_5_cse = and_dcpl_74 | and_dcpl_77 | and_dcpl_259 | and_dcpl_260
      | and_dcpl_263;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse = (z_out_7[5]) & (z_out_7[1]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_208_cse;
  assign COMP_LOOP_tmp_nor_37_cse = ~((z_out_7[4]) | (z_out_7[3]) | (z_out_7[1])
      | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse = (z_out_7[5]) & (z_out_7[2]) & COMP_LOOP_tmp_nor_37_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse = (z_out_7[5]) & (z_out_7[2]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_63_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse = (z_out_7[5]) & (z_out_7[2]) & (z_out_7[1])
      & COMP_LOOP_tmp_nor_64_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse = (z_out_7[5]) & (z_out_7[2]) & (z_out_7[1])
      & (z_out_7[0]) & COMP_LOOP_tmp_nor_65_cse;
  assign COMP_LOOP_tmp_nor_41_cse = ~((z_out_7[4]) | (z_out_7[2]) | (z_out_7[1])
      | (z_out_7[0]));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse = (z_out_7[5]) & (z_out_7[3]) & COMP_LOOP_tmp_nor_41_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse = (z_out_7[5]) & (z_out_7[3]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_67_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse = (z_out_7[5]) & (z_out_7[3]) & (z_out_7[1])
      & COMP_LOOP_tmp_nor_68_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse = (z_out_7[5]) & (z_out_7[3]) & (z_out_7[1])
      & (z_out_7[0]) & COMP_LOOP_tmp_nor_69_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse = (z_out_7[5]) & (z_out_7[3]) & (z_out_7[2])
      & COMP_LOOP_tmp_nor_70_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse = (z_out_7[5]) & (z_out_7[3]) & (z_out_7[2])
      & (z_out_7[0]) & COMP_LOOP_tmp_nor_71_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse = (z_out_7[5]) & (z_out_7[3]) & (z_out_7[2])
      & (z_out_7[1]) & COMP_LOOP_tmp_nor_72_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse = (z_out_7[5:0]==6'b101111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse = (z_out_7[5:4]==2'b11) & COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[0])
      & COMP_LOOP_tmp_nor_140_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[1])
      & COMP_LOOP_tmp_nor_141_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[1])
      & (z_out_7[0]) & COMP_LOOP_tmp_nor_76_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[2])
      & COMP_LOOP_tmp_nor_77_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[2])
      & (z_out_7[0]) & COMP_LOOP_tmp_nor_78_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[2])
      & (z_out_7[1]) & COMP_LOOP_tmp_nor_79_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse = (z_out_7[5:0]==6'b110111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse = (z_out_7[5:3]==3'b111) & COMP_LOOP_tmp_nor_80_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[3])
      & (z_out_7[0]) & COMP_LOOP_tmp_nor_81_cse;
  assign COMP_LOOP_tmp_nor_150_cse = ~((z_out_7[5:1]!=5'b00000));
  assign COMP_LOOP_or_74_cse = and_dcpl_260 | and_dcpl_263;
  assign COMP_LOOP_tmp_nor_10_cse = ~((z_out_7[5]) | (z_out_7[4]) | (z_out_7[2])
      | (z_out_7[1]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_nor_151_cse = ~((z_out_7[5]) | (z_out_7[4]) | (z_out_7[3])
      | (z_out_7[2]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_nor_18_cse = ~((z_out_7[5]) | (z_out_7[3]) | (z_out_7[2])
      | (z_out_7[1]) | (z_out_7[0]));
  assign COMP_LOOP_tmp_nor_153_cse = ~((z_out_7[5]) | (z_out_7[4]) | (z_out_7[3])
      | (z_out_7[1]) | (z_out_7[0]));
  assign COMP_LOOP_or_68_itm = and_dcpl_258 | and_dcpl_343 | and_dcpl_346 | and_dcpl_349
      | and_dcpl_351 | and_dcpl_354 | and_dcpl_357 | and_dcpl_359;
  assign COMP_LOOP_tmp_or_36_cse = and_dcpl_77 | and_dcpl_259 | and_dcpl_260 | and_dcpl_263;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse = (z_out_7[5]) & (z_out_7[4]) & (z_out_7[3])
      & (z_out_7[1]) & COMP_LOOP_tmp_nor_82_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse = (z_out_7[5:0]==6'b111011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse = (z_out_7[5:2]==4'b1111) & COMP_LOOP_tmp_nor_83_cse;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse = (z_out_7[5:0]==6'b111101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse = (z_out_7[5:0]==6'b111110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse = (z_out_7[5:0]==6'b111111);
  assign COMP_LOOP_tmp_or_43_cse = and_dcpl_258 | and_dcpl_261;
  assign or_80_cse = (fsm_output[4:2]!=3'b000);
  assign and_478_m1c = and_dcpl_262 & and_dcpl_73;
  assign mux_3357_nl = MUX_s_1_2_2(not_tmp_868, (fsm_output[7]), fsm_output[6]);
  assign mux_3358_nl = MUX_s_1_2_2(mux_3357_nl, mux_tmp_3288, fsm_output[2]);
  assign mux_3356_nl = MUX_s_1_2_2(mux_tmp_3100, mux_tmp_3288, fsm_output[2]);
  assign mux_3359_nl = MUX_s_1_2_2(mux_3358_nl, mux_3356_nl, fsm_output[1]);
  assign mux_3360_tmp = MUX_s_1_2_2(mux_3359_nl, (fsm_output[7]), fsm_output[5]);
  assign and_735_cse = (fsm_output[4]) & (fsm_output[7]);
  assign nl_COMP_LOOP_1_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b000}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_1_acc_10_nl = nl_COMP_LOOP_1_acc_10_nl[10:0];
  assign COMP_LOOP_1_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_1_acc_10_nl);
  assign nl_COMP_LOOP_acc_psp_sva_mx0w0 = (VEC_LOOP_j_10_0_sva_9_0[9:3]) + COMP_LOOP_k_10_3_sva_6_0;
  assign COMP_LOOP_acc_psp_sva_mx0w0 = nl_COMP_LOOP_acc_psp_sva_mx0w0[6:0];
  assign nl_COMP_LOOP_acc_14_psp_sva_1 = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_3_sva_6_0
      , 2'b11});
  assign COMP_LOOP_acc_14_psp_sva_1 = nl_COMP_LOOP_acc_14_psp_sva_1[8:0];
  assign nl_COMP_LOOP_acc_1_cse_4_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b011});
  assign COMP_LOOP_acc_1_cse_4_sva_1 = nl_COMP_LOOP_acc_1_cse_4_sva_1[9:0];
  assign nl_COMP_LOOP_acc_11_psp_sva_1 = (VEC_LOOP_j_10_0_sva_9_0[9:1]) + ({COMP_LOOP_k_10_3_sva_6_0
      , 2'b01});
  assign COMP_LOOP_acc_11_psp_sva_1 = nl_COMP_LOOP_acc_11_psp_sva_1[8:0];
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[9:0];
  assign nl_COMP_LOOP_2_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b001}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_2_acc_10_nl = nl_COMP_LOOP_2_acc_10_nl[10:0];
  assign COMP_LOOP_2_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_2_acc_10_nl);
  assign nl_COMP_LOOP_3_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b010}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_3_acc_10_nl = nl_COMP_LOOP_3_acc_10_nl[10:0];
  assign COMP_LOOP_3_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_3_acc_10_nl);
  assign nl_COMP_LOOP_4_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b011}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_4_acc_10_nl = nl_COMP_LOOP_4_acc_10_nl[10:0];
  assign COMP_LOOP_4_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_4_acc_10_nl);
  assign nl_COMP_LOOP_5_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b100}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_5_acc_10_nl = nl_COMP_LOOP_5_acc_10_nl[10:0];
  assign COMP_LOOP_5_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_5_acc_10_nl);
  assign nl_COMP_LOOP_6_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b101}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_6_acc_10_nl = nl_COMP_LOOP_6_acc_10_nl[10:0];
  assign COMP_LOOP_6_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_6_acc_10_nl);
  assign nl_COMP_LOOP_7_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b110}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_7_acc_10_nl = nl_COMP_LOOP_7_acc_10_nl[10:0];
  assign COMP_LOOP_7_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_7_acc_10_nl);
  assign nl_COMP_LOOP_8_acc_10_nl = conv_u2u_10_11(VEC_LOOP_j_10_0_sva_9_0) + conv_u2u_10_11({COMP_LOOP_k_10_3_sva_6_0
      , 3'b111}) + STAGE_LOOP_lshift_psp_sva;
  assign COMP_LOOP_8_acc_10_nl = nl_COMP_LOOP_8_acc_10_nl[10:0];
  assign COMP_LOOP_8_acc_10_itm_10_1_1 = readslicef_11_10_1(COMP_LOOP_8_acc_10_nl);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[1])
      & COMP_LOOP_tmp_nor_151_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[2])
      & COMP_LOOP_tmp_nor_153_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[3])
      & COMP_LOOP_tmp_nor_157_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[4])
      & COMP_LOOP_tmp_nor_165_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt = (COMP_LOOP_2_tmp_lshift_ncse_sva[5])
      & COMP_LOOP_tmp_nor_180_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[1])
      & COMP_LOOP_tmp_nor_207_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[2])
      & COMP_LOOP_tmp_nor_209_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[3])
      & COMP_LOOP_tmp_nor_213_itm;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt = (COMP_LOOP_3_tmp_lshift_ncse_sva[4])
      & COMP_LOOP_tmp_nor_220_itm;
  assign nor_tmp_1 = (fsm_output[4]) & (fsm_output[0]) & (fsm_output[3]);
  assign mux_tmp_6 = MUX_s_1_2_2((fsm_output[4]), or_595_cse, fsm_output[2]);
  assign and_dcpl_8 = nor_399_cse & (~ (fsm_output[5]));
  assign and_779_cse = (fsm_output[4:2]==3'b111);
  assign or_150_cse = (fsm_output[0]) | (fsm_output[3]);
  assign and_tmp_10 = (fsm_output[4]) & or_150_cse;
  assign or_tmp_105 = (fsm_output[4]) | and_639_cse;
  assign or_tmp_118 = (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_tmp_119 = (fsm_output[3]) | (fsm_output[7]);
  assign not_tmp_88 = ~((fsm_output[4]) | (fsm_output[7]));
  assign nor_tmp_99 = or_341_cse & (fsm_output[7]);
  assign mux_tmp_206 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_341_cse);
  assign or_4050_cse = and_640_cse | (fsm_output[6]);
  assign mux_tmp_293 = MUX_s_1_2_2(and_640_cse, (fsm_output[4]), fsm_output[2]);
  assign mux_510_nl = MUX_s_1_2_2((~ (fsm_output[7])), or_tmp_118, fsm_output[4]);
  assign mux_tmp_444 = MUX_s_1_2_2(mux_510_nl, (fsm_output[7]), fsm_output[6]);
  assign or_tmp_404 = (fsm_output[4]) | (fsm_output[3]) | (~ (fsm_output[7]));
  assign or_201_nl = (fsm_output[4]) | (~ (fsm_output[7]));
  assign mux_tmp_656 = MUX_s_1_2_2(or_201_nl, (fsm_output[7]), fsm_output[6]);
  assign and_dcpl_55 = ~((fsm_output[1]) | (fsm_output[5]));
  assign and_dcpl_57 = nor_1674_cse & and_dcpl_55;
  assign and_dcpl_58 = ~((fsm_output[0]) | (fsm_output[4]));
  assign and_dcpl_59 = ~((fsm_output[7]) | (fsm_output[3]));
  assign and_dcpl_60 = and_dcpl_59 & and_dcpl_58;
  assign and_dcpl_62 = (~ (fsm_output[1])) & (fsm_output[5]);
  assign and_dcpl_64 = and_808_cse & and_dcpl_62;
  assign and_dcpl_65 = (fsm_output[7]) & (~ (fsm_output[3]));
  assign and_dcpl_66 = and_dcpl_65 & and_dcpl_58;
  assign and_tmp_29 = (fsm_output[6]) & and_655_cse;
  assign mux_tmp_720 = MUX_s_1_2_2(and_tmp_29, and_705_cse, fsm_output[2]);
  assign and_dcpl_72 = (fsm_output[1]) & (~ (fsm_output[5]));
  assign and_dcpl_73 = nor_1674_cse & and_dcpl_72;
  assign and_dcpl_74 = and_dcpl_60 & and_dcpl_73;
  assign and_dcpl_75 = (fsm_output[0]) & (~ (fsm_output[4]));
  assign and_dcpl_76 = and_dcpl_59 & and_dcpl_75;
  assign and_dcpl_77 = and_dcpl_76 & and_dcpl_73;
  assign and_dcpl_78 = (~ (fsm_output[6])) & (fsm_output[2]);
  assign and_dcpl_79 = and_dcpl_78 & and_dcpl_72;
  assign and_dcpl_80 = (~ (fsm_output[0])) & (fsm_output[4]);
  assign and_dcpl_81 = (~ (fsm_output[7])) & (fsm_output[3]);
  assign and_dcpl_82 = and_dcpl_81 & and_dcpl_80;
  assign and_dcpl_84 = (fsm_output[0]) & (fsm_output[4]);
  assign and_dcpl_85 = and_dcpl_81 & and_dcpl_84;
  assign and_dcpl_86 = and_dcpl_85 & and_dcpl_79;
  assign and_dcpl_87 = (fsm_output[1]) & (fsm_output[5]);
  assign and_dcpl_88 = nor_1674_cse & and_dcpl_87;
  assign and_dcpl_90 = and_dcpl_85 & and_dcpl_88;
  assign and_dcpl_91 = and_808_cse & and_dcpl_72;
  assign and_dcpl_92 = and_dcpl_59 & and_dcpl_80;
  assign and_dcpl_94 = and_dcpl_59 & and_dcpl_84;
  assign and_dcpl_95 = and_dcpl_94 & and_dcpl_91;
  assign and_dcpl_96 = (fsm_output[6]) & (~ (fsm_output[2]));
  assign and_dcpl_97 = and_dcpl_96 & and_dcpl_87;
  assign and_dcpl_99 = and_dcpl_94 & and_dcpl_97;
  assign and_dcpl_101 = and_763_cse & and_dcpl_58;
  assign and_dcpl_103 = and_763_cse & and_dcpl_75;
  assign and_dcpl_104 = and_dcpl_103 & and_dcpl_79;
  assign and_dcpl_106 = and_dcpl_103 & and_dcpl_88;
  assign and_dcpl_108 = and_dcpl_65 & and_dcpl_75;
  assign and_dcpl_109 = and_dcpl_108 & and_dcpl_91;
  assign and_dcpl_110 = and_dcpl_78 & and_dcpl_55;
  assign and_dcpl_112 = and_dcpl_85 & and_dcpl_110;
  assign and_dcpl_113 = nor_1674_cse & and_dcpl_62;
  assign and_dcpl_115 = and_dcpl_85 & and_dcpl_113;
  assign and_dcpl_116 = and_808_cse & and_dcpl_55;
  assign and_dcpl_118 = and_dcpl_94 & and_dcpl_116;
  assign and_dcpl_119 = and_dcpl_96 & and_dcpl_62;
  assign or_tmp_491 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_495 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_497 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_501 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000000) | (~ and_763_cse);
  assign or_tmp_535 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_539 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_541 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_545 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000001) | (~ and_763_cse);
  assign not_tmp_321 = ~((VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_579 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_583 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_585 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_589 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000010) | (~ and_763_cse);
  assign or_tmp_623 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_627 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_629 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_633 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000011) | (~ and_763_cse);
  assign not_tmp_330 = ~((VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (fsm_output[3])
      & (fsm_output[7]));
  assign or_tmp_667 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_671 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_673 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_677 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000100) | (~ and_763_cse);
  assign or_tmp_711 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_715 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_717 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_721 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000101) | (~ and_763_cse);
  assign or_tmp_755 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_759 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_761 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_765 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000110) | (~ and_763_cse);
  assign or_tmp_799 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_803 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_805 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b000111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_809 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b000111) | (~ and_763_cse);
  assign not_tmp_347 = ~((COMP_LOOP_acc_13_psp_sva[0]) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
      & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_843 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_847 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_849 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_853 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001000) | (~ and_763_cse);
  assign or_tmp_887 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_891 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_893 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_897 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001001) | (~ and_763_cse);
  assign or_tmp_931 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_935 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_937 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_941 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001010) | (~ and_763_cse);
  assign or_tmp_975 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_979 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_981 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_985 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001011) | (~ and_763_cse);
  assign or_tmp_1019 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1023 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1025 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1029 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001100) | (~ and_763_cse);
  assign or_tmp_1063 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1067 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1069 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1073 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001101) | (~ and_763_cse);
  assign or_tmp_1107 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1111 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1113 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1117 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b001110) | (~ and_763_cse);
  assign or_tmp_1151 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1155 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1157 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b001111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1161 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b001111) & and_763_cse);
  assign or_tmp_1195 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1199 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1201 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1205 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010000) | (~ and_763_cse);
  assign not_tmp_384 = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[4]) & (fsm_output[3]) &
      (fsm_output[7]));
  assign not_tmp_388 = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[4]) & (fsm_output[3]) &
      (fsm_output[7]));
  assign or_tmp_1239 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1243 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1245 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1249 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010001) | (~ and_763_cse);
  assign or_tmp_1283 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1287 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1289 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1293 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010010) | (~ and_763_cse);
  assign or_tmp_1327 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1331 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1333 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1337 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010011) | (~ and_763_cse);
  assign or_tmp_1371 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1375 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1377 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1381 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010100) | (~ and_763_cse);
  assign or_tmp_1415 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1419 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1421 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1425 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010101) | (~ and_763_cse);
  assign or_tmp_1459 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1463 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1465 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1469 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b010110) | (~ and_763_cse);
  assign or_tmp_1503 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1507 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1509 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b010111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1513 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b010111) & and_763_cse);
  assign not_tmp_414 = ~((COMP_LOOP_acc_13_psp_sva[2]) & (COMP_LOOP_acc_13_psp_sva[0])
      & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_1547 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1551 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1553 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1557 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b011000) | (~ and_763_cse);
  assign or_tmp_1591 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1595 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1597 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1601 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b011001) | (~ and_763_cse);
  assign or_tmp_1635 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1639 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1641 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1645 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b011010) | (~ and_763_cse);
  assign or_tmp_1679 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1683 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1685 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1689 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b011011) & and_763_cse);
  assign or_tmp_1723 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1727 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1729 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1733 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]!=6'b011100) | (~ and_763_cse);
  assign or_tmp_1767 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1771 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1773 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1777 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b011101) & and_763_cse);
  assign or_tmp_1811 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1815 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1817 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b011110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1821 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b011110) & and_763_cse);
  assign or_tmp_1855 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b011111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1859 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b011111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_1861 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b011111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign or_tmp_1865 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b011111) & and_763_cse);
  assign or_tmp_1898 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1902 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1904 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_452 = ~((COMP_LOOP_acc_1_cse_6_sva[5]) & (fsm_output[3]) & (fsm_output[7]));
  assign not_tmp_453 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[5]) & (fsm_output[3]) &
      (fsm_output[7]));
  assign or_tmp_1908 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00000) | not_tmp_453;
  assign or_tmp_1942 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1946 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1948 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_458 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_6_sva[5])
      & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_1952 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b0000) | not_tmp_458;
  assign or_tmp_1986 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_1990 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_1992 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_1996 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00010) | not_tmp_453;
  assign or_tmp_2030 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2034 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2036 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_467 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[1]) & (COMP_LOOP_acc_10_cse_10_1_6_sva[0])
      & (COMP_LOOP_acc_10_cse_10_1_6_sva[5]) & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_2040 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:2]!=3'b000) | not_tmp_467;
  assign or_tmp_2074 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2078 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2080 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2084 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00100) | not_tmp_453;
  assign or_tmp_2118 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2122 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2124 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2128 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b0010) | not_tmp_458;
  assign or_tmp_2162 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2166 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2168 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2172 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b00110) | not_tmp_453;
  assign or_tmp_2206 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2210 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2212 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b100111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_484 = ~((COMP_LOOP_acc_10_cse_10_1_6_sva[2]) & (COMP_LOOP_acc_10_cse_10_1_6_sva[1])
      & (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_6_sva[5])
      & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_2216 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:3]!=2'b00) | not_tmp_484;
  assign or_tmp_2250 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2254 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2256 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2260 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01000) | not_tmp_453;
  assign or_tmp_2294 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2298 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2300 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2304 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b0100) | not_tmp_458;
  assign or_tmp_2338 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2342 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2344 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2348 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01010) | not_tmp_453;
  assign or_tmp_2382 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2386 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2388 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2392 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:2]!=3'b010) | not_tmp_467;
  assign or_tmp_2426 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2430 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2432 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2436 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01100) | not_tmp_453;
  assign or_tmp_2470 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2474 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2476 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2480 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b0110) | not_tmp_458;
  assign or_tmp_2514 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2518 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2520 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b101110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2524 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b01110) | not_tmp_453;
  assign or_tmp_2558 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b101111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2562 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b101111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_2564 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b101111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign or_tmp_2567 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4]) | (~((COMP_LOOP_acc_10_cse_10_1_6_sva[3])
      & (COMP_LOOP_acc_10_cse_10_1_6_sva[2]) & (COMP_LOOP_acc_10_cse_10_1_6_sva[1])
      & (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_6_sva[5])
      & (fsm_output[3]) & (fsm_output[7])));
  assign or_tmp_2601 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2605 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2607 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_522 = ~((COMP_LOOP_acc_1_cse_6_sva[5:4]==2'b11) & (fsm_output[3])
      & (fsm_output[7]));
  assign or_tmp_2611 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10000) | not_tmp_453;
  assign not_tmp_523 = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:4]==2'b11) & (fsm_output[3])
      & (fsm_output[7]));
  assign not_tmp_527 = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:4]==2'b11) & (fsm_output[3])
      & (fsm_output[7]));
  assign or_tmp_2645 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2649 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2651 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2655 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b1000) | not_tmp_458;
  assign or_tmp_2689 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2693 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2695 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2699 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10010) | not_tmp_453;
  assign or_tmp_2733 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2737 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2739 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2743 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:2]!=3'b100) | not_tmp_467;
  assign or_tmp_2777 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2781 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2783 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2787 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10100) | not_tmp_453;
  assign not_tmp_544 = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[2]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[5])
      & (COMP_LOOP_acc_10_cse_10_1_7_sva[4]) & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_2821 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2825 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2827 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2831 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b1010) | not_tmp_458;
  assign not_tmp_549 = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      & (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[4])
      & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_2865 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2869 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2871 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b110110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_2875 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b10110) | not_tmp_453;
  assign or_tmp_2909 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b110111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2913 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b110111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_2915 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b110111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign or_tmp_2919 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:3]!=2'b10) | not_tmp_484;
  assign or_tmp_2953 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_2957 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_2959 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b111000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_559 = ~((COMP_LOOP_acc_1_cse_6_sva[5:3]==3'b111) & (fsm_output[3])
      & (fsm_output[7]));
  assign or_tmp_2963 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11000) | not_tmp_453;
  assign not_tmp_560 = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:3]==3'b111) & (fsm_output[3])
      & (fsm_output[7]));
  assign or_tmp_2997 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_3001 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_3003 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b111001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign not_tmp_565 = ~((COMP_LOOP_acc_1_cse_6_sva[0]) & (COMP_LOOP_acc_1_cse_6_sva[3])
      & (COMP_LOOP_acc_1_cse_6_sva[4]) & (COMP_LOOP_acc_1_cse_6_sva[5]) & (fsm_output[3])
      & (fsm_output[7]));
  assign or_tmp_3007 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]!=4'b1100) | not_tmp_458;
  assign or_tmp_3041 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_3045 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_3047 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b111010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_3051 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11010) | not_tmp_453;
  assign not_tmp_570 = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      & (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[4])
      & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_3085 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_3089 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b111011) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_3091 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b111011) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign not_tmp_575 = ~((COMP_LOOP_acc_1_cse_6_sva[1]) & (COMP_LOOP_acc_1_cse_6_sva[0])
      & (COMP_LOOP_acc_1_cse_6_sva[3]) & (COMP_LOOP_acc_1_cse_6_sva[4]) & (COMP_LOOP_acc_1_cse_6_sva[5])
      & (fsm_output[3]) & (fsm_output[7]));
  assign or_tmp_3094 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:2]!=3'b110) | not_tmp_467;
  assign or_tmp_3128 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_3132 = (COMP_LOOP_acc_10_cse_10_1_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign or_tmp_3134 = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]!=6'b111100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign or_tmp_3138 = (COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]!=5'b11100) | not_tmp_453;
  assign or_tmp_3172 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_3176 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b111101) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_3178 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b111101) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign or_tmp_3182 = (~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:1]==4'b1110))) | not_tmp_458;
  assign or_tmp_3215 = (COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]!=6'b111110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_tmp_3219 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b111110) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_3221 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b111110) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign or_tmp_3225 = (~((COMP_LOOP_acc_10_cse_10_1_6_sva[4:0]==5'b11110))) | not_tmp_453;
  assign or_tmp_3258 = ~((COMP_LOOP_acc_10_cse_10_1_4_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (~ (fsm_output[7])));
  assign or_tmp_3262 = ~((COMP_LOOP_acc_10_cse_10_1_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign or_tmp_3264 = ~((COMP_LOOP_acc_10_cse_10_1_2_sva[5:0]==6'b111111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign nor_tmp_306 = (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b111111) & (fsm_output[3])
      & (fsm_output[7]);
  assign nor_tmp_307 = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:0]==6'b111111) & (fsm_output[3])
      & (fsm_output[7]);
  assign and_dcpl_258 = and_dcpl_60 & and_dcpl_110;
  assign and_dcpl_259 = and_dcpl_76 & and_dcpl_110;
  assign and_dcpl_260 = and_dcpl_60 & and_dcpl_79;
  assign and_dcpl_261 = and_dcpl_76 & and_dcpl_79;
  assign and_dcpl_262 = and_dcpl_81 & and_dcpl_58;
  assign and_dcpl_263 = and_dcpl_262 & and_dcpl_57;
  assign and_dcpl_264 = and_dcpl_81 & and_dcpl_75;
  assign and_dcpl_265 = and_dcpl_264 & and_dcpl_57;
  assign and_dcpl_268 = not_tmp_88 & nor_1683_cse;
  assign mux_tmp_2924 = MUX_s_1_2_2((~ and_763_cse), or_tmp_118, fsm_output[4]);
  assign or_tmp_3717 = (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_tmp_2927 = MUX_s_1_2_2(or_tmp_3717, or_tmp_119, fsm_output[4]);
  assign or_tmp_3718 = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]);
  assign and_dcpl_340 = (fsm_output[1:0]==2'b01);
  assign or_tmp_3721 = (~ (fsm_output[4])) | (fsm_output[3]) | (~ (fsm_output[7]));
  assign and_dcpl_343 = and_dcpl_60 & and_dcpl_113;
  assign and_dcpl_344 = and_dcpl_78 & and_dcpl_62;
  assign and_dcpl_346 = and_dcpl_82 & and_dcpl_344;
  assign and_dcpl_347 = and_dcpl_96 & and_dcpl_55;
  assign and_dcpl_349 = and_dcpl_82 & and_dcpl_347;
  assign and_dcpl_351 = and_dcpl_92 & and_dcpl_64;
  assign and_dcpl_353 = and_dcpl_65 & and_dcpl_80;
  assign and_dcpl_354 = and_dcpl_353 & and_dcpl_57;
  assign and_dcpl_355 = and_763_cse & and_dcpl_80;
  assign and_dcpl_357 = and_dcpl_101 & and_dcpl_344;
  assign and_dcpl_359 = and_dcpl_101 & and_dcpl_347;
  assign mux_522_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[4]);
  assign mux_3004_nl = MUX_s_1_2_2(and_735_cse, mux_522_nl, fsm_output[0]);
  assign nand_tmp_142 = ~((fsm_output[3]) & (~ mux_3004_nl));
  assign or_3843_nl = (fsm_output[0]) | (~ and_735_cse);
  assign mux_tmp_2939 = MUX_s_1_2_2(or_364_cse, or_3843_nl, fsm_output[3]);
  assign or_tmp_3734 = (fsm_output[5]) | (~ (fsm_output[1]));
  assign and_dcpl_365 = (~ (fsm_output[3])) & (fsm_output[0]);
  assign or_dcpl_122 = (fsm_output[6]) | (fsm_output[2]) | or_tmp_3734;
  assign or_dcpl_125 = or_tmp_119 | (fsm_output[0]) | (fsm_output[4]) | or_dcpl_122;
  assign mux_tmp_2953 = MUX_s_1_2_2(and_dcpl_60, and_655_cse, fsm_output[6]);
  assign mux_tmp_2955 = MUX_s_1_2_2((~ or_477_cse), and_655_cse, fsm_output[6]);
  assign mux_tmp_2956 = MUX_s_1_2_2(mux_tmp_2955, and_tmp_29, fsm_output[2]);
  assign mux_3021_nl = MUX_s_1_2_2(mux_tmp_2953, and_78_cse, fsm_output[2]);
  assign mux_3024_nl = MUX_s_1_2_2(mux_tmp_2956, mux_3021_nl, fsm_output[1]);
  assign mux_3025_itm = MUX_s_1_2_2(mux_3024_nl, and_705_cse, fsm_output[5]);
  assign mux_tmp_2959 = MUX_s_1_2_2((~ or_595_cse), and_640_cse, fsm_output[6]);
  assign mux_tmp_2960 = MUX_s_1_2_2(mux_tmp_2959, and_677_cse, fsm_output[2]);
  assign mux_tmp_2961 = MUX_s_1_2_2((~ or_4007_cse), and_640_cse, fsm_output[6]);
  assign mux_tmp_2965 = MUX_s_1_2_2((~ or_595_cse), (fsm_output[4]), fsm_output[6]);
  assign mux_tmp_2966 = MUX_s_1_2_2(mux_tmp_2959, mux_tmp_2965, fsm_output[2]);
  assign mux_3034_nl = MUX_s_1_2_2((~ (fsm_output[4])), and_640_cse, fsm_output[6]);
  assign mux_tmp_2968 = MUX_s_1_2_2(mux_3034_nl, mux_tmp_2965, fsm_output[2]);
  assign and_dcpl_370 = and_dcpl_264 & and_dcpl_113;
  assign mux_tmp_2971 = MUX_s_1_2_2(mux_tmp_2959, and_673_cse, fsm_output[2]);
  assign mux_3041_nl = MUX_s_1_2_2(and_dcpl_365, (fsm_output[3]), fsm_output[4]);
  assign or_tmp_3744 = (fsm_output[6]) | mux_3041_nl;
  assign mux_tmp_2975 = MUX_s_1_2_2((fsm_output[6]), or_tmp_3744, fsm_output[2]);
  assign or_tmp_3746 = (fsm_output[6]) | (~((fsm_output[4]) | (~ and_639_cse)));
  assign mux_tmp_2976 = MUX_s_1_2_2(or_tmp_3746, (fsm_output[6]), fsm_output[2]);
  assign and_dcpl_375 = and_dcpl_264 & and_dcpl_88;
  assign or_tmp_3747 = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[3]);
  assign and_dcpl_377 = and_dcpl_78 & and_dcpl_87;
  assign and_dcpl_382 = and_dcpl_94 & and_dcpl_377;
  assign or_3880_nl = (fsm_output[6]) | nor_398_cse;
  assign mux_3057_nl = MUX_s_1_2_2((fsm_output[6]), or_3880_nl, fsm_output[2]);
  assign mux_3058_itm = MUX_s_1_2_2(mux_tmp_2976, mux_3057_nl, fsm_output[1]);
  assign and_dcpl_384 = and_dcpl_85 & and_dcpl_57;
  assign mux_tmp_2993 = MUX_s_1_2_2(or_4050_cse, or_tmp_3744, fsm_output[2]);
  assign mux_tmp_2994 = MUX_s_1_2_2(or_tmp_3746, or_4050_cse, fsm_output[2]);
  assign or_tmp_3757 = (~((~ (fsm_output[0])) | (fsm_output[3]))) | (fsm_output[7]);
  assign or_tmp_3760 = and_639_cse | (fsm_output[7]);
  assign or_3887_nl = (fsm_output[4]) | (~ or_tmp_3760);
  assign mux_tmp_3001 = MUX_s_1_2_2(or_3887_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_3069_nl = MUX_s_1_2_2(mux_tmp_3001, mux_tmp_656, fsm_output[2]);
  assign or_3884_nl = (fsm_output[4]) | (~ or_tmp_3757);
  assign mux_3065_nl = MUX_s_1_2_2(or_3884_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_3067_nl = MUX_s_1_2_2(mux_tmp_656, mux_3065_nl, fsm_output[2]);
  assign mux_tmp_3003 = MUX_s_1_2_2(mux_3069_nl, mux_3067_nl, fsm_output[1]);
  assign mux_3075_nl = MUX_s_1_2_2((~ or_tmp_3757), or_tmp_118, fsm_output[4]);
  assign mux_tmp_3009 = MUX_s_1_2_2(mux_3075_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_tmp_3012 = MUX_s_1_2_2(mux_tmp_444, mux_tmp_3009, fsm_output[2]);
  assign mux_tmp_3013 = MUX_s_1_2_2(mux_tmp_3001, mux_tmp_444, fsm_output[2]);
  assign mux_tmp_3016 = MUX_s_1_2_2(and_dcpl_59, (fsm_output[7]), or_341_cse);
  assign and_dcpl_387 = and_dcpl_264 & and_dcpl_79;
  assign or_tmp_3773 = nor_1744_cse | (fsm_output[7]);
  assign and_dcpl_388 = and_dcpl_94 & and_dcpl_79;
  assign mux_tmp_3042 = MUX_s_1_2_2(mux_tmp_2953, and_705_cse, fsm_output[2]);
  assign and_tmp_31 = (fsm_output[6]) & (fsm_output[4]) & or_150_cse;
  assign or_3906_nl = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0])
      | (fsm_output[3]);
  assign mux_3114_itm = MUX_s_1_2_2(or_tmp_3747, or_3906_nl, fsm_output[1]);
  assign mux_tmp_3049 = MUX_s_1_2_2(mux_tmp_2961, and_673_cse, fsm_output[2]);
  assign mux_3117_nl = MUX_s_1_2_2(mux_tmp_2959, and_tmp_31, fsm_output[2]);
  assign mux_3118_nl = MUX_s_1_2_2(mux_3117_nl, mux_tmp_3049, fsm_output[1]);
  assign mux_3119_nl = MUX_s_1_2_2(mux_3118_nl, (fsm_output[6]), fsm_output[5]);
  assign and_dcpl_390 = ~(mux_3119_nl | (fsm_output[7]));
  assign mux_67_nl = MUX_s_1_2_2(nor_tmp_1, and_640_cse, or_359_cse);
  assign mux_3122_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_67_nl), fsm_output[5]);
  assign and_dcpl_392 = mux_3122_nl & nor_399_cse;
  assign and_dcpl_396 = mux_221_cse & and_dcpl_8;
  assign mux_3129_nl = MUX_s_1_2_2(mux_221_cse, (~ and_779_cse), fsm_output[5]);
  assign and_dcpl_399 = mux_3129_nl & nor_399_cse;
  assign mux_3133_nl = MUX_s_1_2_2(mux_tmp_2961, and_677_cse, fsm_output[2]);
  assign mux_3134_nl = MUX_s_1_2_2(mux_tmp_2960, mux_3133_nl, fsm_output[1]);
  assign mux_3135_nl = MUX_s_1_2_2(mux_3134_nl, (fsm_output[6]), fsm_output[5]);
  assign and_dcpl_402 = ~(mux_3135_nl | (fsm_output[7]));
  assign nor_1425_nl = ~((fsm_output[0]) | (fsm_output[3]) | (fsm_output[7]));
  assign mux_tmp_3069 = MUX_s_1_2_2(nor_1425_nl, (fsm_output[7]), or_341_cse);
  assign mux_tmp_3070 = MUX_s_1_2_2(mux_tmp_3069, and_736_cse, fsm_output[2]);
  assign mux_tmp_3078 = MUX_s_1_2_2(mux_tmp_3016, nor_tmp_99, fsm_output[2]);
  assign mux_3148_nl = MUX_s_1_2_2((~ mux_3114_itm), mux_180_cse, fsm_output[5]);
  assign and_dcpl_403 = ~(mux_3148_nl | (fsm_output[7]));
  assign mux_210_nl = MUX_s_1_2_2(and_640_cse, and_tmp_10, and_507_cse);
  assign mux_3150_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_210_nl), fsm_output[5]);
  assign and_dcpl_404 = mux_3150_nl & nor_399_cse;
  assign mux_214_nl = MUX_s_1_2_2(or_tmp_105, or_595_cse, fsm_output[2]);
  assign mux_215_nl = MUX_s_1_2_2(mux_tmp_6, mux_214_nl, fsm_output[1]);
  assign mux_3156_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_215_nl), fsm_output[5]);
  assign and_dcpl_406 = mux_3156_nl & nor_399_cse;
  assign mux_217_nl = MUX_s_1_2_2(or_tmp_105, or_595_cse, or_359_cse);
  assign mux_3158_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_217_nl), fsm_output[5]);
  assign and_dcpl_407 = mux_3158_nl & nor_399_cse;
  assign mux_tmp_3098 = MUX_s_1_2_2(and_dcpl_60, (fsm_output[7]), fsm_output[6]);
  assign mux_tmp_3100 = MUX_s_1_2_2((~ or_477_cse), (fsm_output[7]), fsm_output[6]);
  assign mux_tmp_3101 = MUX_s_1_2_2(mux_tmp_3100, and_705_cse, fsm_output[2]);
  assign mux_3166_nl = MUX_s_1_2_2(mux_tmp_3098, and_705_cse, fsm_output[2]);
  assign mux_tmp_3102 = MUX_s_1_2_2(mux_tmp_3101, mux_3166_nl, fsm_output[1]);
  assign mux_3173_nl = MUX_s_1_2_2(mux_tmp_3069, nor_tmp_99, fsm_output[2]);
  assign mux_3174_nl = MUX_s_1_2_2(mux_tmp_3078, mux_3173_nl, fsm_output[1]);
  assign mux_3175_itm = MUX_s_1_2_2(mux_3174_nl, (fsm_output[7]), fsm_output[5]);
  assign mux_3176_nl = MUX_s_1_2_2(nor_tmp_1, and_640_cse, fsm_output[2]);
  assign mux_3177_nl = MUX_s_1_2_2(and_779_cse, mux_3176_nl, fsm_output[1]);
  assign mux_3178_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_3177_nl), fsm_output[5]);
  assign and_dcpl_410 = mux_3178_nl & nor_399_cse;
  assign mux_3179_nl = MUX_s_1_2_2(or_4007_cse, (~ nor_tmp_1), fsm_output[2]);
  assign mux_3180_nl = MUX_s_1_2_2(or_80_cse, mux_3179_nl, fsm_output[1]);
  assign and_dcpl_411 = mux_3180_nl & and_dcpl_8;
  assign mux_3184_nl = MUX_s_1_2_2(mux_tmp_2956, mux_tmp_3042, fsm_output[1]);
  assign mux_3185_itm = MUX_s_1_2_2(mux_3184_nl, and_705_cse, fsm_output[5]);
  assign mux_tmp_3119 = MUX_s_1_2_2(nor_tmp_99, and_736_cse, fsm_output[2]);
  assign mux_3187_itm = MUX_s_1_2_2(mux_tmp_3102, mux_tmp_3119, fsm_output[5]);
  assign nor_1524_nl = ~((fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[7]));
  assign nor_409_nl = ~((fsm_output[2]) | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign not_tmp_811 = MUX_s_1_2_2(nor_1524_nl, nor_409_nl, fsm_output[1]);
  assign mux_3199_nl = MUX_s_1_2_2(mux_tmp_2953, and_tmp_29, fsm_output[2]);
  assign mux_tmp_3133 = MUX_s_1_2_2(mux_tmp_2956, mux_3199_nl, fsm_output[1]);
  assign mux_3201_itm = MUX_s_1_2_2(mux_tmp_3133, and_705_cse, fsm_output[5]);
  assign or_tmp_3801 = (fsm_output[6]) | (fsm_output[4]) | (fsm_output[0]) | (fsm_output[3]);
  assign and_tmp_33 = (fsm_output[6]) & or_595_cse;
  assign and_dcpl_421 = and_dcpl_85 & and_dcpl_73;
  assign mux_tmp_3169 = MUX_s_1_2_2(or_tmp_3717, or_tmp_118, fsm_output[4]);
  assign mux_tmp_3193 = MUX_s_1_2_2((~ (fsm_output[7])), and_655_cse, fsm_output[6]);
  assign nor_400_nl = ~((~((~ (fsm_output[0])) | (~ (fsm_output[3])) | (fsm_output[4])))
      | (fsm_output[7]));
  assign mux_3262_nl = MUX_s_1_2_2(nor_400_nl, and_655_cse, fsm_output[6]);
  assign mux_tmp_3196 = MUX_s_1_2_2(mux_3262_nl, mux_tmp_3193, fsm_output[2]);
  assign and_tmp_35 = (fsm_output[5]) & mux_297_cse;
  assign mux_tmp_3210 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_595_cse);
  assign and_tmp_36 = (fsm_output[6]) & mux_tmp_3210;
  assign mux_tmp_3213 = MUX_s_1_2_2(or_tmp_3717, (fsm_output[7]), fsm_output[4]);
  assign mux_tmp_3214 = MUX_s_1_2_2((~ or_477_cse), mux_tmp_3213, fsm_output[6]);
  assign nor_1474_nl = ~(and_640_cse | (fsm_output[7]));
  assign mux_tmp_3218 = MUX_s_1_2_2(nor_1474_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_75_nl = MUX_s_1_2_2(or_595_cse, or_4007_cse, fsm_output[2]);
  assign mux_3305_itm = MUX_s_1_2_2(mux_75_nl, or_80_cse, fsm_output[1]);
  assign or_dcpl_134 = or_tmp_119 | (~ (fsm_output[0])) | (fsm_output[4]);
  assign nor_1709_nl = ~((fsm_output[3:2]!=2'b10));
  assign nor_1710_nl = ~((fsm_output[3:2]!=2'b01));
  assign mux_3314_nl = MUX_s_1_2_2(nor_1709_nl, nor_1710_nl, fsm_output[1]);
  assign and_dcpl_432 = mux_3314_nl & (~ (fsm_output[7])) & and_dcpl_75 & nor_1683_cse;
  assign or_tmp_3833 = (fsm_output[4]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign nor_tmp_391 = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[7]);
  assign mux_tmp_3280 = MUX_s_1_2_2((~ or_477_cse), and_735_cse, fsm_output[6]);
  assign not_tmp_868 = ~((fsm_output[4]) | or_tmp_3760);
  assign or_dcpl_150 = or_dcpl_134 | (fsm_output[6]) | (~ (fsm_output[2])) | or_tmp_3734;
  assign mux_3354_nl = MUX_s_1_2_2(and_dcpl_59, and_763_cse, fsm_output[4]);
  assign mux_tmp_3288 = MUX_s_1_2_2(mux_3354_nl, (fsm_output[7]), fsm_output[6]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_66 & and_dcpl_64;
  assign VEC_LOOP_j_10_0_sva_9_0_mx0c0 = and_dcpl_76 & and_dcpl_57;
  assign mux_3318_nl = MUX_s_1_2_2(mux_tmp_2927, or_tmp_3833, fsm_output[6]);
  assign mux_3317_nl = MUX_s_1_2_2((~ nor_tmp_391), or_tmp_3721, fsm_output[6]);
  assign mux_3319_nl = MUX_s_1_2_2(mux_3318_nl, mux_3317_nl, fsm_output[2]);
  assign or_3973_nl = (fsm_output[6]) | (~ nor_tmp_391);
  assign mux_3315_nl = MUX_s_1_2_2(or_tmp_3833, or_477_cse, fsm_output[6]);
  assign mux_3316_nl = MUX_s_1_2_2(or_3973_nl, mux_3315_nl, fsm_output[2]);
  assign mux_3320_nl = MUX_s_1_2_2(mux_3319_nl, mux_3316_nl, fsm_output[5]);
  assign COMP_LOOP_1_acc_8_itm_mx0c4 = (~ mux_3320_nl) & and_dcpl_340;
  assign mux_3340_nl = MUX_s_1_2_2(mux_3305_itm, (~ mux_tmp_6), fsm_output[5]);
  assign and_474_tmp = mux_3340_nl & nor_399_cse;
  assign mux_104_nl = MUX_s_1_2_2((~ or_595_cse), or_595_cse, fsm_output[6]);
  assign mux_3342_nl = MUX_s_1_2_2(mux_104_nl, and_tmp_33, and_507_cse);
  assign mux_3343_nl = MUX_s_1_2_2(mux_3342_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_1579_tmp = ~(mux_3343_nl | (fsm_output[7]));
  assign mux_3345_nl = MUX_s_1_2_2(or_4057_cse, or_tmp_3801, and_507_cse);
  assign mux_3344_nl = MUX_s_1_2_2(and_tmp_33, (fsm_output[6]), fsm_output[2]);
  assign mux_3346_nl = MUX_s_1_2_2(mux_3345_nl, (~ mux_3344_nl), fsm_output[5]);
  assign and_476_tmp = mux_3346_nl & (~ (fsm_output[7]));
  assign nor_tmp_396 = ~((~(or_595_cse | (fsm_output[6:5]!=2'b00))) | (fsm_output[7]));
  assign and_102_nl = ((fsm_output[7]) ^ (fsm_output[4])) & ((fsm_output[3]) ^ (fsm_output[6]))
      & (~ (fsm_output[1])) & ((fsm_output[2]) ^ (fsm_output[5])) & (fsm_output[0]);
  assign vec_rsc_0_0_i_d_d_pff = MUX_v_64_2_2(COMP_LOOP_1_modulo_dev_cmp_return_rsc_z,
      COMP_LOOP_1_acc_8_itm, and_102_nl);
  assign and_114_nl = and_dcpl_82 & and_dcpl_79;
  assign and_120_nl = and_dcpl_82 & and_dcpl_88;
  assign and_124_nl = and_dcpl_92 & and_dcpl_91;
  assign and_129_nl = and_dcpl_92 & and_dcpl_97;
  assign and_133_nl = and_dcpl_101 & and_dcpl_79;
  assign and_136_nl = and_dcpl_101 & and_dcpl_88;
  assign and_138_nl = and_dcpl_66 & and_dcpl_91;
  assign vec_rsc_0_0_i_radr_d_pff = MUX1HOT_v_4_16_2((COMP_LOOP_1_acc_10_itm_10_1_1[9:6]),
      (COMP_LOOP_acc_psp_sva[6:3]), (COMP_LOOP_acc_1_cse_2_sva[9:6]), (COMP_LOOP_acc_10_cse_10_1_2_sva[9:6]),
      (COMP_LOOP_acc_11_psp_sva[8:5]), (COMP_LOOP_acc_10_cse_10_1_3_sva[9:6]), (COMP_LOOP_acc_1_cse_4_sva[9:6]),
      (COMP_LOOP_acc_10_cse_10_1_4_sva[9:6]), (COMP_LOOP_acc_13_psp_sva[7:4]), (COMP_LOOP_acc_10_cse_10_1_5_sva[9:6]),
      (COMP_LOOP_acc_1_cse_6_sva[9:6]), (COMP_LOOP_acc_10_cse_10_1_6_sva[9:6]), (COMP_LOOP_acc_14_psp_sva[8:5]),
      (COMP_LOOP_acc_10_cse_10_1_7_sva[9:6]), (COMP_LOOP_acc_1_cse_sva[9:6]), (COMP_LOOP_acc_10_cse_10_1_sva[9:6]),
      {and_dcpl_74 , and_dcpl_77 , and_114_nl , and_dcpl_86 , and_120_nl , and_dcpl_90
      , and_124_nl , and_dcpl_95 , and_129_nl , and_dcpl_99 , and_133_nl , and_dcpl_104
      , and_136_nl , and_dcpl_106 , and_138_nl , and_dcpl_109});
  assign and_142_nl = and_dcpl_82 & and_dcpl_110;
  assign and_145_nl = and_dcpl_82 & and_dcpl_113;
  assign and_148_nl = and_dcpl_92 & and_dcpl_116;
  assign and_151_nl = and_dcpl_92 & and_dcpl_119;
  assign and_152_nl = and_dcpl_94 & and_dcpl_119;
  assign and_153_nl = and_dcpl_101 & and_dcpl_110;
  assign and_154_nl = and_dcpl_103 & and_dcpl_110;
  assign and_155_nl = and_dcpl_101 & and_dcpl_113;
  assign and_156_nl = and_dcpl_103 & and_dcpl_113;
  assign and_157_nl = and_dcpl_66 & and_dcpl_116;
  assign and_158_nl = and_dcpl_108 & and_dcpl_116;
  assign and_159_nl = and_dcpl_66 & and_dcpl_119;
  assign and_160_nl = and_dcpl_108 & and_dcpl_119;
  assign vec_rsc_0_0_i_wadr_d_pff = MUX1HOT_v_4_16_2((COMP_LOOP_acc_10_cse_10_1_1_sva[9:6]),
      (COMP_LOOP_acc_psp_sva[6:3]), (COMP_LOOP_acc_10_cse_10_1_2_sva[9:6]), (COMP_LOOP_acc_1_cse_2_sva[9:6]),
      (COMP_LOOP_acc_10_cse_10_1_3_sva[9:6]), (COMP_LOOP_acc_11_psp_sva[8:5]), (COMP_LOOP_acc_10_cse_10_1_4_sva[9:6]),
      (COMP_LOOP_acc_1_cse_4_sva[9:6]), (COMP_LOOP_acc_10_cse_10_1_5_sva[9:6]), (COMP_LOOP_acc_13_psp_sva[7:4]),
      (COMP_LOOP_acc_10_cse_10_1_6_sva[9:6]), (COMP_LOOP_acc_1_cse_6_sva[9:6]), (COMP_LOOP_acc_10_cse_10_1_7_sva[9:6]),
      (COMP_LOOP_acc_14_psp_sva[8:5]), (COMP_LOOP_acc_10_cse_10_1_sva[9:6]), (COMP_LOOP_acc_1_cse_sva[9:6]),
      {and_142_nl , and_dcpl_112 , and_145_nl , and_dcpl_115 , and_148_nl , and_dcpl_118
      , and_151_nl , and_152_nl , and_153_nl , and_154_nl , and_155_nl , and_156_nl
      , and_157_nl , and_158_nl , and_159_nl , and_160_nl});
  assign nor_1414_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000000) | (~ and_763_cse));
  assign nor_1415_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_802_nl = MUX_s_1_2_2(nor_1414_nl, nor_1415_nl, fsm_output[0]);
  assign nor_1416_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1417_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_801_nl = MUX_s_1_2_2(nor_1416_nl, nor_1417_nl, fsm_output[0]);
  assign mux_803_nl = MUX_s_1_2_2(mux_802_nl, mux_801_nl, fsm_output[4]);
  assign nor_1418_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1419_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_799_nl = MUX_s_1_2_2(nor_1418_nl, nor_1419_nl, fsm_output[0]);
  assign nor_1420_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1421_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_798_nl = MUX_s_1_2_2(nor_1420_nl, nor_1421_nl, fsm_output[0]);
  assign mux_800_nl = MUX_s_1_2_2(mux_799_nl, mux_798_nl, fsm_output[4]);
  assign mux_804_nl = MUX_s_1_2_2(mux_803_nl, mux_800_nl, fsm_output[6]);
  assign nand_469_nl = ~((fsm_output[2]) & mux_804_nl);
  assign or_615_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000000) | (~ and_763_cse);
  assign mux_795_nl = MUX_s_1_2_2(or_tmp_501, or_615_nl, fsm_output[0]);
  assign or_612_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_794_nl = MUX_s_1_2_2(or_tmp_497, or_612_nl, fsm_output[0]);
  assign mux_796_nl = MUX_s_1_2_2(mux_795_nl, mux_794_nl, fsm_output[4]);
  assign or_609_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_792_nl = MUX_s_1_2_2(or_tmp_495, or_609_nl, fsm_output[0]);
  assign or_606_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_791_nl = MUX_s_1_2_2(or_tmp_491, or_606_nl, fsm_output[0]);
  assign mux_793_nl = MUX_s_1_2_2(mux_792_nl, mux_791_nl, fsm_output[4]);
  assign mux_797_nl = MUX_s_1_2_2(mux_796_nl, mux_793_nl, fsm_output[6]);
  assign or_4142_nl = (fsm_output[2]) | mux_797_nl;
  assign mux_805_nl = MUX_s_1_2_2(nand_469_nl, or_4142_nl, fsm_output[5]);
  assign vec_rsc_0_0_i_we_d_pff = ~(mux_805_nl | (fsm_output[1]));
  assign or_648_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_647_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_818_nl = MUX_s_1_2_2(or_648_nl, or_647_nl, fsm_output[0]);
  assign or_649_nl = (fsm_output[6]) | (fsm_output[4]) | mux_818_nl;
  assign or_645_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000000)
      | (~ and_763_cse);
  assign mux_815_nl = MUX_s_1_2_2(or_645_nl, or_tmp_501, fsm_output[0]);
  assign or_643_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_814_nl = MUX_s_1_2_2(or_643_nl, or_tmp_497, fsm_output[0]);
  assign mux_816_nl = MUX_s_1_2_2(mux_815_nl, mux_814_nl, fsm_output[4]);
  assign or_642_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_812_nl = MUX_s_1_2_2(or_642_nl, or_tmp_495, fsm_output[0]);
  assign or_640_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_811_nl = MUX_s_1_2_2(or_640_nl, or_tmp_491, fsm_output[0]);
  assign mux_813_nl = MUX_s_1_2_2(mux_812_nl, mux_811_nl, fsm_output[4]);
  assign mux_817_nl = MUX_s_1_2_2(mux_816_nl, mux_813_nl, fsm_output[6]);
  assign mux_819_nl = MUX_s_1_2_2(or_649_nl, mux_817_nl, fsm_output[2]);
  assign or_638_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_636_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000000) | (~ and_763_cse);
  assign mux_808_nl = MUX_s_1_2_2(or_638_nl, or_636_nl, fsm_output[0]);
  assign or_634_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_633_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_807_nl = MUX_s_1_2_2(or_634_nl, or_633_nl, fsm_output[0]);
  assign mux_809_nl = MUX_s_1_2_2(mux_808_nl, mux_807_nl, fsm_output[4]);
  assign nor_1412_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1413_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_806_nl = MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, fsm_output[0]);
  assign nand_15_nl = ~((fsm_output[4]) & mux_806_nl);
  assign mux_810_nl = MUX_s_1_2_2(mux_809_nl, nand_15_nl, fsm_output[6]);
  assign or_639_nl = (fsm_output[2]) | mux_810_nl;
  assign mux_820_nl = MUX_s_1_2_2(mux_819_nl, or_639_nl, fsm_output[5]);
  assign vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_820_nl) & (fsm_output[1]);
  assign nor_1403_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000001) | (~ and_763_cse));
  assign nor_1404_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_832_nl = MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output[0]);
  assign nor_1405_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1406_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_831_nl = MUX_s_1_2_2(nor_1405_nl, nor_1406_nl, fsm_output[0]);
  assign mux_833_nl = MUX_s_1_2_2(mux_832_nl, mux_831_nl, fsm_output[4]);
  assign nor_1407_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1408_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_829_nl = MUX_s_1_2_2(nor_1407_nl, nor_1408_nl, fsm_output[0]);
  assign nor_1409_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1410_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_828_nl = MUX_s_1_2_2(nor_1409_nl, nor_1410_nl, fsm_output[0]);
  assign mux_830_nl = MUX_s_1_2_2(mux_829_nl, mux_828_nl, fsm_output[4]);
  assign mux_834_nl = MUX_s_1_2_2(mux_833_nl, mux_830_nl, fsm_output[6]);
  assign nand_468_nl = ~((fsm_output[2]) & mux_834_nl);
  assign or_659_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000001) | (~ and_763_cse);
  assign mux_825_nl = MUX_s_1_2_2(or_tmp_545, or_659_nl, fsm_output[0]);
  assign or_656_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_824_nl = MUX_s_1_2_2(or_tmp_541, or_656_nl, fsm_output[0]);
  assign mux_826_nl = MUX_s_1_2_2(mux_825_nl, mux_824_nl, fsm_output[4]);
  assign or_653_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_822_nl = MUX_s_1_2_2(or_tmp_539, or_653_nl, fsm_output[0]);
  assign or_650_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_821_nl = MUX_s_1_2_2(or_tmp_535, or_650_nl, fsm_output[0]);
  assign mux_823_nl = MUX_s_1_2_2(mux_822_nl, mux_821_nl, fsm_output[4]);
  assign mux_827_nl = MUX_s_1_2_2(mux_826_nl, mux_823_nl, fsm_output[6]);
  assign or_4141_nl = (fsm_output[2]) | mux_827_nl;
  assign mux_835_nl = MUX_s_1_2_2(nand_468_nl, or_4141_nl, fsm_output[5]);
  assign vec_rsc_0_1_i_we_d_pff = ~(mux_835_nl | (fsm_output[1]));
  assign or_692_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_691_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_848_nl = MUX_s_1_2_2(or_692_nl, or_691_nl, fsm_output[0]);
  assign or_693_nl = (fsm_output[6]) | (fsm_output[4]) | mux_848_nl;
  assign or_689_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000001)
      | (~ and_763_cse);
  assign mux_845_nl = MUX_s_1_2_2(or_689_nl, or_tmp_545, fsm_output[0]);
  assign or_687_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_844_nl = MUX_s_1_2_2(or_687_nl, or_tmp_541, fsm_output[0]);
  assign mux_846_nl = MUX_s_1_2_2(mux_845_nl, mux_844_nl, fsm_output[4]);
  assign or_686_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_842_nl = MUX_s_1_2_2(or_686_nl, or_tmp_539, fsm_output[0]);
  assign or_684_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_841_nl = MUX_s_1_2_2(or_684_nl, or_tmp_535, fsm_output[0]);
  assign mux_843_nl = MUX_s_1_2_2(mux_842_nl, mux_841_nl, fsm_output[4]);
  assign mux_847_nl = MUX_s_1_2_2(mux_846_nl, mux_843_nl, fsm_output[6]);
  assign mux_849_nl = MUX_s_1_2_2(or_693_nl, mux_847_nl, fsm_output[2]);
  assign or_682_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_680_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000001) | (~ and_763_cse);
  assign mux_838_nl = MUX_s_1_2_2(or_682_nl, or_680_nl, fsm_output[0]);
  assign or_678_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_677_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_837_nl = MUX_s_1_2_2(or_678_nl, or_677_nl, fsm_output[0]);
  assign mux_839_nl = MUX_s_1_2_2(mux_838_nl, mux_837_nl, fsm_output[4]);
  assign nor_1401_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1402_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_836_nl = MUX_s_1_2_2(nor_1401_nl, nor_1402_nl, fsm_output[0]);
  assign nand_17_nl = ~((fsm_output[4]) & mux_836_nl);
  assign mux_840_nl = MUX_s_1_2_2(mux_839_nl, nand_17_nl, fsm_output[6]);
  assign or_683_nl = (fsm_output[2]) | mux_840_nl;
  assign mux_850_nl = MUX_s_1_2_2(mux_849_nl, or_683_nl, fsm_output[5]);
  assign vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_850_nl) & (fsm_output[1]);
  assign nor_1392_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000010) | (~ and_763_cse));
  assign nor_1393_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_862_nl = MUX_s_1_2_2(nor_1392_nl, nor_1393_nl, fsm_output[0]);
  assign nor_1394_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1395_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_861_nl = MUX_s_1_2_2(nor_1394_nl, nor_1395_nl, fsm_output[0]);
  assign mux_863_nl = MUX_s_1_2_2(mux_862_nl, mux_861_nl, fsm_output[4]);
  assign nor_1396_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1397_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_859_nl = MUX_s_1_2_2(nor_1396_nl, nor_1397_nl, fsm_output[0]);
  assign nor_1398_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1399_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_858_nl = MUX_s_1_2_2(nor_1398_nl, nor_1399_nl, fsm_output[0]);
  assign mux_860_nl = MUX_s_1_2_2(mux_859_nl, mux_858_nl, fsm_output[4]);
  assign mux_864_nl = MUX_s_1_2_2(mux_863_nl, mux_860_nl, fsm_output[6]);
  assign nand_467_nl = ~((fsm_output[2]) & mux_864_nl);
  assign or_703_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000010) | (~ and_763_cse);
  assign mux_855_nl = MUX_s_1_2_2(or_tmp_589, or_703_nl, fsm_output[0]);
  assign or_700_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_854_nl = MUX_s_1_2_2(or_tmp_585, or_700_nl, fsm_output[0]);
  assign mux_856_nl = MUX_s_1_2_2(mux_855_nl, mux_854_nl, fsm_output[4]);
  assign or_697_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_852_nl = MUX_s_1_2_2(or_tmp_583, or_697_nl, fsm_output[0]);
  assign or_694_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_851_nl = MUX_s_1_2_2(or_tmp_579, or_694_nl, fsm_output[0]);
  assign mux_853_nl = MUX_s_1_2_2(mux_852_nl, mux_851_nl, fsm_output[4]);
  assign mux_857_nl = MUX_s_1_2_2(mux_856_nl, mux_853_nl, fsm_output[6]);
  assign or_4140_nl = (fsm_output[2]) | mux_857_nl;
  assign mux_865_nl = MUX_s_1_2_2(nand_467_nl, or_4140_nl, fsm_output[5]);
  assign vec_rsc_0_2_i_we_d_pff = ~(mux_865_nl | (fsm_output[1]));
  assign or_736_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_735_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_878_nl = MUX_s_1_2_2(or_736_nl, or_735_nl, fsm_output[0]);
  assign or_737_nl = (fsm_output[6]) | (fsm_output[4]) | mux_878_nl;
  assign or_733_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000010)
      | (~ and_763_cse);
  assign mux_875_nl = MUX_s_1_2_2(or_733_nl, or_tmp_589, fsm_output[0]);
  assign or_731_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_874_nl = MUX_s_1_2_2(or_731_nl, or_tmp_585, fsm_output[0]);
  assign mux_876_nl = MUX_s_1_2_2(mux_875_nl, mux_874_nl, fsm_output[4]);
  assign or_730_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_872_nl = MUX_s_1_2_2(or_730_nl, or_tmp_583, fsm_output[0]);
  assign or_728_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_871_nl = MUX_s_1_2_2(or_728_nl, or_tmp_579, fsm_output[0]);
  assign mux_873_nl = MUX_s_1_2_2(mux_872_nl, mux_871_nl, fsm_output[4]);
  assign mux_877_nl = MUX_s_1_2_2(mux_876_nl, mux_873_nl, fsm_output[6]);
  assign mux_879_nl = MUX_s_1_2_2(or_737_nl, mux_877_nl, fsm_output[2]);
  assign or_726_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_724_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000010) | (~ and_763_cse);
  assign mux_868_nl = MUX_s_1_2_2(or_726_nl, or_724_nl, fsm_output[0]);
  assign or_722_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_721_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_867_nl = MUX_s_1_2_2(or_722_nl, or_721_nl, fsm_output[0]);
  assign mux_869_nl = MUX_s_1_2_2(mux_868_nl, mux_867_nl, fsm_output[4]);
  assign nor_1390_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1391_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_866_nl = MUX_s_1_2_2(nor_1390_nl, nor_1391_nl, fsm_output[0]);
  assign nand_19_nl = ~((fsm_output[4]) & mux_866_nl);
  assign mux_870_nl = MUX_s_1_2_2(mux_869_nl, nand_19_nl, fsm_output[6]);
  assign or_727_nl = (fsm_output[2]) | mux_870_nl;
  assign mux_880_nl = MUX_s_1_2_2(mux_879_nl, or_727_nl, fsm_output[5]);
  assign vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_880_nl) & (fsm_output[1]);
  assign nor_1381_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000011) | (~ and_763_cse));
  assign nor_1382_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | not_tmp_330);
  assign mux_892_nl = MUX_s_1_2_2(nor_1381_nl, nor_1382_nl, fsm_output[0]);
  assign nor_1383_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1384_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_891_nl = MUX_s_1_2_2(nor_1383_nl, nor_1384_nl, fsm_output[0]);
  assign mux_893_nl = MUX_s_1_2_2(mux_892_nl, mux_891_nl, fsm_output[4]);
  assign nor_1385_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1386_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_889_nl = MUX_s_1_2_2(nor_1385_nl, nor_1386_nl, fsm_output[0]);
  assign nor_1387_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1388_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_888_nl = MUX_s_1_2_2(nor_1387_nl, nor_1388_nl, fsm_output[0]);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, mux_888_nl, fsm_output[4]);
  assign mux_894_nl = MUX_s_1_2_2(mux_893_nl, mux_890_nl, fsm_output[6]);
  assign nand_466_nl = ~((fsm_output[2]) & mux_894_nl);
  assign or_747_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000011) | (~ and_763_cse);
  assign mux_885_nl = MUX_s_1_2_2(or_tmp_633, or_747_nl, fsm_output[0]);
  assign or_744_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_884_nl = MUX_s_1_2_2(or_tmp_629, or_744_nl, fsm_output[0]);
  assign mux_886_nl = MUX_s_1_2_2(mux_885_nl, mux_884_nl, fsm_output[4]);
  assign or_741_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_882_nl = MUX_s_1_2_2(or_tmp_627, or_741_nl, fsm_output[0]);
  assign or_738_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_881_nl = MUX_s_1_2_2(or_tmp_623, or_738_nl, fsm_output[0]);
  assign mux_883_nl = MUX_s_1_2_2(mux_882_nl, mux_881_nl, fsm_output[4]);
  assign mux_887_nl = MUX_s_1_2_2(mux_886_nl, mux_883_nl, fsm_output[6]);
  assign or_4139_nl = (fsm_output[2]) | mux_887_nl;
  assign mux_895_nl = MUX_s_1_2_2(nand_466_nl, or_4139_nl, fsm_output[5]);
  assign vec_rsc_0_3_i_we_d_pff = ~(mux_895_nl | (fsm_output[1]));
  assign or_780_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_779_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_908_nl = MUX_s_1_2_2(or_780_nl, or_779_nl, fsm_output[0]);
  assign or_781_nl = (fsm_output[6]) | (fsm_output[4]) | mux_908_nl;
  assign or_777_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000011)
      | (~ and_763_cse);
  assign mux_905_nl = MUX_s_1_2_2(or_777_nl, or_tmp_633, fsm_output[0]);
  assign or_775_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_904_nl = MUX_s_1_2_2(or_775_nl, or_tmp_629, fsm_output[0]);
  assign mux_906_nl = MUX_s_1_2_2(mux_905_nl, mux_904_nl, fsm_output[4]);
  assign or_774_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_902_nl = MUX_s_1_2_2(or_774_nl, or_tmp_627, fsm_output[0]);
  assign or_772_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_901_nl = MUX_s_1_2_2(or_772_nl, or_tmp_623, fsm_output[0]);
  assign mux_903_nl = MUX_s_1_2_2(mux_902_nl, mux_901_nl, fsm_output[4]);
  assign mux_907_nl = MUX_s_1_2_2(mux_906_nl, mux_903_nl, fsm_output[6]);
  assign mux_909_nl = MUX_s_1_2_2(or_781_nl, mux_907_nl, fsm_output[2]);
  assign or_770_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_768_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000011) | (~ and_763_cse);
  assign mux_898_nl = MUX_s_1_2_2(or_770_nl, or_768_nl, fsm_output[0]);
  assign or_766_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_765_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_897_nl = MUX_s_1_2_2(or_766_nl, or_765_nl, fsm_output[0]);
  assign mux_899_nl = MUX_s_1_2_2(mux_898_nl, mux_897_nl, fsm_output[4]);
  assign nor_1379_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1380_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_896_nl = MUX_s_1_2_2(nor_1379_nl, nor_1380_nl, fsm_output[0]);
  assign nand_21_nl = ~((fsm_output[4]) & mux_896_nl);
  assign mux_900_nl = MUX_s_1_2_2(mux_899_nl, nand_21_nl, fsm_output[6]);
  assign or_771_nl = (fsm_output[2]) | mux_900_nl;
  assign mux_910_nl = MUX_s_1_2_2(mux_909_nl, or_771_nl, fsm_output[5]);
  assign vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_910_nl) & (fsm_output[1]);
  assign nor_1370_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000100) | (~ and_763_cse));
  assign nor_1371_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_922_nl = MUX_s_1_2_2(nor_1370_nl, nor_1371_nl, fsm_output[0]);
  assign nor_1372_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1373_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_921_nl = MUX_s_1_2_2(nor_1372_nl, nor_1373_nl, fsm_output[0]);
  assign mux_923_nl = MUX_s_1_2_2(mux_922_nl, mux_921_nl, fsm_output[4]);
  assign nor_1374_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1375_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_919_nl = MUX_s_1_2_2(nor_1374_nl, nor_1375_nl, fsm_output[0]);
  assign nor_1376_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1377_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_918_nl = MUX_s_1_2_2(nor_1376_nl, nor_1377_nl, fsm_output[0]);
  assign mux_920_nl = MUX_s_1_2_2(mux_919_nl, mux_918_nl, fsm_output[4]);
  assign mux_924_nl = MUX_s_1_2_2(mux_923_nl, mux_920_nl, fsm_output[6]);
  assign nand_465_nl = ~((fsm_output[2]) & mux_924_nl);
  assign or_791_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000100) | (~ and_763_cse);
  assign mux_915_nl = MUX_s_1_2_2(or_tmp_677, or_791_nl, fsm_output[0]);
  assign or_788_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_914_nl = MUX_s_1_2_2(or_tmp_673, or_788_nl, fsm_output[0]);
  assign mux_916_nl = MUX_s_1_2_2(mux_915_nl, mux_914_nl, fsm_output[4]);
  assign or_785_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_912_nl = MUX_s_1_2_2(or_tmp_671, or_785_nl, fsm_output[0]);
  assign or_782_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_911_nl = MUX_s_1_2_2(or_tmp_667, or_782_nl, fsm_output[0]);
  assign mux_913_nl = MUX_s_1_2_2(mux_912_nl, mux_911_nl, fsm_output[4]);
  assign mux_917_nl = MUX_s_1_2_2(mux_916_nl, mux_913_nl, fsm_output[6]);
  assign or_4138_nl = (fsm_output[2]) | mux_917_nl;
  assign mux_925_nl = MUX_s_1_2_2(nand_465_nl, or_4138_nl, fsm_output[5]);
  assign vec_rsc_0_4_i_we_d_pff = ~(mux_925_nl | (fsm_output[1]));
  assign or_824_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_823_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_938_nl = MUX_s_1_2_2(or_824_nl, or_823_nl, fsm_output[0]);
  assign or_825_nl = (fsm_output[6]) | (fsm_output[4]) | mux_938_nl;
  assign or_821_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000100)
      | (~ and_763_cse);
  assign mux_935_nl = MUX_s_1_2_2(or_821_nl, or_tmp_677, fsm_output[0]);
  assign or_819_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_934_nl = MUX_s_1_2_2(or_819_nl, or_tmp_673, fsm_output[0]);
  assign mux_936_nl = MUX_s_1_2_2(mux_935_nl, mux_934_nl, fsm_output[4]);
  assign or_818_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_932_nl = MUX_s_1_2_2(or_818_nl, or_tmp_671, fsm_output[0]);
  assign or_816_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_931_nl = MUX_s_1_2_2(or_816_nl, or_tmp_667, fsm_output[0]);
  assign mux_933_nl = MUX_s_1_2_2(mux_932_nl, mux_931_nl, fsm_output[4]);
  assign mux_937_nl = MUX_s_1_2_2(mux_936_nl, mux_933_nl, fsm_output[6]);
  assign mux_939_nl = MUX_s_1_2_2(or_825_nl, mux_937_nl, fsm_output[2]);
  assign or_814_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_812_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000100) | (~ and_763_cse);
  assign mux_928_nl = MUX_s_1_2_2(or_814_nl, or_812_nl, fsm_output[0]);
  assign or_810_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_809_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_927_nl = MUX_s_1_2_2(or_810_nl, or_809_nl, fsm_output[0]);
  assign mux_929_nl = MUX_s_1_2_2(mux_928_nl, mux_927_nl, fsm_output[4]);
  assign nor_1368_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1369_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_926_nl = MUX_s_1_2_2(nor_1368_nl, nor_1369_nl, fsm_output[0]);
  assign nand_23_nl = ~((fsm_output[4]) & mux_926_nl);
  assign mux_930_nl = MUX_s_1_2_2(mux_929_nl, nand_23_nl, fsm_output[6]);
  assign or_815_nl = (fsm_output[2]) | mux_930_nl;
  assign mux_940_nl = MUX_s_1_2_2(mux_939_nl, or_815_nl, fsm_output[5]);
  assign vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_940_nl) & (fsm_output[1]);
  assign nor_1359_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000101) | (~ and_763_cse));
  assign nor_1360_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_952_nl = MUX_s_1_2_2(nor_1359_nl, nor_1360_nl, fsm_output[0]);
  assign nor_1361_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1362_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_951_nl = MUX_s_1_2_2(nor_1361_nl, nor_1362_nl, fsm_output[0]);
  assign mux_953_nl = MUX_s_1_2_2(mux_952_nl, mux_951_nl, fsm_output[4]);
  assign nor_1363_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1364_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_949_nl = MUX_s_1_2_2(nor_1363_nl, nor_1364_nl, fsm_output[0]);
  assign nor_1365_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1366_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_948_nl = MUX_s_1_2_2(nor_1365_nl, nor_1366_nl, fsm_output[0]);
  assign mux_950_nl = MUX_s_1_2_2(mux_949_nl, mux_948_nl, fsm_output[4]);
  assign mux_954_nl = MUX_s_1_2_2(mux_953_nl, mux_950_nl, fsm_output[6]);
  assign nand_464_nl = ~((fsm_output[2]) & mux_954_nl);
  assign or_835_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000101) | (~ and_763_cse);
  assign mux_945_nl = MUX_s_1_2_2(or_tmp_721, or_835_nl, fsm_output[0]);
  assign or_832_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_944_nl = MUX_s_1_2_2(or_tmp_717, or_832_nl, fsm_output[0]);
  assign mux_946_nl = MUX_s_1_2_2(mux_945_nl, mux_944_nl, fsm_output[4]);
  assign or_829_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_942_nl = MUX_s_1_2_2(or_tmp_715, or_829_nl, fsm_output[0]);
  assign or_826_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_941_nl = MUX_s_1_2_2(or_tmp_711, or_826_nl, fsm_output[0]);
  assign mux_943_nl = MUX_s_1_2_2(mux_942_nl, mux_941_nl, fsm_output[4]);
  assign mux_947_nl = MUX_s_1_2_2(mux_946_nl, mux_943_nl, fsm_output[6]);
  assign or_4137_nl = (fsm_output[2]) | mux_947_nl;
  assign mux_955_nl = MUX_s_1_2_2(nand_464_nl, or_4137_nl, fsm_output[5]);
  assign vec_rsc_0_5_i_we_d_pff = ~(mux_955_nl | (fsm_output[1]));
  assign or_868_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_867_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_968_nl = MUX_s_1_2_2(or_868_nl, or_867_nl, fsm_output[0]);
  assign or_869_nl = (fsm_output[6]) | (fsm_output[4]) | mux_968_nl;
  assign or_865_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000101)
      | (~ and_763_cse);
  assign mux_965_nl = MUX_s_1_2_2(or_865_nl, or_tmp_721, fsm_output[0]);
  assign or_863_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_964_nl = MUX_s_1_2_2(or_863_nl, or_tmp_717, fsm_output[0]);
  assign mux_966_nl = MUX_s_1_2_2(mux_965_nl, mux_964_nl, fsm_output[4]);
  assign or_862_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_962_nl = MUX_s_1_2_2(or_862_nl, or_tmp_715, fsm_output[0]);
  assign or_860_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_961_nl = MUX_s_1_2_2(or_860_nl, or_tmp_711, fsm_output[0]);
  assign mux_963_nl = MUX_s_1_2_2(mux_962_nl, mux_961_nl, fsm_output[4]);
  assign mux_967_nl = MUX_s_1_2_2(mux_966_nl, mux_963_nl, fsm_output[6]);
  assign mux_969_nl = MUX_s_1_2_2(or_869_nl, mux_967_nl, fsm_output[2]);
  assign or_858_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_856_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000101) | (~ and_763_cse);
  assign mux_958_nl = MUX_s_1_2_2(or_858_nl, or_856_nl, fsm_output[0]);
  assign or_854_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_853_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_957_nl = MUX_s_1_2_2(or_854_nl, or_853_nl, fsm_output[0]);
  assign mux_959_nl = MUX_s_1_2_2(mux_958_nl, mux_957_nl, fsm_output[4]);
  assign nor_1357_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1358_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_956_nl = MUX_s_1_2_2(nor_1357_nl, nor_1358_nl, fsm_output[0]);
  assign nand_25_nl = ~((fsm_output[4]) & mux_956_nl);
  assign mux_960_nl = MUX_s_1_2_2(mux_959_nl, nand_25_nl, fsm_output[6]);
  assign or_859_nl = (fsm_output[2]) | mux_960_nl;
  assign mux_970_nl = MUX_s_1_2_2(mux_969_nl, or_859_nl, fsm_output[5]);
  assign vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_970_nl) & (fsm_output[1]);
  assign nor_1348_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000110) | (~ and_763_cse));
  assign nor_1349_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_982_nl = MUX_s_1_2_2(nor_1348_nl, nor_1349_nl, fsm_output[0]);
  assign nor_1350_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1351_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_981_nl = MUX_s_1_2_2(nor_1350_nl, nor_1351_nl, fsm_output[0]);
  assign mux_983_nl = MUX_s_1_2_2(mux_982_nl, mux_981_nl, fsm_output[4]);
  assign nor_1352_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1353_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_979_nl = MUX_s_1_2_2(nor_1352_nl, nor_1353_nl, fsm_output[0]);
  assign nor_1354_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1355_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_978_nl = MUX_s_1_2_2(nor_1354_nl, nor_1355_nl, fsm_output[0]);
  assign mux_980_nl = MUX_s_1_2_2(mux_979_nl, mux_978_nl, fsm_output[4]);
  assign mux_984_nl = MUX_s_1_2_2(mux_983_nl, mux_980_nl, fsm_output[6]);
  assign nand_463_nl = ~((fsm_output[2]) & mux_984_nl);
  assign or_879_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000110) | (~ and_763_cse);
  assign mux_975_nl = MUX_s_1_2_2(or_tmp_765, or_879_nl, fsm_output[0]);
  assign or_876_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_974_nl = MUX_s_1_2_2(or_tmp_761, or_876_nl, fsm_output[0]);
  assign mux_976_nl = MUX_s_1_2_2(mux_975_nl, mux_974_nl, fsm_output[4]);
  assign or_873_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_972_nl = MUX_s_1_2_2(or_tmp_759, or_873_nl, fsm_output[0]);
  assign or_870_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_971_nl = MUX_s_1_2_2(or_tmp_755, or_870_nl, fsm_output[0]);
  assign mux_973_nl = MUX_s_1_2_2(mux_972_nl, mux_971_nl, fsm_output[4]);
  assign mux_977_nl = MUX_s_1_2_2(mux_976_nl, mux_973_nl, fsm_output[6]);
  assign or_4136_nl = (fsm_output[2]) | mux_977_nl;
  assign mux_985_nl = MUX_s_1_2_2(nand_463_nl, or_4136_nl, fsm_output[5]);
  assign vec_rsc_0_6_i_we_d_pff = ~(mux_985_nl | (fsm_output[1]));
  assign or_912_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_911_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_998_nl = MUX_s_1_2_2(or_912_nl, or_911_nl, fsm_output[0]);
  assign or_913_nl = (fsm_output[6]) | (fsm_output[4]) | mux_998_nl;
  assign or_909_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000110)
      | (~ and_763_cse);
  assign mux_995_nl = MUX_s_1_2_2(or_909_nl, or_tmp_765, fsm_output[0]);
  assign or_907_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_994_nl = MUX_s_1_2_2(or_907_nl, or_tmp_761, fsm_output[0]);
  assign mux_996_nl = MUX_s_1_2_2(mux_995_nl, mux_994_nl, fsm_output[4]);
  assign or_906_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_992_nl = MUX_s_1_2_2(or_906_nl, or_tmp_759, fsm_output[0]);
  assign or_904_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_991_nl = MUX_s_1_2_2(or_904_nl, or_tmp_755, fsm_output[0]);
  assign mux_993_nl = MUX_s_1_2_2(mux_992_nl, mux_991_nl, fsm_output[4]);
  assign mux_997_nl = MUX_s_1_2_2(mux_996_nl, mux_993_nl, fsm_output[6]);
  assign mux_999_nl = MUX_s_1_2_2(or_913_nl, mux_997_nl, fsm_output[2]);
  assign or_902_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_900_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000110) | (~ and_763_cse);
  assign mux_988_nl = MUX_s_1_2_2(or_902_nl, or_900_nl, fsm_output[0]);
  assign or_898_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_897_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_987_nl = MUX_s_1_2_2(or_898_nl, or_897_nl, fsm_output[0]);
  assign mux_989_nl = MUX_s_1_2_2(mux_988_nl, mux_987_nl, fsm_output[4]);
  assign nor_1346_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1347_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_986_nl = MUX_s_1_2_2(nor_1346_nl, nor_1347_nl, fsm_output[0]);
  assign nand_27_nl = ~((fsm_output[4]) & mux_986_nl);
  assign mux_990_nl = MUX_s_1_2_2(mux_989_nl, nand_27_nl, fsm_output[6]);
  assign or_903_nl = (fsm_output[2]) | mux_990_nl;
  assign mux_1000_nl = MUX_s_1_2_2(mux_999_nl, or_903_nl, fsm_output[5]);
  assign vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1000_nl) & (fsm_output[1]);
  assign nor_1337_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000111) | (~ and_763_cse));
  assign nor_1338_nl = ~((COMP_LOOP_acc_13_psp_sva[3:1]!=3'b000) | not_tmp_347);
  assign mux_1012_nl = MUX_s_1_2_2(nor_1337_nl, nor_1338_nl, fsm_output[0]);
  assign nor_1339_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b000111) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1340_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1011_nl = MUX_s_1_2_2(nor_1339_nl, nor_1340_nl, fsm_output[0]);
  assign mux_1013_nl = MUX_s_1_2_2(mux_1012_nl, mux_1011_nl, fsm_output[4]);
  assign nor_1341_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1342_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1009_nl = MUX_s_1_2_2(nor_1341_nl, nor_1342_nl, fsm_output[0]);
  assign nor_1343_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1344_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1008_nl = MUX_s_1_2_2(nor_1343_nl, nor_1344_nl, fsm_output[0]);
  assign mux_1010_nl = MUX_s_1_2_2(mux_1009_nl, mux_1008_nl, fsm_output[4]);
  assign mux_1014_nl = MUX_s_1_2_2(mux_1013_nl, mux_1010_nl, fsm_output[6]);
  assign nand_462_nl = ~((fsm_output[2]) & mux_1014_nl);
  assign or_923_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000111) | (~ and_763_cse);
  assign mux_1005_nl = MUX_s_1_2_2(or_tmp_809, or_923_nl, fsm_output[0]);
  assign or_920_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1004_nl = MUX_s_1_2_2(or_tmp_805, or_920_nl, fsm_output[0]);
  assign mux_1006_nl = MUX_s_1_2_2(mux_1005_nl, mux_1004_nl, fsm_output[4]);
  assign or_917_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1002_nl = MUX_s_1_2_2(or_tmp_803, or_917_nl, fsm_output[0]);
  assign or_914_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1001_nl = MUX_s_1_2_2(or_tmp_799, or_914_nl, fsm_output[0]);
  assign mux_1003_nl = MUX_s_1_2_2(mux_1002_nl, mux_1001_nl, fsm_output[4]);
  assign mux_1007_nl = MUX_s_1_2_2(mux_1006_nl, mux_1003_nl, fsm_output[6]);
  assign or_4135_nl = (fsm_output[2]) | mux_1007_nl;
  assign mux_1015_nl = MUX_s_1_2_2(nand_462_nl, or_4135_nl, fsm_output[5]);
  assign vec_rsc_0_7_i_we_d_pff = ~(mux_1015_nl | (fsm_output[1]));
  assign or_956_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_955_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1028_nl = MUX_s_1_2_2(or_956_nl, or_955_nl, fsm_output[0]);
  assign or_957_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1028_nl;
  assign or_953_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b000111)
      | (~ and_763_cse);
  assign mux_1025_nl = MUX_s_1_2_2(or_953_nl, or_tmp_809, fsm_output[0]);
  assign or_951_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b000111)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1024_nl = MUX_s_1_2_2(or_951_nl, or_tmp_805, fsm_output[0]);
  assign mux_1026_nl = MUX_s_1_2_2(mux_1025_nl, mux_1024_nl, fsm_output[4]);
  assign or_950_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b000111)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1022_nl = MUX_s_1_2_2(or_950_nl, or_tmp_803, fsm_output[0]);
  assign or_948_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b000111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1021_nl = MUX_s_1_2_2(or_948_nl, or_tmp_799, fsm_output[0]);
  assign mux_1023_nl = MUX_s_1_2_2(mux_1022_nl, mux_1021_nl, fsm_output[4]);
  assign mux_1027_nl = MUX_s_1_2_2(mux_1026_nl, mux_1023_nl, fsm_output[6]);
  assign mux_1029_nl = MUX_s_1_2_2(or_957_nl, mux_1027_nl, fsm_output[2]);
  assign or_946_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_944_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b000111) | (~ and_763_cse);
  assign mux_1018_nl = MUX_s_1_2_2(or_946_nl, or_944_nl, fsm_output[0]);
  assign or_942_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_941_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b000111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1017_nl = MUX_s_1_2_2(or_942_nl, or_941_nl, fsm_output[0]);
  assign mux_1019_nl = MUX_s_1_2_2(mux_1018_nl, mux_1017_nl, fsm_output[4]);
  assign nor_1335_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1336_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b000111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1016_nl = MUX_s_1_2_2(nor_1335_nl, nor_1336_nl, fsm_output[0]);
  assign nand_29_nl = ~((fsm_output[4]) & mux_1016_nl);
  assign mux_1020_nl = MUX_s_1_2_2(mux_1019_nl, nand_29_nl, fsm_output[6]);
  assign or_947_nl = (fsm_output[2]) | mux_1020_nl;
  assign mux_1030_nl = MUX_s_1_2_2(mux_1029_nl, or_947_nl, fsm_output[5]);
  assign vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1030_nl) & (fsm_output[1]);
  assign nor_1326_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001000) | (~ and_763_cse));
  assign nor_1327_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1042_nl = MUX_s_1_2_2(nor_1326_nl, nor_1327_nl, fsm_output[0]);
  assign nor_1328_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1329_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1041_nl = MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output[0]);
  assign mux_1043_nl = MUX_s_1_2_2(mux_1042_nl, mux_1041_nl, fsm_output[4]);
  assign nor_1330_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1331_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1039_nl = MUX_s_1_2_2(nor_1330_nl, nor_1331_nl, fsm_output[0]);
  assign nor_1332_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1333_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1038_nl = MUX_s_1_2_2(nor_1332_nl, nor_1333_nl, fsm_output[0]);
  assign mux_1040_nl = MUX_s_1_2_2(mux_1039_nl, mux_1038_nl, fsm_output[4]);
  assign mux_1044_nl = MUX_s_1_2_2(mux_1043_nl, mux_1040_nl, fsm_output[6]);
  assign nand_461_nl = ~((fsm_output[2]) & mux_1044_nl);
  assign or_967_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001000) | (~ and_763_cse);
  assign mux_1035_nl = MUX_s_1_2_2(or_tmp_853, or_967_nl, fsm_output[0]);
  assign or_964_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1034_nl = MUX_s_1_2_2(or_tmp_849, or_964_nl, fsm_output[0]);
  assign mux_1036_nl = MUX_s_1_2_2(mux_1035_nl, mux_1034_nl, fsm_output[4]);
  assign or_961_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1032_nl = MUX_s_1_2_2(or_tmp_847, or_961_nl, fsm_output[0]);
  assign or_958_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1031_nl = MUX_s_1_2_2(or_tmp_843, or_958_nl, fsm_output[0]);
  assign mux_1033_nl = MUX_s_1_2_2(mux_1032_nl, mux_1031_nl, fsm_output[4]);
  assign mux_1037_nl = MUX_s_1_2_2(mux_1036_nl, mux_1033_nl, fsm_output[6]);
  assign or_4134_nl = (fsm_output[2]) | mux_1037_nl;
  assign mux_1045_nl = MUX_s_1_2_2(nand_461_nl, or_4134_nl, fsm_output[5]);
  assign vec_rsc_0_8_i_we_d_pff = ~(mux_1045_nl | (fsm_output[1]));
  assign or_1000_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_999_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1058_nl = MUX_s_1_2_2(or_1000_nl, or_999_nl, fsm_output[0]);
  assign or_1001_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1058_nl;
  assign or_997_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001000)
      | (~ and_763_cse);
  assign mux_1055_nl = MUX_s_1_2_2(or_997_nl, or_tmp_853, fsm_output[0]);
  assign or_995_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1054_nl = MUX_s_1_2_2(or_995_nl, or_tmp_849, fsm_output[0]);
  assign mux_1056_nl = MUX_s_1_2_2(mux_1055_nl, mux_1054_nl, fsm_output[4]);
  assign or_994_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1052_nl = MUX_s_1_2_2(or_994_nl, or_tmp_847, fsm_output[0]);
  assign or_992_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1051_nl = MUX_s_1_2_2(or_992_nl, or_tmp_843, fsm_output[0]);
  assign mux_1053_nl = MUX_s_1_2_2(mux_1052_nl, mux_1051_nl, fsm_output[4]);
  assign mux_1057_nl = MUX_s_1_2_2(mux_1056_nl, mux_1053_nl, fsm_output[6]);
  assign mux_1059_nl = MUX_s_1_2_2(or_1001_nl, mux_1057_nl, fsm_output[2]);
  assign or_990_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_988_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001000) | (~ and_763_cse);
  assign mux_1048_nl = MUX_s_1_2_2(or_990_nl, or_988_nl, fsm_output[0]);
  assign or_986_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_985_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1047_nl = MUX_s_1_2_2(or_986_nl, or_985_nl, fsm_output[0]);
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, mux_1047_nl, fsm_output[4]);
  assign nor_1324_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1325_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1046_nl = MUX_s_1_2_2(nor_1324_nl, nor_1325_nl, fsm_output[0]);
  assign nand_31_nl = ~((fsm_output[4]) & mux_1046_nl);
  assign mux_1050_nl = MUX_s_1_2_2(mux_1049_nl, nand_31_nl, fsm_output[6]);
  assign or_991_nl = (fsm_output[2]) | mux_1050_nl;
  assign mux_1060_nl = MUX_s_1_2_2(mux_1059_nl, or_991_nl, fsm_output[5]);
  assign vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1060_nl) & (fsm_output[1]);
  assign nor_1315_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001001) | (~ and_763_cse));
  assign nor_1316_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1072_nl = MUX_s_1_2_2(nor_1315_nl, nor_1316_nl, fsm_output[0]);
  assign nor_1317_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1318_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1071_nl = MUX_s_1_2_2(nor_1317_nl, nor_1318_nl, fsm_output[0]);
  assign mux_1073_nl = MUX_s_1_2_2(mux_1072_nl, mux_1071_nl, fsm_output[4]);
  assign nor_1319_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1320_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1069_nl = MUX_s_1_2_2(nor_1319_nl, nor_1320_nl, fsm_output[0]);
  assign nor_1321_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1322_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1068_nl = MUX_s_1_2_2(nor_1321_nl, nor_1322_nl, fsm_output[0]);
  assign mux_1070_nl = MUX_s_1_2_2(mux_1069_nl, mux_1068_nl, fsm_output[4]);
  assign mux_1074_nl = MUX_s_1_2_2(mux_1073_nl, mux_1070_nl, fsm_output[6]);
  assign nand_460_nl = ~((fsm_output[2]) & mux_1074_nl);
  assign or_1011_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001001) | (~ and_763_cse);
  assign mux_1065_nl = MUX_s_1_2_2(or_tmp_897, or_1011_nl, fsm_output[0]);
  assign or_1008_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1064_nl = MUX_s_1_2_2(or_tmp_893, or_1008_nl, fsm_output[0]);
  assign mux_1066_nl = MUX_s_1_2_2(mux_1065_nl, mux_1064_nl, fsm_output[4]);
  assign or_1005_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1062_nl = MUX_s_1_2_2(or_tmp_891, or_1005_nl, fsm_output[0]);
  assign or_1002_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1061_nl = MUX_s_1_2_2(or_tmp_887, or_1002_nl, fsm_output[0]);
  assign mux_1063_nl = MUX_s_1_2_2(mux_1062_nl, mux_1061_nl, fsm_output[4]);
  assign mux_1067_nl = MUX_s_1_2_2(mux_1066_nl, mux_1063_nl, fsm_output[6]);
  assign or_4133_nl = (fsm_output[2]) | mux_1067_nl;
  assign mux_1075_nl = MUX_s_1_2_2(nand_460_nl, or_4133_nl, fsm_output[5]);
  assign vec_rsc_0_9_i_we_d_pff = ~(mux_1075_nl | (fsm_output[1]));
  assign or_1044_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1043_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1088_nl = MUX_s_1_2_2(or_1044_nl, or_1043_nl, fsm_output[0]);
  assign or_1045_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1088_nl;
  assign or_1041_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001001)
      | (~ and_763_cse);
  assign mux_1085_nl = MUX_s_1_2_2(or_1041_nl, or_tmp_897, fsm_output[0]);
  assign or_1039_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1084_nl = MUX_s_1_2_2(or_1039_nl, or_tmp_893, fsm_output[0]);
  assign mux_1086_nl = MUX_s_1_2_2(mux_1085_nl, mux_1084_nl, fsm_output[4]);
  assign or_1038_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1082_nl = MUX_s_1_2_2(or_1038_nl, or_tmp_891, fsm_output[0]);
  assign or_1036_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1081_nl = MUX_s_1_2_2(or_1036_nl, or_tmp_887, fsm_output[0]);
  assign mux_1083_nl = MUX_s_1_2_2(mux_1082_nl, mux_1081_nl, fsm_output[4]);
  assign mux_1087_nl = MUX_s_1_2_2(mux_1086_nl, mux_1083_nl, fsm_output[6]);
  assign mux_1089_nl = MUX_s_1_2_2(or_1045_nl, mux_1087_nl, fsm_output[2]);
  assign or_1034_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1032_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001001) | (~ and_763_cse);
  assign mux_1078_nl = MUX_s_1_2_2(or_1034_nl, or_1032_nl, fsm_output[0]);
  assign or_1030_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1029_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1077_nl = MUX_s_1_2_2(or_1030_nl, or_1029_nl, fsm_output[0]);
  assign mux_1079_nl = MUX_s_1_2_2(mux_1078_nl, mux_1077_nl, fsm_output[4]);
  assign nor_1313_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1314_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1076_nl = MUX_s_1_2_2(nor_1313_nl, nor_1314_nl, fsm_output[0]);
  assign nand_33_nl = ~((fsm_output[4]) & mux_1076_nl);
  assign mux_1080_nl = MUX_s_1_2_2(mux_1079_nl, nand_33_nl, fsm_output[6]);
  assign or_1035_nl = (fsm_output[2]) | mux_1080_nl;
  assign mux_1090_nl = MUX_s_1_2_2(mux_1089_nl, or_1035_nl, fsm_output[5]);
  assign vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1090_nl) & (fsm_output[1]);
  assign nor_1304_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001010) | (~ and_763_cse));
  assign nor_1305_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1102_nl = MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output[0]);
  assign nor_1306_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1307_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1101_nl = MUX_s_1_2_2(nor_1306_nl, nor_1307_nl, fsm_output[0]);
  assign mux_1103_nl = MUX_s_1_2_2(mux_1102_nl, mux_1101_nl, fsm_output[4]);
  assign nor_1308_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1309_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1099_nl = MUX_s_1_2_2(nor_1308_nl, nor_1309_nl, fsm_output[0]);
  assign nor_1310_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1311_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1098_nl = MUX_s_1_2_2(nor_1310_nl, nor_1311_nl, fsm_output[0]);
  assign mux_1100_nl = MUX_s_1_2_2(mux_1099_nl, mux_1098_nl, fsm_output[4]);
  assign mux_1104_nl = MUX_s_1_2_2(mux_1103_nl, mux_1100_nl, fsm_output[6]);
  assign nand_459_nl = ~((fsm_output[2]) & mux_1104_nl);
  assign or_1055_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001010) | (~ and_763_cse);
  assign mux_1095_nl = MUX_s_1_2_2(or_tmp_941, or_1055_nl, fsm_output[0]);
  assign or_1052_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1094_nl = MUX_s_1_2_2(or_tmp_937, or_1052_nl, fsm_output[0]);
  assign mux_1096_nl = MUX_s_1_2_2(mux_1095_nl, mux_1094_nl, fsm_output[4]);
  assign or_1049_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1092_nl = MUX_s_1_2_2(or_tmp_935, or_1049_nl, fsm_output[0]);
  assign or_1046_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1091_nl = MUX_s_1_2_2(or_tmp_931, or_1046_nl, fsm_output[0]);
  assign mux_1093_nl = MUX_s_1_2_2(mux_1092_nl, mux_1091_nl, fsm_output[4]);
  assign mux_1097_nl = MUX_s_1_2_2(mux_1096_nl, mux_1093_nl, fsm_output[6]);
  assign or_4132_nl = (fsm_output[2]) | mux_1097_nl;
  assign mux_1105_nl = MUX_s_1_2_2(nand_459_nl, or_4132_nl, fsm_output[5]);
  assign vec_rsc_0_10_i_we_d_pff = ~(mux_1105_nl | (fsm_output[1]));
  assign or_1088_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1087_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1118_nl = MUX_s_1_2_2(or_1088_nl, or_1087_nl, fsm_output[0]);
  assign or_1089_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1118_nl;
  assign or_1085_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001010)
      | (~ and_763_cse);
  assign mux_1115_nl = MUX_s_1_2_2(or_1085_nl, or_tmp_941, fsm_output[0]);
  assign or_1083_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1114_nl = MUX_s_1_2_2(or_1083_nl, or_tmp_937, fsm_output[0]);
  assign mux_1116_nl = MUX_s_1_2_2(mux_1115_nl, mux_1114_nl, fsm_output[4]);
  assign or_1082_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1112_nl = MUX_s_1_2_2(or_1082_nl, or_tmp_935, fsm_output[0]);
  assign or_1080_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1111_nl = MUX_s_1_2_2(or_1080_nl, or_tmp_931, fsm_output[0]);
  assign mux_1113_nl = MUX_s_1_2_2(mux_1112_nl, mux_1111_nl, fsm_output[4]);
  assign mux_1117_nl = MUX_s_1_2_2(mux_1116_nl, mux_1113_nl, fsm_output[6]);
  assign mux_1119_nl = MUX_s_1_2_2(or_1089_nl, mux_1117_nl, fsm_output[2]);
  assign or_1078_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1076_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001010) | (~ and_763_cse);
  assign mux_1108_nl = MUX_s_1_2_2(or_1078_nl, or_1076_nl, fsm_output[0]);
  assign or_1074_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1073_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1107_nl = MUX_s_1_2_2(or_1074_nl, or_1073_nl, fsm_output[0]);
  assign mux_1109_nl = MUX_s_1_2_2(mux_1108_nl, mux_1107_nl, fsm_output[4]);
  assign nor_1302_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1303_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1106_nl = MUX_s_1_2_2(nor_1302_nl, nor_1303_nl, fsm_output[0]);
  assign nand_35_nl = ~((fsm_output[4]) & mux_1106_nl);
  assign mux_1110_nl = MUX_s_1_2_2(mux_1109_nl, nand_35_nl, fsm_output[6]);
  assign or_1079_nl = (fsm_output[2]) | mux_1110_nl;
  assign mux_1120_nl = MUX_s_1_2_2(mux_1119_nl, or_1079_nl, fsm_output[5]);
  assign vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1120_nl) & (fsm_output[1]);
  assign nor_1293_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001011) | (~ and_763_cse));
  assign nor_1294_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | not_tmp_330);
  assign mux_1132_nl = MUX_s_1_2_2(nor_1293_nl, nor_1294_nl, fsm_output[0]);
  assign nor_1295_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1296_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1131_nl = MUX_s_1_2_2(nor_1295_nl, nor_1296_nl, fsm_output[0]);
  assign mux_1133_nl = MUX_s_1_2_2(mux_1132_nl, mux_1131_nl, fsm_output[4]);
  assign nor_1297_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1298_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1129_nl = MUX_s_1_2_2(nor_1297_nl, nor_1298_nl, fsm_output[0]);
  assign nor_1299_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1300_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1128_nl = MUX_s_1_2_2(nor_1299_nl, nor_1300_nl, fsm_output[0]);
  assign mux_1130_nl = MUX_s_1_2_2(mux_1129_nl, mux_1128_nl, fsm_output[4]);
  assign mux_1134_nl = MUX_s_1_2_2(mux_1133_nl, mux_1130_nl, fsm_output[6]);
  assign nand_458_nl = ~((fsm_output[2]) & mux_1134_nl);
  assign or_1099_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001011) | (~ and_763_cse);
  assign mux_1125_nl = MUX_s_1_2_2(or_tmp_985, or_1099_nl, fsm_output[0]);
  assign or_1096_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1124_nl = MUX_s_1_2_2(or_tmp_981, or_1096_nl, fsm_output[0]);
  assign mux_1126_nl = MUX_s_1_2_2(mux_1125_nl, mux_1124_nl, fsm_output[4]);
  assign or_1093_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1122_nl = MUX_s_1_2_2(or_tmp_979, or_1093_nl, fsm_output[0]);
  assign or_1090_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1121_nl = MUX_s_1_2_2(or_tmp_975, or_1090_nl, fsm_output[0]);
  assign mux_1123_nl = MUX_s_1_2_2(mux_1122_nl, mux_1121_nl, fsm_output[4]);
  assign mux_1127_nl = MUX_s_1_2_2(mux_1126_nl, mux_1123_nl, fsm_output[6]);
  assign or_4131_nl = (fsm_output[2]) | mux_1127_nl;
  assign mux_1135_nl = MUX_s_1_2_2(nand_458_nl, or_4131_nl, fsm_output[5]);
  assign vec_rsc_0_11_i_we_d_pff = ~(mux_1135_nl | (fsm_output[1]));
  assign or_1132_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1131_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1148_nl = MUX_s_1_2_2(or_1132_nl, or_1131_nl, fsm_output[0]);
  assign or_1133_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1148_nl;
  assign or_1129_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001011)
      | (~ and_763_cse);
  assign mux_1145_nl = MUX_s_1_2_2(or_1129_nl, or_tmp_985, fsm_output[0]);
  assign or_1127_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1144_nl = MUX_s_1_2_2(or_1127_nl, or_tmp_981, fsm_output[0]);
  assign mux_1146_nl = MUX_s_1_2_2(mux_1145_nl, mux_1144_nl, fsm_output[4]);
  assign or_1126_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1142_nl = MUX_s_1_2_2(or_1126_nl, or_tmp_979, fsm_output[0]);
  assign or_1124_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1141_nl = MUX_s_1_2_2(or_1124_nl, or_tmp_975, fsm_output[0]);
  assign mux_1143_nl = MUX_s_1_2_2(mux_1142_nl, mux_1141_nl, fsm_output[4]);
  assign mux_1147_nl = MUX_s_1_2_2(mux_1146_nl, mux_1143_nl, fsm_output[6]);
  assign mux_1149_nl = MUX_s_1_2_2(or_1133_nl, mux_1147_nl, fsm_output[2]);
  assign or_1122_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1120_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001011) | (~ and_763_cse);
  assign mux_1138_nl = MUX_s_1_2_2(or_1122_nl, or_1120_nl, fsm_output[0]);
  assign or_1118_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1117_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1137_nl = MUX_s_1_2_2(or_1118_nl, or_1117_nl, fsm_output[0]);
  assign mux_1139_nl = MUX_s_1_2_2(mux_1138_nl, mux_1137_nl, fsm_output[4]);
  assign nor_1291_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1292_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1136_nl = MUX_s_1_2_2(nor_1291_nl, nor_1292_nl, fsm_output[0]);
  assign nand_37_nl = ~((fsm_output[4]) & mux_1136_nl);
  assign mux_1140_nl = MUX_s_1_2_2(mux_1139_nl, nand_37_nl, fsm_output[6]);
  assign or_1123_nl = (fsm_output[2]) | mux_1140_nl;
  assign mux_1150_nl = MUX_s_1_2_2(mux_1149_nl, or_1123_nl, fsm_output[5]);
  assign vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1150_nl) & (fsm_output[1]);
  assign nor_1282_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001100) | (~ and_763_cse));
  assign nor_1283_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1162_nl = MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, fsm_output[0]);
  assign nor_1284_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1285_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1161_nl = MUX_s_1_2_2(nor_1284_nl, nor_1285_nl, fsm_output[0]);
  assign mux_1163_nl = MUX_s_1_2_2(mux_1162_nl, mux_1161_nl, fsm_output[4]);
  assign nor_1286_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1287_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1159_nl = MUX_s_1_2_2(nor_1286_nl, nor_1287_nl, fsm_output[0]);
  assign nor_1288_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1289_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1158_nl = MUX_s_1_2_2(nor_1288_nl, nor_1289_nl, fsm_output[0]);
  assign mux_1160_nl = MUX_s_1_2_2(mux_1159_nl, mux_1158_nl, fsm_output[4]);
  assign mux_1164_nl = MUX_s_1_2_2(mux_1163_nl, mux_1160_nl, fsm_output[6]);
  assign nand_457_nl = ~((fsm_output[2]) & mux_1164_nl);
  assign or_1143_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001100) | (~ and_763_cse);
  assign mux_1155_nl = MUX_s_1_2_2(or_tmp_1029, or_1143_nl, fsm_output[0]);
  assign or_1140_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1154_nl = MUX_s_1_2_2(or_tmp_1025, or_1140_nl, fsm_output[0]);
  assign mux_1156_nl = MUX_s_1_2_2(mux_1155_nl, mux_1154_nl, fsm_output[4]);
  assign or_1137_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1152_nl = MUX_s_1_2_2(or_tmp_1023, or_1137_nl, fsm_output[0]);
  assign or_1134_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1151_nl = MUX_s_1_2_2(or_tmp_1019, or_1134_nl, fsm_output[0]);
  assign mux_1153_nl = MUX_s_1_2_2(mux_1152_nl, mux_1151_nl, fsm_output[4]);
  assign mux_1157_nl = MUX_s_1_2_2(mux_1156_nl, mux_1153_nl, fsm_output[6]);
  assign or_4130_nl = (fsm_output[2]) | mux_1157_nl;
  assign mux_1165_nl = MUX_s_1_2_2(nand_457_nl, or_4130_nl, fsm_output[5]);
  assign vec_rsc_0_12_i_we_d_pff = ~(mux_1165_nl | (fsm_output[1]));
  assign or_1176_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1175_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1178_nl = MUX_s_1_2_2(or_1176_nl, or_1175_nl, fsm_output[0]);
  assign or_1177_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1178_nl;
  assign or_1173_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001100)
      | (~ and_763_cse);
  assign mux_1175_nl = MUX_s_1_2_2(or_1173_nl, or_tmp_1029, fsm_output[0]);
  assign or_1171_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1174_nl = MUX_s_1_2_2(or_1171_nl, or_tmp_1025, fsm_output[0]);
  assign mux_1176_nl = MUX_s_1_2_2(mux_1175_nl, mux_1174_nl, fsm_output[4]);
  assign or_1170_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1172_nl = MUX_s_1_2_2(or_1170_nl, or_tmp_1023, fsm_output[0]);
  assign or_1168_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1171_nl = MUX_s_1_2_2(or_1168_nl, or_tmp_1019, fsm_output[0]);
  assign mux_1173_nl = MUX_s_1_2_2(mux_1172_nl, mux_1171_nl, fsm_output[4]);
  assign mux_1177_nl = MUX_s_1_2_2(mux_1176_nl, mux_1173_nl, fsm_output[6]);
  assign mux_1179_nl = MUX_s_1_2_2(or_1177_nl, mux_1177_nl, fsm_output[2]);
  assign or_1166_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1164_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001100) | (~ and_763_cse);
  assign mux_1168_nl = MUX_s_1_2_2(or_1166_nl, or_1164_nl, fsm_output[0]);
  assign or_1162_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1161_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1167_nl = MUX_s_1_2_2(or_1162_nl, or_1161_nl, fsm_output[0]);
  assign mux_1169_nl = MUX_s_1_2_2(mux_1168_nl, mux_1167_nl, fsm_output[4]);
  assign nor_1280_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1281_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1166_nl = MUX_s_1_2_2(nor_1280_nl, nor_1281_nl, fsm_output[0]);
  assign nand_39_nl = ~((fsm_output[4]) & mux_1166_nl);
  assign mux_1170_nl = MUX_s_1_2_2(mux_1169_nl, nand_39_nl, fsm_output[6]);
  assign or_1167_nl = (fsm_output[2]) | mux_1170_nl;
  assign mux_1180_nl = MUX_s_1_2_2(mux_1179_nl, or_1167_nl, fsm_output[5]);
  assign vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1180_nl) & (fsm_output[1]);
  assign nor_1271_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001101) | (~ and_763_cse));
  assign nor_1272_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1192_nl = MUX_s_1_2_2(nor_1271_nl, nor_1272_nl, fsm_output[0]);
  assign nor_1273_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1274_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1191_nl = MUX_s_1_2_2(nor_1273_nl, nor_1274_nl, fsm_output[0]);
  assign mux_1193_nl = MUX_s_1_2_2(mux_1192_nl, mux_1191_nl, fsm_output[4]);
  assign nor_1275_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1276_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1189_nl = MUX_s_1_2_2(nor_1275_nl, nor_1276_nl, fsm_output[0]);
  assign nor_1277_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1278_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1188_nl = MUX_s_1_2_2(nor_1277_nl, nor_1278_nl, fsm_output[0]);
  assign mux_1190_nl = MUX_s_1_2_2(mux_1189_nl, mux_1188_nl, fsm_output[4]);
  assign mux_1194_nl = MUX_s_1_2_2(mux_1193_nl, mux_1190_nl, fsm_output[6]);
  assign nand_456_nl = ~((fsm_output[2]) & mux_1194_nl);
  assign or_1187_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001101) | (~ and_763_cse);
  assign mux_1185_nl = MUX_s_1_2_2(or_tmp_1073, or_1187_nl, fsm_output[0]);
  assign or_1184_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1184_nl = MUX_s_1_2_2(or_tmp_1069, or_1184_nl, fsm_output[0]);
  assign mux_1186_nl = MUX_s_1_2_2(mux_1185_nl, mux_1184_nl, fsm_output[4]);
  assign or_1181_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1182_nl = MUX_s_1_2_2(or_tmp_1067, or_1181_nl, fsm_output[0]);
  assign or_1178_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1181_nl = MUX_s_1_2_2(or_tmp_1063, or_1178_nl, fsm_output[0]);
  assign mux_1183_nl = MUX_s_1_2_2(mux_1182_nl, mux_1181_nl, fsm_output[4]);
  assign mux_1187_nl = MUX_s_1_2_2(mux_1186_nl, mux_1183_nl, fsm_output[6]);
  assign or_4129_nl = (fsm_output[2]) | mux_1187_nl;
  assign mux_1195_nl = MUX_s_1_2_2(nand_456_nl, or_4129_nl, fsm_output[5]);
  assign vec_rsc_0_13_i_we_d_pff = ~(mux_1195_nl | (fsm_output[1]));
  assign or_1220_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1219_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1208_nl = MUX_s_1_2_2(or_1220_nl, or_1219_nl, fsm_output[0]);
  assign or_1221_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1208_nl;
  assign or_1217_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001101)
      | (~ and_763_cse);
  assign mux_1205_nl = MUX_s_1_2_2(or_1217_nl, or_tmp_1073, fsm_output[0]);
  assign or_1215_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1204_nl = MUX_s_1_2_2(or_1215_nl, or_tmp_1069, fsm_output[0]);
  assign mux_1206_nl = MUX_s_1_2_2(mux_1205_nl, mux_1204_nl, fsm_output[4]);
  assign or_1214_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1202_nl = MUX_s_1_2_2(or_1214_nl, or_tmp_1067, fsm_output[0]);
  assign or_1212_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1201_nl = MUX_s_1_2_2(or_1212_nl, or_tmp_1063, fsm_output[0]);
  assign mux_1203_nl = MUX_s_1_2_2(mux_1202_nl, mux_1201_nl, fsm_output[4]);
  assign mux_1207_nl = MUX_s_1_2_2(mux_1206_nl, mux_1203_nl, fsm_output[6]);
  assign mux_1209_nl = MUX_s_1_2_2(or_1221_nl, mux_1207_nl, fsm_output[2]);
  assign or_1210_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1208_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001101) | (~ and_763_cse);
  assign mux_1198_nl = MUX_s_1_2_2(or_1210_nl, or_1208_nl, fsm_output[0]);
  assign or_1206_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1205_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1197_nl = MUX_s_1_2_2(or_1206_nl, or_1205_nl, fsm_output[0]);
  assign mux_1199_nl = MUX_s_1_2_2(mux_1198_nl, mux_1197_nl, fsm_output[4]);
  assign nor_1269_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1270_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1196_nl = MUX_s_1_2_2(nor_1269_nl, nor_1270_nl, fsm_output[0]);
  assign nand_41_nl = ~((fsm_output[4]) & mux_1196_nl);
  assign mux_1200_nl = MUX_s_1_2_2(mux_1199_nl, nand_41_nl, fsm_output[6]);
  assign or_1211_nl = (fsm_output[2]) | mux_1200_nl;
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_nl, or_1211_nl, fsm_output[5]);
  assign vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1210_nl) & (fsm_output[1]);
  assign nor_1260_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001110) | (~ and_763_cse));
  assign nor_1261_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1222_nl = MUX_s_1_2_2(nor_1260_nl, nor_1261_nl, fsm_output[0]);
  assign nor_1262_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1263_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1221_nl = MUX_s_1_2_2(nor_1262_nl, nor_1263_nl, fsm_output[0]);
  assign mux_1223_nl = MUX_s_1_2_2(mux_1222_nl, mux_1221_nl, fsm_output[4]);
  assign nor_1264_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1265_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1219_nl = MUX_s_1_2_2(nor_1264_nl, nor_1265_nl, fsm_output[0]);
  assign nor_1266_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1267_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1218_nl = MUX_s_1_2_2(nor_1266_nl, nor_1267_nl, fsm_output[0]);
  assign mux_1220_nl = MUX_s_1_2_2(mux_1219_nl, mux_1218_nl, fsm_output[4]);
  assign mux_1224_nl = MUX_s_1_2_2(mux_1223_nl, mux_1220_nl, fsm_output[6]);
  assign nand_455_nl = ~((fsm_output[2]) & mux_1224_nl);
  assign or_1231_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001110) | (~ and_763_cse);
  assign mux_1215_nl = MUX_s_1_2_2(or_tmp_1117, or_1231_nl, fsm_output[0]);
  assign or_1228_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1214_nl = MUX_s_1_2_2(or_tmp_1113, or_1228_nl, fsm_output[0]);
  assign mux_1216_nl = MUX_s_1_2_2(mux_1215_nl, mux_1214_nl, fsm_output[4]);
  assign or_1225_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1212_nl = MUX_s_1_2_2(or_tmp_1111, or_1225_nl, fsm_output[0]);
  assign or_1222_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1211_nl = MUX_s_1_2_2(or_tmp_1107, or_1222_nl, fsm_output[0]);
  assign mux_1213_nl = MUX_s_1_2_2(mux_1212_nl, mux_1211_nl, fsm_output[4]);
  assign mux_1217_nl = MUX_s_1_2_2(mux_1216_nl, mux_1213_nl, fsm_output[6]);
  assign or_4128_nl = (fsm_output[2]) | mux_1217_nl;
  assign mux_1225_nl = MUX_s_1_2_2(nand_455_nl, or_4128_nl, fsm_output[5]);
  assign vec_rsc_0_14_i_we_d_pff = ~(mux_1225_nl | (fsm_output[1]));
  assign or_1264_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1263_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1238_nl = MUX_s_1_2_2(or_1264_nl, or_1263_nl, fsm_output[0]);
  assign or_1265_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1238_nl;
  assign or_1261_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b001110)
      | (~ and_763_cse);
  assign mux_1235_nl = MUX_s_1_2_2(or_1261_nl, or_tmp_1117, fsm_output[0]);
  assign or_1259_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1234_nl = MUX_s_1_2_2(or_1259_nl, or_tmp_1113, fsm_output[0]);
  assign mux_1236_nl = MUX_s_1_2_2(mux_1235_nl, mux_1234_nl, fsm_output[4]);
  assign or_1258_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1232_nl = MUX_s_1_2_2(or_1258_nl, or_tmp_1111, fsm_output[0]);
  assign or_1256_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1231_nl = MUX_s_1_2_2(or_1256_nl, or_tmp_1107, fsm_output[0]);
  assign mux_1233_nl = MUX_s_1_2_2(mux_1232_nl, mux_1231_nl, fsm_output[4]);
  assign mux_1237_nl = MUX_s_1_2_2(mux_1236_nl, mux_1233_nl, fsm_output[6]);
  assign mux_1239_nl = MUX_s_1_2_2(or_1265_nl, mux_1237_nl, fsm_output[2]);
  assign or_1254_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00111) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1252_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001110) | (~ and_763_cse);
  assign mux_1228_nl = MUX_s_1_2_2(or_1254_nl, or_1252_nl, fsm_output[0]);
  assign or_1250_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00111) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1249_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1227_nl = MUX_s_1_2_2(or_1250_nl, or_1249_nl, fsm_output[0]);
  assign mux_1229_nl = MUX_s_1_2_2(mux_1228_nl, mux_1227_nl, fsm_output[4]);
  assign nor_1258_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1259_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1226_nl = MUX_s_1_2_2(nor_1258_nl, nor_1259_nl, fsm_output[0]);
  assign nand_43_nl = ~((fsm_output[4]) & mux_1226_nl);
  assign mux_1230_nl = MUX_s_1_2_2(mux_1229_nl, nand_43_nl, fsm_output[6]);
  assign or_1255_nl = (fsm_output[2]) | mux_1230_nl;
  assign mux_1240_nl = MUX_s_1_2_2(mux_1239_nl, or_1255_nl, fsm_output[5]);
  assign vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1240_nl) & (fsm_output[1]);
  assign and_618_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b001111) & and_763_cse;
  assign nor_1250_nl = ~((COMP_LOOP_acc_13_psp_sva[3:1]!=3'b001) | not_tmp_347);
  assign mux_1252_nl = MUX_s_1_2_2(and_618_nl, nor_1250_nl, fsm_output[0]);
  assign nor_1251_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b001111) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1252_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1251_nl = MUX_s_1_2_2(nor_1251_nl, nor_1252_nl, fsm_output[0]);
  assign mux_1253_nl = MUX_s_1_2_2(mux_1252_nl, mux_1251_nl, fsm_output[4]);
  assign nor_1253_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1254_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00111) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1249_nl = MUX_s_1_2_2(nor_1253_nl, nor_1254_nl, fsm_output[0]);
  assign nor_1255_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1256_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00111) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1248_nl = MUX_s_1_2_2(nor_1255_nl, nor_1256_nl, fsm_output[0]);
  assign mux_1250_nl = MUX_s_1_2_2(mux_1249_nl, mux_1248_nl, fsm_output[4]);
  assign mux_1254_nl = MUX_s_1_2_2(mux_1253_nl, mux_1250_nl, fsm_output[6]);
  assign nand_454_nl = ~((fsm_output[2]) & mux_1254_nl);
  assign nand_332_nl = ~((COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b001111) & and_763_cse);
  assign mux_1245_nl = MUX_s_1_2_2(or_tmp_1161, nand_332_nl, fsm_output[0]);
  assign or_1272_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1244_nl = MUX_s_1_2_2(or_tmp_1157, or_1272_nl, fsm_output[0]);
  assign mux_1246_nl = MUX_s_1_2_2(mux_1245_nl, mux_1244_nl, fsm_output[4]);
  assign or_1269_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1242_nl = MUX_s_1_2_2(or_tmp_1155, or_1269_nl, fsm_output[0]);
  assign or_1266_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1241_nl = MUX_s_1_2_2(or_tmp_1151, or_1266_nl, fsm_output[0]);
  assign mux_1243_nl = MUX_s_1_2_2(mux_1242_nl, mux_1241_nl, fsm_output[4]);
  assign mux_1247_nl = MUX_s_1_2_2(mux_1246_nl, mux_1243_nl, fsm_output[6]);
  assign or_4127_nl = (fsm_output[2]) | mux_1247_nl;
  assign mux_1255_nl = MUX_s_1_2_2(nand_454_nl, or_4127_nl, fsm_output[5]);
  assign vec_rsc_0_15_i_we_d_pff = ~(mux_1255_nl | (fsm_output[1]));
  assign or_1308_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b001111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1307_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1268_nl = MUX_s_1_2_2(or_1308_nl, or_1307_nl, fsm_output[0]);
  assign or_1309_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1268_nl;
  assign nand_330_nl = ~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b001111)
      & and_763_cse);
  assign mux_1265_nl = MUX_s_1_2_2(nand_330_nl, or_tmp_1161, fsm_output[0]);
  assign or_1303_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b001111)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1264_nl = MUX_s_1_2_2(or_1303_nl, or_tmp_1157, fsm_output[0]);
  assign mux_1266_nl = MUX_s_1_2_2(mux_1265_nl, mux_1264_nl, fsm_output[4]);
  assign or_1302_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b001111)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1262_nl = MUX_s_1_2_2(or_1302_nl, or_tmp_1155, fsm_output[0]);
  assign or_1300_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b001111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1261_nl = MUX_s_1_2_2(or_1300_nl, or_tmp_1151, fsm_output[0]);
  assign mux_1263_nl = MUX_s_1_2_2(mux_1262_nl, mux_1261_nl, fsm_output[4]);
  assign mux_1267_nl = MUX_s_1_2_2(mux_1266_nl, mux_1263_nl, fsm_output[6]);
  assign mux_1269_nl = MUX_s_1_2_2(or_1309_nl, mux_1267_nl, fsm_output[2]);
  assign or_1298_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b00111) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign nand_331_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b001111) & and_763_cse);
  assign mux_1258_nl = MUX_s_1_2_2(or_1298_nl, nand_331_nl, fsm_output[0]);
  assign or_1294_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b00111) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1293_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b001111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1257_nl = MUX_s_1_2_2(or_1294_nl, or_1293_nl, fsm_output[0]);
  assign mux_1259_nl = MUX_s_1_2_2(mux_1258_nl, mux_1257_nl, fsm_output[4]);
  assign nor_1248_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1249_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b001111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1256_nl = MUX_s_1_2_2(nor_1248_nl, nor_1249_nl, fsm_output[0]);
  assign nand_45_nl = ~((fsm_output[4]) & mux_1256_nl);
  assign mux_1260_nl = MUX_s_1_2_2(mux_1259_nl, nand_45_nl, fsm_output[6]);
  assign or_1299_nl = (fsm_output[2]) | mux_1260_nl;
  assign mux_1270_nl = MUX_s_1_2_2(mux_1269_nl, or_1299_nl, fsm_output[5]);
  assign vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1270_nl) & (fsm_output[1]);
  assign nor_1239_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1240_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1282_nl = MUX_s_1_2_2(nor_1239_nl, nor_1240_nl, fsm_output[0]);
  assign nor_1241_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1242_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1281_nl = MUX_s_1_2_2(nor_1241_nl, nor_1242_nl, fsm_output[0]);
  assign mux_1283_nl = MUX_s_1_2_2(mux_1282_nl, mux_1281_nl, fsm_output[4]);
  assign nor_1243_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1244_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1279_nl = MUX_s_1_2_2(nor_1243_nl, nor_1244_nl, fsm_output[0]);
  assign nor_1245_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1246_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1278_nl = MUX_s_1_2_2(nor_1245_nl, nor_1246_nl, fsm_output[0]);
  assign mux_1280_nl = MUX_s_1_2_2(mux_1279_nl, mux_1278_nl, fsm_output[4]);
  assign mux_1284_nl = MUX_s_1_2_2(mux_1283_nl, mux_1280_nl, fsm_output[6]);
  assign nand_453_nl = ~((fsm_output[2]) & mux_1284_nl);
  assign or_1319_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010000) | (~ and_763_cse);
  assign mux_1275_nl = MUX_s_1_2_2(or_tmp_1205, or_1319_nl, fsm_output[0]);
  assign or_1316_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1274_nl = MUX_s_1_2_2(or_tmp_1201, or_1316_nl, fsm_output[0]);
  assign mux_1276_nl = MUX_s_1_2_2(mux_1275_nl, mux_1274_nl, fsm_output[4]);
  assign or_1313_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1272_nl = MUX_s_1_2_2(or_tmp_1199, or_1313_nl, fsm_output[0]);
  assign or_1310_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1271_nl = MUX_s_1_2_2(or_tmp_1195, or_1310_nl, fsm_output[0]);
  assign mux_1273_nl = MUX_s_1_2_2(mux_1272_nl, mux_1271_nl, fsm_output[4]);
  assign mux_1277_nl = MUX_s_1_2_2(mux_1276_nl, mux_1273_nl, fsm_output[6]);
  assign or_4126_nl = (fsm_output[2]) | mux_1277_nl;
  assign mux_1285_nl = MUX_s_1_2_2(nand_453_nl, or_4126_nl, fsm_output[5]);
  assign vec_rsc_0_16_i_we_d_pff = ~(mux_1285_nl | (fsm_output[1]));
  assign or_1352_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1351_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1298_nl = MUX_s_1_2_2(or_1352_nl, or_1351_nl, fsm_output[0]);
  assign or_1353_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1298_nl;
  assign or_1349_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010000)
      | (~ and_763_cse);
  assign mux_1295_nl = MUX_s_1_2_2(or_1349_nl, or_tmp_1205, fsm_output[0]);
  assign or_1347_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1294_nl = MUX_s_1_2_2(or_1347_nl, or_tmp_1201, fsm_output[0]);
  assign mux_1296_nl = MUX_s_1_2_2(mux_1295_nl, mux_1294_nl, fsm_output[4]);
  assign or_1346_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1292_nl = MUX_s_1_2_2(or_1346_nl, or_tmp_1199, fsm_output[0]);
  assign or_1344_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1291_nl = MUX_s_1_2_2(or_1344_nl, or_tmp_1195, fsm_output[0]);
  assign mux_1293_nl = MUX_s_1_2_2(mux_1292_nl, mux_1291_nl, fsm_output[4]);
  assign mux_1297_nl = MUX_s_1_2_2(mux_1296_nl, mux_1293_nl, fsm_output[6]);
  assign mux_1299_nl = MUX_s_1_2_2(or_1353_nl, mux_1297_nl, fsm_output[2]);
  assign or_1342_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1340_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1288_nl = MUX_s_1_2_2(or_1342_nl, or_1340_nl, fsm_output[0]);
  assign or_1338_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1337_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1287_nl = MUX_s_1_2_2(or_1338_nl, or_1337_nl, fsm_output[0]);
  assign mux_1289_nl = MUX_s_1_2_2(mux_1288_nl, mux_1287_nl, fsm_output[4]);
  assign nor_1237_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1238_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1286_nl = MUX_s_1_2_2(nor_1237_nl, nor_1238_nl, fsm_output[0]);
  assign nand_47_nl = ~((fsm_output[4]) & mux_1286_nl);
  assign mux_1290_nl = MUX_s_1_2_2(mux_1289_nl, nand_47_nl, fsm_output[6]);
  assign or_1343_nl = (fsm_output[2]) | mux_1290_nl;
  assign mux_1300_nl = MUX_s_1_2_2(mux_1299_nl, or_1343_nl, fsm_output[5]);
  assign vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1300_nl) & (fsm_output[1]);
  assign nor_1228_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1229_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1312_nl = MUX_s_1_2_2(nor_1228_nl, nor_1229_nl, fsm_output[0]);
  assign nor_1230_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1231_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1311_nl = MUX_s_1_2_2(nor_1230_nl, nor_1231_nl, fsm_output[0]);
  assign mux_1313_nl = MUX_s_1_2_2(mux_1312_nl, mux_1311_nl, fsm_output[4]);
  assign nor_1232_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1233_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1309_nl = MUX_s_1_2_2(nor_1232_nl, nor_1233_nl, fsm_output[0]);
  assign nor_1234_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1235_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1308_nl = MUX_s_1_2_2(nor_1234_nl, nor_1235_nl, fsm_output[0]);
  assign mux_1310_nl = MUX_s_1_2_2(mux_1309_nl, mux_1308_nl, fsm_output[4]);
  assign mux_1314_nl = MUX_s_1_2_2(mux_1313_nl, mux_1310_nl, fsm_output[6]);
  assign nand_452_nl = ~((fsm_output[2]) & mux_1314_nl);
  assign or_1363_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010001) | (~ and_763_cse);
  assign mux_1305_nl = MUX_s_1_2_2(or_tmp_1249, or_1363_nl, fsm_output[0]);
  assign or_1360_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1304_nl = MUX_s_1_2_2(or_tmp_1245, or_1360_nl, fsm_output[0]);
  assign mux_1306_nl = MUX_s_1_2_2(mux_1305_nl, mux_1304_nl, fsm_output[4]);
  assign or_1357_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1302_nl = MUX_s_1_2_2(or_tmp_1243, or_1357_nl, fsm_output[0]);
  assign or_1354_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1301_nl = MUX_s_1_2_2(or_tmp_1239, or_1354_nl, fsm_output[0]);
  assign mux_1303_nl = MUX_s_1_2_2(mux_1302_nl, mux_1301_nl, fsm_output[4]);
  assign mux_1307_nl = MUX_s_1_2_2(mux_1306_nl, mux_1303_nl, fsm_output[6]);
  assign or_4125_nl = (fsm_output[2]) | mux_1307_nl;
  assign mux_1315_nl = MUX_s_1_2_2(nand_452_nl, or_4125_nl, fsm_output[5]);
  assign vec_rsc_0_17_i_we_d_pff = ~(mux_1315_nl | (fsm_output[1]));
  assign or_1396_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1395_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1328_nl = MUX_s_1_2_2(or_1396_nl, or_1395_nl, fsm_output[0]);
  assign or_1397_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1328_nl;
  assign or_1393_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010001)
      | (~ and_763_cse);
  assign mux_1325_nl = MUX_s_1_2_2(or_1393_nl, or_tmp_1249, fsm_output[0]);
  assign or_1391_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1324_nl = MUX_s_1_2_2(or_1391_nl, or_tmp_1245, fsm_output[0]);
  assign mux_1326_nl = MUX_s_1_2_2(mux_1325_nl, mux_1324_nl, fsm_output[4]);
  assign or_1390_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1322_nl = MUX_s_1_2_2(or_1390_nl, or_tmp_1243, fsm_output[0]);
  assign or_1388_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1321_nl = MUX_s_1_2_2(or_1388_nl, or_tmp_1239, fsm_output[0]);
  assign mux_1323_nl = MUX_s_1_2_2(mux_1322_nl, mux_1321_nl, fsm_output[4]);
  assign mux_1327_nl = MUX_s_1_2_2(mux_1326_nl, mux_1323_nl, fsm_output[6]);
  assign mux_1329_nl = MUX_s_1_2_2(or_1397_nl, mux_1327_nl, fsm_output[2]);
  assign or_1386_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1384_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1318_nl = MUX_s_1_2_2(or_1386_nl, or_1384_nl, fsm_output[0]);
  assign or_1382_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1381_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1317_nl = MUX_s_1_2_2(or_1382_nl, or_1381_nl, fsm_output[0]);
  assign mux_1319_nl = MUX_s_1_2_2(mux_1318_nl, mux_1317_nl, fsm_output[4]);
  assign nor_1226_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1227_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1316_nl = MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, fsm_output[0]);
  assign nand_49_nl = ~((fsm_output[4]) & mux_1316_nl);
  assign mux_1320_nl = MUX_s_1_2_2(mux_1319_nl, nand_49_nl, fsm_output[6]);
  assign or_1387_nl = (fsm_output[2]) | mux_1320_nl;
  assign mux_1330_nl = MUX_s_1_2_2(mux_1329_nl, or_1387_nl, fsm_output[5]);
  assign vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1330_nl) & (fsm_output[1]);
  assign nor_1217_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1218_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1342_nl = MUX_s_1_2_2(nor_1217_nl, nor_1218_nl, fsm_output[0]);
  assign nor_1219_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1220_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1341_nl = MUX_s_1_2_2(nor_1219_nl, nor_1220_nl, fsm_output[0]);
  assign mux_1343_nl = MUX_s_1_2_2(mux_1342_nl, mux_1341_nl, fsm_output[4]);
  assign nor_1221_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1222_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1339_nl = MUX_s_1_2_2(nor_1221_nl, nor_1222_nl, fsm_output[0]);
  assign nor_1223_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1224_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1338_nl = MUX_s_1_2_2(nor_1223_nl, nor_1224_nl, fsm_output[0]);
  assign mux_1340_nl = MUX_s_1_2_2(mux_1339_nl, mux_1338_nl, fsm_output[4]);
  assign mux_1344_nl = MUX_s_1_2_2(mux_1343_nl, mux_1340_nl, fsm_output[6]);
  assign nand_451_nl = ~((fsm_output[2]) & mux_1344_nl);
  assign or_1407_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010010) | (~ and_763_cse);
  assign mux_1335_nl = MUX_s_1_2_2(or_tmp_1293, or_1407_nl, fsm_output[0]);
  assign or_1404_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1334_nl = MUX_s_1_2_2(or_tmp_1289, or_1404_nl, fsm_output[0]);
  assign mux_1336_nl = MUX_s_1_2_2(mux_1335_nl, mux_1334_nl, fsm_output[4]);
  assign or_1401_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1332_nl = MUX_s_1_2_2(or_tmp_1287, or_1401_nl, fsm_output[0]);
  assign or_1398_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1331_nl = MUX_s_1_2_2(or_tmp_1283, or_1398_nl, fsm_output[0]);
  assign mux_1333_nl = MUX_s_1_2_2(mux_1332_nl, mux_1331_nl, fsm_output[4]);
  assign mux_1337_nl = MUX_s_1_2_2(mux_1336_nl, mux_1333_nl, fsm_output[6]);
  assign or_4124_nl = (fsm_output[2]) | mux_1337_nl;
  assign mux_1345_nl = MUX_s_1_2_2(nand_451_nl, or_4124_nl, fsm_output[5]);
  assign vec_rsc_0_18_i_we_d_pff = ~(mux_1345_nl | (fsm_output[1]));
  assign or_1440_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1439_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1358_nl = MUX_s_1_2_2(or_1440_nl, or_1439_nl, fsm_output[0]);
  assign or_1441_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1358_nl;
  assign or_1437_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010010)
      | (~ and_763_cse);
  assign mux_1355_nl = MUX_s_1_2_2(or_1437_nl, or_tmp_1293, fsm_output[0]);
  assign or_1435_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1354_nl = MUX_s_1_2_2(or_1435_nl, or_tmp_1289, fsm_output[0]);
  assign mux_1356_nl = MUX_s_1_2_2(mux_1355_nl, mux_1354_nl, fsm_output[4]);
  assign or_1434_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1352_nl = MUX_s_1_2_2(or_1434_nl, or_tmp_1287, fsm_output[0]);
  assign or_1432_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1351_nl = MUX_s_1_2_2(or_1432_nl, or_tmp_1283, fsm_output[0]);
  assign mux_1353_nl = MUX_s_1_2_2(mux_1352_nl, mux_1351_nl, fsm_output[4]);
  assign mux_1357_nl = MUX_s_1_2_2(mux_1356_nl, mux_1353_nl, fsm_output[6]);
  assign mux_1359_nl = MUX_s_1_2_2(or_1441_nl, mux_1357_nl, fsm_output[2]);
  assign or_1430_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1428_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1348_nl = MUX_s_1_2_2(or_1430_nl, or_1428_nl, fsm_output[0]);
  assign or_1426_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1425_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1347_nl = MUX_s_1_2_2(or_1426_nl, or_1425_nl, fsm_output[0]);
  assign mux_1349_nl = MUX_s_1_2_2(mux_1348_nl, mux_1347_nl, fsm_output[4]);
  assign nor_1215_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1216_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1346_nl = MUX_s_1_2_2(nor_1215_nl, nor_1216_nl, fsm_output[0]);
  assign nand_51_nl = ~((fsm_output[4]) & mux_1346_nl);
  assign mux_1350_nl = MUX_s_1_2_2(mux_1349_nl, nand_51_nl, fsm_output[6]);
  assign or_1431_nl = (fsm_output[2]) | mux_1350_nl;
  assign mux_1360_nl = MUX_s_1_2_2(mux_1359_nl, or_1431_nl, fsm_output[5]);
  assign vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1360_nl) & (fsm_output[1]);
  assign nor_1206_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1207_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | not_tmp_330);
  assign mux_1372_nl = MUX_s_1_2_2(nor_1206_nl, nor_1207_nl, fsm_output[0]);
  assign nor_1208_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1209_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1371_nl = MUX_s_1_2_2(nor_1208_nl, nor_1209_nl, fsm_output[0]);
  assign mux_1373_nl = MUX_s_1_2_2(mux_1372_nl, mux_1371_nl, fsm_output[4]);
  assign nor_1210_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1211_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1369_nl = MUX_s_1_2_2(nor_1210_nl, nor_1211_nl, fsm_output[0]);
  assign nor_1212_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1213_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1368_nl = MUX_s_1_2_2(nor_1212_nl, nor_1213_nl, fsm_output[0]);
  assign mux_1370_nl = MUX_s_1_2_2(mux_1369_nl, mux_1368_nl, fsm_output[4]);
  assign mux_1374_nl = MUX_s_1_2_2(mux_1373_nl, mux_1370_nl, fsm_output[6]);
  assign nand_450_nl = ~((fsm_output[2]) & mux_1374_nl);
  assign or_1451_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010011) | (~ and_763_cse);
  assign mux_1365_nl = MUX_s_1_2_2(or_tmp_1337, or_1451_nl, fsm_output[0]);
  assign or_1448_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1364_nl = MUX_s_1_2_2(or_tmp_1333, or_1448_nl, fsm_output[0]);
  assign mux_1366_nl = MUX_s_1_2_2(mux_1365_nl, mux_1364_nl, fsm_output[4]);
  assign or_1445_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1362_nl = MUX_s_1_2_2(or_tmp_1331, or_1445_nl, fsm_output[0]);
  assign or_1442_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1361_nl = MUX_s_1_2_2(or_tmp_1327, or_1442_nl, fsm_output[0]);
  assign mux_1363_nl = MUX_s_1_2_2(mux_1362_nl, mux_1361_nl, fsm_output[4]);
  assign mux_1367_nl = MUX_s_1_2_2(mux_1366_nl, mux_1363_nl, fsm_output[6]);
  assign or_4123_nl = (fsm_output[2]) | mux_1367_nl;
  assign mux_1375_nl = MUX_s_1_2_2(nand_450_nl, or_4123_nl, fsm_output[5]);
  assign vec_rsc_0_19_i_we_d_pff = ~(mux_1375_nl | (fsm_output[1]));
  assign or_1484_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1483_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1388_nl = MUX_s_1_2_2(or_1484_nl, or_1483_nl, fsm_output[0]);
  assign or_1485_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1388_nl;
  assign or_1481_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010011)
      | (~ and_763_cse);
  assign mux_1385_nl = MUX_s_1_2_2(or_1481_nl, or_tmp_1337, fsm_output[0]);
  assign or_1479_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1384_nl = MUX_s_1_2_2(or_1479_nl, or_tmp_1333, fsm_output[0]);
  assign mux_1386_nl = MUX_s_1_2_2(mux_1385_nl, mux_1384_nl, fsm_output[4]);
  assign or_1478_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1382_nl = MUX_s_1_2_2(or_1478_nl, or_tmp_1331, fsm_output[0]);
  assign or_1476_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1381_nl = MUX_s_1_2_2(or_1476_nl, or_tmp_1327, fsm_output[0]);
  assign mux_1383_nl = MUX_s_1_2_2(mux_1382_nl, mux_1381_nl, fsm_output[4]);
  assign mux_1387_nl = MUX_s_1_2_2(mux_1386_nl, mux_1383_nl, fsm_output[6]);
  assign mux_1389_nl = MUX_s_1_2_2(or_1485_nl, mux_1387_nl, fsm_output[2]);
  assign or_1474_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1472_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1378_nl = MUX_s_1_2_2(or_1474_nl, or_1472_nl, fsm_output[0]);
  assign or_1470_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1469_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1377_nl = MUX_s_1_2_2(or_1470_nl, or_1469_nl, fsm_output[0]);
  assign mux_1379_nl = MUX_s_1_2_2(mux_1378_nl, mux_1377_nl, fsm_output[4]);
  assign nor_1204_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1205_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1376_nl = MUX_s_1_2_2(nor_1204_nl, nor_1205_nl, fsm_output[0]);
  assign nand_53_nl = ~((fsm_output[4]) & mux_1376_nl);
  assign mux_1380_nl = MUX_s_1_2_2(mux_1379_nl, nand_53_nl, fsm_output[6]);
  assign or_1475_nl = (fsm_output[2]) | mux_1380_nl;
  assign mux_1390_nl = MUX_s_1_2_2(mux_1389_nl, or_1475_nl, fsm_output[5]);
  assign vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1390_nl) & (fsm_output[1]);
  assign nor_1195_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1196_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1402_nl = MUX_s_1_2_2(nor_1195_nl, nor_1196_nl, fsm_output[0]);
  assign nor_1197_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1198_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1401_nl = MUX_s_1_2_2(nor_1197_nl, nor_1198_nl, fsm_output[0]);
  assign mux_1403_nl = MUX_s_1_2_2(mux_1402_nl, mux_1401_nl, fsm_output[4]);
  assign nor_1199_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1200_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1399_nl = MUX_s_1_2_2(nor_1199_nl, nor_1200_nl, fsm_output[0]);
  assign nor_1201_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1202_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1398_nl = MUX_s_1_2_2(nor_1201_nl, nor_1202_nl, fsm_output[0]);
  assign mux_1400_nl = MUX_s_1_2_2(mux_1399_nl, mux_1398_nl, fsm_output[4]);
  assign mux_1404_nl = MUX_s_1_2_2(mux_1403_nl, mux_1400_nl, fsm_output[6]);
  assign nand_449_nl = ~((fsm_output[2]) & mux_1404_nl);
  assign or_1495_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010100) | (~ and_763_cse);
  assign mux_1395_nl = MUX_s_1_2_2(or_tmp_1381, or_1495_nl, fsm_output[0]);
  assign or_1492_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1394_nl = MUX_s_1_2_2(or_tmp_1377, or_1492_nl, fsm_output[0]);
  assign mux_1396_nl = MUX_s_1_2_2(mux_1395_nl, mux_1394_nl, fsm_output[4]);
  assign or_1489_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1392_nl = MUX_s_1_2_2(or_tmp_1375, or_1489_nl, fsm_output[0]);
  assign or_1486_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1391_nl = MUX_s_1_2_2(or_tmp_1371, or_1486_nl, fsm_output[0]);
  assign mux_1393_nl = MUX_s_1_2_2(mux_1392_nl, mux_1391_nl, fsm_output[4]);
  assign mux_1397_nl = MUX_s_1_2_2(mux_1396_nl, mux_1393_nl, fsm_output[6]);
  assign or_4122_nl = (fsm_output[2]) | mux_1397_nl;
  assign mux_1405_nl = MUX_s_1_2_2(nand_449_nl, or_4122_nl, fsm_output[5]);
  assign vec_rsc_0_20_i_we_d_pff = ~(mux_1405_nl | (fsm_output[1]));
  assign or_1528_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1527_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1418_nl = MUX_s_1_2_2(or_1528_nl, or_1527_nl, fsm_output[0]);
  assign or_1529_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1418_nl;
  assign or_1525_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010100)
      | (~ and_763_cse);
  assign mux_1415_nl = MUX_s_1_2_2(or_1525_nl, or_tmp_1381, fsm_output[0]);
  assign or_1523_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1414_nl = MUX_s_1_2_2(or_1523_nl, or_tmp_1377, fsm_output[0]);
  assign mux_1416_nl = MUX_s_1_2_2(mux_1415_nl, mux_1414_nl, fsm_output[4]);
  assign or_1522_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1412_nl = MUX_s_1_2_2(or_1522_nl, or_tmp_1375, fsm_output[0]);
  assign or_1520_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1411_nl = MUX_s_1_2_2(or_1520_nl, or_tmp_1371, fsm_output[0]);
  assign mux_1413_nl = MUX_s_1_2_2(mux_1412_nl, mux_1411_nl, fsm_output[4]);
  assign mux_1417_nl = MUX_s_1_2_2(mux_1416_nl, mux_1413_nl, fsm_output[6]);
  assign mux_1419_nl = MUX_s_1_2_2(or_1529_nl, mux_1417_nl, fsm_output[2]);
  assign or_1518_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1516_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1408_nl = MUX_s_1_2_2(or_1518_nl, or_1516_nl, fsm_output[0]);
  assign or_1514_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1513_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1407_nl = MUX_s_1_2_2(or_1514_nl, or_1513_nl, fsm_output[0]);
  assign mux_1409_nl = MUX_s_1_2_2(mux_1408_nl, mux_1407_nl, fsm_output[4]);
  assign nor_1193_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1194_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1406_nl = MUX_s_1_2_2(nor_1193_nl, nor_1194_nl, fsm_output[0]);
  assign nand_55_nl = ~((fsm_output[4]) & mux_1406_nl);
  assign mux_1410_nl = MUX_s_1_2_2(mux_1409_nl, nand_55_nl, fsm_output[6]);
  assign or_1519_nl = (fsm_output[2]) | mux_1410_nl;
  assign mux_1420_nl = MUX_s_1_2_2(mux_1419_nl, or_1519_nl, fsm_output[5]);
  assign vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1420_nl) & (fsm_output[1]);
  assign nor_1184_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1185_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1432_nl = MUX_s_1_2_2(nor_1184_nl, nor_1185_nl, fsm_output[0]);
  assign nor_1186_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1187_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1431_nl = MUX_s_1_2_2(nor_1186_nl, nor_1187_nl, fsm_output[0]);
  assign mux_1433_nl = MUX_s_1_2_2(mux_1432_nl, mux_1431_nl, fsm_output[4]);
  assign nor_1188_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1189_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1429_nl = MUX_s_1_2_2(nor_1188_nl, nor_1189_nl, fsm_output[0]);
  assign nor_1190_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1191_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1428_nl = MUX_s_1_2_2(nor_1190_nl, nor_1191_nl, fsm_output[0]);
  assign mux_1430_nl = MUX_s_1_2_2(mux_1429_nl, mux_1428_nl, fsm_output[4]);
  assign mux_1434_nl = MUX_s_1_2_2(mux_1433_nl, mux_1430_nl, fsm_output[6]);
  assign nand_448_nl = ~((fsm_output[2]) & mux_1434_nl);
  assign or_1539_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010101) | (~ and_763_cse);
  assign mux_1425_nl = MUX_s_1_2_2(or_tmp_1425, or_1539_nl, fsm_output[0]);
  assign or_1536_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1424_nl = MUX_s_1_2_2(or_tmp_1421, or_1536_nl, fsm_output[0]);
  assign mux_1426_nl = MUX_s_1_2_2(mux_1425_nl, mux_1424_nl, fsm_output[4]);
  assign or_1533_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1422_nl = MUX_s_1_2_2(or_tmp_1419, or_1533_nl, fsm_output[0]);
  assign or_1530_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1421_nl = MUX_s_1_2_2(or_tmp_1415, or_1530_nl, fsm_output[0]);
  assign mux_1423_nl = MUX_s_1_2_2(mux_1422_nl, mux_1421_nl, fsm_output[4]);
  assign mux_1427_nl = MUX_s_1_2_2(mux_1426_nl, mux_1423_nl, fsm_output[6]);
  assign or_4121_nl = (fsm_output[2]) | mux_1427_nl;
  assign mux_1435_nl = MUX_s_1_2_2(nand_448_nl, or_4121_nl, fsm_output[5]);
  assign vec_rsc_0_21_i_we_d_pff = ~(mux_1435_nl | (fsm_output[1]));
  assign or_1572_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1571_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1448_nl = MUX_s_1_2_2(or_1572_nl, or_1571_nl, fsm_output[0]);
  assign or_1573_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1448_nl;
  assign or_1569_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010101)
      | (~ and_763_cse);
  assign mux_1445_nl = MUX_s_1_2_2(or_1569_nl, or_tmp_1425, fsm_output[0]);
  assign or_1567_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1444_nl = MUX_s_1_2_2(or_1567_nl, or_tmp_1421, fsm_output[0]);
  assign mux_1446_nl = MUX_s_1_2_2(mux_1445_nl, mux_1444_nl, fsm_output[4]);
  assign or_1566_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1442_nl = MUX_s_1_2_2(or_1566_nl, or_tmp_1419, fsm_output[0]);
  assign or_1564_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1441_nl = MUX_s_1_2_2(or_1564_nl, or_tmp_1415, fsm_output[0]);
  assign mux_1443_nl = MUX_s_1_2_2(mux_1442_nl, mux_1441_nl, fsm_output[4]);
  assign mux_1447_nl = MUX_s_1_2_2(mux_1446_nl, mux_1443_nl, fsm_output[6]);
  assign mux_1449_nl = MUX_s_1_2_2(or_1573_nl, mux_1447_nl, fsm_output[2]);
  assign or_1562_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1560_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1438_nl = MUX_s_1_2_2(or_1562_nl, or_1560_nl, fsm_output[0]);
  assign or_1558_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1557_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1437_nl = MUX_s_1_2_2(or_1558_nl, or_1557_nl, fsm_output[0]);
  assign mux_1439_nl = MUX_s_1_2_2(mux_1438_nl, mux_1437_nl, fsm_output[4]);
  assign nor_1182_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1183_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1436_nl = MUX_s_1_2_2(nor_1182_nl, nor_1183_nl, fsm_output[0]);
  assign nand_57_nl = ~((fsm_output[4]) & mux_1436_nl);
  assign mux_1440_nl = MUX_s_1_2_2(mux_1439_nl, nand_57_nl, fsm_output[6]);
  assign or_1563_nl = (fsm_output[2]) | mux_1440_nl;
  assign mux_1450_nl = MUX_s_1_2_2(mux_1449_nl, or_1563_nl, fsm_output[5]);
  assign vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1450_nl) & (fsm_output[1]);
  assign nor_1173_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1174_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1462_nl = MUX_s_1_2_2(nor_1173_nl, nor_1174_nl, fsm_output[0]);
  assign nor_1175_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1176_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1461_nl = MUX_s_1_2_2(nor_1175_nl, nor_1176_nl, fsm_output[0]);
  assign mux_1463_nl = MUX_s_1_2_2(mux_1462_nl, mux_1461_nl, fsm_output[4]);
  assign nor_1177_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1178_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1459_nl = MUX_s_1_2_2(nor_1177_nl, nor_1178_nl, fsm_output[0]);
  assign nor_1179_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1180_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1458_nl = MUX_s_1_2_2(nor_1179_nl, nor_1180_nl, fsm_output[0]);
  assign mux_1460_nl = MUX_s_1_2_2(mux_1459_nl, mux_1458_nl, fsm_output[4]);
  assign mux_1464_nl = MUX_s_1_2_2(mux_1463_nl, mux_1460_nl, fsm_output[6]);
  assign nand_447_nl = ~((fsm_output[2]) & mux_1464_nl);
  assign or_1583_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010110) | (~ and_763_cse);
  assign mux_1455_nl = MUX_s_1_2_2(or_tmp_1469, or_1583_nl, fsm_output[0]);
  assign or_1580_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1454_nl = MUX_s_1_2_2(or_tmp_1465, or_1580_nl, fsm_output[0]);
  assign mux_1456_nl = MUX_s_1_2_2(mux_1455_nl, mux_1454_nl, fsm_output[4]);
  assign or_1577_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1452_nl = MUX_s_1_2_2(or_tmp_1463, or_1577_nl, fsm_output[0]);
  assign or_1574_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1451_nl = MUX_s_1_2_2(or_tmp_1459, or_1574_nl, fsm_output[0]);
  assign mux_1453_nl = MUX_s_1_2_2(mux_1452_nl, mux_1451_nl, fsm_output[4]);
  assign mux_1457_nl = MUX_s_1_2_2(mux_1456_nl, mux_1453_nl, fsm_output[6]);
  assign or_4120_nl = (fsm_output[2]) | mux_1457_nl;
  assign mux_1465_nl = MUX_s_1_2_2(nand_447_nl, or_4120_nl, fsm_output[5]);
  assign vec_rsc_0_22_i_we_d_pff = ~(mux_1465_nl | (fsm_output[1]));
  assign or_1616_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1615_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1478_nl = MUX_s_1_2_2(or_1616_nl, or_1615_nl, fsm_output[0]);
  assign or_1617_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1478_nl;
  assign or_1613_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b010110)
      | (~ and_763_cse);
  assign mux_1475_nl = MUX_s_1_2_2(or_1613_nl, or_tmp_1469, fsm_output[0]);
  assign or_1611_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1474_nl = MUX_s_1_2_2(or_1611_nl, or_tmp_1465, fsm_output[0]);
  assign mux_1476_nl = MUX_s_1_2_2(mux_1475_nl, mux_1474_nl, fsm_output[4]);
  assign or_1610_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1472_nl = MUX_s_1_2_2(or_1610_nl, or_tmp_1463, fsm_output[0]);
  assign or_1608_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1471_nl = MUX_s_1_2_2(or_1608_nl, or_tmp_1459, fsm_output[0]);
  assign mux_1473_nl = MUX_s_1_2_2(mux_1472_nl, mux_1471_nl, fsm_output[4]);
  assign mux_1477_nl = MUX_s_1_2_2(mux_1476_nl, mux_1473_nl, fsm_output[6]);
  assign mux_1479_nl = MUX_s_1_2_2(or_1617_nl, mux_1477_nl, fsm_output[2]);
  assign or_1606_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1604_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1468_nl = MUX_s_1_2_2(or_1606_nl, or_1604_nl, fsm_output[0]);
  assign or_1602_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1601_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1467_nl = MUX_s_1_2_2(or_1602_nl, or_1601_nl, fsm_output[0]);
  assign mux_1469_nl = MUX_s_1_2_2(mux_1468_nl, mux_1467_nl, fsm_output[4]);
  assign nor_1171_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1172_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1466_nl = MUX_s_1_2_2(nor_1171_nl, nor_1172_nl, fsm_output[0]);
  assign nand_59_nl = ~((fsm_output[4]) & mux_1466_nl);
  assign mux_1470_nl = MUX_s_1_2_2(mux_1469_nl, nand_59_nl, fsm_output[6]);
  assign or_1607_nl = (fsm_output[2]) | mux_1470_nl;
  assign mux_1480_nl = MUX_s_1_2_2(mux_1479_nl, or_1607_nl, fsm_output[5]);
  assign vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1480_nl) & (fsm_output[1]);
  assign nor_1162_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1163_nl = ~((COMP_LOOP_acc_13_psp_sva[3]) | (COMP_LOOP_acc_13_psp_sva[1])
      | not_tmp_414);
  assign mux_1492_nl = MUX_s_1_2_2(nor_1162_nl, nor_1163_nl, fsm_output[0]);
  assign nor_1164_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b010111) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1165_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1491_nl = MUX_s_1_2_2(nor_1164_nl, nor_1165_nl, fsm_output[0]);
  assign mux_1493_nl = MUX_s_1_2_2(mux_1492_nl, mux_1491_nl, fsm_output[4]);
  assign nor_1166_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1167_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1489_nl = MUX_s_1_2_2(nor_1166_nl, nor_1167_nl, fsm_output[0]);
  assign nor_1168_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1169_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1488_nl = MUX_s_1_2_2(nor_1168_nl, nor_1169_nl, fsm_output[0]);
  assign mux_1490_nl = MUX_s_1_2_2(mux_1489_nl, mux_1488_nl, fsm_output[4]);
  assign mux_1494_nl = MUX_s_1_2_2(mux_1493_nl, mux_1490_nl, fsm_output[6]);
  assign nand_446_nl = ~((fsm_output[2]) & mux_1494_nl);
  assign nand_326_nl = ~((COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b010111) & and_763_cse);
  assign mux_1485_nl = MUX_s_1_2_2(or_tmp_1513, nand_326_nl, fsm_output[0]);
  assign or_1624_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1484_nl = MUX_s_1_2_2(or_tmp_1509, or_1624_nl, fsm_output[0]);
  assign mux_1486_nl = MUX_s_1_2_2(mux_1485_nl, mux_1484_nl, fsm_output[4]);
  assign or_1621_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1482_nl = MUX_s_1_2_2(or_tmp_1507, or_1621_nl, fsm_output[0]);
  assign or_1618_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1481_nl = MUX_s_1_2_2(or_tmp_1503, or_1618_nl, fsm_output[0]);
  assign mux_1483_nl = MUX_s_1_2_2(mux_1482_nl, mux_1481_nl, fsm_output[4]);
  assign mux_1487_nl = MUX_s_1_2_2(mux_1486_nl, mux_1483_nl, fsm_output[6]);
  assign or_4119_nl = (fsm_output[2]) | mux_1487_nl;
  assign mux_1495_nl = MUX_s_1_2_2(nand_446_nl, or_4119_nl, fsm_output[5]);
  assign vec_rsc_0_23_i_we_d_pff = ~(mux_1495_nl | (fsm_output[1]));
  assign or_1660_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b010111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1659_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1508_nl = MUX_s_1_2_2(or_1660_nl, or_1659_nl, fsm_output[0]);
  assign or_1661_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1508_nl;
  assign nand_325_nl = ~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b010111)
      & and_763_cse);
  assign mux_1505_nl = MUX_s_1_2_2(nand_325_nl, or_tmp_1513, fsm_output[0]);
  assign or_1655_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b010111)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1504_nl = MUX_s_1_2_2(or_1655_nl, or_tmp_1509, fsm_output[0]);
  assign mux_1506_nl = MUX_s_1_2_2(mux_1505_nl, mux_1504_nl, fsm_output[4]);
  assign or_1654_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b010111)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1502_nl = MUX_s_1_2_2(or_1654_nl, or_tmp_1507, fsm_output[0]);
  assign or_1652_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b010111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1501_nl = MUX_s_1_2_2(or_1652_nl, or_tmp_1503, fsm_output[0]);
  assign mux_1503_nl = MUX_s_1_2_2(mux_1502_nl, mux_1501_nl, fsm_output[4]);
  assign mux_1507_nl = MUX_s_1_2_2(mux_1506_nl, mux_1503_nl, fsm_output[6]);
  assign mux_1509_nl = MUX_s_1_2_2(or_1661_nl, mux_1507_nl, fsm_output[2]);
  assign or_1650_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1648_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1498_nl = MUX_s_1_2_2(or_1650_nl, or_1648_nl, fsm_output[0]);
  assign or_1646_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1645_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b010111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1497_nl = MUX_s_1_2_2(or_1646_nl, or_1645_nl, fsm_output[0]);
  assign mux_1499_nl = MUX_s_1_2_2(mux_1498_nl, mux_1497_nl, fsm_output[4]);
  assign nor_1160_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1161_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b010111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1496_nl = MUX_s_1_2_2(nor_1160_nl, nor_1161_nl, fsm_output[0]);
  assign nand_61_nl = ~((fsm_output[4]) & mux_1496_nl);
  assign mux_1500_nl = MUX_s_1_2_2(mux_1499_nl, nand_61_nl, fsm_output[6]);
  assign or_1651_nl = (fsm_output[2]) | mux_1500_nl;
  assign mux_1510_nl = MUX_s_1_2_2(mux_1509_nl, or_1651_nl, fsm_output[5]);
  assign vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1510_nl) & (fsm_output[1]);
  assign nor_1151_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1152_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1522_nl = MUX_s_1_2_2(nor_1151_nl, nor_1152_nl, fsm_output[0]);
  assign nor_1153_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1154_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1521_nl = MUX_s_1_2_2(nor_1153_nl, nor_1154_nl, fsm_output[0]);
  assign mux_1523_nl = MUX_s_1_2_2(mux_1522_nl, mux_1521_nl, fsm_output[4]);
  assign nor_1155_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1156_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1519_nl = MUX_s_1_2_2(nor_1155_nl, nor_1156_nl, fsm_output[0]);
  assign nor_1157_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1158_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1518_nl = MUX_s_1_2_2(nor_1157_nl, nor_1158_nl, fsm_output[0]);
  assign mux_1520_nl = MUX_s_1_2_2(mux_1519_nl, mux_1518_nl, fsm_output[4]);
  assign mux_1524_nl = MUX_s_1_2_2(mux_1523_nl, mux_1520_nl, fsm_output[6]);
  assign nand_445_nl = ~((fsm_output[2]) & mux_1524_nl);
  assign or_1671_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011000) | (~ and_763_cse);
  assign mux_1515_nl = MUX_s_1_2_2(or_tmp_1557, or_1671_nl, fsm_output[0]);
  assign or_1668_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1514_nl = MUX_s_1_2_2(or_tmp_1553, or_1668_nl, fsm_output[0]);
  assign mux_1516_nl = MUX_s_1_2_2(mux_1515_nl, mux_1514_nl, fsm_output[4]);
  assign or_1665_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1512_nl = MUX_s_1_2_2(or_tmp_1551, or_1665_nl, fsm_output[0]);
  assign or_1662_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1511_nl = MUX_s_1_2_2(or_tmp_1547, or_1662_nl, fsm_output[0]);
  assign mux_1513_nl = MUX_s_1_2_2(mux_1512_nl, mux_1511_nl, fsm_output[4]);
  assign mux_1517_nl = MUX_s_1_2_2(mux_1516_nl, mux_1513_nl, fsm_output[6]);
  assign or_4118_nl = (fsm_output[2]) | mux_1517_nl;
  assign mux_1525_nl = MUX_s_1_2_2(nand_445_nl, or_4118_nl, fsm_output[5]);
  assign vec_rsc_0_24_i_we_d_pff = ~(mux_1525_nl | (fsm_output[1]));
  assign or_1704_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1703_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1538_nl = MUX_s_1_2_2(or_1704_nl, or_1703_nl, fsm_output[0]);
  assign or_1705_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1538_nl;
  assign or_1701_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011000)
      | (~ and_763_cse);
  assign mux_1535_nl = MUX_s_1_2_2(or_1701_nl, or_tmp_1557, fsm_output[0]);
  assign or_1699_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1534_nl = MUX_s_1_2_2(or_1699_nl, or_tmp_1553, fsm_output[0]);
  assign mux_1536_nl = MUX_s_1_2_2(mux_1535_nl, mux_1534_nl, fsm_output[4]);
  assign or_1698_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1532_nl = MUX_s_1_2_2(or_1698_nl, or_tmp_1551, fsm_output[0]);
  assign or_1696_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1531_nl = MUX_s_1_2_2(or_1696_nl, or_tmp_1547, fsm_output[0]);
  assign mux_1533_nl = MUX_s_1_2_2(mux_1532_nl, mux_1531_nl, fsm_output[4]);
  assign mux_1537_nl = MUX_s_1_2_2(mux_1536_nl, mux_1533_nl, fsm_output[6]);
  assign mux_1539_nl = MUX_s_1_2_2(or_1705_nl, mux_1537_nl, fsm_output[2]);
  assign or_1694_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1692_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1528_nl = MUX_s_1_2_2(or_1694_nl, or_1692_nl, fsm_output[0]);
  assign or_1690_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1689_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1527_nl = MUX_s_1_2_2(or_1690_nl, or_1689_nl, fsm_output[0]);
  assign mux_1529_nl = MUX_s_1_2_2(mux_1528_nl, mux_1527_nl, fsm_output[4]);
  assign nor_1149_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1150_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1526_nl = MUX_s_1_2_2(nor_1149_nl, nor_1150_nl, fsm_output[0]);
  assign nand_63_nl = ~((fsm_output[4]) & mux_1526_nl);
  assign mux_1530_nl = MUX_s_1_2_2(mux_1529_nl, nand_63_nl, fsm_output[6]);
  assign or_1695_nl = (fsm_output[2]) | mux_1530_nl;
  assign mux_1540_nl = MUX_s_1_2_2(mux_1539_nl, or_1695_nl, fsm_output[5]);
  assign vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1540_nl) & (fsm_output[1]);
  assign nor_1140_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1141_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1552_nl = MUX_s_1_2_2(nor_1140_nl, nor_1141_nl, fsm_output[0]);
  assign nor_1142_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1143_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1551_nl = MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output[0]);
  assign mux_1553_nl = MUX_s_1_2_2(mux_1552_nl, mux_1551_nl, fsm_output[4]);
  assign nor_1144_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1145_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1549_nl = MUX_s_1_2_2(nor_1144_nl, nor_1145_nl, fsm_output[0]);
  assign nor_1146_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1147_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1548_nl = MUX_s_1_2_2(nor_1146_nl, nor_1147_nl, fsm_output[0]);
  assign mux_1550_nl = MUX_s_1_2_2(mux_1549_nl, mux_1548_nl, fsm_output[4]);
  assign mux_1554_nl = MUX_s_1_2_2(mux_1553_nl, mux_1550_nl, fsm_output[6]);
  assign nand_444_nl = ~((fsm_output[2]) & mux_1554_nl);
  assign or_1715_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011001) | (~ and_763_cse);
  assign mux_1545_nl = MUX_s_1_2_2(or_tmp_1601, or_1715_nl, fsm_output[0]);
  assign or_1712_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1544_nl = MUX_s_1_2_2(or_tmp_1597, or_1712_nl, fsm_output[0]);
  assign mux_1546_nl = MUX_s_1_2_2(mux_1545_nl, mux_1544_nl, fsm_output[4]);
  assign or_1709_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1542_nl = MUX_s_1_2_2(or_tmp_1595, or_1709_nl, fsm_output[0]);
  assign or_1706_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1541_nl = MUX_s_1_2_2(or_tmp_1591, or_1706_nl, fsm_output[0]);
  assign mux_1543_nl = MUX_s_1_2_2(mux_1542_nl, mux_1541_nl, fsm_output[4]);
  assign mux_1547_nl = MUX_s_1_2_2(mux_1546_nl, mux_1543_nl, fsm_output[6]);
  assign or_4117_nl = (fsm_output[2]) | mux_1547_nl;
  assign mux_1555_nl = MUX_s_1_2_2(nand_444_nl, or_4117_nl, fsm_output[5]);
  assign vec_rsc_0_25_i_we_d_pff = ~(mux_1555_nl | (fsm_output[1]));
  assign or_1748_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1747_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1568_nl = MUX_s_1_2_2(or_1748_nl, or_1747_nl, fsm_output[0]);
  assign or_1749_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1568_nl;
  assign or_1745_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011001)
      | (~ and_763_cse);
  assign mux_1565_nl = MUX_s_1_2_2(or_1745_nl, or_tmp_1601, fsm_output[0]);
  assign or_1743_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1564_nl = MUX_s_1_2_2(or_1743_nl, or_tmp_1597, fsm_output[0]);
  assign mux_1566_nl = MUX_s_1_2_2(mux_1565_nl, mux_1564_nl, fsm_output[4]);
  assign or_1742_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1562_nl = MUX_s_1_2_2(or_1742_nl, or_tmp_1595, fsm_output[0]);
  assign or_1740_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1561_nl = MUX_s_1_2_2(or_1740_nl, or_tmp_1591, fsm_output[0]);
  assign mux_1563_nl = MUX_s_1_2_2(mux_1562_nl, mux_1561_nl, fsm_output[4]);
  assign mux_1567_nl = MUX_s_1_2_2(mux_1566_nl, mux_1563_nl, fsm_output[6]);
  assign mux_1569_nl = MUX_s_1_2_2(or_1749_nl, mux_1567_nl, fsm_output[2]);
  assign or_1738_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1736_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1558_nl = MUX_s_1_2_2(or_1738_nl, or_1736_nl, fsm_output[0]);
  assign or_1734_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1733_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1557_nl = MUX_s_1_2_2(or_1734_nl, or_1733_nl, fsm_output[0]);
  assign mux_1559_nl = MUX_s_1_2_2(mux_1558_nl, mux_1557_nl, fsm_output[4]);
  assign nor_1138_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1139_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1556_nl = MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output[0]);
  assign nand_65_nl = ~((fsm_output[4]) & mux_1556_nl);
  assign mux_1560_nl = MUX_s_1_2_2(mux_1559_nl, nand_65_nl, fsm_output[6]);
  assign or_1739_nl = (fsm_output[2]) | mux_1560_nl;
  assign mux_1570_nl = MUX_s_1_2_2(mux_1569_nl, or_1739_nl, fsm_output[5]);
  assign vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1570_nl) & (fsm_output[1]);
  assign nor_1129_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1130_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1582_nl = MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output[0]);
  assign nor_1131_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1132_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1581_nl = MUX_s_1_2_2(nor_1131_nl, nor_1132_nl, fsm_output[0]);
  assign mux_1583_nl = MUX_s_1_2_2(mux_1582_nl, mux_1581_nl, fsm_output[4]);
  assign nor_1133_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1134_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1579_nl = MUX_s_1_2_2(nor_1133_nl, nor_1134_nl, fsm_output[0]);
  assign nor_1135_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1136_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1578_nl = MUX_s_1_2_2(nor_1135_nl, nor_1136_nl, fsm_output[0]);
  assign mux_1580_nl = MUX_s_1_2_2(mux_1579_nl, mux_1578_nl, fsm_output[4]);
  assign mux_1584_nl = MUX_s_1_2_2(mux_1583_nl, mux_1580_nl, fsm_output[6]);
  assign nand_443_nl = ~((fsm_output[2]) & mux_1584_nl);
  assign or_1759_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011010) | (~ and_763_cse);
  assign mux_1575_nl = MUX_s_1_2_2(or_tmp_1645, or_1759_nl, fsm_output[0]);
  assign or_1756_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1574_nl = MUX_s_1_2_2(or_tmp_1641, or_1756_nl, fsm_output[0]);
  assign mux_1576_nl = MUX_s_1_2_2(mux_1575_nl, mux_1574_nl, fsm_output[4]);
  assign or_1753_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1572_nl = MUX_s_1_2_2(or_tmp_1639, or_1753_nl, fsm_output[0]);
  assign or_1750_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1571_nl = MUX_s_1_2_2(or_tmp_1635, or_1750_nl, fsm_output[0]);
  assign mux_1573_nl = MUX_s_1_2_2(mux_1572_nl, mux_1571_nl, fsm_output[4]);
  assign mux_1577_nl = MUX_s_1_2_2(mux_1576_nl, mux_1573_nl, fsm_output[6]);
  assign or_4116_nl = (fsm_output[2]) | mux_1577_nl;
  assign mux_1585_nl = MUX_s_1_2_2(nand_443_nl, or_4116_nl, fsm_output[5]);
  assign vec_rsc_0_26_i_we_d_pff = ~(mux_1585_nl | (fsm_output[1]));
  assign or_1792_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1791_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1598_nl = MUX_s_1_2_2(or_1792_nl, or_1791_nl, fsm_output[0]);
  assign or_1793_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1598_nl;
  assign or_1789_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011010)
      | (~ and_763_cse);
  assign mux_1595_nl = MUX_s_1_2_2(or_1789_nl, or_tmp_1645, fsm_output[0]);
  assign or_1787_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1594_nl = MUX_s_1_2_2(or_1787_nl, or_tmp_1641, fsm_output[0]);
  assign mux_1596_nl = MUX_s_1_2_2(mux_1595_nl, mux_1594_nl, fsm_output[4]);
  assign or_1786_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1592_nl = MUX_s_1_2_2(or_1786_nl, or_tmp_1639, fsm_output[0]);
  assign or_1784_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1591_nl = MUX_s_1_2_2(or_1784_nl, or_tmp_1635, fsm_output[0]);
  assign mux_1593_nl = MUX_s_1_2_2(mux_1592_nl, mux_1591_nl, fsm_output[4]);
  assign mux_1597_nl = MUX_s_1_2_2(mux_1596_nl, mux_1593_nl, fsm_output[6]);
  assign mux_1599_nl = MUX_s_1_2_2(or_1793_nl, mux_1597_nl, fsm_output[2]);
  assign or_1782_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1780_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1588_nl = MUX_s_1_2_2(or_1782_nl, or_1780_nl, fsm_output[0]);
  assign or_1778_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1777_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1587_nl = MUX_s_1_2_2(or_1778_nl, or_1777_nl, fsm_output[0]);
  assign mux_1589_nl = MUX_s_1_2_2(mux_1588_nl, mux_1587_nl, fsm_output[4]);
  assign nor_1127_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1128_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1586_nl = MUX_s_1_2_2(nor_1127_nl, nor_1128_nl, fsm_output[0]);
  assign nand_67_nl = ~((fsm_output[4]) & mux_1586_nl);
  assign mux_1590_nl = MUX_s_1_2_2(mux_1589_nl, nand_67_nl, fsm_output[6]);
  assign or_1783_nl = (fsm_output[2]) | mux_1590_nl;
  assign mux_1600_nl = MUX_s_1_2_2(mux_1599_nl, or_1783_nl, fsm_output[5]);
  assign vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1600_nl) & (fsm_output[1]);
  assign nor_1118_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1119_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | not_tmp_330);
  assign mux_1612_nl = MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, fsm_output[0]);
  assign nor_1120_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1121_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1611_nl = MUX_s_1_2_2(nor_1120_nl, nor_1121_nl, fsm_output[0]);
  assign mux_1613_nl = MUX_s_1_2_2(mux_1612_nl, mux_1611_nl, fsm_output[4]);
  assign nor_1122_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1123_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1609_nl = MUX_s_1_2_2(nor_1122_nl, nor_1123_nl, fsm_output[0]);
  assign nor_1124_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1125_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1608_nl = MUX_s_1_2_2(nor_1124_nl, nor_1125_nl, fsm_output[0]);
  assign mux_1610_nl = MUX_s_1_2_2(mux_1609_nl, mux_1608_nl, fsm_output[4]);
  assign mux_1614_nl = MUX_s_1_2_2(mux_1613_nl, mux_1610_nl, fsm_output[6]);
  assign nand_442_nl = ~((fsm_output[2]) & mux_1614_nl);
  assign nand_324_nl = ~((COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011011) & and_763_cse);
  assign mux_1605_nl = MUX_s_1_2_2(or_tmp_1689, nand_324_nl, fsm_output[0]);
  assign or_1800_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1604_nl = MUX_s_1_2_2(or_tmp_1685, or_1800_nl, fsm_output[0]);
  assign mux_1606_nl = MUX_s_1_2_2(mux_1605_nl, mux_1604_nl, fsm_output[4]);
  assign or_1797_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1602_nl = MUX_s_1_2_2(or_tmp_1683, or_1797_nl, fsm_output[0]);
  assign or_1794_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1601_nl = MUX_s_1_2_2(or_tmp_1679, or_1794_nl, fsm_output[0]);
  assign mux_1603_nl = MUX_s_1_2_2(mux_1602_nl, mux_1601_nl, fsm_output[4]);
  assign mux_1607_nl = MUX_s_1_2_2(mux_1606_nl, mux_1603_nl, fsm_output[6]);
  assign or_4115_nl = (fsm_output[2]) | mux_1607_nl;
  assign mux_1615_nl = MUX_s_1_2_2(nand_442_nl, or_4115_nl, fsm_output[5]);
  assign vec_rsc_0_27_i_we_d_pff = ~(mux_1615_nl | (fsm_output[1]));
  assign or_1836_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1835_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1628_nl = MUX_s_1_2_2(or_1836_nl, or_1835_nl, fsm_output[0]);
  assign or_1837_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1628_nl;
  assign nand_323_nl = ~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011011)
      & and_763_cse);
  assign mux_1625_nl = MUX_s_1_2_2(nand_323_nl, or_tmp_1689, fsm_output[0]);
  assign or_1831_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1624_nl = MUX_s_1_2_2(or_1831_nl, or_tmp_1685, fsm_output[0]);
  assign mux_1626_nl = MUX_s_1_2_2(mux_1625_nl, mux_1624_nl, fsm_output[4]);
  assign or_1830_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1622_nl = MUX_s_1_2_2(or_1830_nl, or_tmp_1683, fsm_output[0]);
  assign or_1828_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1621_nl = MUX_s_1_2_2(or_1828_nl, or_tmp_1679, fsm_output[0]);
  assign mux_1623_nl = MUX_s_1_2_2(mux_1622_nl, mux_1621_nl, fsm_output[4]);
  assign mux_1627_nl = MUX_s_1_2_2(mux_1626_nl, mux_1623_nl, fsm_output[6]);
  assign mux_1629_nl = MUX_s_1_2_2(or_1837_nl, mux_1627_nl, fsm_output[2]);
  assign or_1826_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1824_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1618_nl = MUX_s_1_2_2(or_1826_nl, or_1824_nl, fsm_output[0]);
  assign or_1822_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1821_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1617_nl = MUX_s_1_2_2(or_1822_nl, or_1821_nl, fsm_output[0]);
  assign mux_1619_nl = MUX_s_1_2_2(mux_1618_nl, mux_1617_nl, fsm_output[4]);
  assign nor_1116_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1117_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1616_nl = MUX_s_1_2_2(nor_1116_nl, nor_1117_nl, fsm_output[0]);
  assign nand_69_nl = ~((fsm_output[4]) & mux_1616_nl);
  assign mux_1620_nl = MUX_s_1_2_2(mux_1619_nl, nand_69_nl, fsm_output[6]);
  assign or_1827_nl = (fsm_output[2]) | mux_1620_nl;
  assign mux_1630_nl = MUX_s_1_2_2(mux_1629_nl, or_1827_nl, fsm_output[5]);
  assign vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1630_nl) & (fsm_output[1]);
  assign nor_1107_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1108_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0111) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1642_nl = MUX_s_1_2_2(nor_1107_nl, nor_1108_nl, fsm_output[0]);
  assign nor_1109_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1110_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1641_nl = MUX_s_1_2_2(nor_1109_nl, nor_1110_nl, fsm_output[0]);
  assign mux_1643_nl = MUX_s_1_2_2(mux_1642_nl, mux_1641_nl, fsm_output[4]);
  assign nor_1111_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1112_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1639_nl = MUX_s_1_2_2(nor_1111_nl, nor_1112_nl, fsm_output[0]);
  assign nor_1113_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1114_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1638_nl = MUX_s_1_2_2(nor_1113_nl, nor_1114_nl, fsm_output[0]);
  assign mux_1640_nl = MUX_s_1_2_2(mux_1639_nl, mux_1638_nl, fsm_output[4]);
  assign mux_1644_nl = MUX_s_1_2_2(mux_1643_nl, mux_1640_nl, fsm_output[6]);
  assign nand_441_nl = ~((fsm_output[2]) & mux_1644_nl);
  assign or_1847_nl = (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011100) | (~ and_763_cse);
  assign mux_1635_nl = MUX_s_1_2_2(or_tmp_1733, or_1847_nl, fsm_output[0]);
  assign or_1844_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1634_nl = MUX_s_1_2_2(or_tmp_1729, or_1844_nl, fsm_output[0]);
  assign mux_1636_nl = MUX_s_1_2_2(mux_1635_nl, mux_1634_nl, fsm_output[4]);
  assign or_1841_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1632_nl = MUX_s_1_2_2(or_tmp_1727, or_1841_nl, fsm_output[0]);
  assign or_1838_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1631_nl = MUX_s_1_2_2(or_tmp_1723, or_1838_nl, fsm_output[0]);
  assign mux_1633_nl = MUX_s_1_2_2(mux_1632_nl, mux_1631_nl, fsm_output[4]);
  assign mux_1637_nl = MUX_s_1_2_2(mux_1636_nl, mux_1633_nl, fsm_output[6]);
  assign or_4114_nl = (fsm_output[2]) | mux_1637_nl;
  assign mux_1645_nl = MUX_s_1_2_2(nand_441_nl, or_4114_nl, fsm_output[5]);
  assign vec_rsc_0_28_i_we_d_pff = ~(mux_1645_nl | (fsm_output[1]));
  assign or_1880_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1879_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1658_nl = MUX_s_1_2_2(or_1880_nl, or_1879_nl, fsm_output[0]);
  assign or_1881_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1658_nl;
  assign or_1877_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[5:0]!=6'b011100)
      | (~ and_763_cse);
  assign mux_1655_nl = MUX_s_1_2_2(or_1877_nl, or_tmp_1733, fsm_output[0]);
  assign or_1875_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1654_nl = MUX_s_1_2_2(or_1875_nl, or_tmp_1729, fsm_output[0]);
  assign mux_1656_nl = MUX_s_1_2_2(mux_1655_nl, mux_1654_nl, fsm_output[4]);
  assign or_1874_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1652_nl = MUX_s_1_2_2(or_1874_nl, or_tmp_1727, fsm_output[0]);
  assign or_1872_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1651_nl = MUX_s_1_2_2(or_1872_nl, or_tmp_1723, fsm_output[0]);
  assign mux_1653_nl = MUX_s_1_2_2(mux_1652_nl, mux_1651_nl, fsm_output[4]);
  assign mux_1657_nl = MUX_s_1_2_2(mux_1656_nl, mux_1653_nl, fsm_output[6]);
  assign mux_1659_nl = MUX_s_1_2_2(or_1881_nl, mux_1657_nl, fsm_output[2]);
  assign or_1870_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_1868_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1648_nl = MUX_s_1_2_2(or_1870_nl, or_1868_nl, fsm_output[0]);
  assign or_1866_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1865_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1647_nl = MUX_s_1_2_2(or_1866_nl, or_1865_nl, fsm_output[0]);
  assign mux_1649_nl = MUX_s_1_2_2(mux_1648_nl, mux_1647_nl, fsm_output[4]);
  assign nor_1105_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1106_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1646_nl = MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, fsm_output[0]);
  assign nand_71_nl = ~((fsm_output[4]) & mux_1646_nl);
  assign mux_1650_nl = MUX_s_1_2_2(mux_1649_nl, nand_71_nl, fsm_output[6]);
  assign or_1871_nl = (fsm_output[2]) | mux_1650_nl;
  assign mux_1660_nl = MUX_s_1_2_2(mux_1659_nl, or_1871_nl, fsm_output[5]);
  assign vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1660_nl) & (fsm_output[1]);
  assign nor_1096_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign nor_1097_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0111) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1672_nl = MUX_s_1_2_2(nor_1096_nl, nor_1097_nl, fsm_output[0]);
  assign nor_1098_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1099_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1671_nl = MUX_s_1_2_2(nor_1098_nl, nor_1099_nl, fsm_output[0]);
  assign mux_1673_nl = MUX_s_1_2_2(mux_1672_nl, mux_1671_nl, fsm_output[4]);
  assign nor_1100_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1101_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1669_nl = MUX_s_1_2_2(nor_1100_nl, nor_1101_nl, fsm_output[0]);
  assign nor_1102_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1103_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1668_nl = MUX_s_1_2_2(nor_1102_nl, nor_1103_nl, fsm_output[0]);
  assign mux_1670_nl = MUX_s_1_2_2(mux_1669_nl, mux_1668_nl, fsm_output[4]);
  assign mux_1674_nl = MUX_s_1_2_2(mux_1673_nl, mux_1670_nl, fsm_output[6]);
  assign nand_440_nl = ~((fsm_output[2]) & mux_1674_nl);
  assign nand_322_nl = ~((COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011101) & and_763_cse);
  assign mux_1665_nl = MUX_s_1_2_2(or_tmp_1777, nand_322_nl, fsm_output[0]);
  assign or_1888_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1664_nl = MUX_s_1_2_2(or_tmp_1773, or_1888_nl, fsm_output[0]);
  assign mux_1666_nl = MUX_s_1_2_2(mux_1665_nl, mux_1664_nl, fsm_output[4]);
  assign or_1885_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1662_nl = MUX_s_1_2_2(or_tmp_1771, or_1885_nl, fsm_output[0]);
  assign or_1882_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1661_nl = MUX_s_1_2_2(or_tmp_1767, or_1882_nl, fsm_output[0]);
  assign mux_1663_nl = MUX_s_1_2_2(mux_1662_nl, mux_1661_nl, fsm_output[4]);
  assign mux_1667_nl = MUX_s_1_2_2(mux_1666_nl, mux_1663_nl, fsm_output[6]);
  assign or_4113_nl = (fsm_output[2]) | mux_1667_nl;
  assign mux_1675_nl = MUX_s_1_2_2(nand_440_nl, or_4113_nl, fsm_output[5]);
  assign vec_rsc_0_29_i_we_d_pff = ~(mux_1675_nl | (fsm_output[1]));
  assign or_1924_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1923_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1688_nl = MUX_s_1_2_2(or_1924_nl, or_1923_nl, fsm_output[0]);
  assign or_1925_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1688_nl;
  assign nand_321_nl = ~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011101)
      & and_763_cse);
  assign mux_1685_nl = MUX_s_1_2_2(nand_321_nl, or_tmp_1777, fsm_output[0]);
  assign or_1919_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1684_nl = MUX_s_1_2_2(or_1919_nl, or_tmp_1773, fsm_output[0]);
  assign mux_1686_nl = MUX_s_1_2_2(mux_1685_nl, mux_1684_nl, fsm_output[4]);
  assign or_1918_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1682_nl = MUX_s_1_2_2(or_1918_nl, or_tmp_1771, fsm_output[0]);
  assign or_1916_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1681_nl = MUX_s_1_2_2(or_1916_nl, or_tmp_1767, fsm_output[0]);
  assign mux_1683_nl = MUX_s_1_2_2(mux_1682_nl, mux_1681_nl, fsm_output[4]);
  assign mux_1687_nl = MUX_s_1_2_2(mux_1686_nl, mux_1683_nl, fsm_output[6]);
  assign mux_1689_nl = MUX_s_1_2_2(or_1925_nl, mux_1687_nl, fsm_output[2]);
  assign or_1914_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_1912_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[0])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1678_nl = MUX_s_1_2_2(or_1914_nl, or_1912_nl, fsm_output[0]);
  assign or_1910_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1909_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1677_nl = MUX_s_1_2_2(or_1910_nl, or_1909_nl, fsm_output[0]);
  assign mux_1679_nl = MUX_s_1_2_2(mux_1678_nl, mux_1677_nl, fsm_output[4]);
  assign nor_1094_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1095_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1676_nl = MUX_s_1_2_2(nor_1094_nl, nor_1095_nl, fsm_output[0]);
  assign nand_73_nl = ~((fsm_output[4]) & mux_1676_nl);
  assign mux_1680_nl = MUX_s_1_2_2(mux_1679_nl, nand_73_nl, fsm_output[6]);
  assign or_1915_nl = (fsm_output[2]) | mux_1680_nl;
  assign mux_1690_nl = MUX_s_1_2_2(mux_1689_nl, or_1915_nl, fsm_output[5]);
  assign vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1690_nl) & (fsm_output[1]);
  assign nor_1086_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[2]))
      | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) | not_tmp_384);
  assign and_602_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b0111) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b10)
      & and_763_cse;
  assign mux_1702_nl = MUX_s_1_2_2(nor_1086_nl, and_602_nl, fsm_output[0]);
  assign nor_1087_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b011110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1088_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1701_nl = MUX_s_1_2_2(nor_1087_nl, nor_1088_nl, fsm_output[0]);
  assign mux_1703_nl = MUX_s_1_2_2(mux_1702_nl, mux_1701_nl, fsm_output[4]);
  assign nor_1089_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1090_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b01111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1699_nl = MUX_s_1_2_2(nor_1089_nl, nor_1090_nl, fsm_output[0]);
  assign nor_1091_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1092_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1698_nl = MUX_s_1_2_2(nor_1091_nl, nor_1092_nl, fsm_output[0]);
  assign mux_1700_nl = MUX_s_1_2_2(mux_1699_nl, mux_1698_nl, fsm_output[4]);
  assign mux_1704_nl = MUX_s_1_2_2(mux_1703_nl, mux_1700_nl, fsm_output[6]);
  assign nand_439_nl = ~((fsm_output[2]) & mux_1704_nl);
  assign nand_320_nl = ~((COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011110) & and_763_cse);
  assign mux_1695_nl = MUX_s_1_2_2(or_tmp_1821, nand_320_nl, fsm_output[0]);
  assign or_1932_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1694_nl = MUX_s_1_2_2(or_tmp_1817, or_1932_nl, fsm_output[0]);
  assign mux_1696_nl = MUX_s_1_2_2(mux_1695_nl, mux_1694_nl, fsm_output[4]);
  assign or_1929_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1692_nl = MUX_s_1_2_2(or_tmp_1815, or_1929_nl, fsm_output[0]);
  assign or_1926_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1691_nl = MUX_s_1_2_2(or_tmp_1811, or_1926_nl, fsm_output[0]);
  assign mux_1693_nl = MUX_s_1_2_2(mux_1692_nl, mux_1691_nl, fsm_output[4]);
  assign mux_1697_nl = MUX_s_1_2_2(mux_1696_nl, mux_1693_nl, fsm_output[6]);
  assign or_4112_nl = (fsm_output[2]) | mux_1697_nl;
  assign mux_1705_nl = MUX_s_1_2_2(nand_439_nl, or_4112_nl, fsm_output[5]);
  assign vec_rsc_0_30_i_we_d_pff = ~(mux_1705_nl | (fsm_output[1]));
  assign or_1968_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_1967_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1718_nl = MUX_s_1_2_2(or_1968_nl, or_1967_nl, fsm_output[0]);
  assign or_1969_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1718_nl;
  assign nand_318_nl = ~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011110)
      & and_763_cse);
  assign mux_1715_nl = MUX_s_1_2_2(nand_318_nl, or_tmp_1821, fsm_output[0]);
  assign or_1963_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b011110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1714_nl = MUX_s_1_2_2(or_1963_nl, or_tmp_1817, fsm_output[0]);
  assign mux_1716_nl = MUX_s_1_2_2(mux_1715_nl, mux_1714_nl, fsm_output[4]);
  assign or_1962_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b011110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1712_nl = MUX_s_1_2_2(or_1962_nl, or_tmp_1815, fsm_output[0]);
  assign or_1960_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1711_nl = MUX_s_1_2_2(or_1960_nl, or_tmp_1811, fsm_output[0]);
  assign mux_1713_nl = MUX_s_1_2_2(mux_1712_nl, mux_1711_nl, fsm_output[4]);
  assign mux_1717_nl = MUX_s_1_2_2(mux_1716_nl, mux_1713_nl, fsm_output[6]);
  assign mux_1719_nl = MUX_s_1_2_2(or_1969_nl, mux_1717_nl, fsm_output[2]);
  assign nand_319_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b01111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & and_763_cse);
  assign or_1956_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[2]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) | not_tmp_388;
  assign mux_1708_nl = MUX_s_1_2_2(nand_319_nl, or_1956_nl, fsm_output[0]);
  assign or_1954_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01111) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_1953_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1707_nl = MUX_s_1_2_2(or_1954_nl, or_1953_nl, fsm_output[0]);
  assign mux_1709_nl = MUX_s_1_2_2(mux_1708_nl, mux_1707_nl, fsm_output[4]);
  assign nor_1084_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1085_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1706_nl = MUX_s_1_2_2(nor_1084_nl, nor_1085_nl, fsm_output[0]);
  assign nand_75_nl = ~((fsm_output[4]) & mux_1706_nl);
  assign mux_1710_nl = MUX_s_1_2_2(mux_1709_nl, nand_75_nl, fsm_output[6]);
  assign or_1959_nl = (fsm_output[2]) | mux_1710_nl;
  assign mux_1720_nl = MUX_s_1_2_2(mux_1719_nl, or_1959_nl, fsm_output[5]);
  assign vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1720_nl) & (fsm_output[1]);
  assign nor_1077_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      & (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & (COMP_LOOP_acc_10_cse_10_1_5_sva[3])
      & (~ (COMP_LOOP_acc_10_cse_10_1_5_sva[5])))) | not_tmp_384);
  assign nor_1078_nl = ~((COMP_LOOP_acc_13_psp_sva[3]) | (~((COMP_LOOP_acc_13_psp_sva[2:0]==3'b111)
      & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (fsm_output[3]) & (fsm_output[7]))));
  assign mux_1732_nl = MUX_s_1_2_2(nor_1077_nl, nor_1078_nl, fsm_output[0]);
  assign and_599_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b011111) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_600_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b011) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_1731_nl = MUX_s_1_2_2(and_599_nl, and_600_nl, fsm_output[0]);
  assign mux_1733_nl = MUX_s_1_2_2(mux_1732_nl, mux_1731_nl, fsm_output[4]);
  assign and_811_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b011111) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_818_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b01111) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_1729_nl = MUX_s_1_2_2(and_811_nl, and_818_nl, fsm_output[0]);
  assign nor_1081_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b011111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1082_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b01111) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1728_nl = MUX_s_1_2_2(nor_1081_nl, nor_1082_nl, fsm_output[0]);
  assign mux_1730_nl = MUX_s_1_2_2(mux_1729_nl, mux_1728_nl, fsm_output[4]);
  assign mux_1734_nl = MUX_s_1_2_2(mux_1733_nl, mux_1730_nl, fsm_output[6]);
  assign nand_438_nl = ~((fsm_output[2]) & mux_1734_nl);
  assign nand_313_nl = ~((COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011111) & and_763_cse);
  assign mux_1725_nl = MUX_s_1_2_2(or_tmp_1865, nand_313_nl, fsm_output[0]);
  assign nand_314_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b011111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_1724_nl = MUX_s_1_2_2(or_tmp_1861, nand_314_nl, fsm_output[0]);
  assign mux_1726_nl = MUX_s_1_2_2(mux_1725_nl, mux_1724_nl, fsm_output[4]);
  assign nand_478_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b011111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_1722_nl = MUX_s_1_2_2(or_tmp_1859, nand_478_nl, fsm_output[0]);
  assign or_1970_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1721_nl = MUX_s_1_2_2(or_tmp_1855, or_1970_nl, fsm_output[0]);
  assign mux_1723_nl = MUX_s_1_2_2(mux_1722_nl, mux_1721_nl, fsm_output[4]);
  assign mux_1727_nl = MUX_s_1_2_2(mux_1726_nl, mux_1723_nl, fsm_output[6]);
  assign or_4111_nl = (fsm_output[2]) | mux_1727_nl;
  assign mux_1735_nl = MUX_s_1_2_2(nand_438_nl, or_4111_nl, fsm_output[5]);
  assign vec_rsc_0_31_i_we_d_pff = ~(mux_1735_nl | (fsm_output[1]));
  assign or_2011_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b011111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2010_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1748_nl = MUX_s_1_2_2(or_2011_nl, or_2010_nl, fsm_output[0]);
  assign or_2012_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1748_nl;
  assign nand_302_nl = ~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[5:0]==6'b011111)
      & and_763_cse);
  assign mux_1745_nl = MUX_s_1_2_2(nand_302_nl, or_tmp_1865, fsm_output[0]);
  assign nand_303_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b011111)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_1744_nl = MUX_s_1_2_2(nand_303_nl, or_tmp_1861, fsm_output[0]);
  assign mux_1746_nl = MUX_s_1_2_2(mux_1745_nl, mux_1744_nl, fsm_output[4]);
  assign nand_404_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b011111)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_1742_nl = MUX_s_1_2_2(nand_404_nl, or_tmp_1859, fsm_output[0]);
  assign or_2003_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b011111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1741_nl = MUX_s_1_2_2(or_2003_nl, or_tmp_1855, fsm_output[0]);
  assign mux_1743_nl = MUX_s_1_2_2(mux_1742_nl, mux_1741_nl, fsm_output[4]);
  assign mux_1747_nl = MUX_s_1_2_2(mux_1746_nl, mux_1743_nl, fsm_output[6]);
  assign mux_1749_nl = MUX_s_1_2_2(or_2012_nl, mux_1747_nl, fsm_output[2]);
  assign or_2001_nl = (~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b01111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm))
      | not_tmp_321;
  assign or_1999_nl = (~((COMP_LOOP_acc_10_cse_10_1_7_sva[1]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      & (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      & (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[5])))) | not_tmp_388;
  assign mux_1738_nl = MUX_s_1_2_2(or_2001_nl, or_1999_nl, fsm_output[0]);
  assign nand_307_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b01111) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_308_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b011111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_1737_nl = MUX_s_1_2_2(nand_307_nl, nand_308_nl, fsm_output[0]);
  assign mux_1739_nl = MUX_s_1_2_2(mux_1738_nl, mux_1737_nl, fsm_output[4]);
  assign nor_1075_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b0111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1076_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b011111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1736_nl = MUX_s_1_2_2(nor_1075_nl, nor_1076_nl, fsm_output[0]);
  assign nand_77_nl = ~((fsm_output[4]) & mux_1736_nl);
  assign mux_1740_nl = MUX_s_1_2_2(mux_1739_nl, nand_77_nl, fsm_output[6]);
  assign or_2002_nl = (fsm_output[2]) | mux_1740_nl;
  assign mux_1750_nl = MUX_s_1_2_2(mux_1749_nl, or_2002_nl, fsm_output[5]);
  assign vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1750_nl) & (fsm_output[1]);
  assign nor_1066_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100000) | (~ and_763_cse));
  assign nor_1067_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1762_nl = MUX_s_1_2_2(nor_1066_nl, nor_1067_nl, fsm_output[0]);
  assign nor_1068_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1069_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1761_nl = MUX_s_1_2_2(nor_1068_nl, nor_1069_nl, fsm_output[0]);
  assign mux_1763_nl = MUX_s_1_2_2(mux_1762_nl, mux_1761_nl, fsm_output[4]);
  assign nor_1070_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1071_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1759_nl = MUX_s_1_2_2(nor_1070_nl, nor_1071_nl, fsm_output[0]);
  assign nor_1072_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1073_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1758_nl = MUX_s_1_2_2(nor_1072_nl, nor_1073_nl, fsm_output[0]);
  assign mux_1760_nl = MUX_s_1_2_2(mux_1759_nl, mux_1758_nl, fsm_output[4]);
  assign mux_1764_nl = MUX_s_1_2_2(mux_1763_nl, mux_1760_nl, fsm_output[6]);
  assign nand_437_nl = ~((fsm_output[2]) & mux_1764_nl);
  assign or_2022_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00000) | not_tmp_452;
  assign mux_1755_nl = MUX_s_1_2_2(or_tmp_1908, or_2022_nl, fsm_output[0]);
  assign or_2019_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1754_nl = MUX_s_1_2_2(or_tmp_1904, or_2019_nl, fsm_output[0]);
  assign mux_1756_nl = MUX_s_1_2_2(mux_1755_nl, mux_1754_nl, fsm_output[4]);
  assign or_2016_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1752_nl = MUX_s_1_2_2(or_tmp_1902, or_2016_nl, fsm_output[0]);
  assign or_2013_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1751_nl = MUX_s_1_2_2(or_tmp_1898, or_2013_nl, fsm_output[0]);
  assign mux_1753_nl = MUX_s_1_2_2(mux_1752_nl, mux_1751_nl, fsm_output[4]);
  assign mux_1757_nl = MUX_s_1_2_2(mux_1756_nl, mux_1753_nl, fsm_output[6]);
  assign or_4110_nl = (fsm_output[2]) | mux_1757_nl;
  assign mux_1765_nl = MUX_s_1_2_2(nand_437_nl, or_4110_nl, fsm_output[5]);
  assign vec_rsc_0_32_i_we_d_pff = ~(mux_1765_nl | (fsm_output[1]));
  assign or_2055_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2054_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1778_nl = MUX_s_1_2_2(or_2055_nl, or_2054_nl, fsm_output[0]);
  assign or_2056_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1778_nl;
  assign or_2052_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00000)
      | not_tmp_452;
  assign mux_1775_nl = MUX_s_1_2_2(or_2052_nl, or_tmp_1908, fsm_output[0]);
  assign or_2050_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1774_nl = MUX_s_1_2_2(or_2050_nl, or_tmp_1904, fsm_output[0]);
  assign mux_1776_nl = MUX_s_1_2_2(mux_1775_nl, mux_1774_nl, fsm_output[4]);
  assign or_2049_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1772_nl = MUX_s_1_2_2(or_2049_nl, or_tmp_1902, fsm_output[0]);
  assign or_2047_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1771_nl = MUX_s_1_2_2(or_2047_nl, or_tmp_1898, fsm_output[0]);
  assign mux_1773_nl = MUX_s_1_2_2(mux_1772_nl, mux_1771_nl, fsm_output[4]);
  assign mux_1777_nl = MUX_s_1_2_2(mux_1776_nl, mux_1773_nl, fsm_output[6]);
  assign mux_1779_nl = MUX_s_1_2_2(or_2056_nl, mux_1777_nl, fsm_output[2]);
  assign or_2045_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2043_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100000) | (~ and_763_cse);
  assign mux_1768_nl = MUX_s_1_2_2(or_2045_nl, or_2043_nl, fsm_output[0]);
  assign or_2041_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2040_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1767_nl = MUX_s_1_2_2(or_2041_nl, or_2040_nl, fsm_output[0]);
  assign mux_1769_nl = MUX_s_1_2_2(mux_1768_nl, mux_1767_nl, fsm_output[4]);
  assign nor_1064_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1065_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1766_nl = MUX_s_1_2_2(nor_1064_nl, nor_1065_nl, fsm_output[0]);
  assign nand_79_nl = ~((fsm_output[4]) & mux_1766_nl);
  assign mux_1770_nl = MUX_s_1_2_2(mux_1769_nl, nand_79_nl, fsm_output[6]);
  assign or_2046_nl = (fsm_output[2]) | mux_1770_nl;
  assign mux_1780_nl = MUX_s_1_2_2(mux_1779_nl, or_2046_nl, fsm_output[5]);
  assign vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1780_nl) & (fsm_output[1]);
  assign nor_1055_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100001) | (~ and_763_cse));
  assign nor_1056_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1792_nl = MUX_s_1_2_2(nor_1055_nl, nor_1056_nl, fsm_output[0]);
  assign nor_1057_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1058_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1791_nl = MUX_s_1_2_2(nor_1057_nl, nor_1058_nl, fsm_output[0]);
  assign mux_1793_nl = MUX_s_1_2_2(mux_1792_nl, mux_1791_nl, fsm_output[4]);
  assign nor_1059_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1060_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1789_nl = MUX_s_1_2_2(nor_1059_nl, nor_1060_nl, fsm_output[0]);
  assign nor_1061_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1062_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1788_nl = MUX_s_1_2_2(nor_1061_nl, nor_1062_nl, fsm_output[0]);
  assign mux_1790_nl = MUX_s_1_2_2(mux_1789_nl, mux_1788_nl, fsm_output[4]);
  assign mux_1794_nl = MUX_s_1_2_2(mux_1793_nl, mux_1790_nl, fsm_output[6]);
  assign nand_436_nl = ~((fsm_output[2]) & mux_1794_nl);
  assign or_2066_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00001) | not_tmp_452;
  assign mux_1785_nl = MUX_s_1_2_2(or_tmp_1952, or_2066_nl, fsm_output[0]);
  assign or_2063_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1784_nl = MUX_s_1_2_2(or_tmp_1948, or_2063_nl, fsm_output[0]);
  assign mux_1786_nl = MUX_s_1_2_2(mux_1785_nl, mux_1784_nl, fsm_output[4]);
  assign or_2060_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1782_nl = MUX_s_1_2_2(or_tmp_1946, or_2060_nl, fsm_output[0]);
  assign or_2057_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1781_nl = MUX_s_1_2_2(or_tmp_1942, or_2057_nl, fsm_output[0]);
  assign mux_1783_nl = MUX_s_1_2_2(mux_1782_nl, mux_1781_nl, fsm_output[4]);
  assign mux_1787_nl = MUX_s_1_2_2(mux_1786_nl, mux_1783_nl, fsm_output[6]);
  assign or_4109_nl = (fsm_output[2]) | mux_1787_nl;
  assign mux_1795_nl = MUX_s_1_2_2(nand_436_nl, or_4109_nl, fsm_output[5]);
  assign vec_rsc_0_33_i_we_d_pff = ~(mux_1795_nl | (fsm_output[1]));
  assign or_2099_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2098_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1808_nl = MUX_s_1_2_2(or_2099_nl, or_2098_nl, fsm_output[0]);
  assign or_2100_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1808_nl;
  assign or_2096_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00001)
      | not_tmp_452;
  assign mux_1805_nl = MUX_s_1_2_2(or_2096_nl, or_tmp_1952, fsm_output[0]);
  assign or_2094_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1804_nl = MUX_s_1_2_2(or_2094_nl, or_tmp_1948, fsm_output[0]);
  assign mux_1806_nl = MUX_s_1_2_2(mux_1805_nl, mux_1804_nl, fsm_output[4]);
  assign or_2093_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1802_nl = MUX_s_1_2_2(or_2093_nl, or_tmp_1946, fsm_output[0]);
  assign or_2091_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1801_nl = MUX_s_1_2_2(or_2091_nl, or_tmp_1942, fsm_output[0]);
  assign mux_1803_nl = MUX_s_1_2_2(mux_1802_nl, mux_1801_nl, fsm_output[4]);
  assign mux_1807_nl = MUX_s_1_2_2(mux_1806_nl, mux_1803_nl, fsm_output[6]);
  assign mux_1809_nl = MUX_s_1_2_2(or_2100_nl, mux_1807_nl, fsm_output[2]);
  assign or_2089_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2087_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100001) | (~ and_763_cse);
  assign mux_1798_nl = MUX_s_1_2_2(or_2089_nl, or_2087_nl, fsm_output[0]);
  assign or_2085_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2084_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1797_nl = MUX_s_1_2_2(or_2085_nl, or_2084_nl, fsm_output[0]);
  assign mux_1799_nl = MUX_s_1_2_2(mux_1798_nl, mux_1797_nl, fsm_output[4]);
  assign nor_1053_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1054_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1796_nl = MUX_s_1_2_2(nor_1053_nl, nor_1054_nl, fsm_output[0]);
  assign nand_81_nl = ~((fsm_output[4]) & mux_1796_nl);
  assign mux_1800_nl = MUX_s_1_2_2(mux_1799_nl, nand_81_nl, fsm_output[6]);
  assign or_2090_nl = (fsm_output[2]) | mux_1800_nl;
  assign mux_1810_nl = MUX_s_1_2_2(mux_1809_nl, or_2090_nl, fsm_output[5]);
  assign vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1810_nl) & (fsm_output[1]);
  assign nor_1044_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100010) | (~ and_763_cse));
  assign nor_1045_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1822_nl = MUX_s_1_2_2(nor_1044_nl, nor_1045_nl, fsm_output[0]);
  assign nor_1046_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1047_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1821_nl = MUX_s_1_2_2(nor_1046_nl, nor_1047_nl, fsm_output[0]);
  assign mux_1823_nl = MUX_s_1_2_2(mux_1822_nl, mux_1821_nl, fsm_output[4]);
  assign nor_1048_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1049_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1819_nl = MUX_s_1_2_2(nor_1048_nl, nor_1049_nl, fsm_output[0]);
  assign nor_1050_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1051_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1818_nl = MUX_s_1_2_2(nor_1050_nl, nor_1051_nl, fsm_output[0]);
  assign mux_1820_nl = MUX_s_1_2_2(mux_1819_nl, mux_1818_nl, fsm_output[4]);
  assign mux_1824_nl = MUX_s_1_2_2(mux_1823_nl, mux_1820_nl, fsm_output[6]);
  assign nand_435_nl = ~((fsm_output[2]) & mux_1824_nl);
  assign or_2110_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00010) | not_tmp_452;
  assign mux_1815_nl = MUX_s_1_2_2(or_tmp_1996, or_2110_nl, fsm_output[0]);
  assign or_2107_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1814_nl = MUX_s_1_2_2(or_tmp_1992, or_2107_nl, fsm_output[0]);
  assign mux_1816_nl = MUX_s_1_2_2(mux_1815_nl, mux_1814_nl, fsm_output[4]);
  assign or_2104_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1812_nl = MUX_s_1_2_2(or_tmp_1990, or_2104_nl, fsm_output[0]);
  assign or_2101_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1811_nl = MUX_s_1_2_2(or_tmp_1986, or_2101_nl, fsm_output[0]);
  assign mux_1813_nl = MUX_s_1_2_2(mux_1812_nl, mux_1811_nl, fsm_output[4]);
  assign mux_1817_nl = MUX_s_1_2_2(mux_1816_nl, mux_1813_nl, fsm_output[6]);
  assign or_4108_nl = (fsm_output[2]) | mux_1817_nl;
  assign mux_1825_nl = MUX_s_1_2_2(nand_435_nl, or_4108_nl, fsm_output[5]);
  assign vec_rsc_0_34_i_we_d_pff = ~(mux_1825_nl | (fsm_output[1]));
  assign or_2143_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2142_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1838_nl = MUX_s_1_2_2(or_2143_nl, or_2142_nl, fsm_output[0]);
  assign or_2144_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1838_nl;
  assign or_2140_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00010)
      | not_tmp_452;
  assign mux_1835_nl = MUX_s_1_2_2(or_2140_nl, or_tmp_1996, fsm_output[0]);
  assign or_2138_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1834_nl = MUX_s_1_2_2(or_2138_nl, or_tmp_1992, fsm_output[0]);
  assign mux_1836_nl = MUX_s_1_2_2(mux_1835_nl, mux_1834_nl, fsm_output[4]);
  assign or_2137_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1832_nl = MUX_s_1_2_2(or_2137_nl, or_tmp_1990, fsm_output[0]);
  assign or_2135_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1831_nl = MUX_s_1_2_2(or_2135_nl, or_tmp_1986, fsm_output[0]);
  assign mux_1833_nl = MUX_s_1_2_2(mux_1832_nl, mux_1831_nl, fsm_output[4]);
  assign mux_1837_nl = MUX_s_1_2_2(mux_1836_nl, mux_1833_nl, fsm_output[6]);
  assign mux_1839_nl = MUX_s_1_2_2(or_2144_nl, mux_1837_nl, fsm_output[2]);
  assign or_2133_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2131_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100010) | (~ and_763_cse);
  assign mux_1828_nl = MUX_s_1_2_2(or_2133_nl, or_2131_nl, fsm_output[0]);
  assign or_2129_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2128_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1827_nl = MUX_s_1_2_2(or_2129_nl, or_2128_nl, fsm_output[0]);
  assign mux_1829_nl = MUX_s_1_2_2(mux_1828_nl, mux_1827_nl, fsm_output[4]);
  assign nor_1042_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1043_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1826_nl = MUX_s_1_2_2(nor_1042_nl, nor_1043_nl, fsm_output[0]);
  assign nand_83_nl = ~((fsm_output[4]) & mux_1826_nl);
  assign mux_1830_nl = MUX_s_1_2_2(mux_1829_nl, nand_83_nl, fsm_output[6]);
  assign or_2134_nl = (fsm_output[2]) | mux_1830_nl;
  assign mux_1840_nl = MUX_s_1_2_2(mux_1839_nl, or_2134_nl, fsm_output[5]);
  assign vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1840_nl) & (fsm_output[1]);
  assign nor_1033_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100011) | (~ and_763_cse));
  assign nor_1034_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | not_tmp_330);
  assign mux_1852_nl = MUX_s_1_2_2(nor_1033_nl, nor_1034_nl, fsm_output[0]);
  assign nor_1035_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1036_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1851_nl = MUX_s_1_2_2(nor_1035_nl, nor_1036_nl, fsm_output[0]);
  assign mux_1853_nl = MUX_s_1_2_2(mux_1852_nl, mux_1851_nl, fsm_output[4]);
  assign nor_1037_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1038_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1849_nl = MUX_s_1_2_2(nor_1037_nl, nor_1038_nl, fsm_output[0]);
  assign nor_1039_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1040_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1848_nl = MUX_s_1_2_2(nor_1039_nl, nor_1040_nl, fsm_output[0]);
  assign mux_1850_nl = MUX_s_1_2_2(mux_1849_nl, mux_1848_nl, fsm_output[4]);
  assign mux_1854_nl = MUX_s_1_2_2(mux_1853_nl, mux_1850_nl, fsm_output[6]);
  assign nand_434_nl = ~((fsm_output[2]) & mux_1854_nl);
  assign or_2154_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00011) | not_tmp_452;
  assign mux_1845_nl = MUX_s_1_2_2(or_tmp_2040, or_2154_nl, fsm_output[0]);
  assign or_2151_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1844_nl = MUX_s_1_2_2(or_tmp_2036, or_2151_nl, fsm_output[0]);
  assign mux_1846_nl = MUX_s_1_2_2(mux_1845_nl, mux_1844_nl, fsm_output[4]);
  assign or_2148_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1842_nl = MUX_s_1_2_2(or_tmp_2034, or_2148_nl, fsm_output[0]);
  assign or_2145_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1841_nl = MUX_s_1_2_2(or_tmp_2030, or_2145_nl, fsm_output[0]);
  assign mux_1843_nl = MUX_s_1_2_2(mux_1842_nl, mux_1841_nl, fsm_output[4]);
  assign mux_1847_nl = MUX_s_1_2_2(mux_1846_nl, mux_1843_nl, fsm_output[6]);
  assign or_4107_nl = (fsm_output[2]) | mux_1847_nl;
  assign mux_1855_nl = MUX_s_1_2_2(nand_434_nl, or_4107_nl, fsm_output[5]);
  assign vec_rsc_0_35_i_we_d_pff = ~(mux_1855_nl | (fsm_output[1]));
  assign or_2187_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2186_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1868_nl = MUX_s_1_2_2(or_2187_nl, or_2186_nl, fsm_output[0]);
  assign or_2188_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1868_nl;
  assign or_2184_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00011)
      | not_tmp_452;
  assign mux_1865_nl = MUX_s_1_2_2(or_2184_nl, or_tmp_2040, fsm_output[0]);
  assign or_2182_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1864_nl = MUX_s_1_2_2(or_2182_nl, or_tmp_2036, fsm_output[0]);
  assign mux_1866_nl = MUX_s_1_2_2(mux_1865_nl, mux_1864_nl, fsm_output[4]);
  assign or_2181_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1862_nl = MUX_s_1_2_2(or_2181_nl, or_tmp_2034, fsm_output[0]);
  assign or_2179_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1861_nl = MUX_s_1_2_2(or_2179_nl, or_tmp_2030, fsm_output[0]);
  assign mux_1863_nl = MUX_s_1_2_2(mux_1862_nl, mux_1861_nl, fsm_output[4]);
  assign mux_1867_nl = MUX_s_1_2_2(mux_1866_nl, mux_1863_nl, fsm_output[6]);
  assign mux_1869_nl = MUX_s_1_2_2(or_2188_nl, mux_1867_nl, fsm_output[2]);
  assign or_2177_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2175_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100011) | (~ and_763_cse);
  assign mux_1858_nl = MUX_s_1_2_2(or_2177_nl, or_2175_nl, fsm_output[0]);
  assign or_2173_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2172_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1857_nl = MUX_s_1_2_2(or_2173_nl, or_2172_nl, fsm_output[0]);
  assign mux_1859_nl = MUX_s_1_2_2(mux_1858_nl, mux_1857_nl, fsm_output[4]);
  assign nor_1031_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1000) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1032_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1856_nl = MUX_s_1_2_2(nor_1031_nl, nor_1032_nl, fsm_output[0]);
  assign nand_85_nl = ~((fsm_output[4]) & mux_1856_nl);
  assign mux_1860_nl = MUX_s_1_2_2(mux_1859_nl, nand_85_nl, fsm_output[6]);
  assign or_2178_nl = (fsm_output[2]) | mux_1860_nl;
  assign mux_1870_nl = MUX_s_1_2_2(mux_1869_nl, or_2178_nl, fsm_output[5]);
  assign vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1870_nl) & (fsm_output[1]);
  assign nor_1022_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100100) | (~ and_763_cse));
  assign nor_1023_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_1882_nl = MUX_s_1_2_2(nor_1022_nl, nor_1023_nl, fsm_output[0]);
  assign nor_1024_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1025_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1881_nl = MUX_s_1_2_2(nor_1024_nl, nor_1025_nl, fsm_output[0]);
  assign mux_1883_nl = MUX_s_1_2_2(mux_1882_nl, mux_1881_nl, fsm_output[4]);
  assign nor_1026_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1027_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1879_nl = MUX_s_1_2_2(nor_1026_nl, nor_1027_nl, fsm_output[0]);
  assign nor_1028_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1029_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1878_nl = MUX_s_1_2_2(nor_1028_nl, nor_1029_nl, fsm_output[0]);
  assign mux_1880_nl = MUX_s_1_2_2(mux_1879_nl, mux_1878_nl, fsm_output[4]);
  assign mux_1884_nl = MUX_s_1_2_2(mux_1883_nl, mux_1880_nl, fsm_output[6]);
  assign nand_433_nl = ~((fsm_output[2]) & mux_1884_nl);
  assign or_2198_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00100) | not_tmp_452;
  assign mux_1875_nl = MUX_s_1_2_2(or_tmp_2084, or_2198_nl, fsm_output[0]);
  assign or_2195_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1874_nl = MUX_s_1_2_2(or_tmp_2080, or_2195_nl, fsm_output[0]);
  assign mux_1876_nl = MUX_s_1_2_2(mux_1875_nl, mux_1874_nl, fsm_output[4]);
  assign or_2192_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1872_nl = MUX_s_1_2_2(or_tmp_2078, or_2192_nl, fsm_output[0]);
  assign or_2189_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1871_nl = MUX_s_1_2_2(or_tmp_2074, or_2189_nl, fsm_output[0]);
  assign mux_1873_nl = MUX_s_1_2_2(mux_1872_nl, mux_1871_nl, fsm_output[4]);
  assign mux_1877_nl = MUX_s_1_2_2(mux_1876_nl, mux_1873_nl, fsm_output[6]);
  assign or_4106_nl = (fsm_output[2]) | mux_1877_nl;
  assign mux_1885_nl = MUX_s_1_2_2(nand_433_nl, or_4106_nl, fsm_output[5]);
  assign vec_rsc_0_36_i_we_d_pff = ~(mux_1885_nl | (fsm_output[1]));
  assign or_2231_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2230_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1898_nl = MUX_s_1_2_2(or_2231_nl, or_2230_nl, fsm_output[0]);
  assign or_2232_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1898_nl;
  assign or_2228_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00100)
      | not_tmp_452;
  assign mux_1895_nl = MUX_s_1_2_2(or_2228_nl, or_tmp_2084, fsm_output[0]);
  assign or_2226_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1894_nl = MUX_s_1_2_2(or_2226_nl, or_tmp_2080, fsm_output[0]);
  assign mux_1896_nl = MUX_s_1_2_2(mux_1895_nl, mux_1894_nl, fsm_output[4]);
  assign or_2225_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1892_nl = MUX_s_1_2_2(or_2225_nl, or_tmp_2078, fsm_output[0]);
  assign or_2223_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1891_nl = MUX_s_1_2_2(or_2223_nl, or_tmp_2074, fsm_output[0]);
  assign mux_1893_nl = MUX_s_1_2_2(mux_1892_nl, mux_1891_nl, fsm_output[4]);
  assign mux_1897_nl = MUX_s_1_2_2(mux_1896_nl, mux_1893_nl, fsm_output[6]);
  assign mux_1899_nl = MUX_s_1_2_2(or_2232_nl, mux_1897_nl, fsm_output[2]);
  assign or_2221_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2219_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100100) | (~ and_763_cse);
  assign mux_1888_nl = MUX_s_1_2_2(or_2221_nl, or_2219_nl, fsm_output[0]);
  assign or_2217_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2216_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1887_nl = MUX_s_1_2_2(or_2217_nl, or_2216_nl, fsm_output[0]);
  assign mux_1889_nl = MUX_s_1_2_2(mux_1888_nl, mux_1887_nl, fsm_output[4]);
  assign nor_1020_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1021_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1886_nl = MUX_s_1_2_2(nor_1020_nl, nor_1021_nl, fsm_output[0]);
  assign nand_87_nl = ~((fsm_output[4]) & mux_1886_nl);
  assign mux_1890_nl = MUX_s_1_2_2(mux_1889_nl, nand_87_nl, fsm_output[6]);
  assign or_2222_nl = (fsm_output[2]) | mux_1890_nl;
  assign mux_1900_nl = MUX_s_1_2_2(mux_1899_nl, or_2222_nl, fsm_output[5]);
  assign vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1900_nl) & (fsm_output[1]);
  assign nor_1011_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100101) | (~ and_763_cse));
  assign nor_1012_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_1912_nl = MUX_s_1_2_2(nor_1011_nl, nor_1012_nl, fsm_output[0]);
  assign nor_1013_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1014_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1911_nl = MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output[0]);
  assign mux_1913_nl = MUX_s_1_2_2(mux_1912_nl, mux_1911_nl, fsm_output[4]);
  assign nor_1015_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1016_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1909_nl = MUX_s_1_2_2(nor_1015_nl, nor_1016_nl, fsm_output[0]);
  assign nor_1017_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1018_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1908_nl = MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output[0]);
  assign mux_1910_nl = MUX_s_1_2_2(mux_1909_nl, mux_1908_nl, fsm_output[4]);
  assign mux_1914_nl = MUX_s_1_2_2(mux_1913_nl, mux_1910_nl, fsm_output[6]);
  assign nand_432_nl = ~((fsm_output[2]) & mux_1914_nl);
  assign or_2242_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00101) | not_tmp_452;
  assign mux_1905_nl = MUX_s_1_2_2(or_tmp_2128, or_2242_nl, fsm_output[0]);
  assign or_2239_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1904_nl = MUX_s_1_2_2(or_tmp_2124, or_2239_nl, fsm_output[0]);
  assign mux_1906_nl = MUX_s_1_2_2(mux_1905_nl, mux_1904_nl, fsm_output[4]);
  assign or_2236_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1902_nl = MUX_s_1_2_2(or_tmp_2122, or_2236_nl, fsm_output[0]);
  assign or_2233_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1901_nl = MUX_s_1_2_2(or_tmp_2118, or_2233_nl, fsm_output[0]);
  assign mux_1903_nl = MUX_s_1_2_2(mux_1902_nl, mux_1901_nl, fsm_output[4]);
  assign mux_1907_nl = MUX_s_1_2_2(mux_1906_nl, mux_1903_nl, fsm_output[6]);
  assign or_4105_nl = (fsm_output[2]) | mux_1907_nl;
  assign mux_1915_nl = MUX_s_1_2_2(nand_432_nl, or_4105_nl, fsm_output[5]);
  assign vec_rsc_0_37_i_we_d_pff = ~(mux_1915_nl | (fsm_output[1]));
  assign or_2275_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2274_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1928_nl = MUX_s_1_2_2(or_2275_nl, or_2274_nl, fsm_output[0]);
  assign or_2276_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1928_nl;
  assign or_2272_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00101)
      | not_tmp_452;
  assign mux_1925_nl = MUX_s_1_2_2(or_2272_nl, or_tmp_2128, fsm_output[0]);
  assign or_2270_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1924_nl = MUX_s_1_2_2(or_2270_nl, or_tmp_2124, fsm_output[0]);
  assign mux_1926_nl = MUX_s_1_2_2(mux_1925_nl, mux_1924_nl, fsm_output[4]);
  assign or_2269_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1922_nl = MUX_s_1_2_2(or_2269_nl, or_tmp_2122, fsm_output[0]);
  assign or_2267_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1921_nl = MUX_s_1_2_2(or_2267_nl, or_tmp_2118, fsm_output[0]);
  assign mux_1923_nl = MUX_s_1_2_2(mux_1922_nl, mux_1921_nl, fsm_output[4]);
  assign mux_1927_nl = MUX_s_1_2_2(mux_1926_nl, mux_1923_nl, fsm_output[6]);
  assign mux_1929_nl = MUX_s_1_2_2(or_2276_nl, mux_1927_nl, fsm_output[2]);
  assign or_2265_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2263_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100101) | (~ and_763_cse);
  assign mux_1918_nl = MUX_s_1_2_2(or_2265_nl, or_2263_nl, fsm_output[0]);
  assign or_2261_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2260_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1917_nl = MUX_s_1_2_2(or_2261_nl, or_2260_nl, fsm_output[0]);
  assign mux_1919_nl = MUX_s_1_2_2(mux_1918_nl, mux_1917_nl, fsm_output[4]);
  assign nor_1009_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1010_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1916_nl = MUX_s_1_2_2(nor_1009_nl, nor_1010_nl, fsm_output[0]);
  assign nand_89_nl = ~((fsm_output[4]) & mux_1916_nl);
  assign mux_1920_nl = MUX_s_1_2_2(mux_1919_nl, nand_89_nl, fsm_output[6]);
  assign or_2266_nl = (fsm_output[2]) | mux_1920_nl;
  assign mux_1930_nl = MUX_s_1_2_2(mux_1929_nl, or_2266_nl, fsm_output[5]);
  assign vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1930_nl) & (fsm_output[1]);
  assign nor_1000_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100110) | (~ and_763_cse));
  assign nor_1001_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_1942_nl = MUX_s_1_2_2(nor_1000_nl, nor_1001_nl, fsm_output[0]);
  assign nor_1002_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_1003_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1941_nl = MUX_s_1_2_2(nor_1002_nl, nor_1003_nl, fsm_output[0]);
  assign mux_1943_nl = MUX_s_1_2_2(mux_1942_nl, mux_1941_nl, fsm_output[4]);
  assign nor_1004_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_1005_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1939_nl = MUX_s_1_2_2(nor_1004_nl, nor_1005_nl, fsm_output[0]);
  assign nor_1006_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_1007_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1938_nl = MUX_s_1_2_2(nor_1006_nl, nor_1007_nl, fsm_output[0]);
  assign mux_1940_nl = MUX_s_1_2_2(mux_1939_nl, mux_1938_nl, fsm_output[4]);
  assign mux_1944_nl = MUX_s_1_2_2(mux_1943_nl, mux_1940_nl, fsm_output[6]);
  assign nand_431_nl = ~((fsm_output[2]) & mux_1944_nl);
  assign or_2286_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00110) | not_tmp_452;
  assign mux_1935_nl = MUX_s_1_2_2(or_tmp_2172, or_2286_nl, fsm_output[0]);
  assign or_2283_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1934_nl = MUX_s_1_2_2(or_tmp_2168, or_2283_nl, fsm_output[0]);
  assign mux_1936_nl = MUX_s_1_2_2(mux_1935_nl, mux_1934_nl, fsm_output[4]);
  assign or_2280_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1932_nl = MUX_s_1_2_2(or_tmp_2166, or_2280_nl, fsm_output[0]);
  assign or_2277_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1931_nl = MUX_s_1_2_2(or_tmp_2162, or_2277_nl, fsm_output[0]);
  assign mux_1933_nl = MUX_s_1_2_2(mux_1932_nl, mux_1931_nl, fsm_output[4]);
  assign mux_1937_nl = MUX_s_1_2_2(mux_1936_nl, mux_1933_nl, fsm_output[6]);
  assign or_4104_nl = (fsm_output[2]) | mux_1937_nl;
  assign mux_1945_nl = MUX_s_1_2_2(nand_431_nl, or_4104_nl, fsm_output[5]);
  assign vec_rsc_0_38_i_we_d_pff = ~(mux_1945_nl | (fsm_output[1]));
  assign or_2319_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2318_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1958_nl = MUX_s_1_2_2(or_2319_nl, or_2318_nl, fsm_output[0]);
  assign or_2320_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1958_nl;
  assign or_2316_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00110)
      | not_tmp_452;
  assign mux_1955_nl = MUX_s_1_2_2(or_2316_nl, or_tmp_2172, fsm_output[0]);
  assign or_2314_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1954_nl = MUX_s_1_2_2(or_2314_nl, or_tmp_2168, fsm_output[0]);
  assign mux_1956_nl = MUX_s_1_2_2(mux_1955_nl, mux_1954_nl, fsm_output[4]);
  assign or_2313_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1952_nl = MUX_s_1_2_2(or_2313_nl, or_tmp_2166, fsm_output[0]);
  assign or_2311_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1951_nl = MUX_s_1_2_2(or_2311_nl, or_tmp_2162, fsm_output[0]);
  assign mux_1953_nl = MUX_s_1_2_2(mux_1952_nl, mux_1951_nl, fsm_output[4]);
  assign mux_1957_nl = MUX_s_1_2_2(mux_1956_nl, mux_1953_nl, fsm_output[6]);
  assign mux_1959_nl = MUX_s_1_2_2(or_2320_nl, mux_1957_nl, fsm_output[2]);
  assign or_2309_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2307_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100110) | (~ and_763_cse);
  assign mux_1948_nl = MUX_s_1_2_2(or_2309_nl, or_2307_nl, fsm_output[0]);
  assign or_2305_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2304_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1947_nl = MUX_s_1_2_2(or_2305_nl, or_2304_nl, fsm_output[0]);
  assign mux_1949_nl = MUX_s_1_2_2(mux_1948_nl, mux_1947_nl, fsm_output[4]);
  assign nor_998_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_999_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1946_nl = MUX_s_1_2_2(nor_998_nl, nor_999_nl, fsm_output[0]);
  assign nand_91_nl = ~((fsm_output[4]) & mux_1946_nl);
  assign mux_1950_nl = MUX_s_1_2_2(mux_1949_nl, nand_91_nl, fsm_output[6]);
  assign or_2310_nl = (fsm_output[2]) | mux_1950_nl;
  assign mux_1960_nl = MUX_s_1_2_2(mux_1959_nl, or_2310_nl, fsm_output[5]);
  assign vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1960_nl) & (fsm_output[1]);
  assign and_590_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b100111) & and_763_cse;
  assign nor_990_nl = ~((COMP_LOOP_acc_13_psp_sva[3:1]!=3'b100) | not_tmp_347);
  assign mux_1972_nl = MUX_s_1_2_2(and_590_nl, nor_990_nl, fsm_output[0]);
  assign nor_991_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b100111) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_992_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_1971_nl = MUX_s_1_2_2(nor_991_nl, nor_992_nl, fsm_output[0]);
  assign mux_1973_nl = MUX_s_1_2_2(mux_1972_nl, mux_1971_nl, fsm_output[4]);
  assign nor_993_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_994_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1969_nl = MUX_s_1_2_2(nor_993_nl, nor_994_nl, fsm_output[0]);
  assign nor_995_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_996_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1968_nl = MUX_s_1_2_2(nor_995_nl, nor_996_nl, fsm_output[0]);
  assign mux_1970_nl = MUX_s_1_2_2(mux_1969_nl, mux_1968_nl, fsm_output[4]);
  assign mux_1974_nl = MUX_s_1_2_2(mux_1973_nl, mux_1970_nl, fsm_output[6]);
  assign nand_430_nl = ~((fsm_output[2]) & mux_1974_nl);
  assign or_2330_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00111) | not_tmp_452;
  assign mux_1965_nl = MUX_s_1_2_2(or_tmp_2216, or_2330_nl, fsm_output[0]);
  assign or_2327_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1964_nl = MUX_s_1_2_2(or_tmp_2212, or_2327_nl, fsm_output[0]);
  assign mux_1966_nl = MUX_s_1_2_2(mux_1965_nl, mux_1964_nl, fsm_output[4]);
  assign or_2324_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1962_nl = MUX_s_1_2_2(or_tmp_2210, or_2324_nl, fsm_output[0]);
  assign or_2321_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1961_nl = MUX_s_1_2_2(or_tmp_2206, or_2321_nl, fsm_output[0]);
  assign mux_1963_nl = MUX_s_1_2_2(mux_1962_nl, mux_1961_nl, fsm_output[4]);
  assign mux_1967_nl = MUX_s_1_2_2(mux_1966_nl, mux_1963_nl, fsm_output[6]);
  assign or_4103_nl = (fsm_output[2]) | mux_1967_nl;
  assign mux_1975_nl = MUX_s_1_2_2(nand_430_nl, or_4103_nl, fsm_output[5]);
  assign vec_rsc_0_39_i_we_d_pff = ~(mux_1975_nl | (fsm_output[1]));
  assign or_2363_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b100111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2362_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1988_nl = MUX_s_1_2_2(or_2363_nl, or_2362_nl, fsm_output[0]);
  assign or_2364_nl = (fsm_output[6]) | (fsm_output[4]) | mux_1988_nl;
  assign or_2360_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b00111)
      | not_tmp_452;
  assign mux_1985_nl = MUX_s_1_2_2(or_2360_nl, or_tmp_2216, fsm_output[0]);
  assign or_2358_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b100111)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_1984_nl = MUX_s_1_2_2(or_2358_nl, or_tmp_2212, fsm_output[0]);
  assign mux_1986_nl = MUX_s_1_2_2(mux_1985_nl, mux_1984_nl, fsm_output[4]);
  assign or_2357_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b100111)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_1982_nl = MUX_s_1_2_2(or_2357_nl, or_tmp_2210, fsm_output[0]);
  assign or_2355_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b100111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_1981_nl = MUX_s_1_2_2(or_2355_nl, or_tmp_2206, fsm_output[0]);
  assign mux_1983_nl = MUX_s_1_2_2(mux_1982_nl, mux_1981_nl, fsm_output[4]);
  assign mux_1987_nl = MUX_s_1_2_2(mux_1986_nl, mux_1983_nl, fsm_output[6]);
  assign mux_1989_nl = MUX_s_1_2_2(or_2364_nl, mux_1987_nl, fsm_output[2]);
  assign or_2353_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10011) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign nand_296_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b100111) & and_763_cse);
  assign mux_1978_nl = MUX_s_1_2_2(or_2353_nl, nand_296_nl, fsm_output[0]);
  assign or_2349_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2348_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b100111) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1977_nl = MUX_s_1_2_2(or_2349_nl, or_2348_nl, fsm_output[0]);
  assign mux_1979_nl = MUX_s_1_2_2(mux_1978_nl, mux_1977_nl, fsm_output[4]);
  assign nor_988_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1001) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_989_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b100111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_1976_nl = MUX_s_1_2_2(nor_988_nl, nor_989_nl, fsm_output[0]);
  assign nand_93_nl = ~((fsm_output[4]) & mux_1976_nl);
  assign mux_1980_nl = MUX_s_1_2_2(mux_1979_nl, nand_93_nl, fsm_output[6]);
  assign or_2354_nl = (fsm_output[2]) | mux_1980_nl;
  assign mux_1990_nl = MUX_s_1_2_2(mux_1989_nl, or_2354_nl, fsm_output[5]);
  assign vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_1990_nl) & (fsm_output[1]);
  assign nor_979_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101000) | (~ and_763_cse));
  assign nor_980_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_2002_nl = MUX_s_1_2_2(nor_979_nl, nor_980_nl, fsm_output[0]);
  assign nor_981_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_982_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2001_nl = MUX_s_1_2_2(nor_981_nl, nor_982_nl, fsm_output[0]);
  assign mux_2003_nl = MUX_s_1_2_2(mux_2002_nl, mux_2001_nl, fsm_output[4]);
  assign nor_983_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_984_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_1999_nl = MUX_s_1_2_2(nor_983_nl, nor_984_nl, fsm_output[0]);
  assign nor_985_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_986_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_1998_nl = MUX_s_1_2_2(nor_985_nl, nor_986_nl, fsm_output[0]);
  assign mux_2000_nl = MUX_s_1_2_2(mux_1999_nl, mux_1998_nl, fsm_output[4]);
  assign mux_2004_nl = MUX_s_1_2_2(mux_2003_nl, mux_2000_nl, fsm_output[6]);
  assign nand_429_nl = ~((fsm_output[2]) & mux_2004_nl);
  assign or_2374_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01000) | not_tmp_452;
  assign mux_1995_nl = MUX_s_1_2_2(or_tmp_2260, or_2374_nl, fsm_output[0]);
  assign or_2371_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_1994_nl = MUX_s_1_2_2(or_tmp_2256, or_2371_nl, fsm_output[0]);
  assign mux_1996_nl = MUX_s_1_2_2(mux_1995_nl, mux_1994_nl, fsm_output[4]);
  assign or_2368_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_1992_nl = MUX_s_1_2_2(or_tmp_2254, or_2368_nl, fsm_output[0]);
  assign or_2365_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_1991_nl = MUX_s_1_2_2(or_tmp_2250, or_2365_nl, fsm_output[0]);
  assign mux_1993_nl = MUX_s_1_2_2(mux_1992_nl, mux_1991_nl, fsm_output[4]);
  assign mux_1997_nl = MUX_s_1_2_2(mux_1996_nl, mux_1993_nl, fsm_output[6]);
  assign or_4102_nl = (fsm_output[2]) | mux_1997_nl;
  assign mux_2005_nl = MUX_s_1_2_2(nand_429_nl, or_4102_nl, fsm_output[5]);
  assign vec_rsc_0_40_i_we_d_pff = ~(mux_2005_nl | (fsm_output[1]));
  assign or_2407_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2406_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2018_nl = MUX_s_1_2_2(or_2407_nl, or_2406_nl, fsm_output[0]);
  assign or_2408_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2018_nl;
  assign or_2404_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01000)
      | not_tmp_452;
  assign mux_2015_nl = MUX_s_1_2_2(or_2404_nl, or_tmp_2260, fsm_output[0]);
  assign or_2402_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2014_nl = MUX_s_1_2_2(or_2402_nl, or_tmp_2256, fsm_output[0]);
  assign mux_2016_nl = MUX_s_1_2_2(mux_2015_nl, mux_2014_nl, fsm_output[4]);
  assign or_2401_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2012_nl = MUX_s_1_2_2(or_2401_nl, or_tmp_2254, fsm_output[0]);
  assign or_2399_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2011_nl = MUX_s_1_2_2(or_2399_nl, or_tmp_2250, fsm_output[0]);
  assign mux_2013_nl = MUX_s_1_2_2(mux_2012_nl, mux_2011_nl, fsm_output[4]);
  assign mux_2017_nl = MUX_s_1_2_2(mux_2016_nl, mux_2013_nl, fsm_output[6]);
  assign mux_2019_nl = MUX_s_1_2_2(or_2408_nl, mux_2017_nl, fsm_output[2]);
  assign or_2397_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2395_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101000) | (~ and_763_cse);
  assign mux_2008_nl = MUX_s_1_2_2(or_2397_nl, or_2395_nl, fsm_output[0]);
  assign or_2393_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2392_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2007_nl = MUX_s_1_2_2(or_2393_nl, or_2392_nl, fsm_output[0]);
  assign mux_2009_nl = MUX_s_1_2_2(mux_2008_nl, mux_2007_nl, fsm_output[4]);
  assign nor_977_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_978_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2006_nl = MUX_s_1_2_2(nor_977_nl, nor_978_nl, fsm_output[0]);
  assign nand_95_nl = ~((fsm_output[4]) & mux_2006_nl);
  assign mux_2010_nl = MUX_s_1_2_2(mux_2009_nl, nand_95_nl, fsm_output[6]);
  assign or_2398_nl = (fsm_output[2]) | mux_2010_nl;
  assign mux_2020_nl = MUX_s_1_2_2(mux_2019_nl, or_2398_nl, fsm_output[5]);
  assign vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2020_nl) & (fsm_output[1]);
  assign nor_968_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101001) | (~ and_763_cse));
  assign nor_969_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_2032_nl = MUX_s_1_2_2(nor_968_nl, nor_969_nl, fsm_output[0]);
  assign nor_970_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_971_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2031_nl = MUX_s_1_2_2(nor_970_nl, nor_971_nl, fsm_output[0]);
  assign mux_2033_nl = MUX_s_1_2_2(mux_2032_nl, mux_2031_nl, fsm_output[4]);
  assign nor_972_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_973_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2029_nl = MUX_s_1_2_2(nor_972_nl, nor_973_nl, fsm_output[0]);
  assign nor_974_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_975_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2028_nl = MUX_s_1_2_2(nor_974_nl, nor_975_nl, fsm_output[0]);
  assign mux_2030_nl = MUX_s_1_2_2(mux_2029_nl, mux_2028_nl, fsm_output[4]);
  assign mux_2034_nl = MUX_s_1_2_2(mux_2033_nl, mux_2030_nl, fsm_output[6]);
  assign nand_428_nl = ~((fsm_output[2]) & mux_2034_nl);
  assign or_2418_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01001) | not_tmp_452;
  assign mux_2025_nl = MUX_s_1_2_2(or_tmp_2304, or_2418_nl, fsm_output[0]);
  assign or_2415_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2024_nl = MUX_s_1_2_2(or_tmp_2300, or_2415_nl, fsm_output[0]);
  assign mux_2026_nl = MUX_s_1_2_2(mux_2025_nl, mux_2024_nl, fsm_output[4]);
  assign or_2412_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2022_nl = MUX_s_1_2_2(or_tmp_2298, or_2412_nl, fsm_output[0]);
  assign or_2409_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2021_nl = MUX_s_1_2_2(or_tmp_2294, or_2409_nl, fsm_output[0]);
  assign mux_2023_nl = MUX_s_1_2_2(mux_2022_nl, mux_2021_nl, fsm_output[4]);
  assign mux_2027_nl = MUX_s_1_2_2(mux_2026_nl, mux_2023_nl, fsm_output[6]);
  assign or_4101_nl = (fsm_output[2]) | mux_2027_nl;
  assign mux_2035_nl = MUX_s_1_2_2(nand_428_nl, or_4101_nl, fsm_output[5]);
  assign vec_rsc_0_41_i_we_d_pff = ~(mux_2035_nl | (fsm_output[1]));
  assign or_2451_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2450_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2048_nl = MUX_s_1_2_2(or_2451_nl, or_2450_nl, fsm_output[0]);
  assign or_2452_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2048_nl;
  assign or_2448_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01001)
      | not_tmp_452;
  assign mux_2045_nl = MUX_s_1_2_2(or_2448_nl, or_tmp_2304, fsm_output[0]);
  assign or_2446_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2044_nl = MUX_s_1_2_2(or_2446_nl, or_tmp_2300, fsm_output[0]);
  assign mux_2046_nl = MUX_s_1_2_2(mux_2045_nl, mux_2044_nl, fsm_output[4]);
  assign or_2445_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2042_nl = MUX_s_1_2_2(or_2445_nl, or_tmp_2298, fsm_output[0]);
  assign or_2443_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2041_nl = MUX_s_1_2_2(or_2443_nl, or_tmp_2294, fsm_output[0]);
  assign mux_2043_nl = MUX_s_1_2_2(mux_2042_nl, mux_2041_nl, fsm_output[4]);
  assign mux_2047_nl = MUX_s_1_2_2(mux_2046_nl, mux_2043_nl, fsm_output[6]);
  assign mux_2049_nl = MUX_s_1_2_2(or_2452_nl, mux_2047_nl, fsm_output[2]);
  assign or_2441_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2439_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101001) | (~ and_763_cse);
  assign mux_2038_nl = MUX_s_1_2_2(or_2441_nl, or_2439_nl, fsm_output[0]);
  assign or_2437_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2436_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2037_nl = MUX_s_1_2_2(or_2437_nl, or_2436_nl, fsm_output[0]);
  assign mux_2039_nl = MUX_s_1_2_2(mux_2038_nl, mux_2037_nl, fsm_output[4]);
  assign nor_966_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_967_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2036_nl = MUX_s_1_2_2(nor_966_nl, nor_967_nl, fsm_output[0]);
  assign nand_97_nl = ~((fsm_output[4]) & mux_2036_nl);
  assign mux_2040_nl = MUX_s_1_2_2(mux_2039_nl, nand_97_nl, fsm_output[6]);
  assign or_2442_nl = (fsm_output[2]) | mux_2040_nl;
  assign mux_2050_nl = MUX_s_1_2_2(mux_2049_nl, or_2442_nl, fsm_output[5]);
  assign vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2050_nl) & (fsm_output[1]);
  assign nor_957_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101010) | (~ and_763_cse));
  assign nor_958_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_2062_nl = MUX_s_1_2_2(nor_957_nl, nor_958_nl, fsm_output[0]);
  assign nor_959_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_960_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2061_nl = MUX_s_1_2_2(nor_959_nl, nor_960_nl, fsm_output[0]);
  assign mux_2063_nl = MUX_s_1_2_2(mux_2062_nl, mux_2061_nl, fsm_output[4]);
  assign nor_961_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_962_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2059_nl = MUX_s_1_2_2(nor_961_nl, nor_962_nl, fsm_output[0]);
  assign nor_963_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_964_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2058_nl = MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output[0]);
  assign mux_2060_nl = MUX_s_1_2_2(mux_2059_nl, mux_2058_nl, fsm_output[4]);
  assign mux_2064_nl = MUX_s_1_2_2(mux_2063_nl, mux_2060_nl, fsm_output[6]);
  assign nand_427_nl = ~((fsm_output[2]) & mux_2064_nl);
  assign or_2462_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01010) | not_tmp_452;
  assign mux_2055_nl = MUX_s_1_2_2(or_tmp_2348, or_2462_nl, fsm_output[0]);
  assign or_2459_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2054_nl = MUX_s_1_2_2(or_tmp_2344, or_2459_nl, fsm_output[0]);
  assign mux_2056_nl = MUX_s_1_2_2(mux_2055_nl, mux_2054_nl, fsm_output[4]);
  assign or_2456_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2052_nl = MUX_s_1_2_2(or_tmp_2342, or_2456_nl, fsm_output[0]);
  assign or_2453_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2051_nl = MUX_s_1_2_2(or_tmp_2338, or_2453_nl, fsm_output[0]);
  assign mux_2053_nl = MUX_s_1_2_2(mux_2052_nl, mux_2051_nl, fsm_output[4]);
  assign mux_2057_nl = MUX_s_1_2_2(mux_2056_nl, mux_2053_nl, fsm_output[6]);
  assign or_4100_nl = (fsm_output[2]) | mux_2057_nl;
  assign mux_2065_nl = MUX_s_1_2_2(nand_427_nl, or_4100_nl, fsm_output[5]);
  assign vec_rsc_0_42_i_we_d_pff = ~(mux_2065_nl | (fsm_output[1]));
  assign or_2495_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2494_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2078_nl = MUX_s_1_2_2(or_2495_nl, or_2494_nl, fsm_output[0]);
  assign or_2496_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2078_nl;
  assign or_2492_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01010)
      | not_tmp_452;
  assign mux_2075_nl = MUX_s_1_2_2(or_2492_nl, or_tmp_2348, fsm_output[0]);
  assign or_2490_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2074_nl = MUX_s_1_2_2(or_2490_nl, or_tmp_2344, fsm_output[0]);
  assign mux_2076_nl = MUX_s_1_2_2(mux_2075_nl, mux_2074_nl, fsm_output[4]);
  assign or_2489_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2072_nl = MUX_s_1_2_2(or_2489_nl, or_tmp_2342, fsm_output[0]);
  assign or_2487_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2071_nl = MUX_s_1_2_2(or_2487_nl, or_tmp_2338, fsm_output[0]);
  assign mux_2073_nl = MUX_s_1_2_2(mux_2072_nl, mux_2071_nl, fsm_output[4]);
  assign mux_2077_nl = MUX_s_1_2_2(mux_2076_nl, mux_2073_nl, fsm_output[6]);
  assign mux_2079_nl = MUX_s_1_2_2(or_2496_nl, mux_2077_nl, fsm_output[2]);
  assign or_2485_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2483_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101010) | (~ and_763_cse);
  assign mux_2068_nl = MUX_s_1_2_2(or_2485_nl, or_2483_nl, fsm_output[0]);
  assign or_2481_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2480_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2067_nl = MUX_s_1_2_2(or_2481_nl, or_2480_nl, fsm_output[0]);
  assign mux_2069_nl = MUX_s_1_2_2(mux_2068_nl, mux_2067_nl, fsm_output[4]);
  assign nor_955_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_956_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2066_nl = MUX_s_1_2_2(nor_955_nl, nor_956_nl, fsm_output[0]);
  assign nand_99_nl = ~((fsm_output[4]) & mux_2066_nl);
  assign mux_2070_nl = MUX_s_1_2_2(mux_2069_nl, nand_99_nl, fsm_output[6]);
  assign or_2486_nl = (fsm_output[2]) | mux_2070_nl;
  assign mux_2080_nl = MUX_s_1_2_2(mux_2079_nl, or_2486_nl, fsm_output[5]);
  assign vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2080_nl) & (fsm_output[1]);
  assign and_585_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b101011) & and_763_cse;
  assign nor_947_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | not_tmp_330);
  assign mux_2092_nl = MUX_s_1_2_2(and_585_nl, nor_947_nl, fsm_output[0]);
  assign nor_948_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_949_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2091_nl = MUX_s_1_2_2(nor_948_nl, nor_949_nl, fsm_output[0]);
  assign mux_2093_nl = MUX_s_1_2_2(mux_2092_nl, mux_2091_nl, fsm_output[4]);
  assign nor_950_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_951_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2089_nl = MUX_s_1_2_2(nor_950_nl, nor_951_nl, fsm_output[0]);
  assign nor_952_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_953_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2088_nl = MUX_s_1_2_2(nor_952_nl, nor_953_nl, fsm_output[0]);
  assign mux_2090_nl = MUX_s_1_2_2(mux_2089_nl, mux_2088_nl, fsm_output[4]);
  assign mux_2094_nl = MUX_s_1_2_2(mux_2093_nl, mux_2090_nl, fsm_output[6]);
  assign nand_426_nl = ~((fsm_output[2]) & mux_2094_nl);
  assign or_2506_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01011) | not_tmp_452;
  assign mux_2085_nl = MUX_s_1_2_2(or_tmp_2392, or_2506_nl, fsm_output[0]);
  assign or_2503_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2084_nl = MUX_s_1_2_2(or_tmp_2388, or_2503_nl, fsm_output[0]);
  assign mux_2086_nl = MUX_s_1_2_2(mux_2085_nl, mux_2084_nl, fsm_output[4]);
  assign or_2500_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2082_nl = MUX_s_1_2_2(or_tmp_2386, or_2500_nl, fsm_output[0]);
  assign or_2497_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2081_nl = MUX_s_1_2_2(or_tmp_2382, or_2497_nl, fsm_output[0]);
  assign mux_2083_nl = MUX_s_1_2_2(mux_2082_nl, mux_2081_nl, fsm_output[4]);
  assign mux_2087_nl = MUX_s_1_2_2(mux_2086_nl, mux_2083_nl, fsm_output[6]);
  assign or_4099_nl = (fsm_output[2]) | mux_2087_nl;
  assign mux_2095_nl = MUX_s_1_2_2(nand_426_nl, or_4099_nl, fsm_output[5]);
  assign vec_rsc_0_43_i_we_d_pff = ~(mux_2095_nl | (fsm_output[1]));
  assign or_2539_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2538_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2108_nl = MUX_s_1_2_2(or_2539_nl, or_2538_nl, fsm_output[0]);
  assign or_2540_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2108_nl;
  assign or_2536_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01011)
      | not_tmp_452;
  assign mux_2105_nl = MUX_s_1_2_2(or_2536_nl, or_tmp_2392, fsm_output[0]);
  assign or_2534_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2104_nl = MUX_s_1_2_2(or_2534_nl, or_tmp_2388, fsm_output[0]);
  assign mux_2106_nl = MUX_s_1_2_2(mux_2105_nl, mux_2104_nl, fsm_output[4]);
  assign or_2533_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2102_nl = MUX_s_1_2_2(or_2533_nl, or_tmp_2386, fsm_output[0]);
  assign or_2531_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2101_nl = MUX_s_1_2_2(or_2531_nl, or_tmp_2382, fsm_output[0]);
  assign mux_2103_nl = MUX_s_1_2_2(mux_2102_nl, mux_2101_nl, fsm_output[4]);
  assign mux_2107_nl = MUX_s_1_2_2(mux_2106_nl, mux_2103_nl, fsm_output[6]);
  assign mux_2109_nl = MUX_s_1_2_2(or_2540_nl, mux_2107_nl, fsm_output[2]);
  assign or_2529_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10101) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign nand_295_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b101011) & and_763_cse);
  assign mux_2098_nl = MUX_s_1_2_2(or_2529_nl, nand_295_nl, fsm_output[0]);
  assign or_2525_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2524_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2097_nl = MUX_s_1_2_2(or_2525_nl, or_2524_nl, fsm_output[0]);
  assign mux_2099_nl = MUX_s_1_2_2(mux_2098_nl, mux_2097_nl, fsm_output[4]);
  assign nor_945_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1010) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_946_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2096_nl = MUX_s_1_2_2(nor_945_nl, nor_946_nl, fsm_output[0]);
  assign nand_101_nl = ~((fsm_output[4]) & mux_2096_nl);
  assign mux_2100_nl = MUX_s_1_2_2(mux_2099_nl, nand_101_nl, fsm_output[6]);
  assign or_2530_nl = (fsm_output[2]) | mux_2100_nl;
  assign mux_2110_nl = MUX_s_1_2_2(mux_2109_nl, or_2530_nl, fsm_output[5]);
  assign vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2110_nl) & (fsm_output[1]);
  assign nor_936_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101100) | (~ and_763_cse));
  assign nor_937_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1011) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_2122_nl = MUX_s_1_2_2(nor_936_nl, nor_937_nl, fsm_output[0]);
  assign nor_938_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_939_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2121_nl = MUX_s_1_2_2(nor_938_nl, nor_939_nl, fsm_output[0]);
  assign mux_2123_nl = MUX_s_1_2_2(mux_2122_nl, mux_2121_nl, fsm_output[4]);
  assign nor_940_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_941_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2119_nl = MUX_s_1_2_2(nor_940_nl, nor_941_nl, fsm_output[0]);
  assign nor_942_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_943_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2118_nl = MUX_s_1_2_2(nor_942_nl, nor_943_nl, fsm_output[0]);
  assign mux_2120_nl = MUX_s_1_2_2(mux_2119_nl, mux_2118_nl, fsm_output[4]);
  assign mux_2124_nl = MUX_s_1_2_2(mux_2123_nl, mux_2120_nl, fsm_output[6]);
  assign nand_425_nl = ~((fsm_output[2]) & mux_2124_nl);
  assign or_2550_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01100) | not_tmp_452;
  assign mux_2115_nl = MUX_s_1_2_2(or_tmp_2436, or_2550_nl, fsm_output[0]);
  assign or_2547_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2114_nl = MUX_s_1_2_2(or_tmp_2432, or_2547_nl, fsm_output[0]);
  assign mux_2116_nl = MUX_s_1_2_2(mux_2115_nl, mux_2114_nl, fsm_output[4]);
  assign or_2544_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2112_nl = MUX_s_1_2_2(or_tmp_2430, or_2544_nl, fsm_output[0]);
  assign or_2541_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2111_nl = MUX_s_1_2_2(or_tmp_2426, or_2541_nl, fsm_output[0]);
  assign mux_2113_nl = MUX_s_1_2_2(mux_2112_nl, mux_2111_nl, fsm_output[4]);
  assign mux_2117_nl = MUX_s_1_2_2(mux_2116_nl, mux_2113_nl, fsm_output[6]);
  assign or_4098_nl = (fsm_output[2]) | mux_2117_nl;
  assign mux_2125_nl = MUX_s_1_2_2(nand_425_nl, or_4098_nl, fsm_output[5]);
  assign vec_rsc_0_44_i_we_d_pff = ~(mux_2125_nl | (fsm_output[1]));
  assign or_2583_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2582_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2138_nl = MUX_s_1_2_2(or_2583_nl, or_2582_nl, fsm_output[0]);
  assign or_2584_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2138_nl;
  assign or_2580_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01100)
      | not_tmp_452;
  assign mux_2135_nl = MUX_s_1_2_2(or_2580_nl, or_tmp_2436, fsm_output[0]);
  assign or_2578_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2134_nl = MUX_s_1_2_2(or_2578_nl, or_tmp_2432, fsm_output[0]);
  assign mux_2136_nl = MUX_s_1_2_2(mux_2135_nl, mux_2134_nl, fsm_output[4]);
  assign or_2577_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2132_nl = MUX_s_1_2_2(or_2577_nl, or_tmp_2430, fsm_output[0]);
  assign or_2575_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2131_nl = MUX_s_1_2_2(or_2575_nl, or_tmp_2426, fsm_output[0]);
  assign mux_2133_nl = MUX_s_1_2_2(mux_2132_nl, mux_2131_nl, fsm_output[4]);
  assign mux_2137_nl = MUX_s_1_2_2(mux_2136_nl, mux_2133_nl, fsm_output[6]);
  assign mux_2139_nl = MUX_s_1_2_2(or_2584_nl, mux_2137_nl, fsm_output[2]);
  assign or_2573_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2571_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101100) | (~ and_763_cse);
  assign mux_2128_nl = MUX_s_1_2_2(or_2573_nl, or_2571_nl, fsm_output[0]);
  assign or_2569_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2568_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2127_nl = MUX_s_1_2_2(or_2569_nl, or_2568_nl, fsm_output[0]);
  assign mux_2129_nl = MUX_s_1_2_2(mux_2128_nl, mux_2127_nl, fsm_output[4]);
  assign nor_934_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_935_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2126_nl = MUX_s_1_2_2(nor_934_nl, nor_935_nl, fsm_output[0]);
  assign nand_103_nl = ~((fsm_output[4]) & mux_2126_nl);
  assign mux_2130_nl = MUX_s_1_2_2(mux_2129_nl, nand_103_nl, fsm_output[6]);
  assign or_2574_nl = (fsm_output[2]) | mux_2130_nl;
  assign mux_2140_nl = MUX_s_1_2_2(mux_2139_nl, or_2574_nl, fsm_output[5]);
  assign vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2140_nl) & (fsm_output[1]);
  assign and_582_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b101101) & and_763_cse;
  assign nor_926_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1011) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_2152_nl = MUX_s_1_2_2(and_582_nl, nor_926_nl, fsm_output[0]);
  assign nor_927_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_928_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2151_nl = MUX_s_1_2_2(nor_927_nl, nor_928_nl, fsm_output[0]);
  assign mux_2153_nl = MUX_s_1_2_2(mux_2152_nl, mux_2151_nl, fsm_output[4]);
  assign nor_929_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_930_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2149_nl = MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output[0]);
  assign nor_931_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_932_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2148_nl = MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output[0]);
  assign mux_2150_nl = MUX_s_1_2_2(mux_2149_nl, mux_2148_nl, fsm_output[4]);
  assign mux_2154_nl = MUX_s_1_2_2(mux_2153_nl, mux_2150_nl, fsm_output[6]);
  assign nand_424_nl = ~((fsm_output[2]) & mux_2154_nl);
  assign or_2594_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01101) | not_tmp_452;
  assign mux_2145_nl = MUX_s_1_2_2(or_tmp_2480, or_2594_nl, fsm_output[0]);
  assign or_2591_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2144_nl = MUX_s_1_2_2(or_tmp_2476, or_2591_nl, fsm_output[0]);
  assign mux_2146_nl = MUX_s_1_2_2(mux_2145_nl, mux_2144_nl, fsm_output[4]);
  assign or_2588_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2142_nl = MUX_s_1_2_2(or_tmp_2474, or_2588_nl, fsm_output[0]);
  assign or_2585_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2141_nl = MUX_s_1_2_2(or_tmp_2470, or_2585_nl, fsm_output[0]);
  assign mux_2143_nl = MUX_s_1_2_2(mux_2142_nl, mux_2141_nl, fsm_output[4]);
  assign mux_2147_nl = MUX_s_1_2_2(mux_2146_nl, mux_2143_nl, fsm_output[6]);
  assign or_4097_nl = (fsm_output[2]) | mux_2147_nl;
  assign mux_2155_nl = MUX_s_1_2_2(nand_424_nl, or_4097_nl, fsm_output[5]);
  assign vec_rsc_0_45_i_we_d_pff = ~(mux_2155_nl | (fsm_output[1]));
  assign or_2627_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2626_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2168_nl = MUX_s_1_2_2(or_2627_nl, or_2626_nl, fsm_output[0]);
  assign or_2628_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2168_nl;
  assign or_2624_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01101)
      | not_tmp_452;
  assign mux_2165_nl = MUX_s_1_2_2(or_2624_nl, or_tmp_2480, fsm_output[0]);
  assign or_2622_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2164_nl = MUX_s_1_2_2(or_2622_nl, or_tmp_2476, fsm_output[0]);
  assign mux_2166_nl = MUX_s_1_2_2(mux_2165_nl, mux_2164_nl, fsm_output[4]);
  assign or_2621_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2162_nl = MUX_s_1_2_2(or_2621_nl, or_tmp_2474, fsm_output[0]);
  assign or_2619_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2161_nl = MUX_s_1_2_2(or_2619_nl, or_tmp_2470, fsm_output[0]);
  assign mux_2163_nl = MUX_s_1_2_2(mux_2162_nl, mux_2161_nl, fsm_output[4]);
  assign mux_2167_nl = MUX_s_1_2_2(mux_2166_nl, mux_2163_nl, fsm_output[6]);
  assign mux_2169_nl = MUX_s_1_2_2(or_2628_nl, mux_2167_nl, fsm_output[2]);
  assign or_2617_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10110) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign nand_294_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b101101) & and_763_cse);
  assign mux_2158_nl = MUX_s_1_2_2(or_2617_nl, nand_294_nl, fsm_output[0]);
  assign or_2613_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2612_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2157_nl = MUX_s_1_2_2(or_2613_nl, or_2612_nl, fsm_output[0]);
  assign mux_2159_nl = MUX_s_1_2_2(mux_2158_nl, mux_2157_nl, fsm_output[4]);
  assign nor_924_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_925_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2156_nl = MUX_s_1_2_2(nor_924_nl, nor_925_nl, fsm_output[0]);
  assign nand_105_nl = ~((fsm_output[4]) & mux_2156_nl);
  assign mux_2160_nl = MUX_s_1_2_2(mux_2159_nl, nand_105_nl, fsm_output[6]);
  assign or_2618_nl = (fsm_output[2]) | mux_2160_nl;
  assign mux_2170_nl = MUX_s_1_2_2(mux_2169_nl, or_2618_nl, fsm_output[5]);
  assign vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2170_nl) & (fsm_output[1]);
  assign and_579_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b101110) & and_763_cse;
  assign and_580_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1011) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b10)
      & and_763_cse;
  assign mux_2182_nl = MUX_s_1_2_2(and_579_nl, and_580_nl, fsm_output[0]);
  assign nor_917_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b101110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_918_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2181_nl = MUX_s_1_2_2(nor_917_nl, nor_918_nl, fsm_output[0]);
  assign mux_2183_nl = MUX_s_1_2_2(mux_2182_nl, mux_2181_nl, fsm_output[4]);
  assign nor_919_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_920_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b10111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2179_nl = MUX_s_1_2_2(nor_919_nl, nor_920_nl, fsm_output[0]);
  assign nor_921_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_922_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2178_nl = MUX_s_1_2_2(nor_921_nl, nor_922_nl, fsm_output[0]);
  assign mux_2180_nl = MUX_s_1_2_2(mux_2179_nl, mux_2178_nl, fsm_output[4]);
  assign mux_2184_nl = MUX_s_1_2_2(mux_2183_nl, mux_2180_nl, fsm_output[6]);
  assign nand_423_nl = ~((fsm_output[2]) & mux_2184_nl);
  assign or_2638_nl = (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01110) | not_tmp_452;
  assign mux_2175_nl = MUX_s_1_2_2(or_tmp_2524, or_2638_nl, fsm_output[0]);
  assign or_2635_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2174_nl = MUX_s_1_2_2(or_tmp_2520, or_2635_nl, fsm_output[0]);
  assign mux_2176_nl = MUX_s_1_2_2(mux_2175_nl, mux_2174_nl, fsm_output[4]);
  assign or_2632_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2172_nl = MUX_s_1_2_2(or_tmp_2518, or_2632_nl, fsm_output[0]);
  assign or_2629_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2171_nl = MUX_s_1_2_2(or_tmp_2514, or_2629_nl, fsm_output[0]);
  assign mux_2173_nl = MUX_s_1_2_2(mux_2172_nl, mux_2171_nl, fsm_output[4]);
  assign mux_2177_nl = MUX_s_1_2_2(mux_2176_nl, mux_2173_nl, fsm_output[6]);
  assign or_4096_nl = (fsm_output[2]) | mux_2177_nl;
  assign mux_2185_nl = MUX_s_1_2_2(nand_423_nl, or_4096_nl, fsm_output[5]);
  assign vec_rsc_0_46_i_we_d_pff = ~(mux_2185_nl | (fsm_output[1]));
  assign or_2671_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2670_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2198_nl = MUX_s_1_2_2(or_2671_nl, or_2670_nl, fsm_output[0]);
  assign or_2672_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2198_nl;
  assign or_2668_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[4:0]!=5'b01110)
      | not_tmp_452;
  assign mux_2195_nl = MUX_s_1_2_2(or_2668_nl, or_tmp_2524, fsm_output[0]);
  assign or_2666_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b101110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2194_nl = MUX_s_1_2_2(or_2666_nl, or_tmp_2520, fsm_output[0]);
  assign mux_2196_nl = MUX_s_1_2_2(mux_2195_nl, mux_2194_nl, fsm_output[4]);
  assign or_2665_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b101110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2192_nl = MUX_s_1_2_2(or_2665_nl, or_tmp_2518, fsm_output[0]);
  assign or_2663_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2191_nl = MUX_s_1_2_2(or_2663_nl, or_tmp_2514, fsm_output[0]);
  assign mux_2193_nl = MUX_s_1_2_2(mux_2192_nl, mux_2191_nl, fsm_output[4]);
  assign mux_2197_nl = MUX_s_1_2_2(mux_2196_nl, mux_2193_nl, fsm_output[6]);
  assign mux_2199_nl = MUX_s_1_2_2(or_2672_nl, mux_2197_nl, fsm_output[2]);
  assign nand_292_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b10111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & and_763_cse);
  assign nand_293_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b101110) & and_763_cse);
  assign mux_2188_nl = MUX_s_1_2_2(nand_292_nl, nand_293_nl, fsm_output[0]);
  assign or_2657_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10111) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2656_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2187_nl = MUX_s_1_2_2(or_2657_nl, or_2656_nl, fsm_output[0]);
  assign mux_2189_nl = MUX_s_1_2_2(mux_2188_nl, mux_2187_nl, fsm_output[4]);
  assign nor_915_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_916_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2186_nl = MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output[0]);
  assign nand_107_nl = ~((fsm_output[4]) & mux_2186_nl);
  assign mux_2190_nl = MUX_s_1_2_2(mux_2189_nl, nand_107_nl, fsm_output[6]);
  assign or_2662_nl = (fsm_output[2]) | mux_2190_nl;
  assign mux_2200_nl = MUX_s_1_2_2(mux_2199_nl, or_2662_nl, fsm_output[5]);
  assign vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2200_nl) & (fsm_output[1]);
  assign and_575_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b101111) & and_763_cse;
  assign nor_909_nl = ~((COMP_LOOP_acc_13_psp_sva[3:1]!=3'b101) | not_tmp_347);
  assign mux_2212_nl = MUX_s_1_2_2(and_575_nl, nor_909_nl, fsm_output[0]);
  assign and_576_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b101111) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_577_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b101) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_2211_nl = MUX_s_1_2_2(and_576_nl, and_577_nl, fsm_output[0]);
  assign mux_2213_nl = MUX_s_1_2_2(mux_2212_nl, mux_2211_nl, fsm_output[4]);
  assign and_812_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b101111) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_819_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b10111) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_2209_nl = MUX_s_1_2_2(and_812_nl, and_819_nl, fsm_output[0]);
  assign nor_912_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b101111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_913_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b10111) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2208_nl = MUX_s_1_2_2(nor_912_nl, nor_913_nl, fsm_output[0]);
  assign mux_2210_nl = MUX_s_1_2_2(mux_2209_nl, mux_2208_nl, fsm_output[4]);
  assign mux_2214_nl = MUX_s_1_2_2(mux_2213_nl, mux_2210_nl, fsm_output[6]);
  assign nand_422_nl = ~((fsm_output[2]) & mux_2214_nl);
  assign or_2682_nl = (~((COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b01111))) | not_tmp_452;
  assign mux_2205_nl = MUX_s_1_2_2(or_tmp_2567, or_2682_nl, fsm_output[0]);
  assign nand_287_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b101111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2204_nl = MUX_s_1_2_2(or_tmp_2564, nand_287_nl, fsm_output[0]);
  assign mux_2206_nl = MUX_s_1_2_2(mux_2205_nl, mux_2204_nl, fsm_output[4]);
  assign nand_477_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b101111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_2202_nl = MUX_s_1_2_2(or_tmp_2562, nand_477_nl, fsm_output[0]);
  assign or_2673_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2201_nl = MUX_s_1_2_2(or_tmp_2558, or_2673_nl, fsm_output[0]);
  assign mux_2203_nl = MUX_s_1_2_2(mux_2202_nl, mux_2201_nl, fsm_output[4]);
  assign mux_2207_nl = MUX_s_1_2_2(mux_2206_nl, mux_2203_nl, fsm_output[6]);
  assign or_4095_nl = (fsm_output[2]) | mux_2207_nl;
  assign mux_2215_nl = MUX_s_1_2_2(nand_422_nl, or_4095_nl, fsm_output[5]);
  assign vec_rsc_0_47_i_we_d_pff = ~(mux_2215_nl | (fsm_output[1]));
  assign or_2714_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b101111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2713_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2228_nl = MUX_s_1_2_2(or_2714_nl, or_2713_nl, fsm_output[0]);
  assign or_2715_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2228_nl;
  assign or_2711_nl = (~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[4:0]==5'b01111)))
      | not_tmp_452;
  assign mux_2225_nl = MUX_s_1_2_2(or_2711_nl, or_tmp_2567, fsm_output[0]);
  assign nand_278_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b101111)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_2224_nl = MUX_s_1_2_2(nand_278_nl, or_tmp_2564, fsm_output[0]);
  assign mux_2226_nl = MUX_s_1_2_2(mux_2225_nl, mux_2224_nl, fsm_output[4]);
  assign nand_402_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b101111)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_2222_nl = MUX_s_1_2_2(nand_402_nl, or_tmp_2562, fsm_output[0]);
  assign or_2706_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b101111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2221_nl = MUX_s_1_2_2(or_2706_nl, or_tmp_2558, fsm_output[0]);
  assign mux_2223_nl = MUX_s_1_2_2(mux_2222_nl, mux_2221_nl, fsm_output[4]);
  assign mux_2227_nl = MUX_s_1_2_2(mux_2226_nl, mux_2223_nl, fsm_output[6]);
  assign mux_2229_nl = MUX_s_1_2_2(or_2715_nl, mux_2227_nl, fsm_output[2]);
  assign or_2704_nl = (~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b10111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm))
      | not_tmp_321;
  assign nand_281_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b101111) & and_763_cse);
  assign mux_2218_nl = MUX_s_1_2_2(or_2704_nl, nand_281_nl, fsm_output[0]);
  assign nand_282_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b10111) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_283_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b101111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2217_nl = MUX_s_1_2_2(nand_282_nl, nand_283_nl, fsm_output[0]);
  assign mux_2219_nl = MUX_s_1_2_2(mux_2218_nl, mux_2217_nl, fsm_output[4]);
  assign nor_907_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1011) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_908_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b101111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2216_nl = MUX_s_1_2_2(nor_907_nl, nor_908_nl, fsm_output[0]);
  assign nand_109_nl = ~((fsm_output[4]) & mux_2216_nl);
  assign mux_2220_nl = MUX_s_1_2_2(mux_2219_nl, nand_109_nl, fsm_output[6]);
  assign or_2705_nl = (fsm_output[2]) | mux_2220_nl;
  assign mux_2230_nl = MUX_s_1_2_2(mux_2229_nl, or_2705_nl, fsm_output[5]);
  assign vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2230_nl) & (fsm_output[1]);
  assign nor_898_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0000) | not_tmp_523);
  assign nor_899_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_2242_nl = MUX_s_1_2_2(nor_898_nl, nor_899_nl, fsm_output[0]);
  assign nor_900_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_901_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2241_nl = MUX_s_1_2_2(nor_900_nl, nor_901_nl, fsm_output[0]);
  assign mux_2243_nl = MUX_s_1_2_2(mux_2242_nl, mux_2241_nl, fsm_output[4]);
  assign nor_902_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_903_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2239_nl = MUX_s_1_2_2(nor_902_nl, nor_903_nl, fsm_output[0]);
  assign nor_904_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_905_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11000) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2238_nl = MUX_s_1_2_2(nor_904_nl, nor_905_nl, fsm_output[0]);
  assign mux_2240_nl = MUX_s_1_2_2(mux_2239_nl, mux_2238_nl, fsm_output[4]);
  assign mux_2244_nl = MUX_s_1_2_2(mux_2243_nl, mux_2240_nl, fsm_output[6]);
  assign nand_421_nl = ~((fsm_output[2]) & mux_2244_nl);
  assign or_2725_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | not_tmp_522;
  assign mux_2235_nl = MUX_s_1_2_2(or_tmp_2611, or_2725_nl, fsm_output[0]);
  assign or_2722_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2234_nl = MUX_s_1_2_2(or_tmp_2607, or_2722_nl, fsm_output[0]);
  assign mux_2236_nl = MUX_s_1_2_2(mux_2235_nl, mux_2234_nl, fsm_output[4]);
  assign or_2719_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2232_nl = MUX_s_1_2_2(or_tmp_2605, or_2719_nl, fsm_output[0]);
  assign or_2716_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2231_nl = MUX_s_1_2_2(or_tmp_2601, or_2716_nl, fsm_output[0]);
  assign mux_2233_nl = MUX_s_1_2_2(mux_2232_nl, mux_2231_nl, fsm_output[4]);
  assign mux_2237_nl = MUX_s_1_2_2(mux_2236_nl, mux_2233_nl, fsm_output[6]);
  assign or_4094_nl = (fsm_output[2]) | mux_2237_nl;
  assign mux_2245_nl = MUX_s_1_2_2(nand_421_nl, or_4094_nl, fsm_output[5]);
  assign vec_rsc_0_48_i_we_d_pff = ~(mux_2245_nl | (fsm_output[1]));
  assign or_2758_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2757_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2258_nl = MUX_s_1_2_2(or_2758_nl, or_2757_nl, fsm_output[0]);
  assign or_2759_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2258_nl;
  assign or_2755_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000)
      | not_tmp_522;
  assign mux_2255_nl = MUX_s_1_2_2(or_2755_nl, or_tmp_2611, fsm_output[0]);
  assign or_2753_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2254_nl = MUX_s_1_2_2(or_2753_nl, or_tmp_2607, fsm_output[0]);
  assign mux_2256_nl = MUX_s_1_2_2(mux_2255_nl, mux_2254_nl, fsm_output[4]);
  assign or_2752_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2252_nl = MUX_s_1_2_2(or_2752_nl, or_tmp_2605, fsm_output[0]);
  assign or_2750_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2251_nl = MUX_s_1_2_2(or_2750_nl, or_tmp_2601, fsm_output[0]);
  assign mux_2253_nl = MUX_s_1_2_2(mux_2252_nl, mux_2251_nl, fsm_output[4]);
  assign mux_2257_nl = MUX_s_1_2_2(mux_2256_nl, mux_2253_nl, fsm_output[6]);
  assign mux_2259_nl = MUX_s_1_2_2(or_2759_nl, mux_2257_nl, fsm_output[2]);
  assign or_2748_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2746_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0000) | not_tmp_527;
  assign mux_2248_nl = MUX_s_1_2_2(or_2748_nl, or_2746_nl, fsm_output[0]);
  assign or_2744_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2743_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2247_nl = MUX_s_1_2_2(or_2744_nl, or_2743_nl, fsm_output[0]);
  assign mux_2249_nl = MUX_s_1_2_2(mux_2248_nl, mux_2247_nl, fsm_output[4]);
  assign nor_896_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_897_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2246_nl = MUX_s_1_2_2(nor_896_nl, nor_897_nl, fsm_output[0]);
  assign nand_111_nl = ~((fsm_output[4]) & mux_2246_nl);
  assign mux_2250_nl = MUX_s_1_2_2(mux_2249_nl, nand_111_nl, fsm_output[6]);
  assign or_2749_nl = (fsm_output[2]) | mux_2250_nl;
  assign mux_2260_nl = MUX_s_1_2_2(mux_2259_nl, or_2749_nl, fsm_output[5]);
  assign vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2260_nl) & (fsm_output[1]);
  assign nor_887_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0001) | not_tmp_523);
  assign nor_888_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_2272_nl = MUX_s_1_2_2(nor_887_nl, nor_888_nl, fsm_output[0]);
  assign nor_889_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_890_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2271_nl = MUX_s_1_2_2(nor_889_nl, nor_890_nl, fsm_output[0]);
  assign mux_2273_nl = MUX_s_1_2_2(mux_2272_nl, mux_2271_nl, fsm_output[4]);
  assign nor_891_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_892_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2269_nl = MUX_s_1_2_2(nor_891_nl, nor_892_nl, fsm_output[0]);
  assign nor_893_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_894_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11000) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2268_nl = MUX_s_1_2_2(nor_893_nl, nor_894_nl, fsm_output[0]);
  assign mux_2270_nl = MUX_s_1_2_2(mux_2269_nl, mux_2268_nl, fsm_output[4]);
  assign mux_2274_nl = MUX_s_1_2_2(mux_2273_nl, mux_2270_nl, fsm_output[6]);
  assign nand_420_nl = ~((fsm_output[2]) & mux_2274_nl);
  assign or_2769_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | not_tmp_522;
  assign mux_2265_nl = MUX_s_1_2_2(or_tmp_2655, or_2769_nl, fsm_output[0]);
  assign or_2766_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2264_nl = MUX_s_1_2_2(or_tmp_2651, or_2766_nl, fsm_output[0]);
  assign mux_2266_nl = MUX_s_1_2_2(mux_2265_nl, mux_2264_nl, fsm_output[4]);
  assign or_2763_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2262_nl = MUX_s_1_2_2(or_tmp_2649, or_2763_nl, fsm_output[0]);
  assign or_2760_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2261_nl = MUX_s_1_2_2(or_tmp_2645, or_2760_nl, fsm_output[0]);
  assign mux_2263_nl = MUX_s_1_2_2(mux_2262_nl, mux_2261_nl, fsm_output[4]);
  assign mux_2267_nl = MUX_s_1_2_2(mux_2266_nl, mux_2263_nl, fsm_output[6]);
  assign or_4093_nl = (fsm_output[2]) | mux_2267_nl;
  assign mux_2275_nl = MUX_s_1_2_2(nand_420_nl, or_4093_nl, fsm_output[5]);
  assign vec_rsc_0_49_i_we_d_pff = ~(mux_2275_nl | (fsm_output[1]));
  assign or_2802_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2801_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2288_nl = MUX_s_1_2_2(or_2802_nl, or_2801_nl, fsm_output[0]);
  assign or_2803_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2288_nl;
  assign or_2799_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001)
      | not_tmp_522;
  assign mux_2285_nl = MUX_s_1_2_2(or_2799_nl, or_tmp_2655, fsm_output[0]);
  assign or_2797_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2284_nl = MUX_s_1_2_2(or_2797_nl, or_tmp_2651, fsm_output[0]);
  assign mux_2286_nl = MUX_s_1_2_2(mux_2285_nl, mux_2284_nl, fsm_output[4]);
  assign or_2796_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2282_nl = MUX_s_1_2_2(or_2796_nl, or_tmp_2649, fsm_output[0]);
  assign or_2794_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2281_nl = MUX_s_1_2_2(or_2794_nl, or_tmp_2645, fsm_output[0]);
  assign mux_2283_nl = MUX_s_1_2_2(mux_2282_nl, mux_2281_nl, fsm_output[4]);
  assign mux_2287_nl = MUX_s_1_2_2(mux_2286_nl, mux_2283_nl, fsm_output[6]);
  assign mux_2289_nl = MUX_s_1_2_2(or_2803_nl, mux_2287_nl, fsm_output[2]);
  assign or_2792_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11000) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2790_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0001) | not_tmp_527;
  assign mux_2278_nl = MUX_s_1_2_2(or_2792_nl, or_2790_nl, fsm_output[0]);
  assign or_2788_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11000) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2787_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2277_nl = MUX_s_1_2_2(or_2788_nl, or_2787_nl, fsm_output[0]);
  assign mux_2279_nl = MUX_s_1_2_2(mux_2278_nl, mux_2277_nl, fsm_output[4]);
  assign nor_885_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_886_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2276_nl = MUX_s_1_2_2(nor_885_nl, nor_886_nl, fsm_output[0]);
  assign nand_113_nl = ~((fsm_output[4]) & mux_2276_nl);
  assign mux_2280_nl = MUX_s_1_2_2(mux_2279_nl, nand_113_nl, fsm_output[6]);
  assign or_2793_nl = (fsm_output[2]) | mux_2280_nl;
  assign mux_2290_nl = MUX_s_1_2_2(mux_2289_nl, or_2793_nl, fsm_output[5]);
  assign vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2290_nl) & (fsm_output[1]);
  assign nor_876_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0010) | not_tmp_523);
  assign nor_877_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10)
      | (~ and_763_cse));
  assign mux_2302_nl = MUX_s_1_2_2(nor_876_nl, nor_877_nl, fsm_output[0]);
  assign nor_878_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_879_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2301_nl = MUX_s_1_2_2(nor_878_nl, nor_879_nl, fsm_output[0]);
  assign mux_2303_nl = MUX_s_1_2_2(mux_2302_nl, mux_2301_nl, fsm_output[4]);
  assign nor_880_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_881_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2299_nl = MUX_s_1_2_2(nor_880_nl, nor_881_nl, fsm_output[0]);
  assign nor_882_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_883_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11001) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2298_nl = MUX_s_1_2_2(nor_882_nl, nor_883_nl, fsm_output[0]);
  assign mux_2300_nl = MUX_s_1_2_2(mux_2299_nl, mux_2298_nl, fsm_output[4]);
  assign mux_2304_nl = MUX_s_1_2_2(mux_2303_nl, mux_2300_nl, fsm_output[6]);
  assign nand_419_nl = ~((fsm_output[2]) & mux_2304_nl);
  assign or_2813_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | not_tmp_522;
  assign mux_2295_nl = MUX_s_1_2_2(or_tmp_2699, or_2813_nl, fsm_output[0]);
  assign or_2810_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2294_nl = MUX_s_1_2_2(or_tmp_2695, or_2810_nl, fsm_output[0]);
  assign mux_2296_nl = MUX_s_1_2_2(mux_2295_nl, mux_2294_nl, fsm_output[4]);
  assign or_2807_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2292_nl = MUX_s_1_2_2(or_tmp_2693, or_2807_nl, fsm_output[0]);
  assign or_2804_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2291_nl = MUX_s_1_2_2(or_tmp_2689, or_2804_nl, fsm_output[0]);
  assign mux_2293_nl = MUX_s_1_2_2(mux_2292_nl, mux_2291_nl, fsm_output[4]);
  assign mux_2297_nl = MUX_s_1_2_2(mux_2296_nl, mux_2293_nl, fsm_output[6]);
  assign or_4092_nl = (fsm_output[2]) | mux_2297_nl;
  assign mux_2305_nl = MUX_s_1_2_2(nand_419_nl, or_4092_nl, fsm_output[5]);
  assign vec_rsc_0_50_i_we_d_pff = ~(mux_2305_nl | (fsm_output[1]));
  assign or_2846_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2845_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2318_nl = MUX_s_1_2_2(or_2846_nl, or_2845_nl, fsm_output[0]);
  assign or_2847_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2318_nl;
  assign or_2843_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010)
      | not_tmp_522;
  assign mux_2315_nl = MUX_s_1_2_2(or_2843_nl, or_tmp_2699, fsm_output[0]);
  assign or_2841_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2314_nl = MUX_s_1_2_2(or_2841_nl, or_tmp_2695, fsm_output[0]);
  assign mux_2316_nl = MUX_s_1_2_2(mux_2315_nl, mux_2314_nl, fsm_output[4]);
  assign or_2840_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2312_nl = MUX_s_1_2_2(or_2840_nl, or_tmp_2693, fsm_output[0]);
  assign or_2838_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2311_nl = MUX_s_1_2_2(or_2838_nl, or_tmp_2689, fsm_output[0]);
  assign mux_2313_nl = MUX_s_1_2_2(mux_2312_nl, mux_2311_nl, fsm_output[4]);
  assign mux_2317_nl = MUX_s_1_2_2(mux_2316_nl, mux_2313_nl, fsm_output[6]);
  assign mux_2319_nl = MUX_s_1_2_2(or_2847_nl, mux_2317_nl, fsm_output[2]);
  assign or_2836_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2834_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0010) | not_tmp_527;
  assign mux_2308_nl = MUX_s_1_2_2(or_2836_nl, or_2834_nl, fsm_output[0]);
  assign or_2832_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2831_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2307_nl = MUX_s_1_2_2(or_2832_nl, or_2831_nl, fsm_output[0]);
  assign mux_2309_nl = MUX_s_1_2_2(mux_2308_nl, mux_2307_nl, fsm_output[4]);
  assign nor_874_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_875_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2306_nl = MUX_s_1_2_2(nor_874_nl, nor_875_nl, fsm_output[0]);
  assign nand_115_nl = ~((fsm_output[4]) & mux_2306_nl);
  assign mux_2310_nl = MUX_s_1_2_2(mux_2309_nl, nand_115_nl, fsm_output[6]);
  assign or_2837_nl = (fsm_output[2]) | mux_2310_nl;
  assign mux_2320_nl = MUX_s_1_2_2(mux_2319_nl, or_2837_nl, fsm_output[5]);
  assign vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2320_nl) & (fsm_output[1]);
  assign nor_865_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0011) | not_tmp_523);
  assign nor_866_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | not_tmp_330);
  assign mux_2332_nl = MUX_s_1_2_2(nor_865_nl, nor_866_nl, fsm_output[0]);
  assign nor_867_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110011) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_868_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2331_nl = MUX_s_1_2_2(nor_867_nl, nor_868_nl, fsm_output[0]);
  assign mux_2333_nl = MUX_s_1_2_2(mux_2332_nl, mux_2331_nl, fsm_output[4]);
  assign nor_869_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_870_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2329_nl = MUX_s_1_2_2(nor_869_nl, nor_870_nl, fsm_output[0]);
  assign nor_871_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_872_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11001) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2328_nl = MUX_s_1_2_2(nor_871_nl, nor_872_nl, fsm_output[0]);
  assign mux_2330_nl = MUX_s_1_2_2(mux_2329_nl, mux_2328_nl, fsm_output[4]);
  assign mux_2334_nl = MUX_s_1_2_2(mux_2333_nl, mux_2330_nl, fsm_output[6]);
  assign nand_418_nl = ~((fsm_output[2]) & mux_2334_nl);
  assign or_2857_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | not_tmp_522;
  assign mux_2325_nl = MUX_s_1_2_2(or_tmp_2743, or_2857_nl, fsm_output[0]);
  assign or_2854_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2324_nl = MUX_s_1_2_2(or_tmp_2739, or_2854_nl, fsm_output[0]);
  assign mux_2326_nl = MUX_s_1_2_2(mux_2325_nl, mux_2324_nl, fsm_output[4]);
  assign or_2851_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2322_nl = MUX_s_1_2_2(or_tmp_2737, or_2851_nl, fsm_output[0]);
  assign or_2848_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2321_nl = MUX_s_1_2_2(or_tmp_2733, or_2848_nl, fsm_output[0]);
  assign mux_2323_nl = MUX_s_1_2_2(mux_2322_nl, mux_2321_nl, fsm_output[4]);
  assign mux_2327_nl = MUX_s_1_2_2(mux_2326_nl, mux_2323_nl, fsm_output[6]);
  assign or_4091_nl = (fsm_output[2]) | mux_2327_nl;
  assign mux_2335_nl = MUX_s_1_2_2(nand_418_nl, or_4091_nl, fsm_output[5]);
  assign vec_rsc_0_51_i_we_d_pff = ~(mux_2335_nl | (fsm_output[1]));
  assign or_2890_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2889_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2348_nl = MUX_s_1_2_2(or_2890_nl, or_2889_nl, fsm_output[0]);
  assign or_2891_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2348_nl;
  assign or_2887_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011)
      | not_tmp_522;
  assign mux_2345_nl = MUX_s_1_2_2(or_2887_nl, or_tmp_2743, fsm_output[0]);
  assign or_2885_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110011)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2344_nl = MUX_s_1_2_2(or_2885_nl, or_tmp_2739, fsm_output[0]);
  assign mux_2346_nl = MUX_s_1_2_2(mux_2345_nl, mux_2344_nl, fsm_output[4]);
  assign or_2884_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110011)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2342_nl = MUX_s_1_2_2(or_2884_nl, or_tmp_2737, fsm_output[0]);
  assign or_2882_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2341_nl = MUX_s_1_2_2(or_2882_nl, or_tmp_2733, fsm_output[0]);
  assign mux_2343_nl = MUX_s_1_2_2(mux_2342_nl, mux_2341_nl, fsm_output[4]);
  assign mux_2347_nl = MUX_s_1_2_2(mux_2346_nl, mux_2343_nl, fsm_output[6]);
  assign mux_2349_nl = MUX_s_1_2_2(or_2891_nl, mux_2347_nl, fsm_output[2]);
  assign or_2880_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11001) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2878_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b0011) | not_tmp_527;
  assign mux_2338_nl = MUX_s_1_2_2(or_2880_nl, or_2878_nl, fsm_output[0]);
  assign or_2876_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11001) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2875_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110011) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2337_nl = MUX_s_1_2_2(or_2876_nl, or_2875_nl, fsm_output[0]);
  assign mux_2339_nl = MUX_s_1_2_2(mux_2338_nl, mux_2337_nl, fsm_output[4]);
  assign nor_863_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1100) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_864_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2336_nl = MUX_s_1_2_2(nor_863_nl, nor_864_nl, fsm_output[0]);
  assign nand_117_nl = ~((fsm_output[4]) & mux_2336_nl);
  assign mux_2340_nl = MUX_s_1_2_2(mux_2339_nl, nand_117_nl, fsm_output[6]);
  assign or_2881_nl = (fsm_output[2]) | mux_2340_nl;
  assign mux_2350_nl = MUX_s_1_2_2(mux_2349_nl, or_2881_nl, fsm_output[5]);
  assign vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2350_nl) & (fsm_output[1]);
  assign nor_854_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0100) | not_tmp_523);
  assign nor_855_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1101) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_2362_nl = MUX_s_1_2_2(nor_854_nl, nor_855_nl, fsm_output[0]);
  assign nor_856_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_857_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2361_nl = MUX_s_1_2_2(nor_856_nl, nor_857_nl, fsm_output[0]);
  assign mux_2363_nl = MUX_s_1_2_2(mux_2362_nl, mux_2361_nl, fsm_output[4]);
  assign nor_858_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_859_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2359_nl = MUX_s_1_2_2(nor_858_nl, nor_859_nl, fsm_output[0]);
  assign nor_860_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_861_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11010) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2358_nl = MUX_s_1_2_2(nor_860_nl, nor_861_nl, fsm_output[0]);
  assign mux_2360_nl = MUX_s_1_2_2(mux_2359_nl, mux_2358_nl, fsm_output[4]);
  assign mux_2364_nl = MUX_s_1_2_2(mux_2363_nl, mux_2360_nl, fsm_output[6]);
  assign nand_417_nl = ~((fsm_output[2]) & mux_2364_nl);
  assign or_2901_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | not_tmp_522;
  assign mux_2355_nl = MUX_s_1_2_2(or_tmp_2787, or_2901_nl, fsm_output[0]);
  assign or_2898_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2354_nl = MUX_s_1_2_2(or_tmp_2783, or_2898_nl, fsm_output[0]);
  assign mux_2356_nl = MUX_s_1_2_2(mux_2355_nl, mux_2354_nl, fsm_output[4]);
  assign or_2895_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2352_nl = MUX_s_1_2_2(or_tmp_2781, or_2895_nl, fsm_output[0]);
  assign or_2892_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2351_nl = MUX_s_1_2_2(or_tmp_2777, or_2892_nl, fsm_output[0]);
  assign mux_2353_nl = MUX_s_1_2_2(mux_2352_nl, mux_2351_nl, fsm_output[4]);
  assign mux_2357_nl = MUX_s_1_2_2(mux_2356_nl, mux_2353_nl, fsm_output[6]);
  assign or_4090_nl = (fsm_output[2]) | mux_2357_nl;
  assign mux_2365_nl = MUX_s_1_2_2(nand_417_nl, or_4090_nl, fsm_output[5]);
  assign vec_rsc_0_52_i_we_d_pff = ~(mux_2365_nl | (fsm_output[1]));
  assign or_2934_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2933_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2378_nl = MUX_s_1_2_2(or_2934_nl, or_2933_nl, fsm_output[0]);
  assign or_2935_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2378_nl;
  assign or_2931_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100)
      | not_tmp_522;
  assign mux_2375_nl = MUX_s_1_2_2(or_2931_nl, or_tmp_2787, fsm_output[0]);
  assign or_2929_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2374_nl = MUX_s_1_2_2(or_2929_nl, or_tmp_2783, fsm_output[0]);
  assign mux_2376_nl = MUX_s_1_2_2(mux_2375_nl, mux_2374_nl, fsm_output[4]);
  assign or_2928_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2372_nl = MUX_s_1_2_2(or_2928_nl, or_tmp_2781, fsm_output[0]);
  assign or_2926_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2371_nl = MUX_s_1_2_2(or_2926_nl, or_tmp_2777, fsm_output[0]);
  assign mux_2373_nl = MUX_s_1_2_2(mux_2372_nl, mux_2371_nl, fsm_output[4]);
  assign mux_2377_nl = MUX_s_1_2_2(mux_2376_nl, mux_2373_nl, fsm_output[6]);
  assign mux_2379_nl = MUX_s_1_2_2(or_2935_nl, mux_2377_nl, fsm_output[2]);
  assign or_2924_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_2922_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | not_tmp_544;
  assign mux_2368_nl = MUX_s_1_2_2(or_2924_nl, or_2922_nl, fsm_output[0]);
  assign or_2920_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2919_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2367_nl = MUX_s_1_2_2(or_2920_nl, or_2919_nl, fsm_output[0]);
  assign mux_2369_nl = MUX_s_1_2_2(mux_2368_nl, mux_2367_nl, fsm_output[4]);
  assign nor_852_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_853_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2366_nl = MUX_s_1_2_2(nor_852_nl, nor_853_nl, fsm_output[0]);
  assign nand_119_nl = ~((fsm_output[4]) & mux_2366_nl);
  assign mux_2370_nl = MUX_s_1_2_2(mux_2369_nl, nand_119_nl, fsm_output[6]);
  assign or_2925_nl = (fsm_output[2]) | mux_2370_nl;
  assign mux_2380_nl = MUX_s_1_2_2(mux_2379_nl, or_2925_nl, fsm_output[5]);
  assign vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2380_nl) & (fsm_output[1]);
  assign nor_843_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0101) | not_tmp_523);
  assign nor_844_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1101) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_2392_nl = MUX_s_1_2_2(nor_843_nl, nor_844_nl, fsm_output[0]);
  assign nor_845_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110101) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_846_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2391_nl = MUX_s_1_2_2(nor_845_nl, nor_846_nl, fsm_output[0]);
  assign mux_2393_nl = MUX_s_1_2_2(mux_2392_nl, mux_2391_nl, fsm_output[4]);
  assign nor_847_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_848_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2389_nl = MUX_s_1_2_2(nor_847_nl, nor_848_nl, fsm_output[0]);
  assign nor_849_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_850_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11010) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2388_nl = MUX_s_1_2_2(nor_849_nl, nor_850_nl, fsm_output[0]);
  assign mux_2390_nl = MUX_s_1_2_2(mux_2389_nl, mux_2388_nl, fsm_output[4]);
  assign mux_2394_nl = MUX_s_1_2_2(mux_2393_nl, mux_2390_nl, fsm_output[6]);
  assign nand_416_nl = ~((fsm_output[2]) & mux_2394_nl);
  assign or_2945_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | not_tmp_522;
  assign mux_2385_nl = MUX_s_1_2_2(or_tmp_2831, or_2945_nl, fsm_output[0]);
  assign or_2942_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2384_nl = MUX_s_1_2_2(or_tmp_2827, or_2942_nl, fsm_output[0]);
  assign mux_2386_nl = MUX_s_1_2_2(mux_2385_nl, mux_2384_nl, fsm_output[4]);
  assign or_2939_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2382_nl = MUX_s_1_2_2(or_tmp_2825, or_2939_nl, fsm_output[0]);
  assign or_2936_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2381_nl = MUX_s_1_2_2(or_tmp_2821, or_2936_nl, fsm_output[0]);
  assign mux_2383_nl = MUX_s_1_2_2(mux_2382_nl, mux_2381_nl, fsm_output[4]);
  assign mux_2387_nl = MUX_s_1_2_2(mux_2386_nl, mux_2383_nl, fsm_output[6]);
  assign or_4089_nl = (fsm_output[2]) | mux_2387_nl;
  assign mux_2395_nl = MUX_s_1_2_2(nand_416_nl, or_4089_nl, fsm_output[5]);
  assign vec_rsc_0_53_i_we_d_pff = ~(mux_2395_nl | (fsm_output[1]));
  assign or_2978_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_2977_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2408_nl = MUX_s_1_2_2(or_2978_nl, or_2977_nl, fsm_output[0]);
  assign or_2979_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2408_nl;
  assign or_2975_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101)
      | not_tmp_522;
  assign mux_2405_nl = MUX_s_1_2_2(or_2975_nl, or_tmp_2831, fsm_output[0]);
  assign or_2973_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110101)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2404_nl = MUX_s_1_2_2(or_2973_nl, or_tmp_2827, fsm_output[0]);
  assign mux_2406_nl = MUX_s_1_2_2(mux_2405_nl, mux_2404_nl, fsm_output[4]);
  assign or_2972_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110101)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2402_nl = MUX_s_1_2_2(or_2972_nl, or_tmp_2825, fsm_output[0]);
  assign or_2970_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2401_nl = MUX_s_1_2_2(or_2970_nl, or_tmp_2821, fsm_output[0]);
  assign mux_2403_nl = MUX_s_1_2_2(mux_2402_nl, mux_2401_nl, fsm_output[4]);
  assign mux_2407_nl = MUX_s_1_2_2(mux_2406_nl, mux_2403_nl, fsm_output[6]);
  assign mux_2409_nl = MUX_s_1_2_2(or_2979_nl, mux_2407_nl, fsm_output[2]);
  assign or_2968_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11010) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_2966_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | not_tmp_549;
  assign mux_2398_nl = MUX_s_1_2_2(or_2968_nl, or_2966_nl, fsm_output[0]);
  assign or_2964_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11010) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_2963_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110101) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2397_nl = MUX_s_1_2_2(or_2964_nl, or_2963_nl, fsm_output[0]);
  assign mux_2399_nl = MUX_s_1_2_2(mux_2398_nl, mux_2397_nl, fsm_output[4]);
  assign nor_841_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_842_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2396_nl = MUX_s_1_2_2(nor_841_nl, nor_842_nl, fsm_output[0]);
  assign nand_121_nl = ~((fsm_output[4]) & mux_2396_nl);
  assign mux_2400_nl = MUX_s_1_2_2(mux_2399_nl, nand_121_nl, fsm_output[6]);
  assign or_2969_nl = (fsm_output[2]) | mux_2400_nl;
  assign mux_2410_nl = MUX_s_1_2_2(mux_2409_nl, or_2969_nl, fsm_output[5]);
  assign vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2410_nl) & (fsm_output[1]);
  assign nor_833_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]!=4'b0110) | not_tmp_523);
  assign and_567_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1101) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b10)
      & and_763_cse;
  assign mux_2422_nl = MUX_s_1_2_2(nor_833_nl, and_567_nl, fsm_output[0]);
  assign nor_834_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b110110) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_835_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2421_nl = MUX_s_1_2_2(nor_834_nl, nor_835_nl, fsm_output[0]);
  assign mux_2423_nl = MUX_s_1_2_2(mux_2422_nl, mux_2421_nl, fsm_output[4]);
  assign nor_836_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_837_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2419_nl = MUX_s_1_2_2(nor_836_nl, nor_837_nl, fsm_output[0]);
  assign nor_838_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_839_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11011) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2418_nl = MUX_s_1_2_2(nor_838_nl, nor_839_nl, fsm_output[0]);
  assign mux_2420_nl = MUX_s_1_2_2(mux_2419_nl, mux_2418_nl, fsm_output[4]);
  assign mux_2424_nl = MUX_s_1_2_2(mux_2423_nl, mux_2420_nl, fsm_output[6]);
  assign nand_415_nl = ~((fsm_output[2]) & mux_2424_nl);
  assign or_2989_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | not_tmp_522;
  assign mux_2415_nl = MUX_s_1_2_2(or_tmp_2875, or_2989_nl, fsm_output[0]);
  assign or_2986_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2414_nl = MUX_s_1_2_2(or_tmp_2871, or_2986_nl, fsm_output[0]);
  assign mux_2416_nl = MUX_s_1_2_2(mux_2415_nl, mux_2414_nl, fsm_output[4]);
  assign or_2983_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2412_nl = MUX_s_1_2_2(or_tmp_2869, or_2983_nl, fsm_output[0]);
  assign or_2980_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2411_nl = MUX_s_1_2_2(or_tmp_2865, or_2980_nl, fsm_output[0]);
  assign mux_2413_nl = MUX_s_1_2_2(mux_2412_nl, mux_2411_nl, fsm_output[4]);
  assign mux_2417_nl = MUX_s_1_2_2(mux_2416_nl, mux_2413_nl, fsm_output[6]);
  assign or_4088_nl = (fsm_output[2]) | mux_2417_nl;
  assign mux_2425_nl = MUX_s_1_2_2(nand_415_nl, or_4088_nl, fsm_output[5]);
  assign vec_rsc_0_54_i_we_d_pff = ~(mux_2425_nl | (fsm_output[1]));
  assign or_3022_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3021_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2438_nl = MUX_s_1_2_2(or_3022_nl, or_3021_nl, fsm_output[0]);
  assign or_3023_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2438_nl;
  assign or_3019_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110)
      | not_tmp_522;
  assign mux_2435_nl = MUX_s_1_2_2(or_3019_nl, or_tmp_2875, fsm_output[0]);
  assign or_3017_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b110110)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2434_nl = MUX_s_1_2_2(or_3017_nl, or_tmp_2871, fsm_output[0]);
  assign mux_2436_nl = MUX_s_1_2_2(mux_2435_nl, mux_2434_nl, fsm_output[4]);
  assign or_3016_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b110110)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2432_nl = MUX_s_1_2_2(or_3016_nl, or_tmp_2869, fsm_output[0]);
  assign or_3014_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2431_nl = MUX_s_1_2_2(or_3014_nl, or_tmp_2865, fsm_output[0]);
  assign mux_2433_nl = MUX_s_1_2_2(mux_2432_nl, mux_2431_nl, fsm_output[4]);
  assign mux_2437_nl = MUX_s_1_2_2(mux_2436_nl, mux_2433_nl, fsm_output[6]);
  assign mux_2439_nl = MUX_s_1_2_2(or_3023_nl, mux_2437_nl, fsm_output[2]);
  assign nand_271_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11011) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & and_763_cse);
  assign or_3010_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | not_tmp_544;
  assign mux_2428_nl = MUX_s_1_2_2(nand_271_nl, or_3010_nl, fsm_output[0]);
  assign or_3008_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11011) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_3007_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110110) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2427_nl = MUX_s_1_2_2(or_3008_nl, or_3007_nl, fsm_output[0]);
  assign mux_2429_nl = MUX_s_1_2_2(mux_2428_nl, mux_2427_nl, fsm_output[4]);
  assign nor_831_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_832_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2426_nl = MUX_s_1_2_2(nor_831_nl, nor_832_nl, fsm_output[0]);
  assign nand_123_nl = ~((fsm_output[4]) & mux_2426_nl);
  assign mux_2430_nl = MUX_s_1_2_2(mux_2429_nl, nand_123_nl, fsm_output[6]);
  assign or_3013_nl = (fsm_output[2]) | mux_2430_nl;
  assign mux_2440_nl = MUX_s_1_2_2(mux_2439_nl, or_3013_nl, fsm_output[5]);
  assign vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2440_nl) & (fsm_output[1]);
  assign nor_824_nl = ~((~((COMP_LOOP_acc_10_cse_10_1_5_sva[3:0]==4'b0111))) | not_tmp_523);
  assign nor_825_nl = ~((~ (COMP_LOOP_acc_13_psp_sva[3])) | (COMP_LOOP_acc_13_psp_sva[1])
      | not_tmp_414);
  assign mux_2452_nl = MUX_s_1_2_2(nor_824_nl, nor_825_nl, fsm_output[0]);
  assign and_564_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b110111) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_565_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b110) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_2451_nl = MUX_s_1_2_2(and_564_nl, and_565_nl, fsm_output[0]);
  assign mux_2453_nl = MUX_s_1_2_2(mux_2452_nl, mux_2451_nl, fsm_output[4]);
  assign and_813_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b110111) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_820_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b11011) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_2449_nl = MUX_s_1_2_2(and_813_nl, and_820_nl, fsm_output[0]);
  assign nor_828_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b110111) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_829_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11011) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2448_nl = MUX_s_1_2_2(nor_828_nl, nor_829_nl, fsm_output[0]);
  assign mux_2450_nl = MUX_s_1_2_2(mux_2449_nl, mux_2448_nl, fsm_output[4]);
  assign mux_2454_nl = MUX_s_1_2_2(mux_2453_nl, mux_2450_nl, fsm_output[6]);
  assign nand_414_nl = ~((fsm_output[2]) & mux_2454_nl);
  assign or_3033_nl = (~((COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0111))) | not_tmp_522;
  assign mux_2445_nl = MUX_s_1_2_2(or_tmp_2919, or_3033_nl, fsm_output[0]);
  assign nand_267_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b110111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2444_nl = MUX_s_1_2_2(or_tmp_2915, nand_267_nl, fsm_output[0]);
  assign mux_2446_nl = MUX_s_1_2_2(mux_2445_nl, mux_2444_nl, fsm_output[4]);
  assign nand_476_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b110111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_2442_nl = MUX_s_1_2_2(or_tmp_2913, nand_476_nl, fsm_output[0]);
  assign or_3024_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110111) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2441_nl = MUX_s_1_2_2(or_tmp_2909, or_3024_nl, fsm_output[0]);
  assign mux_2443_nl = MUX_s_1_2_2(mux_2442_nl, mux_2441_nl, fsm_output[4]);
  assign mux_2447_nl = MUX_s_1_2_2(mux_2446_nl, mux_2443_nl, fsm_output[6]);
  assign or_4087_nl = (fsm_output[2]) | mux_2447_nl;
  assign mux_2455_nl = MUX_s_1_2_2(nand_414_nl, or_4087_nl, fsm_output[5]);
  assign vec_rsc_0_55_i_we_d_pff = ~(mux_2455_nl | (fsm_output[1]));
  assign or_3066_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b110111) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3065_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2468_nl = MUX_s_1_2_2(or_3066_nl, or_3065_nl, fsm_output[0]);
  assign or_3067_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2468_nl;
  assign or_3063_nl = (~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b0111)))
      | not_tmp_522;
  assign mux_2465_nl = MUX_s_1_2_2(or_3063_nl, or_tmp_2919, fsm_output[0]);
  assign nand_258_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b110111)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_2464_nl = MUX_s_1_2_2(nand_258_nl, or_tmp_2915, fsm_output[0]);
  assign mux_2466_nl = MUX_s_1_2_2(mux_2465_nl, mux_2464_nl, fsm_output[4]);
  assign nand_400_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b110111)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_2462_nl = MUX_s_1_2_2(nand_400_nl, or_tmp_2913, fsm_output[0]);
  assign or_3058_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b110111)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2461_nl = MUX_s_1_2_2(or_3058_nl, or_tmp_2909, fsm_output[0]);
  assign mux_2463_nl = MUX_s_1_2_2(mux_2462_nl, mux_2461_nl, fsm_output[4]);
  assign mux_2467_nl = MUX_s_1_2_2(mux_2466_nl, mux_2463_nl, fsm_output[6]);
  assign mux_2469_nl = MUX_s_1_2_2(or_3067_nl, mux_2467_nl, fsm_output[2]);
  assign or_3056_nl = (~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11011) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm))
      | not_tmp_321;
  assign or_3054_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      | not_tmp_549;
  assign mux_2458_nl = MUX_s_1_2_2(or_3056_nl, or_3054_nl, fsm_output[0]);
  assign nand_261_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b11011) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_262_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b110111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2457_nl = MUX_s_1_2_2(nand_261_nl, nand_262_nl, fsm_output[0]);
  assign mux_2459_nl = MUX_s_1_2_2(mux_2458_nl, mux_2457_nl, fsm_output[4]);
  assign nor_822_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1101) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_823_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b110111) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2456_nl = MUX_s_1_2_2(nor_822_nl, nor_823_nl, fsm_output[0]);
  assign nand_125_nl = ~((fsm_output[4]) & mux_2456_nl);
  assign mux_2460_nl = MUX_s_1_2_2(mux_2459_nl, nand_125_nl, fsm_output[6]);
  assign or_3057_nl = (fsm_output[2]) | mux_2460_nl;
  assign mux_2470_nl = MUX_s_1_2_2(mux_2469_nl, or_3057_nl, fsm_output[5]);
  assign vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2470_nl) & (fsm_output[1]);
  assign nor_813_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[2:0]!=3'b000) | not_tmp_560);
  assign nor_814_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1110) | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)
      | (~ and_763_cse));
  assign mux_2482_nl = MUX_s_1_2_2(nor_813_nl, nor_814_nl, fsm_output[0]);
  assign nor_815_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b111000) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_816_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2481_nl = MUX_s_1_2_2(nor_815_nl, nor_816_nl, fsm_output[0]);
  assign mux_2483_nl = MUX_s_1_2_2(mux_2482_nl, mux_2481_nl, fsm_output[4]);
  assign nor_817_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_818_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2479_nl = MUX_s_1_2_2(nor_817_nl, nor_818_nl, fsm_output[0]);
  assign nor_819_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_820_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11100) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2478_nl = MUX_s_1_2_2(nor_819_nl, nor_820_nl, fsm_output[0]);
  assign mux_2480_nl = MUX_s_1_2_2(mux_2479_nl, mux_2478_nl, fsm_output[4]);
  assign mux_2484_nl = MUX_s_1_2_2(mux_2483_nl, mux_2480_nl, fsm_output[6]);
  assign nand_413_nl = ~((fsm_output[2]) & mux_2484_nl);
  assign or_3077_nl = (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000) | not_tmp_559;
  assign mux_2475_nl = MUX_s_1_2_2(or_tmp_2963, or_3077_nl, fsm_output[0]);
  assign or_3074_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2474_nl = MUX_s_1_2_2(or_tmp_2959, or_3074_nl, fsm_output[0]);
  assign mux_2476_nl = MUX_s_1_2_2(mux_2475_nl, mux_2474_nl, fsm_output[4]);
  assign or_3071_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2472_nl = MUX_s_1_2_2(or_tmp_2957, or_3071_nl, fsm_output[0]);
  assign or_3068_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2471_nl = MUX_s_1_2_2(or_tmp_2953, or_3068_nl, fsm_output[0]);
  assign mux_2473_nl = MUX_s_1_2_2(mux_2472_nl, mux_2471_nl, fsm_output[4]);
  assign mux_2477_nl = MUX_s_1_2_2(mux_2476_nl, mux_2473_nl, fsm_output[6]);
  assign or_4086_nl = (fsm_output[2]) | mux_2477_nl;
  assign mux_2485_nl = MUX_s_1_2_2(nand_413_nl, or_4086_nl, fsm_output[5]);
  assign vec_rsc_0_56_i_we_d_pff = ~(mux_2485_nl | (fsm_output[1]));
  assign or_3110_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111000) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3109_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2498_nl = MUX_s_1_2_2(or_3110_nl, or_3109_nl, fsm_output[0]);
  assign or_3111_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2498_nl;
  assign or_3107_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b000)
      | not_tmp_559;
  assign mux_2495_nl = MUX_s_1_2_2(or_3107_nl, or_tmp_2963, fsm_output[0]);
  assign or_3105_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111000)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2494_nl = MUX_s_1_2_2(or_3105_nl, or_tmp_2959, fsm_output[0]);
  assign mux_2496_nl = MUX_s_1_2_2(mux_2495_nl, mux_2494_nl, fsm_output[4]);
  assign or_3104_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111000)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2492_nl = MUX_s_1_2_2(or_3104_nl, or_tmp_2957, fsm_output[0]);
  assign or_3102_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111000)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2491_nl = MUX_s_1_2_2(or_3102_nl, or_tmp_2953, fsm_output[0]);
  assign mux_2493_nl = MUX_s_1_2_2(mux_2492_nl, mux_2491_nl, fsm_output[4]);
  assign mux_2497_nl = MUX_s_1_2_2(mux_2496_nl, mux_2493_nl, fsm_output[6]);
  assign mux_2499_nl = MUX_s_1_2_2(or_3111_nl, mux_2497_nl, fsm_output[2]);
  assign or_3100_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ and_763_cse);
  assign or_3098_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1000) | not_tmp_527;
  assign mux_2488_nl = MUX_s_1_2_2(or_3100_nl, or_3098_nl, fsm_output[0]);
  assign or_3096_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_3095_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111000) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2487_nl = MUX_s_1_2_2(or_3096_nl, or_3095_nl, fsm_output[0]);
  assign mux_2489_nl = MUX_s_1_2_2(mux_2488_nl, mux_2487_nl, fsm_output[4]);
  assign nor_811_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_812_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111000) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2486_nl = MUX_s_1_2_2(nor_811_nl, nor_812_nl, fsm_output[0]);
  assign nand_127_nl = ~((fsm_output[4]) & mux_2486_nl);
  assign mux_2490_nl = MUX_s_1_2_2(mux_2489_nl, nand_127_nl, fsm_output[6]);
  assign or_3101_nl = (fsm_output[2]) | mux_2490_nl;
  assign mux_2500_nl = MUX_s_1_2_2(mux_2499_nl, or_3101_nl, fsm_output[5]);
  assign vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2500_nl) & (fsm_output[1]);
  assign nor_802_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[2:0]!=3'b001) | not_tmp_560);
  assign nor_803_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1110) | (VEC_LOOP_j_10_0_sva_9_0[1])
      | not_tmp_321);
  assign mux_2512_nl = MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output[0]);
  assign nor_804_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b111001) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_805_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2511_nl = MUX_s_1_2_2(nor_804_nl, nor_805_nl, fsm_output[0]);
  assign mux_2513_nl = MUX_s_1_2_2(mux_2512_nl, mux_2511_nl, fsm_output[4]);
  assign nor_806_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_807_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2509_nl = MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output[0]);
  assign nor_808_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_809_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11100) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2508_nl = MUX_s_1_2_2(nor_808_nl, nor_809_nl, fsm_output[0]);
  assign mux_2510_nl = MUX_s_1_2_2(mux_2509_nl, mux_2508_nl, fsm_output[4]);
  assign mux_2514_nl = MUX_s_1_2_2(mux_2513_nl, mux_2510_nl, fsm_output[6]);
  assign nand_412_nl = ~((fsm_output[2]) & mux_2514_nl);
  assign or_3121_nl = (COMP_LOOP_acc_1_cse_6_sva[2:1]!=2'b00) | not_tmp_565;
  assign mux_2505_nl = MUX_s_1_2_2(or_tmp_3007, or_3121_nl, fsm_output[0]);
  assign or_3118_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2504_nl = MUX_s_1_2_2(or_tmp_3003, or_3118_nl, fsm_output[0]);
  assign mux_2506_nl = MUX_s_1_2_2(mux_2505_nl, mux_2504_nl, fsm_output[4]);
  assign or_3115_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2502_nl = MUX_s_1_2_2(or_tmp_3001, or_3115_nl, fsm_output[0]);
  assign or_3112_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2501_nl = MUX_s_1_2_2(or_tmp_2997, or_3112_nl, fsm_output[0]);
  assign mux_2503_nl = MUX_s_1_2_2(mux_2502_nl, mux_2501_nl, fsm_output[4]);
  assign mux_2507_nl = MUX_s_1_2_2(mux_2506_nl, mux_2503_nl, fsm_output[6]);
  assign or_4085_nl = (fsm_output[2]) | mux_2507_nl;
  assign mux_2515_nl = MUX_s_1_2_2(nand_412_nl, or_4085_nl, fsm_output[5]);
  assign vec_rsc_0_57_i_we_d_pff = ~(mux_2515_nl | (fsm_output[1]));
  assign or_3154_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111001) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3153_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2528_nl = MUX_s_1_2_2(or_3154_nl, or_3153_nl, fsm_output[0]);
  assign or_3155_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2528_nl;
  assign or_3151_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:1]!=2'b00)
      | not_tmp_565;
  assign mux_2525_nl = MUX_s_1_2_2(or_3151_nl, or_tmp_3007, fsm_output[0]);
  assign or_3149_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111001)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2524_nl = MUX_s_1_2_2(or_3149_nl, or_tmp_3003, fsm_output[0]);
  assign mux_2526_nl = MUX_s_1_2_2(mux_2525_nl, mux_2524_nl, fsm_output[4]);
  assign or_3148_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111001)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2522_nl = MUX_s_1_2_2(or_3148_nl, or_tmp_3001, fsm_output[0]);
  assign or_3146_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111001)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2521_nl = MUX_s_1_2_2(or_3146_nl, or_tmp_2997, fsm_output[0]);
  assign mux_2523_nl = MUX_s_1_2_2(mux_2522_nl, mux_2521_nl, fsm_output[4]);
  assign mux_2527_nl = MUX_s_1_2_2(mux_2526_nl, mux_2523_nl, fsm_output[6]);
  assign mux_2529_nl = MUX_s_1_2_2(or_3155_nl, mux_2527_nl, fsm_output[2]);
  assign or_3144_nl = (COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11100) | (~ COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm)
      | not_tmp_321;
  assign or_3142_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1001) | not_tmp_527;
  assign mux_2518_nl = MUX_s_1_2_2(or_3144_nl, or_3142_nl, fsm_output[0]);
  assign or_3140_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11100) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (~ (VEC_LOOP_j_10_0_sva_9_0[0])) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_3139_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111001) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2517_nl = MUX_s_1_2_2(or_3140_nl, or_3139_nl, fsm_output[0]);
  assign mux_2519_nl = MUX_s_1_2_2(mux_2518_nl, mux_2517_nl, fsm_output[4]);
  assign nor_800_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_801_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111001) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2516_nl = MUX_s_1_2_2(nor_800_nl, nor_801_nl, fsm_output[0]);
  assign nand_129_nl = ~((fsm_output[4]) & mux_2516_nl);
  assign mux_2520_nl = MUX_s_1_2_2(mux_2519_nl, nand_129_nl, fsm_output[6]);
  assign or_3145_nl = (fsm_output[2]) | mux_2520_nl;
  assign mux_2530_nl = MUX_s_1_2_2(mux_2529_nl, or_3145_nl, fsm_output[5]);
  assign vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2530_nl) & (fsm_output[1]);
  assign nor_792_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | not_tmp_570);
  assign and_560_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1110) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b10)
      & and_763_cse;
  assign mux_2542_nl = MUX_s_1_2_2(nor_792_nl, and_560_nl, fsm_output[0]);
  assign nor_793_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b111010) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_794_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2541_nl = MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output[0]);
  assign mux_2543_nl = MUX_s_1_2_2(mux_2542_nl, mux_2541_nl, fsm_output[4]);
  assign nor_795_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_796_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2539_nl = MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output[0]);
  assign nor_797_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_798_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11101) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2538_nl = MUX_s_1_2_2(nor_797_nl, nor_798_nl, fsm_output[0]);
  assign mux_2540_nl = MUX_s_1_2_2(mux_2539_nl, mux_2538_nl, fsm_output[4]);
  assign mux_2544_nl = MUX_s_1_2_2(mux_2543_nl, mux_2540_nl, fsm_output[6]);
  assign nand_411_nl = ~((fsm_output[2]) & mux_2544_nl);
  assign or_3165_nl = (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010) | not_tmp_559;
  assign mux_2535_nl = MUX_s_1_2_2(or_tmp_3051, or_3165_nl, fsm_output[0]);
  assign or_3162_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2534_nl = MUX_s_1_2_2(or_tmp_3047, or_3162_nl, fsm_output[0]);
  assign mux_2536_nl = MUX_s_1_2_2(mux_2535_nl, mux_2534_nl, fsm_output[4]);
  assign or_3159_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2532_nl = MUX_s_1_2_2(or_tmp_3045, or_3159_nl, fsm_output[0]);
  assign or_3156_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2531_nl = MUX_s_1_2_2(or_tmp_3041, or_3156_nl, fsm_output[0]);
  assign mux_2533_nl = MUX_s_1_2_2(mux_2532_nl, mux_2531_nl, fsm_output[4]);
  assign mux_2537_nl = MUX_s_1_2_2(mux_2536_nl, mux_2533_nl, fsm_output[6]);
  assign or_4084_nl = (fsm_output[2]) | mux_2537_nl;
  assign mux_2545_nl = MUX_s_1_2_2(nand_411_nl, or_4084_nl, fsm_output[5]);
  assign vec_rsc_0_58_i_we_d_pff = ~(mux_2545_nl | (fsm_output[1]));
  assign or_3198_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111010) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3197_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2558_nl = MUX_s_1_2_2(or_3198_nl, or_3197_nl, fsm_output[0]);
  assign or_3199_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2558_nl;
  assign or_3195_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b010)
      | not_tmp_559;
  assign mux_2555_nl = MUX_s_1_2_2(or_3195_nl, or_tmp_3051, fsm_output[0]);
  assign or_3193_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111010)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2554_nl = MUX_s_1_2_2(or_3193_nl, or_tmp_3047, fsm_output[0]);
  assign mux_2556_nl = MUX_s_1_2_2(mux_2555_nl, mux_2554_nl, fsm_output[4]);
  assign or_3192_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111010)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2552_nl = MUX_s_1_2_2(or_3192_nl, or_tmp_3045, fsm_output[0]);
  assign or_3190_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111010)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2551_nl = MUX_s_1_2_2(or_3190_nl, or_tmp_3041, fsm_output[0]);
  assign mux_2553_nl = MUX_s_1_2_2(mux_2552_nl, mux_2551_nl, fsm_output[4]);
  assign mux_2557_nl = MUX_s_1_2_2(mux_2556_nl, mux_2553_nl, fsm_output[6]);
  assign mux_2559_nl = MUX_s_1_2_2(or_3199_nl, mux_2557_nl, fsm_output[2]);
  assign nand_252_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11101) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & and_763_cse);
  assign or_3186_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]!=4'b1010) | not_tmp_527;
  assign mux_2548_nl = MUX_s_1_2_2(nand_252_nl, or_3186_nl, fsm_output[0]);
  assign or_3184_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11101) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_3183_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111010) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2547_nl = MUX_s_1_2_2(or_3184_nl, or_3183_nl, fsm_output[0]);
  assign mux_2549_nl = MUX_s_1_2_2(mux_2548_nl, mux_2547_nl, fsm_output[4]);
  assign nor_790_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_791_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111010) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2546_nl = MUX_s_1_2_2(nor_790_nl, nor_791_nl, fsm_output[0]);
  assign nand_131_nl = ~((fsm_output[4]) & mux_2546_nl);
  assign mux_2550_nl = MUX_s_1_2_2(mux_2549_nl, nand_131_nl, fsm_output[6]);
  assign or_3189_nl = (fsm_output[2]) | mux_2550_nl;
  assign mux_2560_nl = MUX_s_1_2_2(mux_2559_nl, or_3189_nl, fsm_output[5]);
  assign vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2560_nl) & (fsm_output[1]);
  assign nor_783_nl = ~((~ (COMP_LOOP_acc_10_cse_10_1_5_sva[0])) | (COMP_LOOP_acc_10_cse_10_1_5_sva[2])
      | not_tmp_570);
  assign nor_784_nl = ~((~((COMP_LOOP_acc_13_psp_sva[3:0]==4'b1110))) | not_tmp_330);
  assign mux_2572_nl = MUX_s_1_2_2(nor_783_nl, nor_784_nl, fsm_output[0]);
  assign and_557_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b111011) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_558_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b011)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_2571_nl = MUX_s_1_2_2(and_557_nl, and_558_nl, fsm_output[0]);
  assign mux_2573_nl = MUX_s_1_2_2(mux_2572_nl, mux_2571_nl, fsm_output[4]);
  assign and_814_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b111011) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_821_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b11101) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_2569_nl = MUX_s_1_2_2(and_814_nl, and_821_nl, fsm_output[0]);
  assign nor_787_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111011) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_788_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11101) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2568_nl = MUX_s_1_2_2(nor_787_nl, nor_788_nl, fsm_output[0]);
  assign mux_2570_nl = MUX_s_1_2_2(mux_2569_nl, mux_2568_nl, fsm_output[4]);
  assign mux_2574_nl = MUX_s_1_2_2(mux_2573_nl, mux_2570_nl, fsm_output[6]);
  assign nand_410_nl = ~((fsm_output[2]) & mux_2574_nl);
  assign or_3208_nl = (COMP_LOOP_acc_1_cse_6_sva[2]) | not_tmp_575;
  assign mux_2565_nl = MUX_s_1_2_2(or_tmp_3094, or_3208_nl, fsm_output[0]);
  assign nand_247_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111011) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2564_nl = MUX_s_1_2_2(or_tmp_3091, nand_247_nl, fsm_output[0]);
  assign mux_2566_nl = MUX_s_1_2_2(mux_2565_nl, mux_2564_nl, fsm_output[4]);
  assign nand_475_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b111011) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_2562_nl = MUX_s_1_2_2(or_tmp_3089, nand_475_nl, fsm_output[0]);
  assign or_3200_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111011) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2561_nl = MUX_s_1_2_2(or_tmp_3085, or_3200_nl, fsm_output[0]);
  assign mux_2563_nl = MUX_s_1_2_2(mux_2562_nl, mux_2561_nl, fsm_output[4]);
  assign mux_2567_nl = MUX_s_1_2_2(mux_2566_nl, mux_2563_nl, fsm_output[6]);
  assign or_4083_nl = (fsm_output[2]) | mux_2567_nl;
  assign mux_2575_nl = MUX_s_1_2_2(nand_410_nl, or_4083_nl, fsm_output[5]);
  assign vec_rsc_0_59_i_we_d_pff = ~(mux_2575_nl | (fsm_output[1]));
  assign or_3241_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111011) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3240_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2588_nl = MUX_s_1_2_2(or_3241_nl, or_3240_nl, fsm_output[0]);
  assign or_3242_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2588_nl;
  assign or_3238_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[2])
      | not_tmp_575;
  assign mux_2585_nl = MUX_s_1_2_2(or_3238_nl, or_tmp_3094, fsm_output[0]);
  assign nand_238_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111011)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_2584_nl = MUX_s_1_2_2(nand_238_nl, or_tmp_3091, fsm_output[0]);
  assign mux_2586_nl = MUX_s_1_2_2(mux_2585_nl, mux_2584_nl, fsm_output[4]);
  assign nand_398_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b111011)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_2582_nl = MUX_s_1_2_2(nand_398_nl, or_tmp_3089, fsm_output[0]);
  assign or_3233_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111011)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2581_nl = MUX_s_1_2_2(or_3233_nl, or_tmp_3085, fsm_output[0]);
  assign mux_2583_nl = MUX_s_1_2_2(mux_2582_nl, mux_2581_nl, fsm_output[4]);
  assign mux_2587_nl = MUX_s_1_2_2(mux_2586_nl, mux_2583_nl, fsm_output[6]);
  assign mux_2589_nl = MUX_s_1_2_2(or_3242_nl, mux_2587_nl, fsm_output[2]);
  assign or_3231_nl = (~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11101) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm))
      | not_tmp_321;
  assign or_3229_nl = (~((COMP_LOOP_acc_10_cse_10_1_7_sva[3:0]==4'b1011))) | not_tmp_527;
  assign mux_2578_nl = MUX_s_1_2_2(or_3231_nl, or_3229_nl, fsm_output[0]);
  assign nand_242_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b11101) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_243_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b111011) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2577_nl = MUX_s_1_2_2(nand_242_nl, nand_243_nl, fsm_output[0]);
  assign mux_2579_nl = MUX_s_1_2_2(mux_2578_nl, mux_2577_nl, fsm_output[4]);
  assign nor_781_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1110) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b11) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_782_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111011) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2576_nl = MUX_s_1_2_2(nor_781_nl, nor_782_nl, fsm_output[0]);
  assign nand_133_nl = ~((fsm_output[4]) & mux_2576_nl);
  assign mux_2580_nl = MUX_s_1_2_2(mux_2579_nl, nand_133_nl, fsm_output[6]);
  assign or_3232_nl = (fsm_output[2]) | mux_2580_nl;
  assign mux_2590_nl = MUX_s_1_2_2(mux_2589_nl, or_3232_nl, fsm_output[5]);
  assign vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2590_nl) & (fsm_output[1]);
  assign nor_773_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[2:0]!=3'b100) | not_tmp_560);
  assign and_555_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1111) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b00)
      & and_763_cse;
  assign mux_2602_nl = MUX_s_1_2_2(nor_773_nl, and_555_nl, fsm_output[0]);
  assign nor_774_nl = ~((COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]!=6'b111100) | (~ (fsm_output[3]))
      | (fsm_output[7]));
  assign nor_775_nl = ~((COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (~ (fsm_output[3])) | (fsm_output[7]));
  assign mux_2601_nl = MUX_s_1_2_2(nor_774_nl, nor_775_nl, fsm_output[0]);
  assign mux_2603_nl = MUX_s_1_2_2(mux_2602_nl, mux_2601_nl, fsm_output[4]);
  assign nor_776_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (~ (fsm_output[7])));
  assign nor_777_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]!=5'b11110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (~ (fsm_output[7])));
  assign mux_2599_nl = MUX_s_1_2_2(nor_776_nl, nor_777_nl, fsm_output[0]);
  assign nor_778_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_779_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11110) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2598_nl = MUX_s_1_2_2(nor_778_nl, nor_779_nl, fsm_output[0]);
  assign mux_2600_nl = MUX_s_1_2_2(mux_2599_nl, mux_2598_nl, fsm_output[4]);
  assign mux_2604_nl = MUX_s_1_2_2(mux_2603_nl, mux_2600_nl, fsm_output[6]);
  assign nand_409_nl = ~((fsm_output[2]) & mux_2604_nl);
  assign or_3252_nl = (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100) | not_tmp_559;
  assign mux_2595_nl = MUX_s_1_2_2(or_tmp_3138, or_3252_nl, fsm_output[0]);
  assign or_3249_nl = (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2594_nl = MUX_s_1_2_2(or_tmp_3134, or_3249_nl, fsm_output[0]);
  assign mux_2596_nl = MUX_s_1_2_2(mux_2595_nl, mux_2594_nl, fsm_output[4]);
  assign or_3246_nl = (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (~ (fsm_output[7]));
  assign mux_2592_nl = MUX_s_1_2_2(or_tmp_3132, or_3246_nl, fsm_output[0]);
  assign or_3243_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2591_nl = MUX_s_1_2_2(or_tmp_3128, or_3243_nl, fsm_output[0]);
  assign mux_2593_nl = MUX_s_1_2_2(mux_2592_nl, mux_2591_nl, fsm_output[4]);
  assign mux_2597_nl = MUX_s_1_2_2(mux_2596_nl, mux_2593_nl, fsm_output[6]);
  assign or_4082_nl = (fsm_output[2]) | mux_2597_nl;
  assign mux_2605_nl = MUX_s_1_2_2(nand_409_nl, or_4082_nl, fsm_output[5]);
  assign vec_rsc_0_60_i_we_d_pff = ~(mux_2605_nl | (fsm_output[1]));
  assign or_3285_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111100) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3284_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2618_nl = MUX_s_1_2_2(or_3285_nl, or_3284_nl, fsm_output[0]);
  assign or_3286_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2618_nl;
  assign or_3282_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b100)
      | not_tmp_559;
  assign mux_2615_nl = MUX_s_1_2_2(or_3282_nl, or_tmp_3138, fsm_output[0]);
  assign or_3280_nl = (~ COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_2_sva[5:0]!=6'b111100)
      | (~ (fsm_output[3])) | (fsm_output[7]);
  assign mux_2614_nl = MUX_s_1_2_2(or_3280_nl, or_tmp_3134, fsm_output[0]);
  assign mux_2616_nl = MUX_s_1_2_2(mux_2615_nl, mux_2614_nl, fsm_output[4]);
  assign or_3279_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm) | (COMP_LOOP_acc_1_cse_sva[5:0]!=6'b111100)
      | (fsm_output[3]) | (~ (fsm_output[7]));
  assign mux_2612_nl = MUX_s_1_2_2(or_3279_nl, or_tmp_3132, fsm_output[0]);
  assign or_3277_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111100)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2611_nl = MUX_s_1_2_2(or_3277_nl, or_tmp_3128, fsm_output[0]);
  assign mux_2613_nl = MUX_s_1_2_2(mux_2612_nl, mux_2611_nl, fsm_output[4]);
  assign mux_2617_nl = MUX_s_1_2_2(mux_2616_nl, mux_2613_nl, fsm_output[6]);
  assign mux_2619_nl = MUX_s_1_2_2(or_3286_nl, mux_2617_nl, fsm_output[2]);
  assign nand_237_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11110) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & and_763_cse);
  assign or_3273_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | not_tmp_544;
  assign mux_2608_nl = MUX_s_1_2_2(nand_237_nl, or_3273_nl, fsm_output[0]);
  assign or_3271_nl = (COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11110) | (~ COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[0]) | (~ (fsm_output[3])) | (fsm_output[7]);
  assign or_3270_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111100) | (~ (fsm_output[3]))
      | (fsm_output[7]);
  assign mux_2607_nl = MUX_s_1_2_2(or_3271_nl, or_3270_nl, fsm_output[0]);
  assign mux_2609_nl = MUX_s_1_2_2(mux_2608_nl, mux_2607_nl, fsm_output[4]);
  assign nor_771_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_772_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111100) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2606_nl = MUX_s_1_2_2(nor_771_nl, nor_772_nl, fsm_output[0]);
  assign nand_135_nl = ~((fsm_output[4]) & mux_2606_nl);
  assign mux_2610_nl = MUX_s_1_2_2(mux_2609_nl, nand_135_nl, fsm_output[6]);
  assign or_3276_nl = (fsm_output[2]) | mux_2610_nl;
  assign mux_2620_nl = MUX_s_1_2_2(mux_2619_nl, or_3276_nl, fsm_output[5]);
  assign vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2620_nl) & (fsm_output[1]);
  assign nor_764_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[2:0]!=3'b101) | not_tmp_560);
  assign nor_765_nl = ~((~((COMP_LOOP_acc_13_psp_sva[3:0]==4'b1111) & (~ (VEC_LOOP_j_10_0_sva_9_0[1]))))
      | not_tmp_321);
  assign mux_2632_nl = MUX_s_1_2_2(nor_764_nl, nor_765_nl, fsm_output[0]);
  assign and_552_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b111101) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_553_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b101)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_2631_nl = MUX_s_1_2_2(and_552_nl, and_553_nl, fsm_output[0]);
  assign mux_2633_nl = MUX_s_1_2_2(mux_2632_nl, mux_2631_nl, fsm_output[4]);
  assign and_815_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b111101) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_822_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b11110) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_2629_nl = MUX_s_1_2_2(and_815_nl, and_822_nl, fsm_output[0]);
  assign nor_768_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111101) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_769_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11110) | (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2628_nl = MUX_s_1_2_2(nor_768_nl, nor_769_nl, fsm_output[0]);
  assign mux_2630_nl = MUX_s_1_2_2(mux_2629_nl, mux_2628_nl, fsm_output[4]);
  assign mux_2634_nl = MUX_s_1_2_2(mux_2633_nl, mux_2630_nl, fsm_output[6]);
  assign nand_408_nl = ~((fsm_output[2]) & mux_2634_nl);
  assign or_3296_nl = (COMP_LOOP_acc_1_cse_6_sva[2:1]!=2'b10) | not_tmp_565;
  assign mux_2625_nl = MUX_s_1_2_2(or_tmp_3182, or_3296_nl, fsm_output[0]);
  assign nand_232_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111101) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2624_nl = MUX_s_1_2_2(or_tmp_3178, nand_232_nl, fsm_output[0]);
  assign mux_2626_nl = MUX_s_1_2_2(mux_2625_nl, mux_2624_nl, fsm_output[4]);
  assign nand_474_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b111101) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_2622_nl = MUX_s_1_2_2(or_tmp_3176, nand_474_nl, fsm_output[0]);
  assign or_3287_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111101) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2621_nl = MUX_s_1_2_2(or_tmp_3172, or_3287_nl, fsm_output[0]);
  assign mux_2623_nl = MUX_s_1_2_2(mux_2622_nl, mux_2621_nl, fsm_output[4]);
  assign mux_2627_nl = MUX_s_1_2_2(mux_2626_nl, mux_2623_nl, fsm_output[6]);
  assign or_4081_nl = (fsm_output[2]) | mux_2627_nl;
  assign mux_2635_nl = MUX_s_1_2_2(nand_408_nl, or_4081_nl, fsm_output[5]);
  assign vec_rsc_0_61_i_we_d_pff = ~(mux_2635_nl | (fsm_output[1]));
  assign or_3328_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111101) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3327_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2648_nl = MUX_s_1_2_2(or_3328_nl, or_3327_nl, fsm_output[0]);
  assign or_3329_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2648_nl;
  assign or_3325_nl = (~ COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm) | (COMP_LOOP_acc_1_cse_6_sva[2:1]!=2'b10)
      | not_tmp_565;
  assign mux_2645_nl = MUX_s_1_2_2(or_3325_nl, or_tmp_3182, fsm_output[0]);
  assign nand_223_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111101)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_2644_nl = MUX_s_1_2_2(nand_223_nl, or_tmp_3178, fsm_output[0]);
  assign mux_2646_nl = MUX_s_1_2_2(mux_2645_nl, mux_2644_nl, fsm_output[4]);
  assign nand_396_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b111101)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_2642_nl = MUX_s_1_2_2(nand_396_nl, or_tmp_3176, fsm_output[0]);
  assign or_3320_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111101)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2641_nl = MUX_s_1_2_2(or_3320_nl, or_tmp_3172, fsm_output[0]);
  assign mux_2643_nl = MUX_s_1_2_2(mux_2642_nl, mux_2641_nl, fsm_output[4]);
  assign mux_2647_nl = MUX_s_1_2_2(mux_2646_nl, mux_2643_nl, fsm_output[6]);
  assign mux_2649_nl = MUX_s_1_2_2(or_3329_nl, mux_2647_nl, fsm_output[2]);
  assign or_3318_nl = (~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11110) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm))
      | not_tmp_321;
  assign or_3316_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) | (~((COMP_LOOP_acc_10_cse_10_1_7_sva[3])
      & (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[2])
      & (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) & (COMP_LOOP_acc_10_cse_10_1_7_sva[4])
      & (fsm_output[3]) & (fsm_output[7])));
  assign mux_2638_nl = MUX_s_1_2_2(or_3318_nl, or_3316_nl, fsm_output[0]);
  assign nand_227_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b11110) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_228_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b111101) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2637_nl = MUX_s_1_2_2(nand_227_nl, nand_228_nl, fsm_output[0]);
  assign mux_2639_nl = MUX_s_1_2_2(mux_2638_nl, mux_2637_nl, fsm_output[4]);
  assign nor_762_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b01) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_763_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111101) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2636_nl = MUX_s_1_2_2(nor_762_nl, nor_763_nl, fsm_output[0]);
  assign nand_137_nl = ~((fsm_output[4]) & mux_2636_nl);
  assign mux_2640_nl = MUX_s_1_2_2(mux_2639_nl, nand_137_nl, fsm_output[6]);
  assign or_3319_nl = (fsm_output[2]) | mux_2640_nl;
  assign mux_2650_nl = MUX_s_1_2_2(mux_2649_nl, or_3319_nl, fsm_output[5]);
  assign vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2650_nl) & (fsm_output[1]);
  assign nor_756_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[0]) | (~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:1]==5'b11111)
      & (fsm_output[3]) & (fsm_output[7]))));
  assign and_548_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1111) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b10)
      & and_763_cse;
  assign mux_2662_nl = MUX_s_1_2_2(nor_756_nl, and_548_nl, fsm_output[0]);
  assign and_549_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b111110) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_550_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b110)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_2661_nl = MUX_s_1_2_2(and_549_nl, and_550_nl, fsm_output[0]);
  assign mux_2663_nl = MUX_s_1_2_2(mux_2662_nl, mux_2661_nl, fsm_output[4]);
  assign and_816_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b111110) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_823_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b11111) & (~ (VEC_LOOP_j_10_0_sva_9_0[0]))
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_2659_nl = MUX_s_1_2_2(and_816_nl, and_823_nl, fsm_output[0]);
  assign nor_759_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]!=6'b111110) | (fsm_output[3])
      | (fsm_output[7]));
  assign nor_760_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]!=5'b11111) | (VEC_LOOP_j_10_0_sva_9_0[0])
      | (fsm_output[3]) | (fsm_output[7]));
  assign mux_2658_nl = MUX_s_1_2_2(nor_759_nl, nor_760_nl, fsm_output[0]);
  assign mux_2660_nl = MUX_s_1_2_2(mux_2659_nl, mux_2658_nl, fsm_output[4]);
  assign mux_2664_nl = MUX_s_1_2_2(mux_2663_nl, mux_2660_nl, fsm_output[6]);
  assign nand_407_nl = ~((fsm_output[2]) & mux_2664_nl);
  assign or_3339_nl = (COMP_LOOP_acc_1_cse_6_sva[2:0]!=3'b110) | not_tmp_559;
  assign mux_2655_nl = MUX_s_1_2_2(or_tmp_3225, or_3339_nl, fsm_output[0]);
  assign nand_218_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111110) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2654_nl = MUX_s_1_2_2(or_tmp_3221, nand_218_nl, fsm_output[0]);
  assign mux_2656_nl = MUX_s_1_2_2(mux_2655_nl, mux_2654_nl, fsm_output[4]);
  assign nand_473_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b111110) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_2652_nl = MUX_s_1_2_2(or_tmp_3219, nand_473_nl, fsm_output[0]);
  assign or_3330_nl = (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111110) | (fsm_output[3])
      | (fsm_output[7]);
  assign mux_2651_nl = MUX_s_1_2_2(or_tmp_3215, or_3330_nl, fsm_output[0]);
  assign mux_2653_nl = MUX_s_1_2_2(mux_2652_nl, mux_2651_nl, fsm_output[4]);
  assign mux_2657_nl = MUX_s_1_2_2(mux_2656_nl, mux_2653_nl, fsm_output[6]);
  assign or_4080_nl = (fsm_output[2]) | mux_2657_nl;
  assign mux_2665_nl = MUX_s_1_2_2(nand_407_nl, or_4080_nl, fsm_output[5]);
  assign vec_rsc_0_62_i_we_d_pff = ~(mux_2665_nl | (fsm_output[1]));
  assign or_3371_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b111110) | (fsm_output[3])
      | (fsm_output[7]);
  assign or_3370_nl = (COMP_LOOP_acc_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2678_nl = MUX_s_1_2_2(or_3371_nl, or_3370_nl, fsm_output[0]);
  assign or_3372_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2678_nl;
  assign or_3368_nl = (~(COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_6_sva[2:0]==3'b110)))
      | not_tmp_559;
  assign mux_2675_nl = MUX_s_1_2_2(or_3368_nl, or_tmp_3225, fsm_output[0]);
  assign nand_210_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111110)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_2674_nl = MUX_s_1_2_2(nand_210_nl, or_tmp_3221, fsm_output[0]);
  assign mux_2676_nl = MUX_s_1_2_2(mux_2675_nl, mux_2674_nl, fsm_output[4]);
  assign nand_394_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b111110)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_2672_nl = MUX_s_1_2_2(nand_394_nl, or_tmp_3219, fsm_output[0]);
  assign or_3363_nl = (~ COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm) | (COMP_LOOP_acc_1_cse_4_sva[5:0]!=6'b111110)
      | (fsm_output[3]) | (fsm_output[7]);
  assign mux_2671_nl = MUX_s_1_2_2(or_3363_nl, or_tmp_3215, fsm_output[0]);
  assign mux_2673_nl = MUX_s_1_2_2(mux_2672_nl, mux_2671_nl, fsm_output[4]);
  assign mux_2677_nl = MUX_s_1_2_2(mux_2676_nl, mux_2673_nl, fsm_output[6]);
  assign mux_2679_nl = MUX_s_1_2_2(or_3372_nl, mux_2677_nl, fsm_output[2]);
  assign nand_212_nl = ~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & and_763_cse);
  assign or_3359_nl = (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[1])) | (~ (COMP_LOOP_acc_10_cse_10_1_7_sva[3]))
      | (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) | not_tmp_544;
  assign mux_2668_nl = MUX_s_1_2_2(nand_212_nl, or_3359_nl, fsm_output[0]);
  assign nand_213_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b11111) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (~ (VEC_LOOP_j_10_0_sva_9_0[0])) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_214_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b111110) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2667_nl = MUX_s_1_2_2(nand_213_nl, nand_214_nl, fsm_output[0]);
  assign mux_2669_nl = MUX_s_1_2_2(mux_2668_nl, mux_2667_nl, fsm_output[4]);
  assign nor_754_nl = ~((COMP_LOOP_acc_13_psp_sva[3:0]!=4'b1111) | (~ COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm)
      | (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b10) | (fsm_output[3]) | (fsm_output[7]));
  assign nor_755_nl = ~((COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]!=6'b111110) | (fsm_output[3])
      | (fsm_output[7]));
  assign mux_2666_nl = MUX_s_1_2_2(nor_754_nl, nor_755_nl, fsm_output[0]);
  assign nand_139_nl = ~((fsm_output[4]) & mux_2666_nl);
  assign mux_2670_nl = MUX_s_1_2_2(mux_2669_nl, nand_139_nl, fsm_output[6]);
  assign or_3362_nl = (fsm_output[2]) | mux_2670_nl;
  assign mux_2680_nl = MUX_s_1_2_2(mux_2679_nl, or_3362_nl, fsm_output[5]);
  assign vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2680_nl) & (fsm_output[1]);
  assign and_539_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b111111) & (fsm_output[3])
      & (fsm_output[7]);
  assign and_540_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1111) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
      & (fsm_output[3]) & (fsm_output[7]);
  assign mux_2692_nl = MUX_s_1_2_2(and_539_nl, and_540_nl, fsm_output[0]);
  assign and_541_nl = (COMP_LOOP_acc_10_cse_10_1_1_sva[5:0]==6'b111111) & (fsm_output[3])
      & (~ (fsm_output[7]));
  assign and_542_nl = (COMP_LOOP_acc_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
      & (fsm_output[3]) & (~ (fsm_output[7]));
  assign mux_2691_nl = MUX_s_1_2_2(and_541_nl, and_542_nl, fsm_output[0]);
  assign mux_2693_nl = MUX_s_1_2_2(mux_2692_nl, mux_2691_nl, fsm_output[4]);
  assign and_817_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (fsm_output[7]);
  assign and_824_nl = (COMP_LOOP_acc_14_psp_sva[4:0]==5'b11111) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (fsm_output[7]);
  assign mux_2689_nl = MUX_s_1_2_2(and_817_nl, and_824_nl, fsm_output[0]);
  assign and_543_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (~ (fsm_output[7]));
  assign and_544_nl = (COMP_LOOP_acc_11_psp_sva[4:0]==5'b11111) & (VEC_LOOP_j_10_0_sva_9_0[0])
      & (~ (fsm_output[3])) & (~ (fsm_output[7]));
  assign mux_2688_nl = MUX_s_1_2_2(and_543_nl, and_544_nl, fsm_output[0]);
  assign mux_2690_nl = MUX_s_1_2_2(mux_2689_nl, mux_2688_nl, fsm_output[4]);
  assign mux_2694_nl = MUX_s_1_2_2(mux_2693_nl, mux_2690_nl, fsm_output[6]);
  assign nand_406_nl = ~((fsm_output[2]) & mux_2694_nl);
  assign mux_2685_nl = MUX_s_1_2_2(nor_tmp_307, nor_tmp_306, fsm_output[0]);
  assign nand_203_nl = ~((COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2684_nl = MUX_s_1_2_2(or_tmp_3264, nand_203_nl, fsm_output[0]);
  assign mux_2686_nl = MUX_s_1_2_2((~ mux_2685_nl), mux_2684_nl, fsm_output[4]);
  assign nand_nl = ~((COMP_LOOP_acc_1_cse_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (fsm_output[7]));
  assign mux_2682_nl = MUX_s_1_2_2(or_tmp_3262, nand_nl, fsm_output[0]);
  assign nand_205_nl = ~((COMP_LOOP_acc_1_cse_4_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (~ (fsm_output[7])));
  assign mux_2681_nl = MUX_s_1_2_2(or_tmp_3258, nand_205_nl, fsm_output[0]);
  assign mux_2683_nl = MUX_s_1_2_2(mux_2682_nl, mux_2681_nl, fsm_output[4]);
  assign mux_2687_nl = MUX_s_1_2_2(mux_2686_nl, mux_2683_nl, fsm_output[6]);
  assign or_4079_nl = (fsm_output[2]) | mux_2687_nl;
  assign mux_2695_nl = MUX_s_1_2_2(nand_406_nl, or_4079_nl, fsm_output[5]);
  assign vec_rsc_0_63_i_we_d_pff = ~(mux_2695_nl | (fsm_output[1]));
  assign nand_192_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (~ (fsm_output[7])));
  assign nand_193_nl = ~((COMP_LOOP_acc_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
      & (~ (fsm_output[3])) & (~ (fsm_output[7])));
  assign mux_2708_nl = MUX_s_1_2_2(nand_192_nl, nand_193_nl, fsm_output[0]);
  assign or_3405_nl = (fsm_output[6]) | (fsm_output[4]) | mux_2708_nl;
  assign and_535_nl = COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm & nor_tmp_306;
  assign mux_2705_nl = MUX_s_1_2_2(and_535_nl, nor_tmp_307, fsm_output[0]);
  assign nand_194_nl = ~(COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm & (COMP_LOOP_acc_1_cse_2_sva[5:0]==6'b111111)
      & (fsm_output[3]) & (~ (fsm_output[7])));
  assign mux_2704_nl = MUX_s_1_2_2(nand_194_nl, or_tmp_3264, fsm_output[0]);
  assign mux_2706_nl = MUX_s_1_2_2((~ mux_2705_nl), mux_2704_nl, fsm_output[4]);
  assign nand_392_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm & (COMP_LOOP_acc_1_cse_sva[5:0]==6'b111111)
      & (~ (fsm_output[3])) & (fsm_output[7]));
  assign mux_2702_nl = MUX_s_1_2_2(nand_392_nl, or_tmp_3262, fsm_output[0]);
  assign nand_196_nl = ~(COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm & (COMP_LOOP_acc_1_cse_4_sva[5:0]==6'b111111)
      & (~ (fsm_output[3])) & (~ (fsm_output[7])));
  assign mux_2701_nl = MUX_s_1_2_2(nand_196_nl, or_tmp_3258, fsm_output[0]);
  assign mux_2703_nl = MUX_s_1_2_2(mux_2702_nl, mux_2701_nl, fsm_output[4]);
  assign mux_2707_nl = MUX_s_1_2_2(mux_2706_nl, mux_2703_nl, fsm_output[6]);
  assign mux_2709_nl = MUX_s_1_2_2(or_3405_nl, mux_2707_nl, fsm_output[2]);
  assign or_4002_nl = (~((COMP_LOOP_acc_14_psp_sva[4:0]==5'b11111) & COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm))
      | not_tmp_321;
  assign nand_198_nl = ~((COMP_LOOP_acc_10_cse_10_1_7_sva[5:0]==6'b111111) & (fsm_output[3])
      & (fsm_output[7]));
  assign mux_2698_nl = MUX_s_1_2_2(or_4002_nl, nand_198_nl, fsm_output[0]);
  assign nand_199_nl = ~((COMP_LOOP_acc_11_psp_sva[4:0]==5'b11111) & COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[0]) & (fsm_output[3]) & (~ (fsm_output[7])));
  assign nand_200_nl = ~((COMP_LOOP_acc_10_cse_10_1_3_sva[5:0]==6'b111111) & (fsm_output[3])
      & (~ (fsm_output[7])));
  assign mux_2697_nl = MUX_s_1_2_2(nand_199_nl, nand_200_nl, fsm_output[0]);
  assign mux_2699_nl = MUX_s_1_2_2(mux_2698_nl, mux_2697_nl, fsm_output[4]);
  assign and_536_nl = (COMP_LOOP_acc_13_psp_sva[3:0]==4'b1111) & COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm
      & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (~ (fsm_output[3])) & (~ (fsm_output[7]));
  assign and_537_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:0]==6'b111111) & (~ (fsm_output[3]))
      & (~ (fsm_output[7]));
  assign mux_2696_nl = MUX_s_1_2_2(and_536_nl, and_537_nl, fsm_output[0]);
  assign nand_141_nl = ~((fsm_output[4]) & mux_2696_nl);
  assign mux_2700_nl = MUX_s_1_2_2(mux_2699_nl, nand_141_nl, fsm_output[6]);
  assign or_3396_nl = (fsm_output[2]) | mux_2700_nl;
  assign mux_2710_nl = MUX_s_1_2_2(mux_2709_nl, or_3396_nl, fsm_output[5]);
  assign vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d = (~ mux_2710_nl) & (fsm_output[1]);
  assign twiddle_rsc_0_0_i_radr_d_pff = MUX1HOT_v_4_7_2((z_out_8[6:3]), (z_out_7[9:6]),
      (z_out_7[8:5]), (COMP_LOOP_5_tmp_mul_idiv_sva[7:4]), (COMP_LOOP_2_tmp_mul_idiv_sva[9:6]),
      (COMP_LOOP_3_tmp_lshift_ncse_sva[8:5]), (COMP_LOOP_2_tmp_lshift_ncse_sva[9:6]),
      {and_dcpl_74 , COMP_LOOP_or_110_rgt , and_dcpl_258 , and_dcpl_260 , and_dcpl_261
      , and_dcpl_263 , and_dcpl_265});
  assign nor_746_cse = ~((z_out_7[5:0]!=6'b000000) | (fsm_output[3]));
  assign nor_743_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b00000) | (~ (fsm_output[3])));
  assign nor_744_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b000000) | (~ (fsm_output[3])));
  assign mux_2715_nl = MUX_s_1_2_2(nor_743_nl, nor_744_nl, fsm_output[0]);
  assign nor_745_nl = ~((z_out_8[2:0]!=3'b000) | (fsm_output[3]));
  assign mux_2714_nl = MUX_s_1_2_2(nor_745_nl, nor_746_cse, fsm_output[0]);
  assign mux_2716_nl = MUX_s_1_2_2(mux_2715_nl, mux_2714_nl, fsm_output[1]);
  assign nor_747_nl = ~((z_out_7[4:0]!=5'b00000) | (fsm_output[3]));
  assign mux_2712_nl = MUX_s_1_2_2(nor_747_nl, nor_746_cse, fsm_output[0]);
  assign nor_749_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0000) | (fsm_output[3]));
  assign nor_750_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b000000) | (fsm_output[3]));
  assign mux_2711_nl = MUX_s_1_2_2(nor_749_nl, nor_750_nl, fsm_output[0]);
  assign mux_2713_nl = MUX_s_1_2_2(mux_2712_nl, mux_2711_nl, fsm_output[1]);
  assign mux_2717_nl = MUX_s_1_2_2(mux_2716_nl, mux_2713_nl, fsm_output[2]);
  assign twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2717_nl & and_dcpl_268;
  assign twiddle_rsc_0_1_i_radr_d_pff = z_out_7[9:6];
  assign nor_740_cse = ~((z_out_7[5:0]!=6'b000001) | (fsm_output[3:2]!=2'b01));
  assign nor_739_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b00000) | nand_191_cse);
  assign mux_2719_nl = MUX_s_1_2_2(nor_739_nl, nor_740_cse, fsm_output[0]);
  assign nor_742_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b000001) | (fsm_output[3]));
  assign mux_2718_nl = MUX_s_1_2_2(nor_740_cse, nor_742_nl, fsm_output[0]);
  assign mux_2720_nl = MUX_s_1_2_2(mux_2719_nl, mux_2718_nl, fsm_output[1]);
  assign twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2720_nl & and_dcpl_268;
  assign twiddle_rsc_0_2_i_radr_d_pff = MUX_v_4_2_2((z_out_7[9:6]), (z_out_7[8:5]),
      COMP_LOOP_tmp_or_43_cse);
  assign nor_735_cse = ~((z_out_7[5:0]!=6'b000010) | (fsm_output[3]));
  assign nor_734_cse = ~((z_out_7[4:0]!=5'b00001) | (fsm_output[3]));
  assign nor_733_nl = ~((z_out_7[5:0]!=6'b000010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2723_nl = MUX_s_1_2_2(nor_734_cse, nor_735_cse, fsm_output[0]);
  assign mux_2724_nl = MUX_s_1_2_2(nor_733_nl, mux_2723_nl, fsm_output[2]);
  assign nor_736_nl = ~((z_out_7[5:0]!=6'b000010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2721_nl = MUX_s_1_2_2(nor_735_cse, nor_734_cse, fsm_output[0]);
  assign mux_2722_nl = MUX_s_1_2_2(nor_736_nl, mux_2721_nl, fsm_output[2]);
  assign mux_2725_nl = MUX_s_1_2_2(mux_2724_nl, mux_2722_nl, fsm_output[1]);
  assign twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2725_nl & and_dcpl_268;
  assign nor_730_cse = ~((z_out_7[5:0]!=6'b000011) | (fsm_output[3:2]!=2'b01));
  assign nor_729_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b0000) | nand_190_cse);
  assign mux_2727_nl = MUX_s_1_2_2(nor_729_nl, nor_730_cse, fsm_output[0]);
  assign nor_732_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b000011) | (fsm_output[3]));
  assign mux_2726_nl = MUX_s_1_2_2(nor_730_cse, nor_732_nl, fsm_output[0]);
  assign mux_2728_nl = MUX_s_1_2_2(mux_2727_nl, mux_2726_nl, fsm_output[1]);
  assign twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2728_nl & and_dcpl_268;
  assign twiddle_rsc_0_4_i_radr_d_pff = MUX1HOT_v_4_6_2((z_out_7[9:6]), (z_out_7[8:5]),
      (COMP_LOOP_5_tmp_mul_idiv_sva[7:4]), (COMP_LOOP_2_tmp_mul_idiv_sva[9:6]), (COMP_LOOP_3_tmp_lshift_ncse_sva[8:5]),
      (COMP_LOOP_2_tmp_lshift_ncse_sva[9:6]), {COMP_LOOP_or_110_rgt , and_dcpl_258
      , and_dcpl_260 , and_dcpl_261 , and_dcpl_263 , and_dcpl_265});
  assign nor_722_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b00010) | (~ (fsm_output[3])));
  assign nor_723_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b000100) | (~ (fsm_output[3])));
  assign mux_2732_nl = MUX_s_1_2_2(nor_722_nl, nor_723_nl, fsm_output[0]);
  assign nor_724_nl = ~((z_out_7[4:0]!=5'b00010) | (fsm_output[3]));
  assign nor_725_nl = ~((z_out_7[5:0]!=6'b000100) | (fsm_output[3]));
  assign mux_2731_nl = MUX_s_1_2_2(nor_724_nl, nor_725_nl, fsm_output[0]);
  assign mux_2733_nl = MUX_s_1_2_2(mux_2732_nl, mux_2731_nl, fsm_output[2]);
  assign nor_726_nl = ~((z_out_7[5:0]!=6'b000100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_727_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0001) | (fsm_output[3]));
  assign nor_728_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b000100) | (fsm_output[3]));
  assign mux_2729_nl = MUX_s_1_2_2(nor_727_nl, nor_728_nl, fsm_output[0]);
  assign mux_2730_nl = MUX_s_1_2_2(nor_726_nl, mux_2729_nl, fsm_output[2]);
  assign mux_2734_nl = MUX_s_1_2_2(mux_2733_nl, mux_2730_nl, fsm_output[1]);
  assign twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2734_nl & and_dcpl_268;
  assign nor_719_cse = ~((z_out_7[5:0]!=6'b000101) | (fsm_output[3:2]!=2'b01));
  assign nor_718_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b00010) | nand_191_cse);
  assign mux_2736_nl = MUX_s_1_2_2(nor_718_nl, nor_719_cse, fsm_output[0]);
  assign nor_721_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b000101) | (fsm_output[3]));
  assign mux_2735_nl = MUX_s_1_2_2(nor_719_cse, nor_721_nl, fsm_output[0]);
  assign mux_2737_nl = MUX_s_1_2_2(mux_2736_nl, mux_2735_nl, fsm_output[1]);
  assign twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2737_nl & and_dcpl_268;
  assign nor_714_cse = ~((z_out_7[5:0]!=6'b000110) | (fsm_output[3]));
  assign nor_713_cse = ~((z_out_7[4:0]!=5'b00011) | (fsm_output[3]));
  assign nor_712_nl = ~((z_out_7[5:0]!=6'b000110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2740_nl = MUX_s_1_2_2(nor_713_cse, nor_714_cse, fsm_output[0]);
  assign mux_2741_nl = MUX_s_1_2_2(nor_712_nl, mux_2740_nl, fsm_output[2]);
  assign nor_715_nl = ~((z_out_7[5:0]!=6'b000110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2738_nl = MUX_s_1_2_2(nor_714_cse, nor_713_cse, fsm_output[0]);
  assign mux_2739_nl = MUX_s_1_2_2(nor_715_nl, mux_2738_nl, fsm_output[2]);
  assign mux_2742_nl = MUX_s_1_2_2(mux_2741_nl, mux_2739_nl, fsm_output[1]);
  assign twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2742_nl & and_dcpl_268;
  assign nor_709_cse = ~((z_out_7[5:0]!=6'b000111) | (fsm_output[3:2]!=2'b01));
  assign nor_708_nl = ~((fsm_output[2]) | (z_out_7[5:3]!=3'b000) | nand_188_cse);
  assign mux_2744_nl = MUX_s_1_2_2(nor_708_nl, nor_709_cse, fsm_output[0]);
  assign nor_711_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b000111) | (fsm_output[3]));
  assign mux_2743_nl = MUX_s_1_2_2(nor_709_cse, nor_711_nl, fsm_output[0]);
  assign mux_2745_nl = MUX_s_1_2_2(mux_2744_nl, mux_2743_nl, fsm_output[1]);
  assign twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2745_nl & and_dcpl_268;
  assign nor_703_cse = ~((z_out_7[5:0]!=6'b001000) | (fsm_output[3]));
  assign nor_700_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b00100) | (~ (fsm_output[3])));
  assign nor_701_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b001000) | (~ (fsm_output[3])));
  assign mux_2750_nl = MUX_s_1_2_2(nor_700_nl, nor_701_nl, fsm_output[0]);
  assign nor_702_nl = ~((z_out_8[2:0]!=3'b001) | (fsm_output[3]));
  assign mux_2749_nl = MUX_s_1_2_2(nor_702_nl, nor_703_cse, fsm_output[0]);
  assign mux_2751_nl = MUX_s_1_2_2(mux_2750_nl, mux_2749_nl, fsm_output[1]);
  assign nor_704_nl = ~((z_out_7[4:0]!=5'b00100) | (fsm_output[3]));
  assign mux_2747_nl = MUX_s_1_2_2(nor_704_nl, nor_703_cse, fsm_output[0]);
  assign nor_706_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0010) | (fsm_output[3]));
  assign nor_707_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b001000) | (fsm_output[3]));
  assign mux_2746_nl = MUX_s_1_2_2(nor_706_nl, nor_707_nl, fsm_output[0]);
  assign mux_2748_nl = MUX_s_1_2_2(mux_2747_nl, mux_2746_nl, fsm_output[1]);
  assign mux_2752_nl = MUX_s_1_2_2(mux_2751_nl, mux_2748_nl, fsm_output[2]);
  assign twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2752_nl & and_dcpl_268;
  assign nor_697_cse = ~((z_out_7[5:0]!=6'b001001) | (fsm_output[3:2]!=2'b01));
  assign nor_696_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b00100) | nand_191_cse);
  assign mux_2754_nl = MUX_s_1_2_2(nor_696_nl, nor_697_cse, fsm_output[0]);
  assign nor_699_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b001001) | (fsm_output[3]));
  assign mux_2753_nl = MUX_s_1_2_2(nor_697_cse, nor_699_nl, fsm_output[0]);
  assign mux_2755_nl = MUX_s_1_2_2(mux_2754_nl, mux_2753_nl, fsm_output[1]);
  assign twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2755_nl & and_dcpl_268;
  assign nor_692_cse = ~((z_out_7[5:0]!=6'b001010) | (fsm_output[3]));
  assign nor_691_cse = ~((z_out_7[4:0]!=5'b00101) | (fsm_output[3]));
  assign nor_690_nl = ~((z_out_7[5:0]!=6'b001010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2758_nl = MUX_s_1_2_2(nor_691_cse, nor_692_cse, fsm_output[0]);
  assign mux_2759_nl = MUX_s_1_2_2(nor_690_nl, mux_2758_nl, fsm_output[2]);
  assign nor_693_nl = ~((z_out_7[5:0]!=6'b001010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2756_nl = MUX_s_1_2_2(nor_692_cse, nor_691_cse, fsm_output[0]);
  assign mux_2757_nl = MUX_s_1_2_2(nor_693_nl, mux_2756_nl, fsm_output[2]);
  assign mux_2760_nl = MUX_s_1_2_2(mux_2759_nl, mux_2757_nl, fsm_output[1]);
  assign twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2760_nl & and_dcpl_268;
  assign nor_687_cse = ~((z_out_7[5:0]!=6'b001011) | (fsm_output[3:2]!=2'b01));
  assign nor_686_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b0010) | nand_190_cse);
  assign mux_2762_nl = MUX_s_1_2_2(nor_686_nl, nor_687_cse, fsm_output[0]);
  assign nor_689_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b001011) | (fsm_output[3]));
  assign mux_2761_nl = MUX_s_1_2_2(nor_687_cse, nor_689_nl, fsm_output[0]);
  assign mux_2763_nl = MUX_s_1_2_2(mux_2762_nl, mux_2761_nl, fsm_output[1]);
  assign twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2763_nl & and_dcpl_268;
  assign nor_679_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b00110) | (~ (fsm_output[3])));
  assign nor_680_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b001100) | (~ (fsm_output[3])));
  assign mux_2767_nl = MUX_s_1_2_2(nor_679_nl, nor_680_nl, fsm_output[0]);
  assign nor_681_nl = ~((z_out_7[4:0]!=5'b00110) | (fsm_output[3]));
  assign nor_682_nl = ~((z_out_7[5:0]!=6'b001100) | (fsm_output[3]));
  assign mux_2766_nl = MUX_s_1_2_2(nor_681_nl, nor_682_nl, fsm_output[0]);
  assign mux_2768_nl = MUX_s_1_2_2(mux_2767_nl, mux_2766_nl, fsm_output[2]);
  assign nor_683_nl = ~((z_out_7[5:0]!=6'b001100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_684_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0011) | (fsm_output[3]));
  assign nor_685_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b001100) | (fsm_output[3]));
  assign mux_2764_nl = MUX_s_1_2_2(nor_684_nl, nor_685_nl, fsm_output[0]);
  assign mux_2765_nl = MUX_s_1_2_2(nor_683_nl, mux_2764_nl, fsm_output[2]);
  assign mux_2769_nl = MUX_s_1_2_2(mux_2768_nl, mux_2765_nl, fsm_output[1]);
  assign twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2769_nl & and_dcpl_268;
  assign nor_676_cse = ~((z_out_7[5:0]!=6'b001101) | (fsm_output[3:2]!=2'b01));
  assign nor_675_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b00110) | nand_191_cse);
  assign mux_2771_nl = MUX_s_1_2_2(nor_675_nl, nor_676_cse, fsm_output[0]);
  assign nor_678_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b001101) | (fsm_output[3]));
  assign mux_2770_nl = MUX_s_1_2_2(nor_676_cse, nor_678_nl, fsm_output[0]);
  assign mux_2772_nl = MUX_s_1_2_2(mux_2771_nl, mux_2770_nl, fsm_output[1]);
  assign twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2772_nl & and_dcpl_268;
  assign nor_671_cse = ~((z_out_7[5:0]!=6'b001110) | (fsm_output[3]));
  assign nor_670_cse = ~((z_out_7[4:0]!=5'b00111) | (fsm_output[3]));
  assign nor_669_nl = ~((z_out_7[5:0]!=6'b001110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2775_nl = MUX_s_1_2_2(nor_670_cse, nor_671_cse, fsm_output[0]);
  assign mux_2776_nl = MUX_s_1_2_2(nor_669_nl, mux_2775_nl, fsm_output[2]);
  assign nor_672_nl = ~((z_out_7[5:0]!=6'b001110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2773_nl = MUX_s_1_2_2(nor_671_cse, nor_670_cse, fsm_output[0]);
  assign mux_2774_nl = MUX_s_1_2_2(nor_672_nl, mux_2773_nl, fsm_output[2]);
  assign mux_2777_nl = MUX_s_1_2_2(mux_2776_nl, mux_2774_nl, fsm_output[1]);
  assign twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2777_nl & and_dcpl_268;
  assign nor_666_cse = ~((z_out_7[5:0]!=6'b001111) | (fsm_output[3:2]!=2'b01));
  assign nor_665_nl = ~((fsm_output[2]) | (z_out_7[5:4]!=2'b00) | nand_184_cse);
  assign mux_2779_nl = MUX_s_1_2_2(nor_665_nl, nor_666_cse, fsm_output[0]);
  assign nor_668_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b001111) | (fsm_output[3]));
  assign mux_2778_nl = MUX_s_1_2_2(nor_666_cse, nor_668_nl, fsm_output[0]);
  assign mux_2780_nl = MUX_s_1_2_2(mux_2779_nl, mux_2778_nl, fsm_output[1]);
  assign twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2780_nl & and_dcpl_268;
  assign nor_660_cse = ~((z_out_7[5:0]!=6'b010000) | (fsm_output[3]));
  assign nor_657_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b01000) | (~ (fsm_output[3])));
  assign nor_658_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b010000) | (~ (fsm_output[3])));
  assign mux_2785_nl = MUX_s_1_2_2(nor_657_nl, nor_658_nl, fsm_output[0]);
  assign nor_659_nl = ~((z_out_8[2:0]!=3'b010) | (fsm_output[3]));
  assign mux_2784_nl = MUX_s_1_2_2(nor_659_nl, nor_660_cse, fsm_output[0]);
  assign mux_2786_nl = MUX_s_1_2_2(mux_2785_nl, mux_2784_nl, fsm_output[1]);
  assign nor_661_nl = ~((z_out_7[4:0]!=5'b01000) | (fsm_output[3]));
  assign mux_2782_nl = MUX_s_1_2_2(nor_661_nl, nor_660_cse, fsm_output[0]);
  assign nor_663_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0100) | (fsm_output[3]));
  assign nor_664_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b010000) | (fsm_output[3]));
  assign mux_2781_nl = MUX_s_1_2_2(nor_663_nl, nor_664_nl, fsm_output[0]);
  assign mux_2783_nl = MUX_s_1_2_2(mux_2782_nl, mux_2781_nl, fsm_output[1]);
  assign mux_2787_nl = MUX_s_1_2_2(mux_2786_nl, mux_2783_nl, fsm_output[2]);
  assign twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2787_nl & and_dcpl_268;
  assign nor_654_cse = ~((z_out_7[5:0]!=6'b010001) | (fsm_output[3:2]!=2'b01));
  assign nor_653_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b01000) | nand_191_cse);
  assign mux_2789_nl = MUX_s_1_2_2(nor_653_nl, nor_654_cse, fsm_output[0]);
  assign nor_656_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b010001) | (fsm_output[3]));
  assign mux_2788_nl = MUX_s_1_2_2(nor_654_cse, nor_656_nl, fsm_output[0]);
  assign mux_2790_nl = MUX_s_1_2_2(mux_2789_nl, mux_2788_nl, fsm_output[1]);
  assign twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2790_nl & and_dcpl_268;
  assign nor_649_cse = ~((z_out_7[5:0]!=6'b010010) | (fsm_output[3]));
  assign nor_648_cse = ~((z_out_7[4:0]!=5'b01001) | (fsm_output[3]));
  assign nor_647_nl = ~((z_out_7[5:0]!=6'b010010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2793_nl = MUX_s_1_2_2(nor_648_cse, nor_649_cse, fsm_output[0]);
  assign mux_2794_nl = MUX_s_1_2_2(nor_647_nl, mux_2793_nl, fsm_output[2]);
  assign nor_650_nl = ~((z_out_7[5:0]!=6'b010010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2791_nl = MUX_s_1_2_2(nor_649_cse, nor_648_cse, fsm_output[0]);
  assign mux_2792_nl = MUX_s_1_2_2(nor_650_nl, mux_2791_nl, fsm_output[2]);
  assign mux_2795_nl = MUX_s_1_2_2(mux_2794_nl, mux_2792_nl, fsm_output[1]);
  assign twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2795_nl & and_dcpl_268;
  assign nor_644_cse = ~((z_out_7[5:0]!=6'b010011) | (fsm_output[3:2]!=2'b01));
  assign nor_643_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b0100) | nand_190_cse);
  assign mux_2797_nl = MUX_s_1_2_2(nor_643_nl, nor_644_cse, fsm_output[0]);
  assign nor_646_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b010011) | (fsm_output[3]));
  assign mux_2796_nl = MUX_s_1_2_2(nor_644_cse, nor_646_nl, fsm_output[0]);
  assign mux_2798_nl = MUX_s_1_2_2(mux_2797_nl, mux_2796_nl, fsm_output[1]);
  assign twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2798_nl & and_dcpl_268;
  assign nor_636_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b01010) | (~ (fsm_output[3])));
  assign nor_637_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b010100) | (~ (fsm_output[3])));
  assign mux_2802_nl = MUX_s_1_2_2(nor_636_nl, nor_637_nl, fsm_output[0]);
  assign nor_638_nl = ~((z_out_7[4:0]!=5'b01010) | (fsm_output[3]));
  assign nor_639_nl = ~((z_out_7[5:0]!=6'b010100) | (fsm_output[3]));
  assign mux_2801_nl = MUX_s_1_2_2(nor_638_nl, nor_639_nl, fsm_output[0]);
  assign mux_2803_nl = MUX_s_1_2_2(mux_2802_nl, mux_2801_nl, fsm_output[2]);
  assign nor_640_nl = ~((z_out_7[5:0]!=6'b010100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_641_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0101) | (fsm_output[3]));
  assign nor_642_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b010100) | (fsm_output[3]));
  assign mux_2799_nl = MUX_s_1_2_2(nor_641_nl, nor_642_nl, fsm_output[0]);
  assign mux_2800_nl = MUX_s_1_2_2(nor_640_nl, mux_2799_nl, fsm_output[2]);
  assign mux_2804_nl = MUX_s_1_2_2(mux_2803_nl, mux_2800_nl, fsm_output[1]);
  assign twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2804_nl & and_dcpl_268;
  assign nor_633_cse = ~((z_out_7[5:0]!=6'b010101) | (fsm_output[3:2]!=2'b01));
  assign nor_632_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b01010) | nand_191_cse);
  assign mux_2806_nl = MUX_s_1_2_2(nor_632_nl, nor_633_cse, fsm_output[0]);
  assign nor_635_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b010101) | (fsm_output[3]));
  assign mux_2805_nl = MUX_s_1_2_2(nor_633_cse, nor_635_nl, fsm_output[0]);
  assign mux_2807_nl = MUX_s_1_2_2(mux_2806_nl, mux_2805_nl, fsm_output[1]);
  assign twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2807_nl & and_dcpl_268;
  assign nor_628_cse = ~((z_out_7[5:0]!=6'b010110) | (fsm_output[3]));
  assign nor_627_cse = ~((z_out_7[4:0]!=5'b01011) | (fsm_output[3]));
  assign nor_626_nl = ~((z_out_7[5:0]!=6'b010110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2810_nl = MUX_s_1_2_2(nor_627_cse, nor_628_cse, fsm_output[0]);
  assign mux_2811_nl = MUX_s_1_2_2(nor_626_nl, mux_2810_nl, fsm_output[2]);
  assign nor_629_nl = ~((z_out_7[5:0]!=6'b010110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2808_nl = MUX_s_1_2_2(nor_628_cse, nor_627_cse, fsm_output[0]);
  assign mux_2809_nl = MUX_s_1_2_2(nor_629_nl, mux_2808_nl, fsm_output[2]);
  assign mux_2812_nl = MUX_s_1_2_2(mux_2811_nl, mux_2809_nl, fsm_output[1]);
  assign twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2812_nl & and_dcpl_268;
  assign nor_623_cse = ~((z_out_7[5:0]!=6'b010111) | (fsm_output[3:2]!=2'b01));
  assign nor_622_nl = ~((fsm_output[2]) | (z_out_7[5:3]!=3'b010) | nand_188_cse);
  assign mux_2814_nl = MUX_s_1_2_2(nor_622_nl, nor_623_cse, fsm_output[0]);
  assign nor_625_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b010111) | (fsm_output[3]));
  assign mux_2813_nl = MUX_s_1_2_2(nor_623_cse, nor_625_nl, fsm_output[0]);
  assign mux_2815_nl = MUX_s_1_2_2(mux_2814_nl, mux_2813_nl, fsm_output[1]);
  assign twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2815_nl & and_dcpl_268;
  assign nor_617_cse = ~((z_out_7[5:0]!=6'b011000) | (fsm_output[3]));
  assign nor_614_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b01100) | (~ (fsm_output[3])));
  assign nor_615_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b011000) | (~ (fsm_output[3])));
  assign mux_2820_nl = MUX_s_1_2_2(nor_614_nl, nor_615_nl, fsm_output[0]);
  assign nor_616_nl = ~((z_out_8[2:0]!=3'b011) | (fsm_output[3]));
  assign mux_2819_nl = MUX_s_1_2_2(nor_616_nl, nor_617_cse, fsm_output[0]);
  assign mux_2821_nl = MUX_s_1_2_2(mux_2820_nl, mux_2819_nl, fsm_output[1]);
  assign nor_618_nl = ~((z_out_7[4:0]!=5'b01100) | (fsm_output[3]));
  assign mux_2817_nl = MUX_s_1_2_2(nor_618_nl, nor_617_cse, fsm_output[0]);
  assign nor_620_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0110) | (fsm_output[3]));
  assign nor_621_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b011000) | (fsm_output[3]));
  assign mux_2816_nl = MUX_s_1_2_2(nor_620_nl, nor_621_nl, fsm_output[0]);
  assign mux_2818_nl = MUX_s_1_2_2(mux_2817_nl, mux_2816_nl, fsm_output[1]);
  assign mux_2822_nl = MUX_s_1_2_2(mux_2821_nl, mux_2818_nl, fsm_output[2]);
  assign twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2822_nl & and_dcpl_268;
  assign nor_611_cse = ~((z_out_7[5:0]!=6'b011001) | (fsm_output[3:2]!=2'b01));
  assign nor_610_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b01100) | nand_191_cse);
  assign mux_2824_nl = MUX_s_1_2_2(nor_610_nl, nor_611_cse, fsm_output[0]);
  assign nor_613_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b011001) | (fsm_output[3]));
  assign mux_2823_nl = MUX_s_1_2_2(nor_611_cse, nor_613_nl, fsm_output[0]);
  assign mux_2825_nl = MUX_s_1_2_2(mux_2824_nl, mux_2823_nl, fsm_output[1]);
  assign twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2825_nl & and_dcpl_268;
  assign nor_606_cse = ~((z_out_7[5:0]!=6'b011010) | (fsm_output[3]));
  assign nor_605_cse = ~((z_out_7[4:0]!=5'b01101) | (fsm_output[3]));
  assign nor_604_nl = ~((z_out_7[5:0]!=6'b011010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2828_nl = MUX_s_1_2_2(nor_605_cse, nor_606_cse, fsm_output[0]);
  assign mux_2829_nl = MUX_s_1_2_2(nor_604_nl, mux_2828_nl, fsm_output[2]);
  assign nor_607_nl = ~((z_out_7[5:0]!=6'b011010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2826_nl = MUX_s_1_2_2(nor_606_cse, nor_605_cse, fsm_output[0]);
  assign mux_2827_nl = MUX_s_1_2_2(nor_607_nl, mux_2826_nl, fsm_output[2]);
  assign mux_2830_nl = MUX_s_1_2_2(mux_2829_nl, mux_2827_nl, fsm_output[1]);
  assign twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2830_nl & and_dcpl_268;
  assign nor_601_cse = ~((z_out_7[5:0]!=6'b011011) | (fsm_output[3:2]!=2'b01));
  assign nor_600_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b0110) | nand_190_cse);
  assign mux_2832_nl = MUX_s_1_2_2(nor_600_nl, nor_601_cse, fsm_output[0]);
  assign nor_603_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b011011) | (fsm_output[3]));
  assign mux_2831_nl = MUX_s_1_2_2(nor_601_cse, nor_603_nl, fsm_output[0]);
  assign mux_2833_nl = MUX_s_1_2_2(mux_2832_nl, mux_2831_nl, fsm_output[1]);
  assign twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2833_nl & and_dcpl_268;
  assign nor_593_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b01110) | (~ (fsm_output[3])));
  assign nor_594_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b011100) | (~ (fsm_output[3])));
  assign mux_2837_nl = MUX_s_1_2_2(nor_593_nl, nor_594_nl, fsm_output[0]);
  assign nor_595_nl = ~((z_out_7[4:0]!=5'b01110) | (fsm_output[3]));
  assign nor_596_nl = ~((z_out_7[5:0]!=6'b011100) | (fsm_output[3]));
  assign mux_2836_nl = MUX_s_1_2_2(nor_595_nl, nor_596_nl, fsm_output[0]);
  assign mux_2838_nl = MUX_s_1_2_2(mux_2837_nl, mux_2836_nl, fsm_output[2]);
  assign nor_597_nl = ~((z_out_7[5:0]!=6'b011100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_598_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b0111) | (fsm_output[3]));
  assign nor_599_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b011100) | (fsm_output[3]));
  assign mux_2834_nl = MUX_s_1_2_2(nor_598_nl, nor_599_nl, fsm_output[0]);
  assign mux_2835_nl = MUX_s_1_2_2(nor_597_nl, mux_2834_nl, fsm_output[2]);
  assign mux_2839_nl = MUX_s_1_2_2(mux_2838_nl, mux_2835_nl, fsm_output[1]);
  assign twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2839_nl & and_dcpl_268;
  assign nor_590_cse = ~((z_out_7[5:0]!=6'b011101) | (fsm_output[3:2]!=2'b01));
  assign nor_589_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b01110) | nand_191_cse);
  assign mux_2841_nl = MUX_s_1_2_2(nor_589_nl, nor_590_cse, fsm_output[0]);
  assign nor_592_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b011101) | (fsm_output[3]));
  assign mux_2840_nl = MUX_s_1_2_2(nor_590_cse, nor_592_nl, fsm_output[0]);
  assign mux_2842_nl = MUX_s_1_2_2(mux_2841_nl, mux_2840_nl, fsm_output[1]);
  assign twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2842_nl & and_dcpl_268;
  assign nor_585_cse = ~((z_out_7[5:0]!=6'b011110) | (fsm_output[3]));
  assign nor_584_cse = ~((z_out_7[4:0]!=5'b01111) | (fsm_output[3]));
  assign nor_583_nl = ~((z_out_7[5:0]!=6'b011110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2845_nl = MUX_s_1_2_2(nor_584_cse, nor_585_cse, fsm_output[0]);
  assign mux_2846_nl = MUX_s_1_2_2(nor_583_nl, mux_2845_nl, fsm_output[2]);
  assign nor_586_nl = ~((z_out_7[5:0]!=6'b011110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2843_nl = MUX_s_1_2_2(nor_585_cse, nor_584_cse, fsm_output[0]);
  assign mux_2844_nl = MUX_s_1_2_2(nor_586_nl, mux_2843_nl, fsm_output[2]);
  assign mux_2847_nl = MUX_s_1_2_2(mux_2846_nl, mux_2844_nl, fsm_output[1]);
  assign twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2847_nl & and_dcpl_268;
  assign and_533_cse = (z_out_7[5:0]==6'b011111) & (fsm_output[3:2]==2'b01);
  assign nor_581_nl = ~((fsm_output[2]) | (z_out_7[5]) | (~((z_out_7[4:0]==5'b11111)
      & (fsm_output[3]))));
  assign mux_2849_nl = MUX_s_1_2_2(nor_581_nl, and_533_cse, fsm_output[0]);
  assign nor_582_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b011111) | (fsm_output[3]));
  assign mux_2848_nl = MUX_s_1_2_2(and_533_cse, nor_582_nl, fsm_output[0]);
  assign mux_2850_nl = MUX_s_1_2_2(mux_2849_nl, mux_2848_nl, fsm_output[1]);
  assign twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2850_nl & and_dcpl_268;
  assign nor_576_cse = ~((z_out_7[5:0]!=6'b100000) | (fsm_output[3]));
  assign nor_573_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:0]!=4'b0000) | nand_174_cse);
  assign nor_574_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:0]!=5'b00000) | nand_175_cse);
  assign mux_2855_nl = MUX_s_1_2_2(nor_573_nl, nor_574_nl, fsm_output[0]);
  assign nor_575_nl = ~((z_out_8[2:0]!=3'b100) | (fsm_output[3]));
  assign mux_2854_nl = MUX_s_1_2_2(nor_575_nl, nor_576_cse, fsm_output[0]);
  assign mux_2856_nl = MUX_s_1_2_2(mux_2855_nl, mux_2854_nl, fsm_output[1]);
  assign nor_577_nl = ~((z_out_7[4:0]!=5'b10000) | (fsm_output[3]));
  assign mux_2852_nl = MUX_s_1_2_2(nor_577_nl, nor_576_cse, fsm_output[0]);
  assign nor_579_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1000) | (fsm_output[3]));
  assign nor_580_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b100000) | (fsm_output[3]));
  assign mux_2851_nl = MUX_s_1_2_2(nor_579_nl, nor_580_nl, fsm_output[0]);
  assign mux_2853_nl = MUX_s_1_2_2(mux_2852_nl, mux_2851_nl, fsm_output[1]);
  assign mux_2857_nl = MUX_s_1_2_2(mux_2856_nl, mux_2853_nl, fsm_output[2]);
  assign twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2857_nl & and_dcpl_268;
  assign nor_570_cse = ~((z_out_7[5:0]!=6'b100001) | (fsm_output[3:2]!=2'b01));
  assign nor_569_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b10000) | nand_191_cse);
  assign mux_2859_nl = MUX_s_1_2_2(nor_569_nl, nor_570_cse, fsm_output[0]);
  assign nor_572_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b100001) | (fsm_output[3]));
  assign mux_2858_nl = MUX_s_1_2_2(nor_570_cse, nor_572_nl, fsm_output[0]);
  assign mux_2860_nl = MUX_s_1_2_2(mux_2859_nl, mux_2858_nl, fsm_output[1]);
  assign twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2860_nl & and_dcpl_268;
  assign nor_565_cse = ~((z_out_7[5:0]!=6'b100010) | (fsm_output[3]));
  assign nor_564_cse = ~((z_out_7[4:0]!=5'b10001) | (fsm_output[3]));
  assign nor_563_nl = ~((z_out_7[5:0]!=6'b100010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2863_nl = MUX_s_1_2_2(nor_564_cse, nor_565_cse, fsm_output[0]);
  assign mux_2864_nl = MUX_s_1_2_2(nor_563_nl, mux_2863_nl, fsm_output[2]);
  assign nor_566_nl = ~((z_out_7[5:0]!=6'b100010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2861_nl = MUX_s_1_2_2(nor_565_cse, nor_564_cse, fsm_output[0]);
  assign mux_2862_nl = MUX_s_1_2_2(nor_566_nl, mux_2861_nl, fsm_output[2]);
  assign mux_2865_nl = MUX_s_1_2_2(mux_2864_nl, mux_2862_nl, fsm_output[1]);
  assign twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2865_nl & and_dcpl_268;
  assign nor_560_cse = ~((z_out_7[5:0]!=6'b100011) | (fsm_output[3:2]!=2'b01));
  assign nor_559_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b1000) | nand_190_cse);
  assign mux_2867_nl = MUX_s_1_2_2(nor_559_nl, nor_560_cse, fsm_output[0]);
  assign nor_562_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b100011) | (fsm_output[3]));
  assign mux_2866_nl = MUX_s_1_2_2(nor_560_cse, nor_562_nl, fsm_output[0]);
  assign mux_2868_nl = MUX_s_1_2_2(mux_2867_nl, mux_2866_nl, fsm_output[1]);
  assign twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2868_nl & and_dcpl_268;
  assign nor_552_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b10010) | (~ (fsm_output[3])));
  assign nor_553_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b100100) | (~ (fsm_output[3])));
  assign mux_2872_nl = MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output[0]);
  assign nor_554_nl = ~((z_out_7[4:0]!=5'b10010) | (fsm_output[3]));
  assign nor_555_nl = ~((z_out_7[5:0]!=6'b100100) | (fsm_output[3]));
  assign mux_2871_nl = MUX_s_1_2_2(nor_554_nl, nor_555_nl, fsm_output[0]);
  assign mux_2873_nl = MUX_s_1_2_2(mux_2872_nl, mux_2871_nl, fsm_output[2]);
  assign nor_556_nl = ~((z_out_7[5:0]!=6'b100100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_557_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1001) | (fsm_output[3]));
  assign nor_558_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b100100) | (fsm_output[3]));
  assign mux_2869_nl = MUX_s_1_2_2(nor_557_nl, nor_558_nl, fsm_output[0]);
  assign mux_2870_nl = MUX_s_1_2_2(nor_556_nl, mux_2869_nl, fsm_output[2]);
  assign mux_2874_nl = MUX_s_1_2_2(mux_2873_nl, mux_2870_nl, fsm_output[1]);
  assign twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2874_nl & and_dcpl_268;
  assign nor_549_cse = ~((z_out_7[5:0]!=6'b100101) | (fsm_output[3:2]!=2'b01));
  assign nor_548_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b10010) | nand_191_cse);
  assign mux_2876_nl = MUX_s_1_2_2(nor_548_nl, nor_549_cse, fsm_output[0]);
  assign nor_551_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b100101) | (fsm_output[3]));
  assign mux_2875_nl = MUX_s_1_2_2(nor_549_cse, nor_551_nl, fsm_output[0]);
  assign mux_2877_nl = MUX_s_1_2_2(mux_2876_nl, mux_2875_nl, fsm_output[1]);
  assign twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2877_nl & and_dcpl_268;
  assign nor_544_cse = ~((z_out_7[5:0]!=6'b100110) | (fsm_output[3]));
  assign nor_543_cse = ~((z_out_7[4:0]!=5'b10011) | (fsm_output[3]));
  assign nor_542_nl = ~((z_out_7[5:0]!=6'b100110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2880_nl = MUX_s_1_2_2(nor_543_cse, nor_544_cse, fsm_output[0]);
  assign mux_2881_nl = MUX_s_1_2_2(nor_542_nl, mux_2880_nl, fsm_output[2]);
  assign nor_545_nl = ~((z_out_7[5:0]!=6'b100110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2878_nl = MUX_s_1_2_2(nor_544_cse, nor_543_cse, fsm_output[0]);
  assign mux_2879_nl = MUX_s_1_2_2(nor_545_nl, mux_2878_nl, fsm_output[2]);
  assign mux_2882_nl = MUX_s_1_2_2(mux_2881_nl, mux_2879_nl, fsm_output[1]);
  assign twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2882_nl & and_dcpl_268;
  assign nor_539_cse = ~((z_out_7[5:0]!=6'b100111) | (fsm_output[3:2]!=2'b01));
  assign nor_538_nl = ~((fsm_output[2]) | (z_out_7[5:3]!=3'b100) | nand_188_cse);
  assign mux_2884_nl = MUX_s_1_2_2(nor_538_nl, nor_539_cse, fsm_output[0]);
  assign nor_541_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b100111) | (fsm_output[3]));
  assign mux_2883_nl = MUX_s_1_2_2(nor_539_cse, nor_541_nl, fsm_output[0]);
  assign mux_2885_nl = MUX_s_1_2_2(mux_2884_nl, mux_2883_nl, fsm_output[1]);
  assign twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2885_nl & and_dcpl_268;
  assign nor_533_cse = ~((z_out_7[5:0]!=6'b101000) | (fsm_output[3]));
  assign nor_530_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[3:0]!=4'b0100) | nand_174_cse);
  assign nor_531_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[4:0]!=5'b01000) | nand_175_cse);
  assign mux_2890_nl = MUX_s_1_2_2(nor_530_nl, nor_531_nl, fsm_output[0]);
  assign nor_532_nl = ~((z_out_8[2:0]!=3'b101) | (fsm_output[3]));
  assign mux_2889_nl = MUX_s_1_2_2(nor_532_nl, nor_533_cse, fsm_output[0]);
  assign mux_2891_nl = MUX_s_1_2_2(mux_2890_nl, mux_2889_nl, fsm_output[1]);
  assign nor_534_nl = ~((z_out_7[4:0]!=5'b10100) | (fsm_output[3]));
  assign mux_2887_nl = MUX_s_1_2_2(nor_534_nl, nor_533_cse, fsm_output[0]);
  assign nor_536_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1010) | (fsm_output[3]));
  assign nor_537_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b101000) | (fsm_output[3]));
  assign mux_2886_nl = MUX_s_1_2_2(nor_536_nl, nor_537_nl, fsm_output[0]);
  assign mux_2888_nl = MUX_s_1_2_2(mux_2887_nl, mux_2886_nl, fsm_output[1]);
  assign mux_2892_nl = MUX_s_1_2_2(mux_2891_nl, mux_2888_nl, fsm_output[2]);
  assign twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2892_nl & and_dcpl_268;
  assign nor_527_cse = ~((z_out_7[5:0]!=6'b101001) | (fsm_output[3:2]!=2'b01));
  assign nor_526_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b10100) | nand_191_cse);
  assign mux_2894_nl = MUX_s_1_2_2(nor_526_nl, nor_527_cse, fsm_output[0]);
  assign nor_529_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b101001) | (fsm_output[3]));
  assign mux_2893_nl = MUX_s_1_2_2(nor_527_cse, nor_529_nl, fsm_output[0]);
  assign mux_2895_nl = MUX_s_1_2_2(mux_2894_nl, mux_2893_nl, fsm_output[1]);
  assign twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2895_nl & and_dcpl_268;
  assign nor_522_cse = ~((z_out_7[5:0]!=6'b101010) | (fsm_output[3]));
  assign nor_521_cse = ~((z_out_7[4:0]!=5'b10101) | (fsm_output[3]));
  assign nor_520_nl = ~((z_out_7[5:0]!=6'b101010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2898_nl = MUX_s_1_2_2(nor_521_cse, nor_522_cse, fsm_output[0]);
  assign mux_2899_nl = MUX_s_1_2_2(nor_520_nl, mux_2898_nl, fsm_output[2]);
  assign nor_523_nl = ~((z_out_7[5:0]!=6'b101010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2896_nl = MUX_s_1_2_2(nor_522_cse, nor_521_cse, fsm_output[0]);
  assign mux_2897_nl = MUX_s_1_2_2(nor_523_nl, mux_2896_nl, fsm_output[2]);
  assign mux_2900_nl = MUX_s_1_2_2(mux_2899_nl, mux_2897_nl, fsm_output[1]);
  assign twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2900_nl & and_dcpl_268;
  assign nor_517_cse = ~((z_out_7[5:0]!=6'b101011) | (fsm_output[3:2]!=2'b01));
  assign nor_516_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b1010) | nand_190_cse);
  assign mux_2902_nl = MUX_s_1_2_2(nor_516_nl, nor_517_cse, fsm_output[0]);
  assign nor_519_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b101011) | (fsm_output[3]));
  assign mux_2901_nl = MUX_s_1_2_2(nor_517_cse, nor_519_nl, fsm_output[0]);
  assign mux_2903_nl = MUX_s_1_2_2(mux_2902_nl, mux_2901_nl, fsm_output[1]);
  assign twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2903_nl & and_dcpl_268;
  assign nor_509_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b10110) | (~ (fsm_output[3])));
  assign nor_510_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b101100) | (~ (fsm_output[3])));
  assign mux_2907_nl = MUX_s_1_2_2(nor_509_nl, nor_510_nl, fsm_output[0]);
  assign nor_511_nl = ~((z_out_7[4:0]!=5'b10110) | (fsm_output[3]));
  assign nor_512_nl = ~((z_out_7[5:0]!=6'b101100) | (fsm_output[3]));
  assign mux_2906_nl = MUX_s_1_2_2(nor_511_nl, nor_512_nl, fsm_output[0]);
  assign mux_2908_nl = MUX_s_1_2_2(mux_2907_nl, mux_2906_nl, fsm_output[2]);
  assign nor_513_nl = ~((z_out_7[5:0]!=6'b101100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_514_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1011) | (fsm_output[3]));
  assign nor_515_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b101100) | (fsm_output[3]));
  assign mux_2904_nl = MUX_s_1_2_2(nor_514_nl, nor_515_nl, fsm_output[0]);
  assign mux_2905_nl = MUX_s_1_2_2(nor_513_nl, mux_2904_nl, fsm_output[2]);
  assign mux_2909_nl = MUX_s_1_2_2(mux_2908_nl, mux_2905_nl, fsm_output[1]);
  assign twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2909_nl & and_dcpl_268;
  assign nor_506_cse = ~((z_out_7[5:0]!=6'b101101) | (fsm_output[3:2]!=2'b01));
  assign nor_505_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b10110) | nand_191_cse);
  assign mux_2911_nl = MUX_s_1_2_2(nor_505_nl, nor_506_cse, fsm_output[0]);
  assign nor_508_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b101101) | (fsm_output[3]));
  assign mux_2910_nl = MUX_s_1_2_2(nor_506_cse, nor_508_nl, fsm_output[0]);
  assign mux_2912_nl = MUX_s_1_2_2(mux_2911_nl, mux_2910_nl, fsm_output[1]);
  assign twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2912_nl & and_dcpl_268;
  assign nor_501_cse = ~((z_out_7[5:0]!=6'b101110) | (fsm_output[3]));
  assign nor_500_cse = ~((z_out_7[4:0]!=5'b10111) | (fsm_output[3]));
  assign nor_499_nl = ~((z_out_7[5:0]!=6'b101110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2915_nl = MUX_s_1_2_2(nor_500_cse, nor_501_cse, fsm_output[0]);
  assign mux_2916_nl = MUX_s_1_2_2(nor_499_nl, mux_2915_nl, fsm_output[2]);
  assign nor_502_nl = ~((z_out_7[5:0]!=6'b101110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2913_nl = MUX_s_1_2_2(nor_501_cse, nor_500_cse, fsm_output[0]);
  assign mux_2914_nl = MUX_s_1_2_2(nor_502_nl, mux_2913_nl, fsm_output[2]);
  assign mux_2917_nl = MUX_s_1_2_2(mux_2916_nl, mux_2914_nl, fsm_output[1]);
  assign twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2917_nl & and_dcpl_268;
  assign and_531_cse = (z_out_7[5:0]==6'b101111) & (fsm_output[3:2]==2'b01);
  assign nor_497_nl = ~((fsm_output[2]) | (z_out_7[5:4]!=2'b10) | nand_184_cse);
  assign mux_2919_nl = MUX_s_1_2_2(nor_497_nl, and_531_cse, fsm_output[0]);
  assign nor_498_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b101111) | (fsm_output[3]));
  assign mux_2918_nl = MUX_s_1_2_2(and_531_cse, nor_498_nl, fsm_output[0]);
  assign mux_2920_nl = MUX_s_1_2_2(mux_2919_nl, mux_2918_nl, fsm_output[1]);
  assign twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2920_nl & and_dcpl_268;
  assign nor_492_cse = ~((z_out_7[5:0]!=6'b110000) | (fsm_output[3]));
  assign nor_489_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[2:0]!=3'b000) | (~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:3]==2'b11)
      & (fsm_output[3]))));
  assign nor_490_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[3:0]!=4'b0000) | (~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:4]==2'b11)
      & (fsm_output[3]))));
  assign mux_2925_nl = MUX_s_1_2_2(nor_489_nl, nor_490_nl, fsm_output[0]);
  assign nor_491_nl = ~((z_out_8[2:0]!=3'b110) | (fsm_output[3]));
  assign mux_2924_nl = MUX_s_1_2_2(nor_491_nl, nor_492_cse, fsm_output[0]);
  assign mux_2926_nl = MUX_s_1_2_2(mux_2925_nl, mux_2924_nl, fsm_output[1]);
  assign nor_493_nl = ~((z_out_7[4:0]!=5'b11000) | (fsm_output[3]));
  assign mux_2922_nl = MUX_s_1_2_2(nor_493_nl, nor_492_cse, fsm_output[0]);
  assign nor_495_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1100) | (fsm_output[3]));
  assign nor_496_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b110000) | (fsm_output[3]));
  assign mux_2921_nl = MUX_s_1_2_2(nor_495_nl, nor_496_nl, fsm_output[0]);
  assign mux_2923_nl = MUX_s_1_2_2(mux_2922_nl, mux_2921_nl, fsm_output[1]);
  assign mux_2927_nl = MUX_s_1_2_2(mux_2926_nl, mux_2923_nl, fsm_output[2]);
  assign twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2927_nl & and_dcpl_268;
  assign nor_486_cse = ~((z_out_7[5:0]!=6'b110001) | (fsm_output[3:2]!=2'b01));
  assign nor_485_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b11000) | nand_191_cse);
  assign mux_2929_nl = MUX_s_1_2_2(nor_485_nl, nor_486_cse, fsm_output[0]);
  assign nor_488_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b110001) | (fsm_output[3]));
  assign mux_2928_nl = MUX_s_1_2_2(nor_486_cse, nor_488_nl, fsm_output[0]);
  assign mux_2930_nl = MUX_s_1_2_2(mux_2929_nl, mux_2928_nl, fsm_output[1]);
  assign twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2930_nl & and_dcpl_268;
  assign nor_481_cse = ~((z_out_7[5:0]!=6'b110010) | (fsm_output[3]));
  assign nor_480_cse = ~((z_out_7[4:0]!=5'b11001) | (fsm_output[3]));
  assign nor_479_nl = ~((z_out_7[5:0]!=6'b110010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2933_nl = MUX_s_1_2_2(nor_480_cse, nor_481_cse, fsm_output[0]);
  assign mux_2934_nl = MUX_s_1_2_2(nor_479_nl, mux_2933_nl, fsm_output[2]);
  assign nor_482_nl = ~((z_out_7[5:0]!=6'b110010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2931_nl = MUX_s_1_2_2(nor_481_cse, nor_480_cse, fsm_output[0]);
  assign mux_2932_nl = MUX_s_1_2_2(nor_482_nl, mux_2931_nl, fsm_output[2]);
  assign mux_2935_nl = MUX_s_1_2_2(mux_2934_nl, mux_2932_nl, fsm_output[1]);
  assign twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2935_nl & and_dcpl_268;
  assign nor_476_cse = ~((z_out_7[5:0]!=6'b110011) | (fsm_output[3:2]!=2'b01));
  assign nor_475_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b1100) | nand_190_cse);
  assign mux_2937_nl = MUX_s_1_2_2(nor_475_nl, nor_476_cse, fsm_output[0]);
  assign nor_478_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b110011) | (fsm_output[3]));
  assign mux_2936_nl = MUX_s_1_2_2(nor_476_cse, nor_478_nl, fsm_output[0]);
  assign mux_2938_nl = MUX_s_1_2_2(mux_2937_nl, mux_2936_nl, fsm_output[1]);
  assign twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2938_nl & and_dcpl_268;
  assign nor_468_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]!=5'b11010) | (~ (fsm_output[3])));
  assign nor_469_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]!=6'b110100) | (~ (fsm_output[3])));
  assign mux_2942_nl = MUX_s_1_2_2(nor_468_nl, nor_469_nl, fsm_output[0]);
  assign nor_470_nl = ~((z_out_7[4:0]!=5'b11010) | (fsm_output[3]));
  assign nor_471_nl = ~((z_out_7[5:0]!=6'b110100) | (fsm_output[3]));
  assign mux_2941_nl = MUX_s_1_2_2(nor_470_nl, nor_471_nl, fsm_output[0]);
  assign mux_2943_nl = MUX_s_1_2_2(mux_2942_nl, mux_2941_nl, fsm_output[2]);
  assign nor_472_nl = ~((z_out_7[5:0]!=6'b110100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign nor_473_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1101) | (fsm_output[3]));
  assign nor_474_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b110100) | (fsm_output[3]));
  assign mux_2939_nl = MUX_s_1_2_2(nor_473_nl, nor_474_nl, fsm_output[0]);
  assign mux_2940_nl = MUX_s_1_2_2(nor_472_nl, mux_2939_nl, fsm_output[2]);
  assign mux_2944_nl = MUX_s_1_2_2(mux_2943_nl, mux_2940_nl, fsm_output[1]);
  assign twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2944_nl & and_dcpl_268;
  assign nor_465_cse = ~((z_out_7[5:0]!=6'b110101) | (fsm_output[3:2]!=2'b01));
  assign nor_464_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b11010) | nand_191_cse);
  assign mux_2946_nl = MUX_s_1_2_2(nor_464_nl, nor_465_cse, fsm_output[0]);
  assign nor_467_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b110101) | (fsm_output[3]));
  assign mux_2945_nl = MUX_s_1_2_2(nor_465_cse, nor_467_nl, fsm_output[0]);
  assign mux_2947_nl = MUX_s_1_2_2(mux_2946_nl, mux_2945_nl, fsm_output[1]);
  assign twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2947_nl & and_dcpl_268;
  assign nor_460_cse = ~((z_out_7[5:0]!=6'b110110) | (fsm_output[3]));
  assign nor_459_cse = ~((z_out_7[4:0]!=5'b11011) | (fsm_output[3]));
  assign nor_458_nl = ~((z_out_7[5:0]!=6'b110110) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2950_nl = MUX_s_1_2_2(nor_459_cse, nor_460_cse, fsm_output[0]);
  assign mux_2951_nl = MUX_s_1_2_2(nor_458_nl, mux_2950_nl, fsm_output[2]);
  assign nor_461_nl = ~((z_out_7[5:0]!=6'b110110) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2948_nl = MUX_s_1_2_2(nor_460_cse, nor_459_cse, fsm_output[0]);
  assign mux_2949_nl = MUX_s_1_2_2(nor_461_nl, mux_2948_nl, fsm_output[2]);
  assign mux_2952_nl = MUX_s_1_2_2(mux_2951_nl, mux_2949_nl, fsm_output[1]);
  assign twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2952_nl & and_dcpl_268;
  assign and_529_cse = (z_out_7[5:0]==6'b110111) & (fsm_output[3:2]==2'b01);
  assign nor_456_nl = ~((fsm_output[2]) | (z_out_7[5:3]!=3'b110) | nand_188_cse);
  assign mux_2954_nl = MUX_s_1_2_2(nor_456_nl, and_529_cse, fsm_output[0]);
  assign nor_457_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b110111) | (fsm_output[3]));
  assign mux_2953_nl = MUX_s_1_2_2(and_529_cse, nor_457_nl, fsm_output[0]);
  assign mux_2955_nl = MUX_s_1_2_2(mux_2954_nl, mux_2953_nl, fsm_output[1]);
  assign twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2955_nl & and_dcpl_268;
  assign nor_451_cse = ~((z_out_7[5:0]!=6'b111000) | (fsm_output[3]));
  assign nor_449_nl = ~((COMP_LOOP_3_tmp_lshift_ncse_sva[1:0]!=2'b00) | (~((COMP_LOOP_3_tmp_lshift_ncse_sva[4:2]==3'b111)
      & (fsm_output[3]))));
  assign nor_450_nl = ~((COMP_LOOP_2_tmp_lshift_ncse_sva[2:0]!=3'b000) | (~((COMP_LOOP_2_tmp_lshift_ncse_sva[5:3]==3'b111)
      & (fsm_output[3]))));
  assign mux_2960_nl = MUX_s_1_2_2(nor_449_nl, nor_450_nl, fsm_output[0]);
  assign and_528_nl = (z_out_8[2:0]==3'b111) & (~ (fsm_output[3]));
  assign mux_2959_nl = MUX_s_1_2_2(and_528_nl, nor_451_cse, fsm_output[0]);
  assign mux_2961_nl = MUX_s_1_2_2(mux_2960_nl, mux_2959_nl, fsm_output[1]);
  assign nor_452_nl = ~((z_out_7[4:0]!=5'b11100) | (fsm_output[3]));
  assign mux_2957_nl = MUX_s_1_2_2(nor_452_nl, nor_451_cse, fsm_output[0]);
  assign nor_454_nl = ~((COMP_LOOP_5_tmp_mul_idiv_sva[3:0]!=4'b1110) | (fsm_output[3]));
  assign nor_455_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b111000) | (fsm_output[3]));
  assign mux_2956_nl = MUX_s_1_2_2(nor_454_nl, nor_455_nl, fsm_output[0]);
  assign mux_2958_nl = MUX_s_1_2_2(mux_2957_nl, mux_2956_nl, fsm_output[1]);
  assign mux_2962_nl = MUX_s_1_2_2(mux_2961_nl, mux_2958_nl, fsm_output[2]);
  assign twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2962_nl & and_dcpl_268;
  assign nor_446_cse = ~((z_out_7[5:0]!=6'b111001) | (fsm_output[3:2]!=2'b01));
  assign nor_445_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b11100) | nand_191_cse);
  assign mux_2964_nl = MUX_s_1_2_2(nor_445_nl, nor_446_cse, fsm_output[0]);
  assign nor_448_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b111001) | (fsm_output[3]));
  assign mux_2963_nl = MUX_s_1_2_2(nor_446_cse, nor_448_nl, fsm_output[0]);
  assign mux_2965_nl = MUX_s_1_2_2(mux_2964_nl, mux_2963_nl, fsm_output[1]);
  assign twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2965_nl & and_dcpl_268;
  assign nor_441_cse = ~((z_out_7[5:0]!=6'b111010) | (fsm_output[3]));
  assign nor_440_cse = ~((z_out_7[4:0]!=5'b11101) | (fsm_output[3]));
  assign nor_439_nl = ~((z_out_7[5:0]!=6'b111010) | (fsm_output[0]) | (~ (fsm_output[3])));
  assign mux_2968_nl = MUX_s_1_2_2(nor_440_cse, nor_441_cse, fsm_output[0]);
  assign mux_2969_nl = MUX_s_1_2_2(nor_439_nl, mux_2968_nl, fsm_output[2]);
  assign nor_442_nl = ~((z_out_7[5:0]!=6'b111010) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign mux_2966_nl = MUX_s_1_2_2(nor_441_cse, nor_440_cse, fsm_output[0]);
  assign mux_2967_nl = MUX_s_1_2_2(nor_442_nl, mux_2966_nl, fsm_output[2]);
  assign mux_2970_nl = MUX_s_1_2_2(mux_2969_nl, mux_2967_nl, fsm_output[1]);
  assign twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2970_nl & and_dcpl_268;
  assign and_526_cse = (z_out_7[5:0]==6'b111011) & (fsm_output[3:2]==2'b01);
  assign nor_437_nl = ~((fsm_output[2]) | (z_out_7[5:2]!=4'b1110) | nand_190_cse);
  assign mux_2972_nl = MUX_s_1_2_2(nor_437_nl, and_526_cse, fsm_output[0]);
  assign nor_438_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b111011) | (fsm_output[3]));
  assign mux_2971_nl = MUX_s_1_2_2(and_526_cse, nor_438_nl, fsm_output[0]);
  assign mux_2973_nl = MUX_s_1_2_2(mux_2972_nl, mux_2971_nl, fsm_output[1]);
  assign twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2973_nl & and_dcpl_268;
  assign and_789_nl = (COMP_LOOP_3_tmp_lshift_ncse_sva[4:0]==5'b11110) & (fsm_output[3]);
  assign and_810_nl = (COMP_LOOP_2_tmp_lshift_ncse_sva[5:0]==6'b111100) & (fsm_output[3]);
  assign mux_2977_nl = MUX_s_1_2_2(and_789_nl, and_810_nl, fsm_output[0]);
  assign nor_433_nl = ~((z_out_7[4:0]!=5'b11110) | (fsm_output[3]));
  assign nor_434_nl = ~((z_out_7[5:0]!=6'b111100) | (fsm_output[3]));
  assign mux_2976_nl = MUX_s_1_2_2(nor_433_nl, nor_434_nl, fsm_output[0]);
  assign mux_2978_nl = MUX_s_1_2_2(mux_2977_nl, mux_2976_nl, fsm_output[2]);
  assign nor_435_nl = ~((z_out_7[5:0]!=6'b111100) | (~ (fsm_output[0])) | (fsm_output[3]));
  assign and_525_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[3:0]==4'b1111) & (~ (fsm_output[3]));
  assign nor_436_nl = ~((COMP_LOOP_2_tmp_mul_idiv_sva[5:0]!=6'b111100) | (fsm_output[3]));
  assign mux_2974_nl = MUX_s_1_2_2(and_525_nl, nor_436_nl, fsm_output[0]);
  assign mux_2975_nl = MUX_s_1_2_2(nor_435_nl, mux_2974_nl, fsm_output[2]);
  assign mux_2979_nl = MUX_s_1_2_2(mux_2978_nl, mux_2975_nl, fsm_output[1]);
  assign twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2979_nl & and_dcpl_268;
  assign and_523_cse = (z_out_7[5:0]==6'b111101) & (fsm_output[3:2]==2'b01);
  assign nor_429_nl = ~((fsm_output[2]) | (z_out_7[5:1]!=5'b11110) | nand_191_cse);
  assign mux_2981_nl = MUX_s_1_2_2(nor_429_nl, and_523_cse, fsm_output[0]);
  assign nor_430_nl = ~((fsm_output[2]) | (z_out_7[5:0]!=6'b111101) | (fsm_output[3]));
  assign mux_2980_nl = MUX_s_1_2_2(and_523_cse, nor_430_nl, fsm_output[0]);
  assign mux_2982_nl = MUX_s_1_2_2(mux_2981_nl, mux_2980_nl, fsm_output[1]);
  assign twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2982_nl & and_dcpl_268;
  assign and_519_cse = (z_out_7[5:0]==6'b111110) & (~ (fsm_output[3]));
  assign and_518_cse = (z_out_7[4:0]==5'b11111) & (~ (fsm_output[3]));
  assign and_790_nl = (z_out_7[5:0]==6'b111110) & (~ (fsm_output[0])) & (fsm_output[3]);
  assign mux_2985_nl = MUX_s_1_2_2(and_518_cse, and_519_cse, fsm_output[0]);
  assign mux_2986_nl = MUX_s_1_2_2(and_790_nl, mux_2985_nl, fsm_output[2]);
  assign and_520_nl = (z_out_7[5:0]==6'b111110) & (fsm_output[0]) & (~ (fsm_output[3]));
  assign mux_2983_nl = MUX_s_1_2_2(and_519_cse, and_518_cse, fsm_output[0]);
  assign mux_2984_nl = MUX_s_1_2_2(and_520_nl, mux_2983_nl, fsm_output[2]);
  assign mux_2987_nl = MUX_s_1_2_2(mux_2986_nl, mux_2984_nl, fsm_output[1]);
  assign twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2987_nl & and_dcpl_268;
  assign and_515_cse = (z_out_7[5:0]==6'b111111) & (fsm_output[3:2]==2'b01);
  assign nor_427_nl = ~((fsm_output[2]) | (~((z_out_7[5:0]==6'b111111) & (fsm_output[3]))));
  assign mux_2989_nl = MUX_s_1_2_2(nor_427_nl, and_515_cse, fsm_output[0]);
  assign and_517_nl = (~ (fsm_output[2])) & (z_out_7[5:0]==6'b111111) & (~ (fsm_output[3]));
  assign mux_2988_nl = MUX_s_1_2_2(and_515_cse, and_517_nl, fsm_output[0]);
  assign mux_2990_nl = MUX_s_1_2_2(mux_2989_nl, mux_2988_nl, fsm_output[1]);
  assign twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d = mux_2990_nl & and_dcpl_268;
  assign nor_1716_cse = ~((fsm_output[7]) | (fsm_output[5]));
  assign nor_1715_cse = ~((fsm_output[3]) | (fsm_output[6]));
  assign and_dcpl_477 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_488 = (~ (fsm_output[4])) & (fsm_output[0]) & (~ (fsm_output[3]))
      & (fsm_output[6]) & and_dcpl_477 & (fsm_output[7]) & (fsm_output[5]);
  assign and_dcpl_501 = ~((fsm_output!=8'b00000010));
  assign and_dcpl_503 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_509 = (~ (fsm_output[7])) & (fsm_output[5]);
  assign and_dcpl_513 = and_dcpl_503 & and_dcpl_509;
  assign and_dcpl_514 = (fsm_output[3]) & (~ (fsm_output[6]));
  assign and_903_cse = and_dcpl_80 & and_dcpl_514 & and_dcpl_513;
  assign and_dcpl_519 = (fsm_output[3]) & (fsm_output[6]);
  assign and_907_cse = and_dcpl_80 & and_dcpl_519 & nor_1744_cse & nor_1716_cse;
  assign and_910_cse = and_dcpl_80 & (~ (fsm_output[3])) & (fsm_output[6]) & and_dcpl_513;
  assign and_dcpl_526 = nor_1744_cse & (fsm_output[7]) & (~ (fsm_output[5]));
  assign and_914_cse = and_dcpl_80 & nor_1715_cse & and_dcpl_526;
  assign and_918_cse = and_dcpl_58 & and_dcpl_514 & and_dcpl_503 & (fsm_output[7])
      & (fsm_output[5]);
  assign and_920_cse = and_dcpl_58 & and_dcpl_519 & and_dcpl_526;
  assign and_dcpl_570 = (fsm_output[2:1]==2'b01) & nor_1716_cse;
  assign and_dcpl_573 = and_dcpl_58 & nor_1715_cse;
  assign and_dcpl_574 = and_dcpl_573 & and_dcpl_570;
  assign and_dcpl_576 = (~ (fsm_output[4])) & (fsm_output[0]) & nor_1715_cse;
  assign and_dcpl_577 = and_dcpl_576 & and_dcpl_570;
  assign and_dcpl_579 = (fsm_output[2:1]==2'b10) & nor_1716_cse;
  assign and_dcpl_580 = and_dcpl_576 & and_dcpl_579;
  assign and_dcpl_582 = (fsm_output[2:1]==2'b11) & nor_1716_cse;
  assign and_dcpl_583 = and_dcpl_573 & and_dcpl_582;
  assign and_dcpl_588 = and_dcpl_58 & (fsm_output[3]) & (~ (fsm_output[6])) & (~
      (fsm_output[2])) & (~ (fsm_output[1])) & nor_1716_cse;
  assign and_dcpl_589 = and_dcpl_573 & and_dcpl_579;
  assign and_dcpl_590 = and_dcpl_576 & and_dcpl_582;
  assign and_dcpl_599 = nor_1744_cse & nor_1716_cse;
  assign and_dcpl_602 = and_dcpl_80 & nor_1715_cse & and_dcpl_599;
  assign and_dcpl_605 = and_dcpl_503 & (~ (fsm_output[7])) & (fsm_output[5]);
  assign and_dcpl_608 = and_dcpl_58 & and_dcpl_514 & and_dcpl_605;
  assign and_dcpl_611 = and_dcpl_58 & (fsm_output[3]) & (fsm_output[6]) & and_dcpl_599;
  assign and_dcpl_612 = (~ (fsm_output[3])) & (fsm_output[6]);
  assign and_dcpl_614 = and_dcpl_58 & and_dcpl_612 & and_dcpl_605;
  assign and_dcpl_615 = (fsm_output[7]) & (~ (fsm_output[5]));
  assign and_dcpl_617 = and_dcpl_573 & nor_1744_cse & and_dcpl_615;
  assign and_dcpl_618 = and_dcpl_503 & and_dcpl_615;
  assign and_dcpl_619 = and_dcpl_80 & and_dcpl_514;
  assign and_dcpl_620 = and_dcpl_619 & and_dcpl_618;
  assign and_dcpl_623 = and_dcpl_619 & nor_1744_cse & (fsm_output[7]) & (fsm_output[5]);
  assign and_dcpl_625 = and_dcpl_80 & and_dcpl_612 & and_dcpl_618;
  assign and_dcpl_632 = and_dcpl_573 & and_dcpl_503 & nor_1716_cse;
  assign and_dcpl_636 = and_dcpl_573 & nor_1744_cse & and_dcpl_509;
  assign COMP_LOOP_or_65_itm = (and_dcpl_58 & nor_1715_cse & nor_1744_cse & and_dcpl_509)
      | and_903_cse | and_907_cse | and_910_cse | and_914_cse | and_918_cse | and_920_cse;
  assign COMP_LOOP_tmp_or_83_itm = and_dcpl_589 | and_dcpl_590;
  assign COMP_LOOP_tmp_or_54_ssc = and_dcpl_580 | and_dcpl_583 | and_dcpl_588;
  always @(posedge clk) begin
    if ( (and_dcpl_60 & and_dcpl_57) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b1010, z_out_4, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_1423_nl, mux_789_nl, fsm_output[5]) ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_63_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      COMP_LOOP_1_tmp_mul_idiv_sva_2_0 <= 3'b000;
      COMP_LOOP_nor_326_itm <= 1'b0;
      COMP_LOOP_nor_319_itm <= 1'b0;
      COMP_LOOP_3_tmp_mul_idiv_sva_4_0 <= 5'b00000;
    end
    else begin
      reg_vec_rsc_triosy_0_63_obj_ld_cse <= and_dcpl_65 & (~ (fsm_output[0])) & (~
          (fsm_output[4])) & (fsm_output[6]) & (fsm_output[2]) & (~ (fsm_output[1]))
          & (fsm_output[5]) & (~ (z_out_2[4]));
      reg_ensig_cgo_cse <= mux_2997_rmff;
      COMP_LOOP_1_tmp_mul_idiv_sva_2_0 <= z_out_8[2:0];
      COMP_LOOP_nor_326_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[3:0]!=4'b0000));
      COMP_LOOP_nor_319_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4]) | (COMP_LOOP_2_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[1]) | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
      COMP_LOOP_3_tmp_mul_idiv_sva_4_0 <= z_out_7[4:0];
    end
  end
  always @(posedge clk) begin
    tmp_21_sva_2 <= MUX_v_64_2_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_58_i_q_d, and_dcpl_263);
    tmp_21_sva_6 <= twiddle_rsc_0_6_i_q_d;
    tmp_21_sva_11 <= MUX_v_64_2_2(twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_30_i_q_d,
        and_dcpl_263);
    tmp_21_sva_13 <= MUX_v_64_2_2(twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_34_i_q_d,
        and_dcpl_263);
    tmp_21_sva_14 <= MUX_v_64_2_2(twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_38_i_q_d,
        and_dcpl_263);
    tmp_21_sva_15 <= MUX_v_64_2_2(twiddle_rsc_0_15_i_q_d, twiddle_rsc_0_42_i_q_d,
        and_dcpl_263);
    tmp_21_sva_17 <= MUX_v_64_2_2(twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_46_i_q_d,
        and_dcpl_263);
    tmp_21_sva_18 <= MUX_v_64_2_2(twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_50_i_q_d,
        and_dcpl_263);
    tmp_21_sva_19 <= MUX_v_64_2_2(twiddle_rsc_0_19_i_q_d, twiddle_rsc_0_54_i_q_d,
        and_dcpl_263);
    tmp_21_sva_21 <= MUX_v_64_2_2(twiddle_rsc_0_21_i_q_d, twiddle_rsc_0_6_i_q_d,
        and_dcpl_263);
    tmp_21_sva_22 <= MUX_v_64_2_2(twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_62_i_q_d,
        and_dcpl_263);
    tmp_21_sva_23 <= MUX_v_64_2_2(twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_10_i_q_d,
        and_dcpl_263);
    tmp_21_sva_25 <= MUX_v_64_2_2(twiddle_rsc_0_25_i_q_d, twiddle_rsc_0_14_i_q_d,
        and_dcpl_263);
    tmp_21_sva_26 <= MUX_v_64_2_2(twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_18_i_q_d,
        and_dcpl_263);
    tmp_21_sva_30 <= twiddle_rsc_0_30_i_q_d;
    tmp_21_sva_34 <= twiddle_rsc_0_34_i_q_d;
    tmp_21_sva_38 <= twiddle_rsc_0_38_i_q_d;
    tmp_21_sva_42 <= twiddle_rsc_0_42_i_q_d;
    tmp_21_sva_46 <= twiddle_rsc_0_46_i_q_d;
    tmp_21_sva_50 <= twiddle_rsc_0_50_i_q_d;
    tmp_21_sva_54 <= twiddle_rsc_0_54_i_q_d;
    tmp_21_sva_58 <= twiddle_rsc_0_58_i_q_d;
    tmp_21_sva_62 <= twiddle_rsc_0_62_i_q_d;
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_10_0_sva_9_0 <= 10'b0000000000;
    end
    else if ( VEC_LOOP_j_10_0_sva_9_0_mx0c0 | (and_dcpl_108 & and_dcpl_97) ) begin
      VEC_LOOP_j_10_0_sva_9_0 <= MUX_v_10_2_2(10'b0000000000, (z_out_3[9:0]), VEC_LOOP_j_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(nor_422_nl, mux_tmp_720, fsm_output[5]) ) begin
      STAGE_LOOP_lshift_psp_sva <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(or_4159_nl, nand_493_nl, fsm_output[7]) ) begin
      COMP_LOOP_k_10_3_sva_6_0 <= MUX_v_7_2_2(7'b0000000, reg_COMP_LOOP_k_10_3_ftd,
          nand_480_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva <= 10'b0000000000;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_acc_10_cse_10_1_1_sva <= COMP_LOOP_1_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_psp_sva <= 7'b0000000;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_5_tmp_mul_idiv_sva <= 8'b00000000;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_5_tmp_mul_idiv_sva <= z_out_7[7:0];
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_2_slc_COMP_LOOP_acc_10_itm <= z_out_3[10];
    end
  end
  always @(posedge clk) begin
    if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_1_tmp_acc_cse_sva <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1518_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_760_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_761_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_509_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_510_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_258_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_260_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_261_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_262_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_264_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_268_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_522_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_270_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_18_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_272_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_20_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_21_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_22_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_23_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_24_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_25_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_26_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_27_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_28_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_29_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_30_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_284_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_285_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_286_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_34_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_288_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_36_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_37_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_38_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_39_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_40_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_41_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_42_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_43_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_44_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_45_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_46_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_47_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_48_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_49_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_50_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_51_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_52_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_53_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_54_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_55_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_56_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_57_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_58_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_59_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_60_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_61_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_62_itm <= 1'b0;
    end
    else if ( mux_3025_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((COMP_LOOP_acc_psp_sva_mx0w0[2:0]!=3'b000)
          | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000));
      COMP_LOOP_COMP_LOOP_and_1518_itm <= (COMP_LOOP_acc_14_psp_sva_1[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (COMP_LOOP_acc_14_psp_sva_1[4:2]==3'b000);
      COMP_LOOP_COMP_LOOP_and_760_itm <= (COMP_LOOP_acc_1_cse_4_sva_1[5:0]==6'b000101);
      COMP_LOOP_COMP_LOOP_and_761_itm <= (COMP_LOOP_acc_1_cse_4_sva_1[5:0]==6'b000110);
      COMP_LOOP_COMP_LOOP_and_509_itm <= (COMP_LOOP_acc_11_psp_sva_1[1:0]==2'b11)
          & (~((COMP_LOOP_acc_11_psp_sva_1[4:2]!=3'b000) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_510_itm <= (COMP_LOOP_acc_11_psp_sva_1[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (COMP_LOOP_acc_11_psp_sva_1[4:2]==3'b000);
      COMP_LOOP_COMP_LOOP_and_258_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b000111);
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111) & (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b000);
      COMP_LOOP_COMP_LOOP_and_260_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b001001);
      COMP_LOOP_COMP_LOOP_and_261_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b001010);
      COMP_LOOP_COMP_LOOP_and_262_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b001011);
      COMP_LOOP_COMP_LOOP_and_10_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[2:1]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_264_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b001101);
      COMP_LOOP_COMP_LOOP_and_12_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[2])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2:1]!=2'b00)
          | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_13_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[2:1]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_14_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[0]) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
          & (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b00);
      COMP_LOOP_COMP_LOOP_and_268_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b010001);
      COMP_LOOP_COMP_LOOP_and_522_itm <= (COMP_LOOP_acc_11_psp_sva_1[3]) & (COMP_LOOP_acc_11_psp_sva_1[0])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_11_psp_sva_1[4]) | (COMP_LOOP_acc_11_psp_sva_1[2])
          | (COMP_LOOP_acc_11_psp_sva_1[1])));
      COMP_LOOP_COMP_LOOP_and_270_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b010011);
      COMP_LOOP_COMP_LOOP_and_18_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) | (COMP_LOOP_acc_psp_sva_mx0w0[0])
          | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_272_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b010101);
      COMP_LOOP_COMP_LOOP_and_20_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[2])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) |
          (COMP_LOOP_acc_psp_sva_mx0w0[0]) | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_21_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) | (COMP_LOOP_acc_psp_sva_mx0w0[0])
          | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_22_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1]) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) | (COMP_LOOP_acc_psp_sva_mx0w0[0])));
      COMP_LOOP_COMP_LOOP_and_23_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)));
      COMP_LOOP_COMP_LOOP_and_24_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) |
          (VEC_LOOP_j_10_0_sva_9_0[2:1]!=2'b00)));
      COMP_LOOP_COMP_LOOP_and_25_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[1]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) |
          (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_26_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2])
          | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_27_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2]) |
          (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)));
      COMP_LOOP_COMP_LOOP_and_28_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2]) & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2])
          | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_29_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11) & (~((COMP_LOOP_acc_psp_sva_mx0w0[2])
          | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_30_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111) & (~ (COMP_LOOP_acc_psp_sva_mx0w0[2]));
      COMP_LOOP_COMP_LOOP_and_284_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b100001);
      COMP_LOOP_COMP_LOOP_and_285_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b100010);
      COMP_LOOP_COMP_LOOP_and_286_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b100011);
      COMP_LOOP_COMP_LOOP_and_34_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_288_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[5:0]==6'b100101);
      COMP_LOOP_COMP_LOOP_and_36_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (VEC_LOOP_j_10_0_sva_9_0[2])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1:0]!=2'b00)
          | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_37_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[1:0]!=2'b00) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_38_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111)
          & (COMP_LOOP_acc_psp_sva_mx0w0[1:0]==2'b00);
      COMP_LOOP_COMP_LOOP_and_39_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)));
      COMP_LOOP_COMP_LOOP_and_40_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) |
          (VEC_LOOP_j_10_0_sva_9_0[2:1]!=2'b00)));
      COMP_LOOP_COMP_LOOP_and_41_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[1]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) |
          (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_42_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1])
          | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_43_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[2]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1]) |
          (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)));
      COMP_LOOP_COMP_LOOP_and_44_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[2]) & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1])
          | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_45_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11) & (~((COMP_LOOP_acc_psp_sva_mx0w0[1])
          | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_46_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2]) & (COMP_LOOP_acc_psp_sva_mx0w0[0])
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111) & (~ (COMP_LOOP_acc_psp_sva_mx0w0[1]));
      COMP_LOOP_COMP_LOOP_and_47_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) | (VEC_LOOP_j_10_0_sva_9_0[2:0]!=3'b000)));
      COMP_LOOP_COMP_LOOP_and_48_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) |
          (VEC_LOOP_j_10_0_sva_9_0[2:1]!=2'b00)));
      COMP_LOOP_COMP_LOOP_and_49_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[1]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) |
          (VEC_LOOP_j_10_0_sva_9_0[2]) | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_50_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[1:0]==2'b11) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0])
          | (VEC_LOOP_j_10_0_sva_9_0[2])));
      COMP_LOOP_COMP_LOOP_and_51_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0]) |
          (VEC_LOOP_j_10_0_sva_9_0[1:0]!=2'b00)));
      COMP_LOOP_COMP_LOOP_and_52_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2]) & (VEC_LOOP_j_10_0_sva_9_0[0]) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0])
          | (VEC_LOOP_j_10_0_sva_9_0[1])));
      COMP_LOOP_COMP_LOOP_and_53_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:1]==2'b11) & (~((COMP_LOOP_acc_psp_sva_mx0w0[0])
          | (VEC_LOOP_j_10_0_sva_9_0[0])));
      COMP_LOOP_COMP_LOOP_and_54_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:1]==2'b11)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111) & (~ (COMP_LOOP_acc_psp_sva_mx0w0[0]));
      COMP_LOOP_COMP_LOOP_and_55_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b000);
      COMP_LOOP_COMP_LOOP_and_56_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b001);
      COMP_LOOP_COMP_LOOP_and_57_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b010);
      COMP_LOOP_COMP_LOOP_and_58_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b011);
      COMP_LOOP_COMP_LOOP_and_59_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b100);
      COMP_LOOP_COMP_LOOP_and_60_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b101);
      COMP_LOOP_COMP_LOOP_and_61_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b110);
      COMP_LOOP_COMP_LOOP_and_62_itm <= (COMP_LOOP_acc_psp_sva_mx0w0[2:0]==3'b111)
          & (VEC_LOOP_j_10_0_sva_9_0[2:0]==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_73_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_74_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_75_itm <= 1'b0;
    end
    else if ( COMP_LOOP_or_121_cse ) begin
      COMP_LOOP_COMP_LOOP_and_73_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_73_nl,
          COMP_LOOP_COMP_LOOP_and_824_nl, and_dcpl_258);
      COMP_LOOP_COMP_LOOP_and_74_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_74_nl,
          COMP_LOOP_COMP_LOOP_and_851_nl, and_dcpl_258);
      COMP_LOOP_COMP_LOOP_and_75_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_75_nl,
          COMP_LOOP_COMP_LOOP_and_858_nl, and_dcpl_258);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_100_itm <= 1'b0;
    end
    else if ( ~(mux_3037_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_100_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_100_nl,
          COMP_LOOP_COMP_LOOP_and_323_nl, COMP_LOOP_COMP_LOOP_and_1073_nl, {and_dcpl_74
          , and_dcpl_261 , and_dcpl_370});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_101_itm <= 1'b0;
    end
    else if ( mux_3039_nl | (fsm_output[7]) ) begin
      COMP_LOOP_COMP_LOOP_and_101_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_101_nl,
          COMP_LOOP_COMP_LOOP_and_348_nl, COMP_LOOP_COMP_LOOP_and_1075_nl, {and_dcpl_74
          , and_dcpl_259 , and_403_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_102_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_109_itm <= 1'b0;
    end
    else if ( COMP_LOOP_or_126_cse ) begin
      COMP_LOOP_COMP_LOOP_and_102_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_102_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, COMP_LOOP_COMP_LOOP_and_1076_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_112});
      COMP_LOOP_COMP_LOOP_and_109_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_109_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_COMP_LOOP_and_1094_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_112});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_103_itm <= 1'b0;
    end
    else if ( ~(mux_3046_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_103_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_103_nl,
          COMP_LOOP_COMP_LOOP_and_350_nl, COMP_LOOP_COMP_LOOP_and_1079_nl, {and_dcpl_74
          , and_dcpl_261 , and_dcpl_375});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_104_itm <= 1'b0;
    end
    else if ( ~(mux_3047_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_104_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_104_nl,
          COMP_LOOP_COMP_LOOP_and_354_nl, COMP_LOOP_COMP_LOOP_and_1080_nl, {and_dcpl_74
          , and_dcpl_77 , and_409_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_105_itm <= 1'b0;
    end
    else if ( ~(mux_3048_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_105_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_105_nl,
          COMP_LOOP_COMP_LOOP_and_362_nl, COMP_LOOP_COMP_LOOP_and_1082_nl, {and_dcpl_74
          , and_dcpl_77 , and_dcpl_375});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_106_itm <= 1'b0;
    end
    else if ( ~(mux_3053_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_106_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_106_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_17_cse, COMP_LOOP_COMP_LOOP_and_1087_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_411_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_107_itm <= 1'b0;
    end
    else if ( mux_3059_nl | (fsm_output[7]) ) begin
      COMP_LOOP_COMP_LOOP_and_107_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_107_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_18_cse, COMP_LOOP_COMP_LOOP_and_1088_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_382});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_108_itm <= 1'b0;
    end
    else if ( ~(mux_3063_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_108_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_108_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_20_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_19_cse, COMP_LOOP_COMP_LOOP_and_1090_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_384});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_110_itm <= 1'b0;
    end
    else if ( mux_3064_nl | (fsm_output[7]) ) begin
      COMP_LOOP_COMP_LOOP_and_110_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_110_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_21_cse, COMP_LOOP_COMP_LOOP_and_1103_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_375});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_115_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_117_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_122_itm <= 1'b0;
    end
    else if ( COMP_LOOP_or_135_cse ) begin
      COMP_LOOP_COMP_LOOP_and_115_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_115_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse, COMP_LOOP_COMP_LOOP_and_1328_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_86});
      COMP_LOOP_COMP_LOOP_and_117_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_117_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse, COMP_LOOP_COMP_LOOP_and_1332_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_86});
      COMP_LOOP_COMP_LOOP_and_122_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_122_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse, COMP_LOOP_COMP_LOOP_and_1355_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_86});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_116_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3003, mux_3073_nl, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_116_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_116_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_28_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_27_cse, COMP_LOOP_COMP_LOOP_and_1331_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_90});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_118_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3081_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_118_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_118_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_29_cse, COMP_LOOP_COMP_LOOP_and_1334_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_384});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_119_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3085_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_119_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_COMP_LOOP_and_119_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse,
          COMP_LOOP_COMP_LOOP_and_1339_nl, {and_dcpl_74 , COMP_LOOP_or_110_rgt ,
          and_dcpl_261 , and_dcpl_265});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_120_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3092_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_120_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_120_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_30_cse, COMP_LOOP_COMP_LOOP_and_1340_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_387});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_121_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2((~ mux_3097_nl), (fsm_output[7]), fsm_output[6]) ) begin
      COMP_LOOP_COMP_LOOP_and_121_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_121_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_32_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_31_cse, COMP_LOOP_COMP_LOOP_and_1342_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_370});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_123_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3003, mux_742_cse, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_123_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_123_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_33_cse, COMP_LOOP_COMP_LOOP_and_1356_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_382});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_124_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3102_nl, (fsm_output[7]), fsm_output[6]) ) begin
      COMP_LOOP_COMP_LOOP_and_124_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_124_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_34_cse, COMP_LOOP_COMP_LOOP_and_1358_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_115});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_125_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3107_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_125_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_125_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_35_cse, COMP_LOOP_COMP_LOOP_and_1362_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_388});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 9'b000000000;
    end
    else if ( MUX_s_1_2_2(mux_3111_nl, and_705_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_14_psp_sva <= COMP_LOOP_acc_14_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 10'b0000000000;
    end
    else if ( mux_3115_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= COMP_LOOP_acc_1_cse_4_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 9'b000000000;
    end
    else if ( ~ and_dcpl_390 ) begin
      COMP_LOOP_acc_11_psp_sva <= COMP_LOOP_acc_11_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 10'b0000000000;
    end
    else if ( ~ and_dcpl_392 ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_2_sva <= 10'b0000000000;
    end
    else if ( ~(mux_3123_nl & nor_399_cse) ) begin
      COMP_LOOP_acc_10_cse_10_1_2_sva <= COMP_LOOP_2_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( ~(mux_3124_nl & nor_399_cse) ) begin
      COMP_LOOP_3_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_3_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_nor_5_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5:0]!=6'b000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_281_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_nor_281_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5:1]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_282_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_nor_282_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5]) | (COMP_LOOP_2_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[3]) | (COMP_LOOP_2_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_284_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_nor_284_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5]) | (COMP_LOOP_2_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[3]) | (COMP_LOOP_2_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_288_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_nor_288_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5]) | (COMP_LOOP_2_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[2]) | (COMP_LOOP_2_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_296_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_nor_296_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5]) | (COMP_LOOP_2_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[2]) | (COMP_LOOP_2_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_333_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_333_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_334_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_334_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_335_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_335_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_336_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_336_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_337_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_337_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_338_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_338_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_339_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_339_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_340_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_340_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_341_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_341_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_342_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_342_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_343_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_343_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_344_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_344_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_345_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_345_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b011111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_311_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_nor_311_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_347_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_347_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b100001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_349_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_349_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b100011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_351_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_351_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b100101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_352_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_352_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b100110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_353_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_353_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b100111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_355_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_355_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_356_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_356_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_357_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_357_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_358_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_358_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_359_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_359_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_360_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_360_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_361_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_361_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b101111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_363_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_363_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_364_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_364_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_365_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_365_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_366_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_366_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_367_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_367_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_368_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_368_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_369_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_369_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b110111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_370_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_370_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_371_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_371_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_372_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_372_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_373_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_373_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_374_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_374_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_375_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_375_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_376_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_376_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_377_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_396 ) begin
      COMP_LOOP_COMP_LOOP_and_377_itm <= (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_315_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_315_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4]) | (COMP_LOOP_2_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[1]) | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_289_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_289_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[5]) | (COMP_LOOP_2_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[2]) | (COMP_LOOP_2_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_313_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_313_itm <= ~((COMP_LOOP_2_acc_10_itm_10_1_1[4]) | (COMP_LOOP_2_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_2_acc_10_itm_10_1_1[2]) | (COMP_LOOP_2_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_3_sva <= 10'b0000000000;
    end
    else if ( mux_3126_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_10_cse_10_1_3_sva <= COMP_LOOP_3_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_3128_nl | (fsm_output[7]) ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_12_8_itm <= readslicef_9_1_8(COMP_LOOP_acc_12_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_nor_9_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5:0]!=6'b000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_505_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_nor_505_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5:1]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_506_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_nor_506_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5]) | (COMP_LOOP_3_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[3]) | (COMP_LOOP_3_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_569_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_569_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b000011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_508_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_nor_508_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5]) | (COMP_LOOP_3_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[3]) | (COMP_LOOP_3_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_571_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_571_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b000101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_572_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_572_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b000110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_573_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_573_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b000111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_512_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_nor_512_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5]) | (COMP_LOOP_3_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[2]) | (COMP_LOOP_3_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_575_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_575_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_576_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_576_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_577_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_577_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_578_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_578_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_579_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_579_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_580_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_580_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_581_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_581_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b001111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_520_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_nor_520_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5]) | (COMP_LOOP_3_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[2]) | (COMP_LOOP_3_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_584_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_584_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b010010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_585_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_585_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b010011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_586_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_586_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b010100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_587_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_587_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b010101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_588_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_588_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b010110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_589_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_589_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b010111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_590_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_590_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_591_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_591_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_592_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_592_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_593_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_593_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_594_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_594_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_595_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_595_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_596_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_596_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_597_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_597_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b011111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_535_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_nor_535_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_599_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_599_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_600_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_600_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_601_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_601_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_602_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_602_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_603_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_603_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_604_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_604_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_605_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_605_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b100111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_606_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_606_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_607_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_607_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_608_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_608_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_609_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_609_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_610_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_610_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_611_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_611_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_612_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_612_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_613_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_613_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b101111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_614_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_614_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_615_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_615_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_616_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_616_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_617_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_617_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_618_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_618_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_619_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_619_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_620_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_620_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_621_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_621_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b110111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_622_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_622_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_623_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_623_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_624_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_624_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_625_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_625_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_626_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_626_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_627_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_627_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_628_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_628_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_629_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_399 ) begin
      COMP_LOOP_COMP_LOOP_and_629_itm <= (COMP_LOOP_3_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_521_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_521_itm <= ~((COMP_LOOP_3_acc_10_itm_10_1_1[5]) | (COMP_LOOP_3_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_3_acc_10_itm_10_1_1[2]) | (COMP_LOOP_3_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_4_sva <= 10'b0000000000;
    end
    else if ( mux_3130_nl | (fsm_output[7]) ) begin
      COMP_LOOP_acc_10_cse_10_1_4_sva <= COMP_LOOP_4_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_3132_nl | (fsm_output[7]) ) begin
      COMP_LOOP_5_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_5_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_nor_13_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5:0]!=6'b000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_729_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_nor_729_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5:1]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_730_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_nor_730_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5]) | (COMP_LOOP_4_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[3]) | (COMP_LOOP_4_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_821_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_821_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b000011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_732_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_nor_732_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5]) | (COMP_LOOP_4_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[3]) | (COMP_LOOP_4_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_823_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_823_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b000101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_825_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_825_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b000111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_736_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_nor_736_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5]) | (COMP_LOOP_4_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[2]) | (COMP_LOOP_4_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_827_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_827_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_828_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_828_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_829_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_829_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_830_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_830_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_831_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_831_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_832_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_832_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_833_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_833_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b001111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_744_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_nor_744_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5]) | (COMP_LOOP_4_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[2]) | (COMP_LOOP_4_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_835_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_835_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_836_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_836_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_837_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_837_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_838_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_838_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_839_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_839_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_840_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_840_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_841_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_841_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b010111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_842_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_842_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_843_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_843_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_844_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_844_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_845_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_845_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_846_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_846_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_847_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_847_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_848_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_848_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_849_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_849_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b011111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_759_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_nor_759_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_852_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_852_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b100010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_853_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_853_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b100011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_854_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_854_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b100100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_855_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_855_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b100101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_856_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_856_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b100110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_857_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_857_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b100111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_859_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_859_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_860_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_860_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_861_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_861_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_862_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_862_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_863_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_863_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_864_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_864_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_865_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_865_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b101111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_866_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_866_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_867_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_867_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_868_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_868_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_869_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_869_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_870_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_870_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_871_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_871_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_872_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_872_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_873_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_873_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b110111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_874_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_874_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_875_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_875_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_876_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_876_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_877_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_877_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_878_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_878_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_879_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_879_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_880_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_880_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_881_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_402 ) begin
      COMP_LOOP_COMP_LOOP_and_881_itm <= (COMP_LOOP_4_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_767_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_767_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4]) | (COMP_LOOP_4_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[1]) | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_760_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_760_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_734_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_734_itm <= ~((COMP_LOOP_4_acc_10_itm_10_1_1[5]) | (COMP_LOOP_4_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_4_acc_10_itm_10_1_1[3]) | (COMP_LOOP_4_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 8'b00000000;
    end
    else if ( MUX_s_1_2_2(mux_3140_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_acc_13_psp_sva <= nl_COMP_LOOP_acc_13_psp_sva[7:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_5_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_3143_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_5_sva <= COMP_LOOP_5_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_3146_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_6_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_6_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_nor_17_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5:0]!=6'b000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_953_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_nor_953_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5:1]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_954_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_nor_954_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[3]) | (COMP_LOOP_5_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_956_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_nor_956_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[3]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1077_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1077_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b000111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_960_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_nor_960_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1081_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1081_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b001011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1083_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1083_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b001101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1084_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1084_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b001110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1085_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1085_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b001111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_968_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_nor_968_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1089_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1089_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b010011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1091_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1091_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b010101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1092_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1092_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b010110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1093_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1093_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b010111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1095_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1095_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1096_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1096_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1097_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1097_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1098_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1098_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1099_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1099_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1100_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1100_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1101_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1101_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b011111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_983_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_nor_983_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4:0]!=5'b00000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1105_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1105_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b100011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1107_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1107_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b100101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1108_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1108_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b100110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1109_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1109_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b100111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1111_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1111_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1112_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1112_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1113_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1113_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1114_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1114_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1115_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1115_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1116_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1116_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1117_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1117_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b101111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1119_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1119_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1120_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1120_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1121_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1121_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1122_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1122_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1123_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1123_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1124_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1124_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1125_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1125_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b110111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1126_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1126_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111000);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1127_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1127_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1128_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1128_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1129_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1129_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1130_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1130_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1131_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1131_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1132_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1132_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1133_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_403 ) begin
      COMP_LOOP_COMP_LOOP_and_1133_itm <= (COMP_LOOP_5_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_970_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_404 ) begin
      COMP_LOOP_nor_970_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_969_itm <= 1'b0;
    end
    else if ( ~(mux_3152_nl & nor_399_cse) ) begin
      COMP_LOOP_nor_969_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_984_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_406 ) begin
      COMP_LOOP_nor_984_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_964_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_406 ) begin
      COMP_LOOP_nor_964_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_961_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_406 ) begin
      COMP_LOOP_nor_961_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_955_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      COMP_LOOP_nor_955_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5:2]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_962_itm <= 1'b0;
    end
    else if ( ~(mux_3160_nl & nor_399_cse) ) begin
      COMP_LOOP_nor_962_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_957_itm <= 1'b0;
    end
    else if ( ~((mux_221_cse ^ (fsm_output[5])) & nor_399_cse) ) begin
      COMP_LOOP_nor_957_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[3]) | (COMP_LOOP_5_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_976_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_976_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_958_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_958_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[3]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_998_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_998_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_972_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_972_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[5]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_987_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_987_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_985_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_985_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4]) | (COMP_LOOP_5_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[2]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_140_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_nor_140_itm <= COMP_LOOP_tmp_nor_140_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_141_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_nor_141_itm <= COMP_LOOP_tmp_nor_141_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm <= (z_out_7[1:0]==2'b11) & COMP_LOOP_tmp_nor_76_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_143_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_nor_143_itm <= COMP_LOOP_tmp_nor_77_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm <= (z_out_7[2]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_78_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm <= (z_out_7[2:1]==2'b11) & COMP_LOOP_tmp_nor_79_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm <= (z_out_7[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_nor_146_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_nor_146_itm <= COMP_LOOP_tmp_nor_80_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm <= (z_out_7[3]) & (z_out_7[0]) & COMP_LOOP_tmp_nor_81_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm <= (z_out_7[3]) & (z_out_7[1]) & COMP_LOOP_tmp_nor_82_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm <= (z_out_7[3:0]==4'b1011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm <= (z_out_7[3:2]==2'b11) & COMP_LOOP_tmp_nor_83_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm <= (z_out_7[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm <= (z_out_7[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm <= (z_out_7[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_991_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_991_itm <= ~((COMP_LOOP_5_acc_10_itm_10_1_1[4]) | (COMP_LOOP_5_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_5_acc_10_itm_10_1_1[1]) | (COMP_LOOP_5_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_3163_nl, (fsm_output[7]), fsm_output[6]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= nl_COMP_LOOP_acc_1_cse_6_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_6_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3102, and_736_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_6_sva <= COMP_LOOP_6_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_tmp_3102, mux_3171_nl, fsm_output[5]) ) begin
      COMP_LOOP_7_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_7_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= 1'b0;
      COMP_LOOP_nor_1177_itm <= 1'b0;
      COMP_LOOP_nor_1178_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1325_itm <= 1'b0;
      COMP_LOOP_nor_1180_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1327_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1329_itm <= 1'b0;
      COMP_LOOP_nor_1184_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1333_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1335_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1336_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1337_itm <= 1'b0;
      COMP_LOOP_nor_1192_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1341_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1343_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1344_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1345_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1346_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1347_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1348_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1349_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1350_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1351_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1352_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1353_itm <= 1'b0;
      COMP_LOOP_nor_1207_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1357_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1359_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1360_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1361_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1363_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1364_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1365_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1366_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1367_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1368_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1369_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1371_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1372_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1373_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1374_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1375_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1376_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1377_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1378_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1379_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1380_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1381_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1382_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1383_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1384_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1385_itm <= 1'b0;
    end
    else if ( mux_3175_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_21_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5:0]!=6'b000000));
      COMP_LOOP_nor_1177_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5:1]!=5'b00000));
      COMP_LOOP_nor_1178_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[3]) | (COMP_LOOP_6_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1325_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b000011);
      COMP_LOOP_nor_1180_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[3]) | (COMP_LOOP_6_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1327_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b000101);
      COMP_LOOP_COMP_LOOP_and_1329_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b000111);
      COMP_LOOP_nor_1184_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1333_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b001011);
      COMP_LOOP_COMP_LOOP_and_1335_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b001101);
      COMP_LOOP_COMP_LOOP_and_1336_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b001110);
      COMP_LOOP_COMP_LOOP_and_1337_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b001111);
      COMP_LOOP_nor_1192_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1341_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b010011);
      COMP_LOOP_COMP_LOOP_and_1343_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b010101);
      COMP_LOOP_COMP_LOOP_and_1344_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b010110);
      COMP_LOOP_COMP_LOOP_and_1345_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b010111);
      COMP_LOOP_COMP_LOOP_and_1346_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011000);
      COMP_LOOP_COMP_LOOP_and_1347_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011001);
      COMP_LOOP_COMP_LOOP_and_1348_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011010);
      COMP_LOOP_COMP_LOOP_and_1349_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011011);
      COMP_LOOP_COMP_LOOP_and_1350_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011100);
      COMP_LOOP_COMP_LOOP_and_1351_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011101);
      COMP_LOOP_COMP_LOOP_and_1352_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011110);
      COMP_LOOP_COMP_LOOP_and_1353_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b011111);
      COMP_LOOP_nor_1207_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4:0]!=5'b00000));
      COMP_LOOP_COMP_LOOP_and_1357_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b100011);
      COMP_LOOP_COMP_LOOP_and_1359_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b100101);
      COMP_LOOP_COMP_LOOP_and_1360_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b100110);
      COMP_LOOP_COMP_LOOP_and_1361_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b100111);
      COMP_LOOP_COMP_LOOP_and_1363_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101001);
      COMP_LOOP_COMP_LOOP_and_1364_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101010);
      COMP_LOOP_COMP_LOOP_and_1365_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101011);
      COMP_LOOP_COMP_LOOP_and_1366_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101100);
      COMP_LOOP_COMP_LOOP_and_1367_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101101);
      COMP_LOOP_COMP_LOOP_and_1368_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101110);
      COMP_LOOP_COMP_LOOP_and_1369_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b101111);
      COMP_LOOP_COMP_LOOP_and_1371_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110001);
      COMP_LOOP_COMP_LOOP_and_1372_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110010);
      COMP_LOOP_COMP_LOOP_and_1373_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110011);
      COMP_LOOP_COMP_LOOP_and_1374_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110100);
      COMP_LOOP_COMP_LOOP_and_1375_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110101);
      COMP_LOOP_COMP_LOOP_and_1376_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110110);
      COMP_LOOP_COMP_LOOP_and_1377_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b110111);
      COMP_LOOP_COMP_LOOP_and_1378_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111000);
      COMP_LOOP_COMP_LOOP_and_1379_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111001);
      COMP_LOOP_COMP_LOOP_and_1380_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111010);
      COMP_LOOP_COMP_LOOP_and_1381_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111011);
      COMP_LOOP_COMP_LOOP_and_1382_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111100);
      COMP_LOOP_COMP_LOOP_and_1383_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111101);
      COMP_LOOP_COMP_LOOP_and_1384_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111110);
      COMP_LOOP_COMP_LOOP_and_1385_itm <= (COMP_LOOP_6_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1185_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_410 ) begin
      COMP_LOOP_nor_1185_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1211_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_392 ) begin
      COMP_LOOP_nor_1211_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[1]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1209_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_404 ) begin
      COMP_LOOP_nor_1209_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1196_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      COMP_LOOP_nor_1196_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[1]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1208_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_411 ) begin
      COMP_LOOP_nor_1208_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1186_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_411 ) begin
      COMP_LOOP_nor_1186_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1182_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_411 ) begin
      COMP_LOOP_nor_1182_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[3]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1222_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1222_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1188_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1188_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[1]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1215_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1215_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[4]) | (COMP_LOOP_6_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[1]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1194_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1194_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1193_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1193_itm <= ~((COMP_LOOP_6_acc_10_itm_10_1_1[5]) | (COMP_LOOP_6_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_6_acc_10_itm_10_1_1[2]) | (COMP_LOOP_6_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_7_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_3182_nl, and_705_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_7_sva <= COMP_LOOP_7_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( mux_3185_itm ) begin
      COMP_LOOP_slc_COMP_LOOP_acc_15_7_itm <= readslicef_8_1_7(COMP_LOOP_acc_15_nl);
      reg_COMP_LOOP_k_10_3_ftd <= z_out_2[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= 1'b0;
      COMP_LOOP_nor_1401_itm <= 1'b0;
      COMP_LOOP_nor_1402_itm <= 1'b0;
      COMP_LOOP_nor_1404_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1579_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1580_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1581_itm <= 1'b0;
      COMP_LOOP_nor_1408_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1583_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1585_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1586_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1587_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1588_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1589_itm <= 1'b0;
      COMP_LOOP_nor_1416_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1591_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1592_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1593_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1595_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1596_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1597_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1599_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1600_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1601_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1602_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1603_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1604_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1605_itm <= 1'b0;
      COMP_LOOP_nor_1431_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1608_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1609_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1611_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1612_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1613_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1615_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1616_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1617_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1618_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1619_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1620_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1621_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1623_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1624_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1625_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1626_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1627_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1628_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1629_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1630_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1631_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1632_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1633_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1634_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1635_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1636_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1637_itm <= 1'b0;
    end
    else if ( mux_3187_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_25_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5:0]!=6'b000000));
      COMP_LOOP_nor_1401_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5:1]!=5'b00000));
      COMP_LOOP_nor_1402_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[3]) | (COMP_LOOP_7_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_nor_1404_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[3]) | (COMP_LOOP_7_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1579_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b000101);
      COMP_LOOP_COMP_LOOP_and_1580_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b000110);
      COMP_LOOP_COMP_LOOP_and_1581_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b000111);
      COMP_LOOP_nor_1408_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[2]) | (COMP_LOOP_7_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1583_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b001001);
      COMP_LOOP_COMP_LOOP_and_1585_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b001011);
      COMP_LOOP_COMP_LOOP_and_1586_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b001100);
      COMP_LOOP_COMP_LOOP_and_1587_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b001101);
      COMP_LOOP_COMP_LOOP_and_1588_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b001110);
      COMP_LOOP_COMP_LOOP_and_1589_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b001111);
      COMP_LOOP_nor_1416_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[2]) | (COMP_LOOP_7_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1591_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b010001);
      COMP_LOOP_COMP_LOOP_and_1592_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b010010);
      COMP_LOOP_COMP_LOOP_and_1593_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b010011);
      COMP_LOOP_COMP_LOOP_and_1595_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b010101);
      COMP_LOOP_COMP_LOOP_and_1596_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b010110);
      COMP_LOOP_COMP_LOOP_and_1597_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b010111);
      COMP_LOOP_COMP_LOOP_and_1599_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011001);
      COMP_LOOP_COMP_LOOP_and_1600_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011010);
      COMP_LOOP_COMP_LOOP_and_1601_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011011);
      COMP_LOOP_COMP_LOOP_and_1602_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011100);
      COMP_LOOP_COMP_LOOP_and_1603_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011101);
      COMP_LOOP_COMP_LOOP_and_1604_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011110);
      COMP_LOOP_COMP_LOOP_and_1605_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b011111);
      COMP_LOOP_nor_1431_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4:0]!=5'b00000));
      COMP_LOOP_COMP_LOOP_and_1608_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b100010);
      COMP_LOOP_COMP_LOOP_and_1609_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b100011);
      COMP_LOOP_COMP_LOOP_and_1611_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b100101);
      COMP_LOOP_COMP_LOOP_and_1612_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b100110);
      COMP_LOOP_COMP_LOOP_and_1613_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b100111);
      COMP_LOOP_COMP_LOOP_and_1615_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101001);
      COMP_LOOP_COMP_LOOP_and_1616_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101010);
      COMP_LOOP_COMP_LOOP_and_1617_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101011);
      COMP_LOOP_COMP_LOOP_and_1618_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101100);
      COMP_LOOP_COMP_LOOP_and_1619_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101101);
      COMP_LOOP_COMP_LOOP_and_1620_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101110);
      COMP_LOOP_COMP_LOOP_and_1621_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b101111);
      COMP_LOOP_COMP_LOOP_and_1623_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110001);
      COMP_LOOP_COMP_LOOP_and_1624_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110010);
      COMP_LOOP_COMP_LOOP_and_1625_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110011);
      COMP_LOOP_COMP_LOOP_and_1626_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110100);
      COMP_LOOP_COMP_LOOP_and_1627_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110101);
      COMP_LOOP_COMP_LOOP_and_1628_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110110);
      COMP_LOOP_COMP_LOOP_and_1629_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b110111);
      COMP_LOOP_COMP_LOOP_and_1630_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111000);
      COMP_LOOP_COMP_LOOP_and_1631_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111001);
      COMP_LOOP_COMP_LOOP_and_1632_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111010);
      COMP_LOOP_COMP_LOOP_and_1633_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111011);
      COMP_LOOP_COMP_LOOP_and_1634_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111100);
      COMP_LOOP_COMP_LOOP_and_1635_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111101);
      COMP_LOOP_COMP_LOOP_and_1636_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111110);
      COMP_LOOP_COMP_LOOP_and_1637_itm <= (COMP_LOOP_7_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1435_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_390 ) begin
      COMP_LOOP_nor_1435_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4]) | (COMP_LOOP_7_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[1]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1446_itm <= 1'b0;
    end
    else if ( ~(mux_3188_nl & nor_399_cse) ) begin
      COMP_LOOP_nor_1446_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1439_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_410 ) begin
      COMP_LOOP_nor_1439_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4]) | (COMP_LOOP_7_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[1]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1420_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_410 ) begin
      COMP_LOOP_nor_1420_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[1]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1432_itm <= 1'b0;
    end
    else if ( ~(mux_3192_nl & nor_399_cse) ) begin
      COMP_LOOP_nor_1432_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[4:1]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1424_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_407 ) begin
      COMP_LOOP_nor_1424_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[1]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1410_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1410_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5]) | (COMP_LOOP_7_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_7_acc_10_itm_10_1_1[2]) | (COMP_LOOP_7_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1403_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1403_itm <= ~((COMP_LOOP_7_acc_10_itm_10_1_1[5:2]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_811, mux_3193_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[9:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_10_1_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(not_tmp_811, and_705_cse, fsm_output[5]) ) begin
      COMP_LOOP_acc_10_cse_10_1_sva <= COMP_LOOP_8_acc_10_itm_10_1_1;
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(not_tmp_811, mux_3197_nl, fsm_output[5]) ) begin
      COMP_LOOP_1_slc_COMP_LOOP_acc_10_itm <= readslicef_11_1_10(COMP_LOOP_1_acc_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= 1'b0;
      COMP_LOOP_nor_1625_itm <= 1'b0;
      COMP_LOOP_nor_1626_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1829_itm <= 1'b0;
      COMP_LOOP_nor_1628_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1833_itm <= 1'b0;
      COMP_LOOP_nor_1632_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1836_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1837_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1838_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1839_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1840_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1841_itm <= 1'b0;
      COMP_LOOP_nor_1640_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1843_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1845_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1846_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1847_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1848_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1849_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1851_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1852_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1853_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1854_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1855_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1856_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1857_itm <= 1'b0;
      COMP_LOOP_nor_1655_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1859_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1860_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1861_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1863_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1864_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1865_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1867_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1868_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1869_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1870_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1871_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1872_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1873_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1875_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1876_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1877_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1878_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1879_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1880_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1881_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1882_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1883_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1884_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1885_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1886_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1887_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1888_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1889_itm <= 1'b0;
    end
    else if ( mux_3201_itm ) begin
      COMP_LOOP_COMP_LOOP_nor_29_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5:0]!=6'b000000));
      COMP_LOOP_nor_1625_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5:1]!=5'b00000));
      COMP_LOOP_nor_1626_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[3]) | (COMP_LOOP_8_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1829_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b000011);
      COMP_LOOP_nor_1628_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[3]) | (COMP_LOOP_8_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1833_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b000111);
      COMP_LOOP_nor_1632_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[2]) | (COMP_LOOP_8_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1836_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b001010);
      COMP_LOOP_COMP_LOOP_and_1837_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b001011);
      COMP_LOOP_COMP_LOOP_and_1838_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b001100);
      COMP_LOOP_COMP_LOOP_and_1839_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b001101);
      COMP_LOOP_COMP_LOOP_and_1840_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b001110);
      COMP_LOOP_COMP_LOOP_and_1841_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b001111);
      COMP_LOOP_nor_1640_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[2]) | (COMP_LOOP_8_acc_10_itm_10_1_1[1])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
      COMP_LOOP_COMP_LOOP_and_1843_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b010001);
      COMP_LOOP_COMP_LOOP_and_1845_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b010011);
      COMP_LOOP_COMP_LOOP_and_1846_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b010100);
      COMP_LOOP_COMP_LOOP_and_1847_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b010101);
      COMP_LOOP_COMP_LOOP_and_1848_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b010110);
      COMP_LOOP_COMP_LOOP_and_1849_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b010111);
      COMP_LOOP_COMP_LOOP_and_1851_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011001);
      COMP_LOOP_COMP_LOOP_and_1852_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011010);
      COMP_LOOP_COMP_LOOP_and_1853_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011011);
      COMP_LOOP_COMP_LOOP_and_1854_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011100);
      COMP_LOOP_COMP_LOOP_and_1855_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011101);
      COMP_LOOP_COMP_LOOP_and_1856_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011110);
      COMP_LOOP_COMP_LOOP_and_1857_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b011111);
      COMP_LOOP_nor_1655_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4:0]!=5'b00000));
      COMP_LOOP_COMP_LOOP_and_1859_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b100001);
      COMP_LOOP_COMP_LOOP_and_1860_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b100010);
      COMP_LOOP_COMP_LOOP_and_1861_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b100011);
      COMP_LOOP_COMP_LOOP_and_1863_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b100101);
      COMP_LOOP_COMP_LOOP_and_1864_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b100110);
      COMP_LOOP_COMP_LOOP_and_1865_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b100111);
      COMP_LOOP_COMP_LOOP_and_1867_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101001);
      COMP_LOOP_COMP_LOOP_and_1868_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101010);
      COMP_LOOP_COMP_LOOP_and_1869_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101011);
      COMP_LOOP_COMP_LOOP_and_1870_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101100);
      COMP_LOOP_COMP_LOOP_and_1871_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101101);
      COMP_LOOP_COMP_LOOP_and_1872_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101110);
      COMP_LOOP_COMP_LOOP_and_1873_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b101111);
      COMP_LOOP_COMP_LOOP_and_1875_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110001);
      COMP_LOOP_COMP_LOOP_and_1876_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110010);
      COMP_LOOP_COMP_LOOP_and_1877_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110011);
      COMP_LOOP_COMP_LOOP_and_1878_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110100);
      COMP_LOOP_COMP_LOOP_and_1879_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110101);
      COMP_LOOP_COMP_LOOP_and_1880_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110110);
      COMP_LOOP_COMP_LOOP_and_1881_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b110111);
      COMP_LOOP_COMP_LOOP_and_1882_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111000);
      COMP_LOOP_COMP_LOOP_and_1883_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111001);
      COMP_LOOP_COMP_LOOP_and_1884_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111010);
      COMP_LOOP_COMP_LOOP_and_1885_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111011);
      COMP_LOOP_COMP_LOOP_and_1886_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111100);
      COMP_LOOP_COMP_LOOP_and_1887_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111101);
      COMP_LOOP_COMP_LOOP_and_1888_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111110);
      COMP_LOOP_COMP_LOOP_and_1889_itm <= (COMP_LOOP_8_acc_10_itm_10_1_1[5:0]==6'b111111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1663_itm <= 1'b0;
    end
    else if ( mux_3205_nl | (fsm_output[7]) ) begin
      COMP_LOOP_nor_1663_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4]) | (COMP_LOOP_8_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[1]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1659_itm <= 1'b0;
    end
    else if ( mux_3210_nl | (fsm_output[7]) ) begin
      COMP_LOOP_nor_1659_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[4]) | (COMP_LOOP_8_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[1]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1633_itm <= 1'b0;
    end
    else if ( mux_3216_nl | (fsm_output[7]) ) begin
      COMP_LOOP_nor_1633_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[2]) | (COMP_LOOP_8_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1642_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_410 ) begin
      COMP_LOOP_nor_1642_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[3])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[2]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1648_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_404 ) begin
      COMP_LOOP_nor_1648_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[2])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[1]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1630_itm <= 1'b0;
    end
    else if ( ~(mux_3219_nl & nor_399_cse) ) begin
      COMP_LOOP_nor_1630_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[3]) | (COMP_LOOP_8_acc_10_itm_10_1_1[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1670_itm <= 1'b0;
    end
    else if ( ~ and_dcpl_411 ) begin
      COMP_LOOP_nor_1670_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_nor_1629_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_125 ) begin
      COMP_LOOP_nor_1629_itm <= ~((COMP_LOOP_8_acc_10_itm_10_1_1[5]) | (COMP_LOOP_8_acc_10_itm_10_1_1[4])
          | (COMP_LOOP_8_acc_10_itm_10_1_1[3]) | (COMP_LOOP_8_acc_10_itm_10_1_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1104_itm <= 1'b0;
    end
    else if ( ~(mux_3223_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_1104_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_111_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_23_cse, COMP_LOOP_COMP_LOOP_and_1104_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_387});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1106_itm <= 1'b0;
    end
    else if ( ~(mux_3226_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_1106_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_112_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_24_cse, COMP_LOOP_COMP_LOOP_and_1106_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_388});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1110_itm <= 1'b0;
    end
    else if ( ~(mux_3227_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_1110_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_113_nl,
          COMP_LOOP_COMP_LOOP_and_1110_nl, and_dcpl_261);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1118_itm <= 1'b0;
    end
    else if ( ~(mux_3229_nl & (~ (fsm_output[7]))) ) begin
      COMP_LOOP_COMP_LOOP_and_1118_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_114_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_120_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_25_cse, COMP_LOOP_COMP_LOOP_and_1118_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_421});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1370_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3231_nl, (fsm_output[7]), fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1370_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_65_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_36_cse, COMP_LOOP_COMP_LOOP_and_1370_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_421});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1577_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1584_itm <= 1'b0;
    end
    else if ( COMP_LOOP_or_151_cse ) begin
      COMP_LOOP_COMP_LOOP_and_1577_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_67_nl,
          COMP_LOOP_COMP_LOOP_and_1577_nl, and_dcpl_258);
      COMP_LOOP_COMP_LOOP_and_1584_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_68_nl,
          COMP_LOOP_COMP_LOOP_and_1584_nl, and_dcpl_258);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1594_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_1614_itm <= 1'b0;
    end
    else if ( COMP_LOOP_or_153_cse ) begin
      COMP_LOOP_COMP_LOOP_and_1594_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_317_nl,
          COMP_LOOP_COMP_LOOP_and_1594_nl, and_dcpl_90);
      COMP_LOOP_COMP_LOOP_and_1614_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_324_nl,
          COMP_LOOP_COMP_LOOP_and_1614_nl, and_dcpl_90);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1598_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3243_nl, (fsm_output[7]), fsm_output[6]) ) begin
      COMP_LOOP_COMP_LOOP_and_1598_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_319_nl,
          COMP_LOOP_COMP_LOOP_and_1598_nl, and_dcpl_370);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1607_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3102, mux_3246_nl, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1607_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_320_nl,
          COMP_LOOP_COMP_LOOP_and_1607_nl, and_458_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1610_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3253_nl, mux_3249_nl, fsm_output[6]) ) begin
      COMP_LOOP_COMP_LOOP_and_1610_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_321_nl,
          COMP_LOOP_COMP_LOOP_and_1610_nl, and_dcpl_118);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1622_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3102, mux_3256_nl, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1622_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_325_nl,
          COMP_LOOP_COMP_LOOP_and_1622_nl, and_459_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1831_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3264_nl, and_705_cse, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1831_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_69_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_37_cse, COMP_LOOP_COMP_LOOP_and_1831_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_112});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1832_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3274_nl, mux_3267_nl, fsm_output[3]) ) begin
      COMP_LOOP_COMP_LOOP_and_1832_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_326_nl,
          COMP_LOOP_COMP_LOOP_and_1832_nl, and_461_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1835_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3283_nl, mux_297_cse, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1835_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_327_nl,
          COMP_LOOP_COMP_LOOP_and_1835_nl, and_463_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1844_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3133, mux_3286_nl, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1844_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_328_nl,
          COMP_LOOP_COMP_LOOP_and_1844_nl, and_dcpl_90);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1850_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3133, mux_tmp_3218, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1850_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_329_nl,
          COMP_LOOP_COMP_LOOP_and_1850_nl, and_dcpl_382);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1862_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3292_nl, mux_297_cse, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1862_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_331_nl,
          COMP_LOOP_COMP_LOOP_and_1862_nl, and_465_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1866_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3298_nl, mux_297_cse, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1866_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_332_nl,
          COMP_LOOP_COMP_LOOP_and_1866_nl, and_468_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_1874_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3302_nl, and_705_cse, fsm_output[5]) ) begin
      COMP_LOOP_COMP_LOOP_and_1874_itm <= MUX1HOT_s_1_5_2(COMP_LOOP_COMP_LOOP_and_71_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_39_cse, COMP_LOOP_COMP_LOOP_and_1874_nl,
          {and_dcpl_74 , and_dcpl_77 , and_dcpl_258 , COMP_LOOP_or_120_rgt , and_dcpl_86});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_583_itm <= 1'b0;
    end
    else if ( ~(mux_3306_nl & nor_399_cse) ) begin
      COMP_LOOP_COMP_LOOP_and_583_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_72_nl,
          COMP_LOOP_COMP_LOOP_and_583_nl, and_dcpl_258);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse, {and_dcpl_74 , and_dcpl_77 , and_dcpl_258
          , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_244_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_11_cse, {and_dcpl_74 , and_dcpl_77 , and_dcpl_258
          , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_12_cse, {and_dcpl_74 , and_dcpl_77 , and_dcpl_258
          , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_13_cse, {and_dcpl_74 , and_dcpl_77 , and_dcpl_258
          , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_tmp_COMP_LOOP_tmp_nor_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_110_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_15_cse, {and_dcpl_74 , and_dcpl_77 , and_dcpl_258
          , COMP_LOOP_or_120_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= 1'b0;
      COMP_LOOP_tmp_nor_10_itm <= 1'b0;
      COMP_LOOP_tmp_nor_151_itm <= 1'b0;
      COMP_LOOP_tmp_nor_153_itm <= 1'b0;
      COMP_LOOP_tmp_nor_157_itm <= 1'b0;
      COMP_LOOP_tmp_nor_165_itm <= 1'b0;
      COMP_LOOP_tmp_nor_180_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_5_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_76_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_40_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_77_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_41_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_79_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_42_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_80_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_43_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_81_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_44_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_82_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_45_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_83_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_46_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_84_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_47_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_85_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_48_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_86_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_49_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_87_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_50_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_88_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_51_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_89_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_52_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_90_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_53_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_91_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_54_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_92_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_55_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_93_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_56_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_95_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_57_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_96_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_58_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_97_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_59_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_98_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_60_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_and_99_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_61_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm <= MUX1HOT_s_1_3_2(COMP_LOOP_COMP_LOOP_nor_1_nl,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_and_62_cse,
          {and_dcpl_74 , and_dcpl_77 , COMP_LOOP_or_120_rgt});
      COMP_LOOP_tmp_nor_10_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_57_nl, COMP_LOOP_tmp_nor_10_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, COMP_LOOP_tmp_nor_150_cse, {and_dcpl_74
          , and_dcpl_77 , and_dcpl_259 , COMP_LOOP_or_74_cse});
      COMP_LOOP_tmp_nor_151_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_58_nl, COMP_LOOP_tmp_nor_18_cse,
          COMP_LOOP_tmp_nor_150_cse, COMP_LOOP_tmp_nor_151_cse, {and_dcpl_74 , and_dcpl_77
          , and_dcpl_259 , COMP_LOOP_or_74_cse});
      COMP_LOOP_tmp_nor_153_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_60_nl, COMP_LOOP_tmp_nor_150_cse,
          COMP_LOOP_tmp_nor_151_cse, COMP_LOOP_tmp_nor_153_cse, {and_dcpl_74 , and_dcpl_77
          , and_dcpl_259 , COMP_LOOP_or_74_cse});
      COMP_LOOP_tmp_nor_157_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_64_nl, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse,
          COMP_LOOP_tmp_nor_153_cse, COMP_LOOP_tmp_nor_10_cse, {and_dcpl_74 , and_dcpl_77
          , and_dcpl_259 , COMP_LOOP_or_74_cse});
      COMP_LOOP_tmp_nor_165_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_72_nl, COMP_LOOP_tmp_nor_151_cse,
          COMP_LOOP_tmp_nor_10_cse, COMP_LOOP_tmp_nor_18_cse, {and_dcpl_74 , and_dcpl_77
          , and_dcpl_259 , COMP_LOOP_or_74_cse});
      COMP_LOOP_tmp_nor_180_itm <= MUX1HOT_s_1_4_2(COMP_LOOP_nor_87_nl, COMP_LOOP_tmp_nor_153_cse,
          COMP_LOOP_tmp_nor_18_cse, COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse, {and_dcpl_74
          , and_dcpl_77 , and_dcpl_259 , COMP_LOOP_or_74_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_2_tmp_mul_idiv_sva <= 10'b0000000000;
    end
    else if ( and_dcpl_77 | and_dcpl_259 | and_dcpl_260 ) begin
      COMP_LOOP_2_tmp_mul_idiv_sva <= z_out_7;
    end
  end
  always @(posedge clk) begin
    if ( ~(or_dcpl_134 | or_dcpl_122) ) begin
      COMP_LOOP_tmp_mux1h_itm <= MUX1HOT_v_64_8_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_8_i_q_d,
          twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_32_i_q_d,
          twiddle_rsc_0_40_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_56_i_q_d,
          {COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm , COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_2_tmp_lshift_ncse_sva <= 10'b0000000000;
    end
    else if ( and_dcpl_77 | and_dcpl_263 ) begin
      COMP_LOOP_2_tmp_lshift_ncse_sva <= MUX_v_10_2_2(z_out_1, z_out_7, and_dcpl_263);
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_77 | and_dcpl_258 | and_dcpl_432 | and_dcpl_263 | COMP_LOOP_1_acc_8_itm_mx0c4
        | and_dcpl_86 | and_dcpl_343 | and_dcpl_90 | and_dcpl_346 | and_dcpl_95 |
        and_dcpl_349 | and_dcpl_99 | and_dcpl_351 | and_dcpl_104 | and_dcpl_354 |
        and_dcpl_106 | and_dcpl_357 | and_dcpl_109 | and_dcpl_359 ) begin
      COMP_LOOP_1_acc_8_itm <= MUX1HOT_v_64_68_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d,
          vec_rsc_0_2_i_q_d, vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d,
          vec_rsc_0_6_i_q_d, vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d,
          vec_rsc_0_10_i_q_d, vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d,
          vec_rsc_0_14_i_q_d, vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d,
          vec_rsc_0_18_i_q_d, vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d,
          vec_rsc_0_22_i_q_d, vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d,
          vec_rsc_0_26_i_q_d, vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d,
          vec_rsc_0_30_i_q_d, vec_rsc_0_31_i_q_d, vec_rsc_0_32_i_q_d, vec_rsc_0_33_i_q_d,
          vec_rsc_0_34_i_q_d, vec_rsc_0_35_i_q_d, vec_rsc_0_36_i_q_d, vec_rsc_0_37_i_q_d,
          vec_rsc_0_38_i_q_d, vec_rsc_0_39_i_q_d, vec_rsc_0_40_i_q_d, vec_rsc_0_41_i_q_d,
          vec_rsc_0_42_i_q_d, vec_rsc_0_43_i_q_d, vec_rsc_0_44_i_q_d, vec_rsc_0_45_i_q_d,
          vec_rsc_0_46_i_q_d, vec_rsc_0_47_i_q_d, vec_rsc_0_48_i_q_d, vec_rsc_0_49_i_q_d,
          vec_rsc_0_50_i_q_d, vec_rsc_0_51_i_q_d, vec_rsc_0_52_i_q_d, vec_rsc_0_53_i_q_d,
          vec_rsc_0_54_i_q_d, vec_rsc_0_55_i_q_d, vec_rsc_0_56_i_q_d, vec_rsc_0_57_i_q_d,
          vec_rsc_0_58_i_q_d, vec_rsc_0_59_i_q_d, vec_rsc_0_60_i_q_d, vec_rsc_0_61_i_q_d,
          vec_rsc_0_62_i_q_d, vec_rsc_0_63_i_q_d, COMP_LOOP_acc_17_nl, twiddle_rsc_0_10_i_q_d,
          twiddle_rsc_0_26_i_q_d, COMP_LOOP_1_modulo_dev_cmp_return_rsc_z, {COMP_LOOP_or_nl
          , COMP_LOOP_or_1_nl , COMP_LOOP_or_2_nl , COMP_LOOP_or_3_nl , COMP_LOOP_or_4_nl
          , COMP_LOOP_or_5_nl , COMP_LOOP_or_6_nl , COMP_LOOP_or_7_nl , COMP_LOOP_or_8_nl
          , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl
          , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl , COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl
          , COMP_LOOP_or_17_nl , COMP_LOOP_or_18_nl , COMP_LOOP_or_19_nl , COMP_LOOP_or_20_nl
          , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl , COMP_LOOP_or_23_nl , COMP_LOOP_or_24_nl
          , COMP_LOOP_or_25_nl , COMP_LOOP_or_26_nl , COMP_LOOP_or_27_nl , COMP_LOOP_or_28_nl
          , COMP_LOOP_or_29_nl , COMP_LOOP_or_30_nl , COMP_LOOP_or_31_nl , COMP_LOOP_or_32_nl
          , COMP_LOOP_or_33_nl , COMP_LOOP_or_34_nl , COMP_LOOP_or_35_nl , COMP_LOOP_or_36_nl
          , COMP_LOOP_or_37_nl , COMP_LOOP_or_38_nl , COMP_LOOP_or_39_nl , COMP_LOOP_or_40_nl
          , COMP_LOOP_or_41_nl , COMP_LOOP_or_42_nl , COMP_LOOP_or_43_nl , COMP_LOOP_or_44_nl
          , COMP_LOOP_or_45_nl , COMP_LOOP_or_46_nl , COMP_LOOP_or_47_nl , COMP_LOOP_or_48_nl
          , COMP_LOOP_or_49_nl , COMP_LOOP_or_50_nl , COMP_LOOP_or_51_nl , COMP_LOOP_or_52_nl
          , COMP_LOOP_or_53_nl , COMP_LOOP_or_54_nl , COMP_LOOP_or_55_nl , COMP_LOOP_or_56_nl
          , COMP_LOOP_or_57_nl , COMP_LOOP_or_58_nl , COMP_LOOP_or_59_nl , COMP_LOOP_or_60_nl
          , COMP_LOOP_or_61_nl , COMP_LOOP_or_62_nl , COMP_LOOP_or_63_nl , COMP_LOOP_or_68_itm
          , and_dcpl_432 , and_dcpl_263 , COMP_LOOP_1_acc_8_itm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= 1'b0;
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_36_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_63_cse, COMP_LOOP_or_120_rgt);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_64_cse, COMP_LOOP_or_120_rgt);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_65_cse, COMP_LOOP_or_120_rgt);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_66_cse, COMP_LOOP_or_120_rgt);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_67_cse, COMP_LOOP_or_120_rgt);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_68_cse, COMP_LOOP_or_120_rgt);
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm <= MUX_s_1_2_2(COMP_LOOP_tmp_COMP_LOOP_tmp_and_103_cse,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_69_cse, COMP_LOOP_or_120_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_3_tmp_lshift_ncse_sva <= 9'b000000000;
      COMP_LOOP_tmp_nor_206_itm <= 1'b0;
      COMP_LOOP_tmp_nor_207_itm <= 1'b0;
      COMP_LOOP_tmp_nor_209_itm <= 1'b0;
      COMP_LOOP_tmp_nor_213_itm <= 1'b0;
      COMP_LOOP_tmp_nor_220_itm <= 1'b0;
    end
    else if ( COMP_LOOP_tmp_or_43_cse ) begin
      COMP_LOOP_3_tmp_lshift_ncse_sva <= MUX_v_9_2_2((z_out_1[8:0]), (z_out_7[8:0]),
          and_dcpl_261);
      COMP_LOOP_tmp_nor_206_itm <= COMP_LOOP_tmp_nor_34_cse;
      COMP_LOOP_tmp_nor_207_itm <= COMP_LOOP_tmp_nor_35_cse;
      COMP_LOOP_tmp_nor_209_itm <= COMP_LOOP_tmp_nor_37_cse;
      COMP_LOOP_tmp_nor_213_itm <= COMP_LOOP_tmp_nor_41_cse;
      COMP_LOOP_tmp_nor_220_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_474_tmp ) begin
      COMP_LOOP_tmp_mux1h_1_itm <= MUX1HOT_v_64_64_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
          twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_5_i_q_d,
          twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d, twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d,
          twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d,
          twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d,
          twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d,
          twiddle_rsc_0_19_i_q_d, twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d,
          twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d,
          twiddle_rsc_0_25_i_q_d, twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d,
          twiddle_rsc_0_28_i_q_d, twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d,
          twiddle_rsc_0_31_i_q_d, twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_33_i_q_d,
          twiddle_rsc_0_34_i_q_d, twiddle_rsc_0_35_i_q_d, twiddle_rsc_0_36_i_q_d,
          twiddle_rsc_0_37_i_q_d, twiddle_rsc_0_38_i_q_d, twiddle_rsc_0_39_i_q_d,
          twiddle_rsc_0_40_i_q_d, twiddle_rsc_0_41_i_q_d, twiddle_rsc_0_42_i_q_d,
          twiddle_rsc_0_43_i_q_d, twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_45_i_q_d,
          twiddle_rsc_0_46_i_q_d, twiddle_rsc_0_47_i_q_d, twiddle_rsc_0_48_i_q_d,
          twiddle_rsc_0_49_i_q_d, twiddle_rsc_0_50_i_q_d, twiddle_rsc_0_51_i_q_d,
          twiddle_rsc_0_52_i_q_d, twiddle_rsc_0_53_i_q_d, twiddle_rsc_0_54_i_q_d,
          twiddle_rsc_0_55_i_q_d, twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_57_i_q_d,
          twiddle_rsc_0_58_i_q_d, twiddle_rsc_0_59_i_q_d, twiddle_rsc_0_60_i_q_d,
          twiddle_rsc_0_61_i_q_d, twiddle_rsc_0_62_i_q_d, twiddle_rsc_0_63_i_q_d,
          {COMP_LOOP_tmp_and_249_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_nl
          , COMP_LOOP_tmp_and_250_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_nl , COMP_LOOP_tmp_and_251_nl
          , COMP_LOOP_tmp_and_252_nl , COMP_LOOP_tmp_and_253_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_nl
          , COMP_LOOP_tmp_and_254_nl , COMP_LOOP_tmp_and_255_nl , COMP_LOOP_tmp_and_256_nl
          , COMP_LOOP_tmp_and_257_nl , COMP_LOOP_tmp_and_258_nl , COMP_LOOP_tmp_and_259_nl
          , COMP_LOOP_tmp_and_260_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_22_nl , COMP_LOOP_tmp_and_261_nl
          , COMP_LOOP_tmp_and_262_nl , COMP_LOOP_tmp_and_263_nl , COMP_LOOP_tmp_and_264_nl
          , COMP_LOOP_tmp_and_265_nl , COMP_LOOP_tmp_and_266_nl , COMP_LOOP_tmp_and_267_nl
          , COMP_LOOP_tmp_and_268_nl , COMP_LOOP_tmp_and_269_nl , COMP_LOOP_tmp_and_270_nl
          , COMP_LOOP_tmp_and_271_nl , COMP_LOOP_tmp_and_272_nl , COMP_LOOP_tmp_and_273_nl
          , COMP_LOOP_tmp_and_274_nl , COMP_LOOP_tmp_and_275_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_nl
          , COMP_LOOP_tmp_and_276_nl , COMP_LOOP_tmp_and_277_nl , COMP_LOOP_tmp_and_278_nl
          , COMP_LOOP_tmp_and_279_nl , COMP_LOOP_tmp_and_280_nl , COMP_LOOP_tmp_and_281_nl
          , COMP_LOOP_tmp_and_282_nl , COMP_LOOP_tmp_and_283_nl , COMP_LOOP_tmp_and_284_nl
          , COMP_LOOP_tmp_and_285_nl , COMP_LOOP_tmp_and_286_nl , COMP_LOOP_tmp_and_287_nl
          , COMP_LOOP_tmp_and_288_nl , COMP_LOOP_tmp_and_289_nl , COMP_LOOP_tmp_and_290_nl
          , COMP_LOOP_tmp_and_291_nl , COMP_LOOP_tmp_and_292_nl , COMP_LOOP_tmp_and_293_nl
          , COMP_LOOP_tmp_and_294_nl , COMP_LOOP_tmp_and_295_nl , COMP_LOOP_tmp_and_296_nl
          , COMP_LOOP_tmp_and_297_nl , COMP_LOOP_tmp_and_298_nl , COMP_LOOP_tmp_and_299_nl
          , COMP_LOOP_tmp_and_300_nl , COMP_LOOP_tmp_and_301_nl , COMP_LOOP_tmp_and_302_nl
          , COMP_LOOP_tmp_and_303_nl , COMP_LOOP_tmp_and_304_nl , COMP_LOOP_tmp_and_305_nl
          , COMP_LOOP_tmp_and_306_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ nor_1579_tmp ) begin
      COMP_LOOP_tmp_mux1h_2_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_2_i_q_d,
          twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_10_i_q_d,
          twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_16_i_q_d,
          twiddle_rsc_0_18_i_q_d, twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_22_i_q_d,
          twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_28_i_q_d,
          twiddle_rsc_0_30_i_q_d, twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_34_i_q_d,
          twiddle_rsc_0_36_i_q_d, twiddle_rsc_0_38_i_q_d, twiddle_rsc_0_40_i_q_d,
          twiddle_rsc_0_42_i_q_d, twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_46_i_q_d,
          twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_50_i_q_d, twiddle_rsc_0_52_i_q_d,
          twiddle_rsc_0_54_i_q_d, twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_58_i_q_d,
          twiddle_rsc_0_60_i_q_d, twiddle_rsc_0_62_i_q_d, {COMP_LOOP_tmp_and_222_nl
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_70_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_71_nl
          , COMP_LOOP_tmp_and_223_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_73_nl , COMP_LOOP_tmp_and_224_nl
          , COMP_LOOP_tmp_and_225_nl , COMP_LOOP_tmp_and_226_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_77_nl
          , COMP_LOOP_tmp_and_227_nl , COMP_LOOP_tmp_and_228_nl , COMP_LOOP_tmp_and_229_nl
          , COMP_LOOP_tmp_and_230_nl , COMP_LOOP_tmp_and_231_nl , COMP_LOOP_tmp_and_232_nl
          , COMP_LOOP_tmp_and_233_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_nl , COMP_LOOP_tmp_and_234_nl
          , COMP_LOOP_tmp_and_235_nl , COMP_LOOP_tmp_and_236_nl , COMP_LOOP_tmp_and_237_nl
          , COMP_LOOP_tmp_and_238_nl , COMP_LOOP_tmp_and_239_nl , COMP_LOOP_tmp_and_240_nl
          , COMP_LOOP_tmp_and_241_nl , COMP_LOOP_tmp_and_242_nl , COMP_LOOP_tmp_and_243_nl
          , COMP_LOOP_tmp_and_244_nl , COMP_LOOP_tmp_and_245_nl , COMP_LOOP_tmp_and_246_nl
          , COMP_LOOP_tmp_and_247_nl , COMP_LOOP_tmp_and_248_nl});
    end
  end
  always @(posedge clk) begin
    if ( ~ and_476_tmp ) begin
      COMP_LOOP_tmp_mux1h_3_itm <= MUX1HOT_v_64_64_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_1_i_q_d,
          twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_3_i_q_d, twiddle_rsc_0_4_i_q_d, twiddle_rsc_0_5_i_q_d,
          twiddle_rsc_0_6_i_q_d, twiddle_rsc_0_7_i_q_d, twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_9_i_q_d,
          twiddle_rsc_0_10_i_q_d, twiddle_rsc_0_11_i_q_d, twiddle_rsc_0_12_i_q_d,
          twiddle_rsc_0_13_i_q_d, twiddle_rsc_0_14_i_q_d, twiddle_rsc_0_15_i_q_d,
          twiddle_rsc_0_16_i_q_d, twiddle_rsc_0_17_i_q_d, twiddle_rsc_0_18_i_q_d,
          twiddle_rsc_0_19_i_q_d, twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_21_i_q_d,
          twiddle_rsc_0_22_i_q_d, twiddle_rsc_0_23_i_q_d, twiddle_rsc_0_24_i_q_d,
          twiddle_rsc_0_25_i_q_d, twiddle_rsc_0_26_i_q_d, twiddle_rsc_0_27_i_q_d,
          twiddle_rsc_0_28_i_q_d, twiddle_rsc_0_29_i_q_d, twiddle_rsc_0_30_i_q_d,
          twiddle_rsc_0_31_i_q_d, twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_33_i_q_d,
          twiddle_rsc_0_34_i_q_d, twiddle_rsc_0_35_i_q_d, twiddle_rsc_0_36_i_q_d,
          twiddle_rsc_0_37_i_q_d, twiddle_rsc_0_38_i_q_d, twiddle_rsc_0_39_i_q_d,
          twiddle_rsc_0_40_i_q_d, twiddle_rsc_0_41_i_q_d, twiddle_rsc_0_42_i_q_d,
          twiddle_rsc_0_43_i_q_d, twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_45_i_q_d,
          twiddle_rsc_0_46_i_q_d, twiddle_rsc_0_47_i_q_d, twiddle_rsc_0_48_i_q_d,
          twiddle_rsc_0_49_i_q_d, twiddle_rsc_0_50_i_q_d, twiddle_rsc_0_51_i_q_d,
          twiddle_rsc_0_52_i_q_d, twiddle_rsc_0_53_i_q_d, twiddle_rsc_0_54_i_q_d,
          twiddle_rsc_0_55_i_q_d, twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_57_i_q_d,
          twiddle_rsc_0_58_i_q_d, twiddle_rsc_0_59_i_q_d, twiddle_rsc_0_60_i_q_d,
          twiddle_rsc_0_61_i_q_d, twiddle_rsc_0_62_i_q_d, twiddle_rsc_0_63_i_q_d,
          {COMP_LOOP_tmp_and_164_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_102_nl
          , COMP_LOOP_tmp_and_165_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_nl , COMP_LOOP_tmp_and_166_nl
          , COMP_LOOP_tmp_and_167_nl , COMP_LOOP_tmp_and_168_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_nl
          , COMP_LOOP_tmp_and_169_nl , COMP_LOOP_tmp_and_170_nl , COMP_LOOP_tmp_and_171_nl
          , COMP_LOOP_tmp_and_172_nl , COMP_LOOP_tmp_and_173_nl , COMP_LOOP_tmp_and_174_nl
          , COMP_LOOP_tmp_and_175_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_nl , COMP_LOOP_tmp_and_176_nl
          , COMP_LOOP_tmp_and_177_nl , COMP_LOOP_tmp_and_178_nl , COMP_LOOP_tmp_and_179_nl
          , COMP_LOOP_tmp_and_180_nl , COMP_LOOP_tmp_and_181_nl , COMP_LOOP_tmp_and_182_nl
          , COMP_LOOP_tmp_and_183_nl , COMP_LOOP_tmp_and_184_nl , COMP_LOOP_tmp_and_185_nl
          , COMP_LOOP_tmp_and_186_nl , COMP_LOOP_tmp_and_187_nl , COMP_LOOP_tmp_and_188_nl
          , COMP_LOOP_tmp_and_189_nl , COMP_LOOP_tmp_and_190_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_nl
          , COMP_LOOP_tmp_and_191_nl , COMP_LOOP_tmp_and_192_nl , COMP_LOOP_tmp_and_193_nl
          , COMP_LOOP_tmp_and_194_nl , COMP_LOOP_tmp_and_195_nl , COMP_LOOP_tmp_and_196_nl
          , COMP_LOOP_tmp_and_197_nl , COMP_LOOP_tmp_and_198_nl , COMP_LOOP_tmp_and_199_nl
          , COMP_LOOP_tmp_and_200_nl , COMP_LOOP_tmp_and_201_nl , COMP_LOOP_tmp_and_202_nl
          , COMP_LOOP_tmp_and_203_nl , COMP_LOOP_tmp_and_204_nl , COMP_LOOP_tmp_and_205_nl
          , COMP_LOOP_tmp_and_206_nl , COMP_LOOP_tmp_and_207_nl , COMP_LOOP_tmp_and_208_nl
          , COMP_LOOP_tmp_and_209_nl , COMP_LOOP_tmp_and_210_nl , COMP_LOOP_tmp_and_211_nl
          , COMP_LOOP_tmp_and_212_nl , COMP_LOOP_tmp_and_213_nl , COMP_LOOP_tmp_and_214_nl
          , COMP_LOOP_tmp_and_215_nl , COMP_LOOP_tmp_and_216_nl , COMP_LOOP_tmp_and_217_nl
          , COMP_LOOP_tmp_and_218_nl , COMP_LOOP_tmp_and_219_nl , COMP_LOOP_tmp_and_220_nl
          , COMP_LOOP_tmp_and_221_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= 1'b0;
    end
    else if ( COMP_LOOP_or_74_cse ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_1_cse;
    end
  end
  always @(posedge clk) begin
    if ( ~ nor_tmp_396 ) begin
      COMP_LOOP_tmp_mux1h_4_itm <= MUX1HOT_v_64_16_2(twiddle_rsc_0_0_i_q_d, twiddle_rsc_0_4_i_q_d,
          twiddle_rsc_0_8_i_q_d, twiddle_rsc_0_12_i_q_d, twiddle_rsc_0_16_i_q_d,
          twiddle_rsc_0_20_i_q_d, twiddle_rsc_0_24_i_q_d, twiddle_rsc_0_28_i_q_d,
          twiddle_rsc_0_32_i_q_d, twiddle_rsc_0_36_i_q_d, twiddle_rsc_0_40_i_q_d,
          twiddle_rsc_0_44_i_q_d, twiddle_rsc_0_48_i_q_d, twiddle_rsc_0_52_i_q_d,
          twiddle_rsc_0_56_i_q_d, twiddle_rsc_0_60_i_q_d, {COMP_LOOP_tmp_and_152_nl
          , COMP_LOOP_tmp_COMP_LOOP_tmp_and_164_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_165_nl
          , COMP_LOOP_tmp_and_153_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_167_nl , COMP_LOOP_tmp_and_154_nl
          , COMP_LOOP_tmp_and_155_nl , COMP_LOOP_tmp_and_156_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_171_nl
          , COMP_LOOP_tmp_and_157_nl , COMP_LOOP_tmp_and_158_nl , COMP_LOOP_tmp_and_159_nl
          , COMP_LOOP_tmp_and_160_nl , COMP_LOOP_tmp_and_161_nl , COMP_LOOP_tmp_and_162_nl
          , COMP_LOOP_tmp_and_163_nl});
    end
  end
  always @(posedge clk) begin
    if ( ((~((COMP_LOOP_2_tmp_lshift_ncse_sva[0]) & COMP_LOOP_tmp_nor_10_itm)) |
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm | COMP_LOOP_COMP_LOOP_and_102_itm
        | COMP_LOOP_COMP_LOOP_and_106_itm | COMP_LOOP_COMP_LOOP_and_107_itm | COMP_LOOP_COMP_LOOP_and_108_itm
        | COMP_LOOP_COMP_LOOP_and_109_itm | COMP_LOOP_COMP_LOOP_and_110_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt
        | COMP_LOOP_COMP_LOOP_and_1104_itm | COMP_LOOP_COMP_LOOP_and_1106_itm | COMP_LOOP_COMP_LOOP_and_1118_itm
        | COMP_LOOP_COMP_LOOP_and_115_itm | COMP_LOOP_COMP_LOOP_and_116_itm | COMP_LOOP_COMP_LOOP_and_117_itm
        | COMP_LOOP_COMP_LOOP_and_118_itm | COMP_LOOP_COMP_LOOP_and_120_itm | COMP_LOOP_COMP_LOOP_and_121_itm
        | COMP_LOOP_COMP_LOOP_and_122_itm | COMP_LOOP_COMP_LOOP_and_123_itm | COMP_LOOP_COMP_LOOP_and_124_itm
        | COMP_LOOP_COMP_LOOP_and_125_itm | COMP_LOOP_COMP_LOOP_and_1370_itm | COMP_LOOP_COMP_LOOP_and_1831_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt | COMP_LOOP_COMP_LOOP_and_1874_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm
        | and_dcpl_432 | and_dcpl_263) & mux_3353_nl ) begin
      tmp_21_sva_1 <= MUX1HOT_v_64_65_2(twiddle_rsc_0_1_i_q_d, twiddle_rsc_0_22_i_q_d,
          twiddle_rsc_0_0_i_q_d, tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d,
          tmp_21_sva_5, tmp_21_sva_6, tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9,
          COMP_LOOP_1_acc_8_itm, tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13,
          tmp_21_sva_14, tmp_21_sva_15, twiddle_rsc_0_16_i_q_d, tmp_21_sva_17, tmp_21_sva_18,
          tmp_21_sva_19, twiddle_rsc_0_20_i_q_d, tmp_21_sva_21, tmp_21_sva_22, tmp_21_sva_23,
          twiddle_rsc_0_24_i_q_d, tmp_21_sva_25, tmp_21_sva_26, tmp_21_sva_27, twiddle_rsc_0_28_i_q_d,
          tmp_21_sva_29, tmp_21_sva_30, tmp_21_sva_31, twiddle_rsc_0_32_i_q_d, tmp_21_sva_33,
          tmp_21_sva_34, tmp_21_sva_35, twiddle_rsc_0_36_i_q_d, tmp_21_sva_37, tmp_21_sva_38,
          tmp_21_sva_39, twiddle_rsc_0_40_i_q_d, tmp_21_sva_41, tmp_21_sva_42, tmp_21_sva_43,
          twiddle_rsc_0_44_i_q_d, tmp_21_sva_45, tmp_21_sva_46, tmp_21_sva_47, twiddle_rsc_0_48_i_q_d,
          tmp_21_sva_49, tmp_21_sva_50, tmp_21_sva_51, twiddle_rsc_0_52_i_q_d, tmp_21_sva_53,
          tmp_21_sva_54, tmp_21_sva_55, twiddle_rsc_0_56_i_q_d, tmp_21_sva_57, tmp_21_sva_58,
          tmp_21_sva_59, twiddle_rsc_0_60_i_q_d, tmp_21_sva_61, tmp_21_sva_62, tmp_21_sva_63,
          {and_dcpl_432 , and_dcpl_263 , COMP_LOOP_tmp_and_89_nl , COMP_LOOP_tmp_and_90_nl
          , COMP_LOOP_tmp_and_91_nl , COMP_LOOP_tmp_and_92_nl , COMP_LOOP_tmp_and_93_nl
          , COMP_LOOP_tmp_and_94_nl , COMP_LOOP_tmp_and_95_nl , COMP_LOOP_tmp_and_96_nl
          , COMP_LOOP_tmp_and_97_nl , COMP_LOOP_tmp_and_98_nl , COMP_LOOP_tmp_and_99_nl
          , COMP_LOOP_tmp_and_100_nl , COMP_LOOP_tmp_and_101_nl , COMP_LOOP_tmp_and_102_nl
          , COMP_LOOP_tmp_and_103_nl , COMP_LOOP_tmp_and_104_nl , COMP_LOOP_tmp_and_105_nl
          , COMP_LOOP_tmp_and_106_nl , COMP_LOOP_tmp_and_107_nl , COMP_LOOP_tmp_and_108_nl
          , COMP_LOOP_tmp_and_109_nl , COMP_LOOP_tmp_and_110_nl , COMP_LOOP_tmp_and_111_nl
          , COMP_LOOP_tmp_and_112_nl , COMP_LOOP_tmp_and_113_nl , COMP_LOOP_tmp_and_114_nl
          , COMP_LOOP_tmp_and_115_nl , COMP_LOOP_tmp_and_116_nl , COMP_LOOP_tmp_and_117_nl
          , COMP_LOOP_tmp_and_118_nl , COMP_LOOP_tmp_and_119_nl , COMP_LOOP_tmp_and_120_nl
          , COMP_LOOP_tmp_and_121_nl , COMP_LOOP_tmp_and_122_nl , COMP_LOOP_tmp_and_123_nl
          , COMP_LOOP_tmp_and_124_nl , COMP_LOOP_tmp_and_125_nl , COMP_LOOP_tmp_and_126_nl
          , COMP_LOOP_tmp_and_127_nl , COMP_LOOP_tmp_and_128_nl , COMP_LOOP_tmp_and_129_nl
          , COMP_LOOP_tmp_and_130_nl , COMP_LOOP_tmp_and_131_nl , COMP_LOOP_tmp_and_132_nl
          , COMP_LOOP_tmp_and_133_nl , COMP_LOOP_tmp_and_134_nl , COMP_LOOP_tmp_and_135_nl
          , COMP_LOOP_tmp_and_136_nl , COMP_LOOP_tmp_and_137_nl , COMP_LOOP_tmp_and_138_nl
          , COMP_LOOP_tmp_and_139_nl , COMP_LOOP_tmp_and_140_nl , COMP_LOOP_tmp_and_141_nl
          , COMP_LOOP_tmp_and_142_nl , COMP_LOOP_tmp_and_143_nl , COMP_LOOP_tmp_and_144_nl
          , COMP_LOOP_tmp_and_145_nl , COMP_LOOP_tmp_and_146_nl , COMP_LOOP_tmp_and_147_nl
          , COMP_LOOP_tmp_and_148_nl , COMP_LOOP_tmp_and_149_nl , COMP_LOOP_tmp_and_150_nl
          , COMP_LOOP_tmp_and_151_nl});
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm ) begin
      tmp_21_sva_3 <= twiddle_rsc_0_3_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm ) begin
      tmp_21_sva_5 <= twiddle_rsc_0_5_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm ) begin
      tmp_21_sva_7 <= twiddle_rsc_0_7_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm ) begin
      tmp_21_sva_9 <= twiddle_rsc_0_9_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_COMP_LOOP_and_123_itm ) begin
      tmp_21_sva_27 <= twiddle_rsc_0_27_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_COMP_LOOP_and_125_itm ) begin
      tmp_21_sva_29 <= twiddle_rsc_0_29_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_COMP_LOOP_and_1831_itm ) begin
      tmp_21_sva_31 <= twiddle_rsc_0_31_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_COMP_LOOP_and_1874_itm ) begin
      tmp_21_sva_33 <= twiddle_rsc_0_33_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm ) begin
      tmp_21_sva_35 <= twiddle_rsc_0_35_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm ) begin
      tmp_21_sva_37 <= twiddle_rsc_0_37_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm ) begin
      tmp_21_sva_39 <= twiddle_rsc_0_39_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm ) begin
      tmp_21_sva_41 <= twiddle_rsc_0_41_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm ) begin
      tmp_21_sva_43 <= twiddle_rsc_0_43_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm ) begin
      tmp_21_sva_45 <= twiddle_rsc_0_45_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm ) begin
      tmp_21_sva_47 <= twiddle_rsc_0_47_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm ) begin
      tmp_21_sva_49 <= twiddle_rsc_0_49_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm ) begin
      tmp_21_sva_51 <= twiddle_rsc_0_51_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm ) begin
      tmp_21_sva_53 <= twiddle_rsc_0_53_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm ) begin
      tmp_21_sva_55 <= twiddle_rsc_0_55_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm ) begin
      tmp_21_sva_57 <= twiddle_rsc_0_57_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm ) begin
      tmp_21_sva_59 <= twiddle_rsc_0_59_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm ) begin
      tmp_21_sva_61 <= twiddle_rsc_0_61_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm ) begin
      tmp_21_sva_63 <= twiddle_rsc_0_63_i_q_d;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_nor_2_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_74_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_75_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_76_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_78_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_79_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_80_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_81_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_82_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_83_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_84_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_86_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_87_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_88_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_89_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_90_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_91_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_92_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_93_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_94_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_95_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_96_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_97_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_98_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_99_cse;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm <= 1'b0;
    end
    else if ( ~ or_dcpl_150 ) begin
      COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm <= COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_cse;
    end
  end
  always @(posedge clk) begin
    if ( mux_3360_tmp ) begin
      COMP_LOOP_tmp_mux1h_5_itm <= MUX1HOT_v_64_64_2(twiddle_rsc_0_0_i_q_d, tmp_21_sva_1,
          tmp_21_sva_2, tmp_21_sva_3, twiddle_rsc_0_4_i_q_d, tmp_21_sva_5, tmp_21_sva_6,
          tmp_21_sva_7, twiddle_rsc_0_8_i_q_d, tmp_21_sva_9, COMP_LOOP_1_acc_8_itm,
          tmp_21_sva_11, twiddle_rsc_0_12_i_q_d, tmp_21_sva_13, tmp_21_sva_14, tmp_21_sva_15,
          twiddle_rsc_0_16_i_q_d, tmp_21_sva_17, tmp_21_sva_18, tmp_21_sva_19, twiddle_rsc_0_20_i_q_d,
          tmp_21_sva_21, tmp_21_sva_22, tmp_21_sva_23, twiddle_rsc_0_24_i_q_d, tmp_21_sva_25,
          tmp_21_sva_26, tmp_21_sva_27, twiddle_rsc_0_28_i_q_d, tmp_21_sva_29, tmp_21_sva_30,
          tmp_21_sva_31, twiddle_rsc_0_32_i_q_d, tmp_21_sva_33, tmp_21_sva_34, tmp_21_sva_35,
          twiddle_rsc_0_36_i_q_d, tmp_21_sva_37, tmp_21_sva_38, tmp_21_sva_39, twiddle_rsc_0_40_i_q_d,
          tmp_21_sva_41, tmp_21_sva_42, tmp_21_sva_43, twiddle_rsc_0_44_i_q_d, tmp_21_sva_45,
          tmp_21_sva_46, tmp_21_sva_47, twiddle_rsc_0_48_i_q_d, tmp_21_sva_49, tmp_21_sva_50,
          tmp_21_sva_51, twiddle_rsc_0_52_i_q_d, tmp_21_sva_53, tmp_21_sva_54, tmp_21_sva_55,
          twiddle_rsc_0_56_i_q_d, tmp_21_sva_57, tmp_21_sva_58, tmp_21_sva_59, twiddle_rsc_0_60_i_q_d,
          tmp_21_sva_61, tmp_21_sva_62, tmp_21_sva_63, {COMP_LOOP_tmp_and_31_nl ,
          COMP_LOOP_tmp_COMP_LOOP_tmp_and_179_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_180_nl
          , COMP_LOOP_tmp_and_32_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_182_nl , COMP_LOOP_tmp_and_33_nl
          , COMP_LOOP_tmp_and_34_nl , COMP_LOOP_tmp_and_35_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_186_nl
          , COMP_LOOP_tmp_and_36_nl , COMP_LOOP_tmp_and_37_nl , COMP_LOOP_tmp_and_38_nl
          , COMP_LOOP_tmp_and_39_nl , COMP_LOOP_tmp_and_40_nl , COMP_LOOP_tmp_and_41_nl
          , COMP_LOOP_tmp_and_42_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_194_nl , COMP_LOOP_tmp_and_43_nl
          , COMP_LOOP_tmp_and_44_nl , COMP_LOOP_tmp_and_45_nl , COMP_LOOP_tmp_and_46_nl
          , COMP_LOOP_tmp_and_47_nl , COMP_LOOP_tmp_and_48_nl , COMP_LOOP_tmp_and_49_nl
          , COMP_LOOP_tmp_and_50_nl , COMP_LOOP_tmp_and_51_nl , COMP_LOOP_tmp_and_52_nl
          , COMP_LOOP_tmp_and_53_nl , COMP_LOOP_tmp_and_54_nl , COMP_LOOP_tmp_and_55_nl
          , COMP_LOOP_tmp_and_56_nl , COMP_LOOP_tmp_and_57_nl , COMP_LOOP_tmp_COMP_LOOP_tmp_and_210_nl
          , COMP_LOOP_tmp_and_58_nl , COMP_LOOP_tmp_and_59_nl , COMP_LOOP_tmp_and_60_nl
          , COMP_LOOP_tmp_and_61_nl , COMP_LOOP_tmp_and_62_nl , COMP_LOOP_tmp_and_63_nl
          , COMP_LOOP_tmp_and_64_nl , COMP_LOOP_tmp_and_65_nl , COMP_LOOP_tmp_and_66_nl
          , COMP_LOOP_tmp_and_67_nl , COMP_LOOP_tmp_and_68_nl , COMP_LOOP_tmp_and_69_nl
          , COMP_LOOP_tmp_and_70_nl , COMP_LOOP_tmp_and_71_nl , COMP_LOOP_tmp_and_72_nl
          , COMP_LOOP_tmp_and_73_nl , COMP_LOOP_tmp_and_74_nl , COMP_LOOP_tmp_and_75_nl
          , COMP_LOOP_tmp_and_76_nl , COMP_LOOP_tmp_and_77_nl , COMP_LOOP_tmp_and_78_nl
          , COMP_LOOP_tmp_and_79_nl , COMP_LOOP_tmp_and_80_nl , COMP_LOOP_tmp_and_81_nl
          , COMP_LOOP_tmp_and_82_nl , COMP_LOOP_tmp_and_83_nl , COMP_LOOP_tmp_and_84_nl
          , COMP_LOOP_tmp_and_85_nl , COMP_LOOP_tmp_and_86_nl , COMP_LOOP_tmp_and_87_nl
          , COMP_LOOP_tmp_and_88_nl});
    end
  end
  always @(posedge clk) begin
    if ( ((~(COMP_LOOP_tmp_nor_206_itm & (COMP_LOOP_3_tmp_lshift_ncse_sva[0]))) |
        COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt
        | COMP_LOOP_COMP_LOOP_and_119_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm | COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm
        | COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm | and_dcpl_263) & mux_3364_nl )
        begin
      COMP_LOOP_tmp_mux1h_6_itm <= MUX1HOT_v_64_32_2(twiddle_rsc_0_2_i_q_d, twiddle_rsc_0_0_i_q_d,
          twiddle_rsc_0_4_i_q_d, tmp_21_sva_21, twiddle_rsc_0_8_i_q_d, tmp_21_sva_23,
          twiddle_rsc_0_12_i_q_d, tmp_21_sva_25, twiddle_rsc_0_16_i_q_d, tmp_21_sva_26,
          twiddle_rsc_0_20_i_q_d, tmp_21_sva_1, twiddle_rsc_0_24_i_q_d, COMP_LOOP_1_acc_8_itm,
          twiddle_rsc_0_28_i_q_d, tmp_21_sva_11, twiddle_rsc_0_32_i_q_d, tmp_21_sva_13,
          twiddle_rsc_0_36_i_q_d, tmp_21_sva_14, twiddle_rsc_0_40_i_q_d, tmp_21_sva_15,
          twiddle_rsc_0_44_i_q_d, tmp_21_sva_17, twiddle_rsc_0_48_i_q_d, tmp_21_sva_18,
          twiddle_rsc_0_52_i_q_d, tmp_21_sva_19, twiddle_rsc_0_56_i_q_d, tmp_21_sva_2,
          twiddle_rsc_0_60_i_q_d, tmp_21_sva_22, {and_dcpl_263 , COMP_LOOP_tmp_and_nl
          , COMP_LOOP_tmp_and_1_nl , COMP_LOOP_tmp_and_2_nl , COMP_LOOP_tmp_and_3_nl
          , COMP_LOOP_tmp_and_4_nl , COMP_LOOP_tmp_and_5_nl , COMP_LOOP_tmp_and_6_nl
          , COMP_LOOP_tmp_and_7_nl , COMP_LOOP_tmp_and_8_nl , COMP_LOOP_tmp_and_9_nl
          , COMP_LOOP_tmp_and_10_nl , COMP_LOOP_tmp_and_11_nl , COMP_LOOP_tmp_and_12_nl
          , COMP_LOOP_tmp_and_13_nl , COMP_LOOP_tmp_and_14_nl , COMP_LOOP_tmp_and_15_nl
          , COMP_LOOP_tmp_and_16_nl , COMP_LOOP_tmp_and_17_nl , COMP_LOOP_tmp_and_18_nl
          , COMP_LOOP_tmp_and_19_nl , COMP_LOOP_tmp_and_20_nl , COMP_LOOP_tmp_and_21_nl
          , COMP_LOOP_tmp_and_22_nl , COMP_LOOP_tmp_and_23_nl , COMP_LOOP_tmp_and_24_nl
          , COMP_LOOP_tmp_and_25_nl , COMP_LOOP_tmp_and_26_nl , COMP_LOOP_tmp_and_27_nl
          , COMP_LOOP_tmp_and_28_nl , COMP_LOOP_tmp_and_29_nl , COMP_LOOP_tmp_and_30_nl});
    end
  end
  assign nor_1423_nl = ~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[4])
      | (fsm_output[0]) | (fsm_output[3]) | (fsm_output[7]));
  assign mux_788_nl = MUX_s_1_2_2(and_tmp_29, and_78_cse, fsm_output[2]);
  assign mux_789_nl = MUX_s_1_2_2(mux_788_nl, mux_tmp_720, fsm_output[1]);
  assign VEC_LOOP_j_not_1_nl = ~ VEC_LOOP_j_10_0_sva_9_0_mx0c0;
  assign nor_422_nl = ~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[4])
      | (fsm_output[3]) | (fsm_output[7]));
  assign nor_1426_nl = ~((fsm_output[1]) | (fsm_output[6]) | (fsm_output[7]));
  assign and_637_nl = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[7]);
  assign mux_781_nl = MUX_s_1_2_2(nor_1426_nl, and_637_nl, fsm_output[5]);
  assign nand_480_nl = ~(mux_781_nl & and_dcpl_365 & (~ (fsm_output[4])) & (~ (fsm_output[2])));
  assign or_4159_nl = (fsm_output[6:4]!=3'b000) | nor_1744_cse | (fsm_output[3]);
  assign nor_1745_nl = ~(((fsm_output[2:0]==3'b111)) | (fsm_output[3]));
  assign or_4154_nl = (fsm_output[2]) | and_1046_cse | (fsm_output[3]);
  assign mux_nl = MUX_s_1_2_2(nor_1745_nl, or_4154_nl, fsm_output[5]);
  assign mux_3365_nl = MUX_s_1_2_2(mux_nl, (fsm_output[5]), fsm_output[4]);
  assign nand_493_nl = ~((fsm_output[6]) & (~ mux_3365_nl));
  assign COMP_LOOP_COMP_LOOP_and_73_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001011);
  assign COMP_LOOP_COMP_LOOP_and_824_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[2:1]==2'b11)
      & COMP_LOOP_nor_734_itm;
  assign COMP_LOOP_COMP_LOOP_and_74_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001100);
  assign COMP_LOOP_COMP_LOOP_and_851_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_4_sva[0]) & COMP_LOOP_nor_760_itm;
  assign COMP_LOOP_COMP_LOOP_and_75_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001101);
  assign COMP_LOOP_COMP_LOOP_and_858_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_4_sva[3]) & COMP_LOOP_nor_767_itm;
  assign COMP_LOOP_COMP_LOOP_and_100_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100110);
  assign COMP_LOOP_COMP_LOOP_and_323_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[3]) &
      (COMP_LOOP_acc_10_cse_10_1_2_sva[0]) & COMP_LOOP_nor_289_itm;
  assign COMP_LOOP_COMP_LOOP_and_1073_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[1:0]==2'b11)
      & COMP_LOOP_nor_955_itm;
  assign mux_3036_nl = MUX_s_1_2_2(mux_tmp_2968, mux_tmp_2966, fsm_output[1]);
  assign mux_3037_nl = MUX_s_1_2_2(or_4057_cse, (~ mux_3036_nl), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_101_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100111);
  assign COMP_LOOP_COMP_LOOP_and_348_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_2_sva[1]) & COMP_LOOP_nor_313_itm;
  assign COMP_LOOP_COMP_LOOP_and_1075_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[2]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) & COMP_LOOP_nor_957_itm;
  assign and_403_nl = and_dcpl_76 & and_dcpl_88;
  assign nor_420_nl = ~(and_507_cse | (fsm_output[6]) | (fsm_output[4]) | (fsm_output[3]));
  assign mux_3039_nl = MUX_s_1_2_2(nor_420_nl, mux_tmp_2971, fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_102_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101000);
  assign COMP_LOOP_COMP_LOOP_and_1076_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[2:1]==2'b11)
      & COMP_LOOP_nor_958_itm;
  assign COMP_LOOP_COMP_LOOP_and_109_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101111);
  assign COMP_LOOP_COMP_LOOP_and_1094_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4:3]==2'b11)
      & COMP_LOOP_nor_976_itm;
  assign COMP_LOOP_COMP_LOOP_and_103_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101001);
  assign COMP_LOOP_COMP_LOOP_and_350_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_2_sva[2]) & COMP_LOOP_nor_315_itm;
  assign COMP_LOOP_COMP_LOOP_and_1079_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) & COMP_LOOP_nor_961_itm;
  assign mux_3046_nl = MUX_s_1_2_2(or_4057_cse, (~ mux_tmp_2968), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_104_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101010);
  assign COMP_LOOP_COMP_LOOP_and_354_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_2_sva[3]) & COMP_LOOP_nor_319_itm;
  assign COMP_LOOP_COMP_LOOP_and_1080_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & COMP_LOOP_nor_962_itm;
  assign and_409_nl = and_dcpl_76 & and_dcpl_377;
  assign mux_3047_nl = MUX_s_1_2_2(or_tmp_3747, (~ mux_tmp_2966), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_105_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101011);
  assign COMP_LOOP_COMP_LOOP_and_362_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[5:4]==2'b11)
      & COMP_LOOP_nor_326_itm;
  assign COMP_LOOP_COMP_LOOP_and_1082_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3:2]==2'b11)
      & COMP_LOOP_nor_964_itm;
  assign mux_3048_nl = MUX_s_1_2_2(or_tmp_3747, (~ mux_tmp_2968), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_106_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101100);
  assign COMP_LOOP_COMP_LOOP_and_1087_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) & COMP_LOOP_nor_969_itm;
  assign and_411_nl = and_dcpl_94 & and_dcpl_113;
  assign or_3878_nl = and_507_cse | (fsm_output[6]);
  assign or_3877_nl = nor_1744_cse | (fsm_output[6]);
  assign mux_3051_nl = MUX_s_1_2_2(or_3878_nl, or_3877_nl, fsm_output[3]);
  assign mux_3052_nl = MUX_s_1_2_2((fsm_output[6]), mux_3051_nl, nor_358_cse);
  assign nor_418_nl = ~((fsm_output[1]) | (fsm_output[6]));
  assign or_3874_nl = (fsm_output[3:2]!=2'b00);
  assign mux_3049_nl = MUX_s_1_2_2(nor_418_nl, (fsm_output[6]), or_3874_nl);
  assign mux_3050_nl = MUX_s_1_2_2((fsm_output[6]), (~ mux_3049_nl), fsm_output[5]);
  assign mux_3053_nl = MUX_s_1_2_2(mux_3052_nl, mux_3050_nl, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_and_107_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101101);
  assign COMP_LOOP_COMP_LOOP_and_1088_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & COMP_LOOP_nor_970_itm;
  assign mux_3055_nl = MUX_s_1_2_2((~ and_640_cse), and_640_cse, fsm_output[6]);
  assign mux_3054_nl = MUX_s_1_2_2((~ and_640_cse), (fsm_output[4]), fsm_output[6]);
  assign mux_3056_nl = MUX_s_1_2_2(mux_3055_nl, mux_3054_nl, fsm_output[2]);
  assign mux_3059_nl = MUX_s_1_2_2((~ mux_3058_itm), mux_3056_nl, fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_108_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b101110);
  assign COMP_LOOP_COMP_LOOP_and_1090_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[2]) & COMP_LOOP_nor_972_itm;
  assign mux_3062_nl = MUX_s_1_2_2(mux_tmp_2994, mux_tmp_2993, fsm_output[1]);
  assign mux_3063_nl = MUX_s_1_2_2(mux_3062_nl, (~ mux_180_cse), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_110_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110000);
  assign COMP_LOOP_COMP_LOOP_and_1103_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) & COMP_LOOP_nor_984_itm;
  assign mux_3064_nl = MUX_s_1_2_2((~ mux_3058_itm), mux_tmp_2968, fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_115_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110101);
  assign COMP_LOOP_COMP_LOOP_and_1328_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2:1]==2'b11)
      & COMP_LOOP_nor_1182_itm;
  assign COMP_LOOP_COMP_LOOP_and_117_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110111);
  assign COMP_LOOP_COMP_LOOP_and_1332_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[1]) & COMP_LOOP_nor_1186_itm;
  assign COMP_LOOP_COMP_LOOP_and_122_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111100);
  assign COMP_LOOP_COMP_LOOP_and_1355_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) & COMP_LOOP_nor_1208_itm;
  assign COMP_LOOP_COMP_LOOP_and_116_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110110);
  assign COMP_LOOP_COMP_LOOP_and_1331_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) & COMP_LOOP_nor_1185_itm;
  assign or_3889_nl = (fsm_output[7:6]!=2'b01);
  assign mux_3073_nl = MUX_s_1_2_2(or_3889_nl, mux_742_cse, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_118_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111000);
  assign COMP_LOOP_COMP_LOOP_and_1334_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3:2]==2'b11)
      & COMP_LOOP_nor_1188_itm;
  assign mux_3081_nl = MUX_s_1_2_2(mux_tmp_3013, mux_tmp_3012, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_119_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111001);
  assign COMP_LOOP_COMP_LOOP_and_1339_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) & COMP_LOOP_nor_1193_itm;
  assign nor_414_nl = ~((~((fsm_output[0]) | (~ (fsm_output[3])))) | (fsm_output[7]));
  assign mux_3084_nl = MUX_s_1_2_2(nor_414_nl, (fsm_output[7]), or_341_cse);
  assign mux_3085_nl = MUX_s_1_2_2(mux_3084_nl, mux_tmp_3016, or_359_cse);
  assign COMP_LOOP_COMP_LOOP_and_120_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111010);
  assign COMP_LOOP_COMP_LOOP_and_1340_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[1]) & COMP_LOOP_nor_1194_itm;
  assign mux_3090_nl = MUX_s_1_2_2((~ or_tmp_3760), (fsm_output[7]), or_341_cse);
  assign mux_3091_nl = MUX_s_1_2_2(mux_3090_nl, mux_tmp_206, fsm_output[2]);
  assign mux_3087_nl = MUX_s_1_2_2((~ or_tmp_3757), (fsm_output[7]), or_341_cse);
  assign mux_3089_nl = MUX_s_1_2_2(mux_tmp_206, mux_3087_nl, fsm_output[2]);
  assign mux_3092_nl = MUX_s_1_2_2(mux_3091_nl, mux_3089_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_121_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111011);
  assign COMP_LOOP_COMP_LOOP_and_1342_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[2]) & COMP_LOOP_nor_1196_itm;
  assign and_503_nl = (fsm_output[3]) & (~ or_tmp_3773);
  assign mux_3096_nl = MUX_s_1_2_2(mux_3095_cse, and_503_nl, fsm_output[5]);
  assign mux_3097_nl = MUX_s_1_2_2(mux_3096_nl, nor_412_cse, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_and_123_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111101);
  assign COMP_LOOP_COMP_LOOP_and_1356_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[1]) & COMP_LOOP_nor_1209_itm;
  assign COMP_LOOP_COMP_LOOP_and_124_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111110);
  assign COMP_LOOP_COMP_LOOP_and_1358_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[2]) & COMP_LOOP_nor_1211_itm;
  assign or_3904_nl = (fsm_output[5]) | (~ mux_3095_cse);
  assign nand_145_nl = ~((fsm_output[5]) & (fsm_output[3]) & (~ or_tmp_3773));
  assign mux_3102_nl = MUX_s_1_2_2(or_3904_nl, nand_145_nl, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_and_125_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b111111);
  assign COMP_LOOP_COMP_LOOP_and_1362_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_6_sva[3]) & COMP_LOOP_nor_1215_itm;
  assign mux_3104_nl = MUX_s_1_2_2((~ or_tmp_3760), or_tmp_118, fsm_output[4]);
  assign mux_3105_nl = MUX_s_1_2_2(mux_3104_nl, (fsm_output[7]), fsm_output[6]);
  assign mux_3106_nl = MUX_s_1_2_2(mux_3105_nl, mux_tmp_444, fsm_output[2]);
  assign mux_3107_nl = MUX_s_1_2_2(mux_3106_nl, mux_tmp_3012, fsm_output[1]);
  assign mux_3110_nl = MUX_s_1_2_2(mux_tmp_2955, and_78_cse, fsm_output[2]);
  assign mux_3111_nl = MUX_s_1_2_2(mux_3110_nl, mux_tmp_3042, fsm_output[1]);
  assign mux_3113_nl = MUX_s_1_2_2(and_tmp_31, and_673_cse, or_359_cse);
  assign mux_3115_nl = MUX_s_1_2_2((~ mux_3114_itm), mux_3113_nl, fsm_output[5]);
  assign mux_3123_nl = MUX_s_1_2_2(mux_221_cse, (~ and_640_cse), fsm_output[5]);
  assign nl_COMP_LOOP_3_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b010}) + 11'b00000000001;
  assign COMP_LOOP_3_acc_nl = nl_COMP_LOOP_3_acc_nl[10:0];
  assign nand_149_nl = ~(or_359_cse & (fsm_output[4:3]==2'b11));
  assign mux_3124_nl = MUX_s_1_2_2(mux_221_cse, nand_149_nl, fsm_output[5]);
  assign mux_3125_nl = MUX_s_1_2_2(mux_tmp_2971, mux_tmp_3049, fsm_output[1]);
  assign mux_3126_nl = MUX_s_1_2_2(mux_3125_nl, (fsm_output[6]), fsm_output[5]);
  assign nl_COMP_LOOP_acc_12_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:3]))})
      + conv_u2u_8_9({COMP_LOOP_k_10_3_sva_6_0 , 1'b0}) + 9'b000000001;
  assign COMP_LOOP_acc_12_nl = nl_COMP_LOOP_acc_12_nl[8:0];
  assign mux_3127_nl = MUX_s_1_2_2(mux_tmp_2960, mux_tmp_3049, fsm_output[1]);
  assign mux_3128_nl = MUX_s_1_2_2(mux_3127_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_3130_nl = MUX_s_1_2_2((~ mux_3114_itm), and_673_cse, fsm_output[5]);
  assign nl_COMP_LOOP_5_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b100}) + 11'b00000000001;
  assign COMP_LOOP_5_acc_nl = nl_COMP_LOOP_5_acc_nl[10:0];
  assign mux_3131_nl = MUX_s_1_2_2(and_677_cse, and_673_cse, or_359_cse);
  assign mux_3132_nl = MUX_s_1_2_2((~ mux_3114_itm), mux_3131_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_13_psp_sva  = (VEC_LOOP_j_10_0_sva_9_0[9:2]) + ({COMP_LOOP_k_10_3_sva_6_0
      , 1'b1});
  assign and_497_nl = (fsm_output[0]) & (fsm_output[3]) & (fsm_output[7]);
  assign mux_3138_nl = MUX_s_1_2_2(and_497_nl, (fsm_output[7]), or_341_cse);
  assign mux_3139_nl = MUX_s_1_2_2(mux_tmp_3016, mux_3138_nl, fsm_output[2]);
  assign mux_3140_nl = MUX_s_1_2_2(mux_3139_nl, mux_tmp_3070, fsm_output[1]);
  assign mux_3142_nl = MUX_s_1_2_2(mux_tmp_3016, and_736_cse, fsm_output[2]);
  assign mux_3143_nl = MUX_s_1_2_2(mux_3142_nl, mux_tmp_3070, fsm_output[1]);
  assign nl_COMP_LOOP_6_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b101}) + 11'b00000000001;
  assign COMP_LOOP_6_acc_nl = nl_COMP_LOOP_6_acc_nl[10:0];
  assign mux_3146_nl = MUX_s_1_2_2(mux_tmp_3078, mux_tmp_3070, fsm_output[1]);
  assign mux_212_nl = MUX_s_1_2_2(and_tmp_10, (fsm_output[4]), or_359_cse);
  assign mux_3152_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_212_nl), fsm_output[5]);
  assign mux_219_nl = MUX_s_1_2_2(or_595_cse, or_4007_cse, and_507_cse);
  assign mux_3160_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_219_nl), fsm_output[5]);
  assign nl_COMP_LOOP_acc_1_cse_6_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b101});
  assign nor_410_nl = ~(and_1046_cse | (fsm_output[5]) | (fsm_output[7]));
  assign and_491_nl = ((fsm_output[1:0]!=2'b00)) & (fsm_output[5]) & (fsm_output[7]);
  assign mux_3161_nl = MUX_s_1_2_2(nor_410_nl, and_491_nl, fsm_output[3]);
  assign and_492_nl = (fsm_output[3]) & (fsm_output[5]) & (fsm_output[7]);
  assign mux_3162_nl = MUX_s_1_2_2(mux_3161_nl, and_492_nl, fsm_output[2]);
  assign mux_3163_nl = MUX_s_1_2_2(mux_3162_nl, and_493_cse, fsm_output[4]);
  assign nl_COMP_LOOP_7_acc_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + conv_u2s_10_11({COMP_LOOP_k_10_3_sva_6_0 , 3'b110}) + 11'b00000000001;
  assign COMP_LOOP_7_acc_nl = nl_COMP_LOOP_7_acc_nl[10:0];
  assign mux_3171_nl = MUX_s_1_2_2(nor_tmp_99, and_736_cse, or_359_cse);
  assign mux_3181_nl = MUX_s_1_2_2(mux_tmp_2955, and_705_cse, fsm_output[2]);
  assign mux_3182_nl = MUX_s_1_2_2(mux_3181_nl, mux_tmp_3042, fsm_output[1]);
  assign nl_COMP_LOOP_acc_15_nl = ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:4]))})
      + conv_u2u_7_8(COMP_LOOP_k_10_3_sva_6_0) + 8'b00000001;
  assign COMP_LOOP_acc_15_nl = nl_COMP_LOOP_acc_15_nl[7:0];
  assign nand_148_nl = ~((fsm_output[4:0]==5'b11111));
  assign mux_3188_nl = MUX_s_1_2_2(mux_221_cse, nand_148_nl, fsm_output[5]);
  assign mux_359_nl = MUX_s_1_2_2(and_tmp_10, (fsm_output[4]), fsm_output[2]);
  assign mux_361_nl = MUX_s_1_2_2(mux_tmp_293, mux_359_nl, fsm_output[1]);
  assign mux_3192_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_361_nl), fsm_output[5]);
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_10_0_sva_9_0 + ({COMP_LOOP_k_10_3_sva_6_0
      , 3'b111});
  assign mux_3193_nl = MUX_s_1_2_2(and_78_cse, and_705_cse, or_359_cse);
  assign nl_COMP_LOOP_1_acc_nl = ({z_out_2 , 3'b000}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))})
      + 11'b00000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[10:0];
  assign mux_3197_nl = MUX_s_1_2_2(and_tmp_29, and_705_cse, or_359_cse);
  assign and_489_nl = (fsm_output[6]) & (fsm_output[4]) & (fsm_output[0]) & (fsm_output[3]);
  assign mux_3203_nl = MUX_s_1_2_2((~ or_4057_cse), and_489_nl, fsm_output[2]);
  assign mux_3202_nl = MUX_s_1_2_2((~ or_tmp_3801), and_677_cse, fsm_output[2]);
  assign mux_3204_nl = MUX_s_1_2_2(mux_3203_nl, mux_3202_nl, fsm_output[1]);
  assign mux_3205_nl = MUX_s_1_2_2(mux_3204_nl, (fsm_output[6]), fsm_output[5]);
  assign and_449_nl = (fsm_output[6]) & or_tmp_105;
  assign mux_3208_nl = MUX_s_1_2_2(mux_tmp_2965, and_449_nl, fsm_output[2]);
  assign mux_3206_nl = MUX_s_1_2_2((~ or_4007_cse), (fsm_output[4]), fsm_output[6]);
  assign mux_3207_nl = MUX_s_1_2_2(mux_3206_nl, and_tmp_33, fsm_output[2]);
  assign mux_3209_nl = MUX_s_1_2_2(mux_3208_nl, mux_3207_nl, fsm_output[1]);
  assign mux_3210_nl = MUX_s_1_2_2(mux_3209_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_3213_nl = MUX_s_1_2_2((~ or_595_cse), or_tmp_105, fsm_output[6]);
  assign mux_3214_nl = MUX_s_1_2_2(mux_3213_nl, and_tmp_33, fsm_output[2]);
  assign mux_3211_nl = MUX_s_1_2_2((~ or_4007_cse), or_595_cse, fsm_output[6]);
  assign mux_3212_nl = MUX_s_1_2_2(mux_3211_nl, and_tmp_33, fsm_output[2]);
  assign mux_3215_nl = MUX_s_1_2_2(mux_3214_nl, mux_3212_nl, fsm_output[1]);
  assign mux_3216_nl = MUX_s_1_2_2(mux_3215_nl, (fsm_output[6]), fsm_output[5]);
  assign mux_434_nl = MUX_s_1_2_2(and_640_cse, and_tmp_10, fsm_output[2]);
  assign mux_435_nl = MUX_s_1_2_2(mux_434_nl, mux_tmp_293, fsm_output[1]);
  assign mux_3219_nl = MUX_s_1_2_2(mux_221_cse, (~ mux_435_nl), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_111_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110001);
  assign COMP_LOOP_COMP_LOOP_and_1104_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) & COMP_LOOP_nor_985_itm;
  assign or_3932_nl = (fsm_output[6]) | (fsm_output[4]) | and_639_cse;
  assign mux_3221_nl = MUX_s_1_2_2(or_3932_nl, or_341_cse, fsm_output[2]);
  assign or_3929_nl = (fsm_output[6]) | (fsm_output[4]) | and_dcpl_365;
  assign mux_3220_nl = MUX_s_1_2_2(or_341_cse, or_3929_nl, fsm_output[2]);
  assign mux_3222_nl = MUX_s_1_2_2(mux_3221_nl, mux_3220_nl, fsm_output[1]);
  assign mux_3223_nl = MUX_s_1_2_2(mux_3222_nl, (~ mux_180_cse), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_112_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110010);
  assign COMP_LOOP_COMP_LOOP_and_1106_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[2]) & COMP_LOOP_nor_987_itm;
  assign or_3934_nl = (fsm_output[6]) | (((fsm_output[4]) | (fsm_output[0])) & (fsm_output[3]));
  assign mux_3224_nl = MUX_s_1_2_2(or_3934_nl, or_4050_cse, fsm_output[2]);
  assign mux_3225_nl = MUX_s_1_2_2(mux_3224_nl, mux_tmp_2993, fsm_output[1]);
  assign mux_3226_nl = MUX_s_1_2_2(mux_3225_nl, (~ mux_180_cse), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_113_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110011);
  assign COMP_LOOP_COMP_LOOP_and_1110_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) & COMP_LOOP_nor_991_itm;
  assign mux_3227_nl = MUX_s_1_2_2(or_4057_cse, (~ mux_180_cse), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_114_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b110100);
  assign COMP_LOOP_COMP_LOOP_and_1118_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5:4]==2'b11)
      & COMP_LOOP_nor_998_itm;
  assign mux_3228_nl = MUX_s_1_2_2(mux_tmp_2994, mux_tmp_2975, fsm_output[1]);
  assign mux_3229_nl = MUX_s_1_2_2(mux_3228_nl, (~ mux_180_cse), fsm_output[5]);
  assign COMP_LOOP_COMP_LOOP_and_65_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b000011);
  assign COMP_LOOP_COMP_LOOP_and_1370_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[5:4]==2'b11)
      & COMP_LOOP_nor_1222_itm;
  assign mux_3230_nl = MUX_s_1_2_2(mux_tmp_656, mux_tmp_3009, fsm_output[2]);
  assign mux_3231_nl = MUX_s_1_2_2(mux_tmp_3013, mux_3230_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_67_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b000101);
  assign COMP_LOOP_COMP_LOOP_and_1577_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1:0]==2'b11)
      & COMP_LOOP_nor_1403_itm;
  assign COMP_LOOP_COMP_LOOP_and_68_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b000110);
  assign COMP_LOOP_COMP_LOOP_and_1584_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3]) &
      (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) & COMP_LOOP_nor_1410_itm;
  assign COMP_LOOP_COMP_LOOP_and_317_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b000011);
  assign COMP_LOOP_COMP_LOOP_and_1594_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_7_sva[2]) & COMP_LOOP_nor_1420_itm;
  assign COMP_LOOP_COMP_LOOP_and_324_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b001010);
  assign COMP_LOOP_COMP_LOOP_and_1614_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_7_sva[3]) & COMP_LOOP_nor_1439_itm;
  assign COMP_LOOP_COMP_LOOP_and_319_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b000101);
  assign COMP_LOOP_COMP_LOOP_and_1598_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4:3]==2'b11)
      & COMP_LOOP_nor_1424_itm;
  assign nor_403_nl = ~((~((~ (fsm_output[3])) | (fsm_output[5]))) | (fsm_output[7]));
  assign nor_405_nl = ~((fsm_output[3]) | nor_358_cse | (fsm_output[7]));
  assign mux_3241_nl = MUX_s_1_2_2(nor_403_nl, nor_405_nl, fsm_output[1]);
  assign mux_3240_nl = MUX_s_1_2_2(nor_412_cse, and_493_cse, fsm_output[3]);
  assign mux_3242_nl = MUX_s_1_2_2(mux_3241_nl, mux_3240_nl, fsm_output[2]);
  assign mux_3243_nl = MUX_s_1_2_2(mux_3242_nl, and_493_cse, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_and_320_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b000110);
  assign COMP_LOOP_COMP_LOOP_and_1607_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) & COMP_LOOP_nor_1432_itm;
  assign and_458_nl = and_dcpl_94 & and_dcpl_88;
  assign mux_3245_nl = MUX_s_1_2_2(or_tmp_3717, (fsm_output[7]), or_341_cse);
  assign mux_3246_nl = MUX_s_1_2_2(mux_tmp_444, mux_3245_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_321_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b000111);
  assign COMP_LOOP_COMP_LOOP_and_1610_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) &
      (COMP_LOOP_acc_10_cse_10_1_7_sva[2]) & COMP_LOOP_nor_1435_itm;
  assign or_3946_nl = (~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[5])))
      | (fsm_output[7]);
  assign mux_3251_nl = MUX_s_1_2_2(or_3946_nl, or_564_cse, fsm_output[2]);
  assign mux_582_nl = MUX_s_1_2_2((~ or_564_cse), (fsm_output[5]), fsm_output[2]);
  assign mux_3252_nl = MUX_s_1_2_2((~ mux_3251_nl), mux_582_nl, fsm_output[3]);
  assign mux_3253_nl = MUX_s_1_2_2(mux_3252_nl, (fsm_output[5]), fsm_output[4]);
  assign or_3943_nl = (~(and_507_cse | (fsm_output[5]))) | (fsm_output[7]);
  assign mux_3248_nl = MUX_s_1_2_2(or_3943_nl, (fsm_output[7]), fsm_output[3]);
  assign mux_3249_nl = MUX_s_1_2_2(or_564_cse, mux_3248_nl, fsm_output[4]);
  assign COMP_LOOP_COMP_LOOP_and_325_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b001011);
  assign COMP_LOOP_COMP_LOOP_and_1622_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5:4]==2'b11)
      & COMP_LOOP_nor_1446_itm;
  assign and_459_nl = and_dcpl_85 & and_dcpl_377;
  assign mux_3255_nl = MUX_s_1_2_2(or_tmp_404, (fsm_output[7]), fsm_output[6]);
  assign mux_3256_nl = MUX_s_1_2_2(mux_tmp_656, mux_3255_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_69_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b000111);
  assign COMP_LOOP_COMP_LOOP_and_1831_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2]) & (COMP_LOOP_acc_10_cse_10_1_sva[0])
      & COMP_LOOP_nor_1629_itm;
  assign mux_3258_nl = MUX_s_1_2_2(or_tmp_3757, or_tmp_119, fsm_output[4]);
  assign mux_3259_nl = MUX_s_1_2_2((~ mux_3258_nl), and_655_cse, fsm_output[6]);
  assign mux_3261_nl = MUX_s_1_2_2(mux_tmp_3193, mux_3259_nl, fsm_output[2]);
  assign mux_3264_nl = MUX_s_1_2_2(mux_tmp_3196, mux_3261_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_326_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b001100);
  assign COMP_LOOP_COMP_LOOP_and_1832_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2:1]==2'b11)
      & COMP_LOOP_nor_1630_itm;
  assign and_461_nl = and_dcpl_94 & and_dcpl_344;
  assign mux_3271_nl = MUX_s_1_2_2(nor_399_cse, mux_297_cse, fsm_output[5]);
  assign mux_3272_nl = MUX_s_1_2_2(mux_3271_nl, and_tmp_35, and_1046_cse);
  assign mux_3270_nl = MUX_s_1_2_2(and_705_cse, mux_297_cse, fsm_output[5]);
  assign mux_3273_nl = MUX_s_1_2_2(mux_3272_nl, mux_3270_nl, fsm_output[4]);
  assign nor_386_nl = ~((fsm_output[1]) | (~ (fsm_output[5])));
  assign mux_3268_nl = MUX_s_1_2_2(and_705_cse, mux_297_cse, nor_386_nl);
  assign mux_3269_nl = MUX_s_1_2_2(and_tmp_35, mux_3268_nl, fsm_output[4]);
  assign mux_3274_nl = MUX_s_1_2_2(mux_3273_nl, mux_3269_nl, fsm_output[2]);
  assign nor_384_nl = ~((fsm_output[5:4]!=2'b10));
  assign mux_3267_nl = MUX_s_1_2_2(and_705_cse, mux_297_cse, nor_384_nl);
  assign COMP_LOOP_COMP_LOOP_and_327_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b001101);
  assign COMP_LOOP_COMP_LOOP_and_1835_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3]) & (COMP_LOOP_acc_10_cse_10_1_sva[0])
      & COMP_LOOP_nor_1633_itm;
  assign and_463_nl = and_dcpl_264 & and_dcpl_347;
  assign mux_3282_nl = MUX_s_1_2_2(mux_tmp_3214, and_tmp_36, fsm_output[2]);
  assign mux_3278_nl = MUX_s_1_2_2(and_dcpl_60, mux_tmp_3210, fsm_output[6]);
  assign mux_3279_nl = MUX_s_1_2_2(mux_3278_nl, and_tmp_36, fsm_output[2]);
  assign mux_3283_nl = MUX_s_1_2_2(mux_3282_nl, mux_3279_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_328_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b001110);
  assign COMP_LOOP_COMP_LOOP_and_1844_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4]) & (COMP_LOOP_acc_10_cse_10_1_sva[1])
      & COMP_LOOP_nor_1642_itm;
  assign mux_3286_nl = MUX_s_1_2_2(mux_297_cse, mux_tmp_3218, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_329_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b001111);
  assign COMP_LOOP_COMP_LOOP_and_1850_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4:3]==2'b11)
      & COMP_LOOP_nor_1648_itm;
  assign COMP_LOOP_COMP_LOOP_and_331_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010001);
  assign COMP_LOOP_COMP_LOOP_and_1862_nl = (COMP_LOOP_acc_10_cse_10_1_sva[5]) & (COMP_LOOP_acc_10_cse_10_1_sva[2])
      & COMP_LOOP_nor_1659_itm;
  assign and_465_nl = and_dcpl_264 & and_dcpl_116;
  assign and_464_nl = (fsm_output[6]) & mux_tmp_3213;
  assign mux_3291_nl = MUX_s_1_2_2(mux_tmp_3214, and_464_nl, fsm_output[2]);
  assign mux_3289_nl = MUX_s_1_2_2(and_dcpl_60, mux_tmp_3213, fsm_output[6]);
  assign mux_3290_nl = MUX_s_1_2_2(mux_3289_nl, and_tmp_36, fsm_output[2]);
  assign mux_3292_nl = MUX_s_1_2_2(mux_3291_nl, mux_3290_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_332_nl = (COMP_LOOP_2_acc_10_itm_10_1_1[5:0]==6'b010010);
  assign COMP_LOOP_COMP_LOOP_and_1866_nl = (COMP_LOOP_acc_10_cse_10_1_sva[5]) & (COMP_LOOP_acc_10_cse_10_1_sva[3])
      & COMP_LOOP_nor_1663_itm;
  assign and_468_nl = and_dcpl_85 & and_dcpl_116;
  assign mux_3296_nl = MUX_s_1_2_2((~ or_477_cse), or_tmp_404, fsm_output[6]);
  assign and_73_nl = (fsm_output[6]) & or_tmp_404;
  assign mux_3297_nl = MUX_s_1_2_2(mux_3296_nl, and_73_nl, fsm_output[2]);
  assign mux_3294_nl = MUX_s_1_2_2(and_dcpl_60, or_tmp_404, fsm_output[6]);
  assign and_466_nl = (fsm_output[6]) & mux_tmp_3169;
  assign mux_3295_nl = MUX_s_1_2_2(mux_3294_nl, and_466_nl, fsm_output[2]);
  assign mux_3298_nl = MUX_s_1_2_2(mux_3297_nl, mux_3295_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_71_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001001);
  assign COMP_LOOP_COMP_LOOP_and_1874_nl = (COMP_LOOP_acc_10_cse_10_1_sva[5:4]==2'b11)
      & COMP_LOOP_nor_1670_itm;
  assign nor_397_nl = ~(nor_398_cse | (fsm_output[7]));
  assign mux_3300_nl = MUX_s_1_2_2(nor_397_nl, and_655_cse, fsm_output[6]);
  assign mux_3301_nl = MUX_s_1_2_2(mux_tmp_3193, mux_3300_nl, fsm_output[2]);
  assign mux_3302_nl = MUX_s_1_2_2(mux_tmp_3196, mux_3301_nl, fsm_output[1]);
  assign COMP_LOOP_COMP_LOOP_and_72_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001010);
  assign COMP_LOOP_COMP_LOOP_and_583_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[4]) &
      (COMP_LOOP_acc_10_cse_10_1_3_sva[0]) & COMP_LOOP_nor_521_itm;
  assign mux_3306_nl = MUX_s_1_2_2(mux_3305_itm, (~ and_779_cse), fsm_output[5]);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_2_nl = (z_out_8[2:0]==3'b011);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_4_nl = (z_out_8[2:0]==3'b101);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_5_nl = (z_out_8[2:0]==3'b110);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_6_nl = (z_out_8[2:0]==3'b111);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_nor_nl = ~((z_out_8[2:0]!=3'b000));
  assign COMP_LOOP_COMP_LOOP_and_76_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001110);
  assign COMP_LOOP_COMP_LOOP_and_77_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b001111);
  assign COMP_LOOP_COMP_LOOP_and_79_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010001);
  assign COMP_LOOP_COMP_LOOP_and_80_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010010);
  assign COMP_LOOP_COMP_LOOP_and_81_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010011);
  assign COMP_LOOP_COMP_LOOP_and_82_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010100);
  assign COMP_LOOP_COMP_LOOP_and_83_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010101);
  assign COMP_LOOP_COMP_LOOP_and_84_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010110);
  assign COMP_LOOP_COMP_LOOP_and_85_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b010111);
  assign COMP_LOOP_COMP_LOOP_and_86_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011000);
  assign COMP_LOOP_COMP_LOOP_and_87_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011001);
  assign COMP_LOOP_COMP_LOOP_and_88_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011010);
  assign COMP_LOOP_COMP_LOOP_and_89_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011011);
  assign COMP_LOOP_COMP_LOOP_and_90_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011100);
  assign COMP_LOOP_COMP_LOOP_and_91_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011101);
  assign COMP_LOOP_COMP_LOOP_and_92_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011110);
  assign COMP_LOOP_COMP_LOOP_and_93_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b011111);
  assign COMP_LOOP_COMP_LOOP_and_95_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100001);
  assign COMP_LOOP_COMP_LOOP_and_96_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100010);
  assign COMP_LOOP_COMP_LOOP_and_97_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100011);
  assign COMP_LOOP_COMP_LOOP_and_98_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100100);
  assign COMP_LOOP_COMP_LOOP_and_99_nl = (COMP_LOOP_1_acc_10_itm_10_1_1[5:0]==6'b100101);
  assign COMP_LOOP_COMP_LOOP_nor_1_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5:0]!=6'b000000));
  assign COMP_LOOP_nor_57_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5:1]!=5'b00000));
  assign COMP_LOOP_nor_58_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5]) | (COMP_LOOP_1_acc_10_itm_10_1_1[4])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[3]) | (COMP_LOOP_1_acc_10_itm_10_1_1[2]) |
      (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_60_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5]) | (COMP_LOOP_1_acc_10_itm_10_1_1[4])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[3]) | (COMP_LOOP_1_acc_10_itm_10_1_1[1]) |
      (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_64_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5]) | (COMP_LOOP_1_acc_10_itm_10_1_1[4])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[2]) | (COMP_LOOP_1_acc_10_itm_10_1_1[1]) |
      (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_72_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[5]) | (COMP_LOOP_1_acc_10_itm_10_1_1[3])
      | (COMP_LOOP_1_acc_10_itm_10_1_1[2]) | (COMP_LOOP_1_acc_10_itm_10_1_1[1]) |
      (COMP_LOOP_1_acc_10_itm_10_1_1[0]));
  assign COMP_LOOP_nor_87_nl = ~((COMP_LOOP_1_acc_10_itm_10_1_1[4:0]!=5'b00000));
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_nl = (COMP_LOOP_1_tmp_mul_idiv_sva_2_0==3'b001);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_1_nl = (COMP_LOOP_1_tmp_mul_idiv_sva_2_0==3'b010);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_3_nl = (COMP_LOOP_1_tmp_mul_idiv_sva_2_0==3'b100);
  assign COMP_LOOP_COMP_LOOP_mux_21_nl = MUX_v_64_2_2(COMP_LOOP_1_acc_8_itm, z_out_9,
      COMP_LOOP_or_65_itm);
  assign nl_COMP_LOOP_acc_17_nl = COMP_LOOP_mux_724_cse + COMP_LOOP_COMP_LOOP_mux_21_nl;
  assign COMP_LOOP_acc_17_nl = nl_COMP_LOOP_acc_17_nl[63:0];
  assign COMP_LOOP_or_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_61_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_60_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_59_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_58_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_57_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_56_itm & and_dcpl_109);
  assign COMP_LOOP_or_1_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[0]) & COMP_LOOP_tmp_nor_10_itm
      & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_61_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_60_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_59_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_58_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_57_itm & and_dcpl_109);
  assign COMP_LOOP_or_2_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[1]) & COMP_LOOP_tmp_nor_151_itm
      & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_1518_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_61_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_60_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_59_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_58_itm & and_dcpl_109);
  assign COMP_LOOP_or_3_nl = (COMP_LOOP_COMP_LOOP_and_1370_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_760_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_1518_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_61_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_60_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_59_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_4_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[2]) & COMP_LOOP_tmp_nor_153_itm
      & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_761_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_760_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_1518_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_61_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_60_itm & and_dcpl_109);
  assign COMP_LOOP_or_5_nl = (COMP_LOOP_COMP_LOOP_and_1577_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_509_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_761_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_760_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_1518_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_61_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_6_nl = (COMP_LOOP_COMP_LOOP_and_1584_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_510_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_509_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_761_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_760_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_1518_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_7_nl = (COMP_LOOP_COMP_LOOP_and_1831_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_258_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_510_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_509_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_761_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_760_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_1518_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_8_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[3]) & COMP_LOOP_tmp_nor_157_itm
      & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_258_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_510_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_509_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_761_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_760_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_1518_itm & and_dcpl_109);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_1874_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_260_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_258_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_510_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_509_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_761_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_760_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_583_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_261_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_260_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_258_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_510_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_509_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_761_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_73_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_262_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_261_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_260_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_258_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_510_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_509_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_74_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_262_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_261_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_260_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_258_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_510_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_75_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_264_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_262_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_261_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_260_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_258_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_264_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_262_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_261_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_260_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_109);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_264_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_262_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_261_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_260_itm & and_dcpl_109);
  assign COMP_LOOP_or_16_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[4]) & COMP_LOOP_tmp_nor_165_itm
      & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_264_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_262_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_261_itm & and_dcpl_109);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_268_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_264_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_262_itm & and_dcpl_109);
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_522_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_268_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_264_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_109);
  assign COMP_LOOP_or_19_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_270_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_522_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_268_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_264_itm & and_dcpl_109);
  assign COMP_LOOP_or_20_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_270_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_522_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_268_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_109);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_272_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_18_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_270_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_522_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_268_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_109);
  assign COMP_LOOP_or_22_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_272_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_270_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_522_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_268_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_109);
  assign COMP_LOOP_or_23_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_20_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_272_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_18_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_270_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_522_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_268_itm & and_dcpl_109);
  assign COMP_LOOP_or_24_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_21_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_272_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_270_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_522_itm & and_dcpl_109);
  assign COMP_LOOP_or_25_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_22_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_20_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_272_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_18_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_270_itm & and_dcpl_109);
  assign COMP_LOOP_or_26_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_23_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_21_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_272_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_18_itm & and_dcpl_109);
  assign COMP_LOOP_or_27_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_24_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_22_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_20_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_272_itm & and_dcpl_109);
  assign COMP_LOOP_or_28_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_25_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_23_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_21_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_20_itm & and_dcpl_109);
  assign COMP_LOOP_or_29_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_26_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_24_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_22_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_21_itm & and_dcpl_109);
  assign COMP_LOOP_or_30_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_27_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_25_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_23_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_22_itm & and_dcpl_109);
  assign COMP_LOOP_or_31_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_28_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_26_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_24_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_23_itm & and_dcpl_109);
  assign COMP_LOOP_or_32_nl = ((COMP_LOOP_acc_10_cse_10_1_1_sva[5]) & COMP_LOOP_tmp_nor_180_itm
      & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_29_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_27_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_25_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_24_itm & and_dcpl_109);
  assign COMP_LOOP_or_33_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_284_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_28_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_26_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_25_itm & and_dcpl_109);
  assign COMP_LOOP_or_34_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_285_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_284_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_29_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_27_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_26_itm & and_dcpl_109);
  assign COMP_LOOP_or_35_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_286_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_285_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_284_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_28_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_27_itm & and_dcpl_109);
  assign COMP_LOOP_or_36_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_34_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_286_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_285_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_284_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_30_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_29_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_28_itm & and_dcpl_109);
  assign COMP_LOOP_or_37_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & and_dcpl_77)
      | (COMP_LOOP_COMP_LOOP_and_288_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_286_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_285_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_284_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_29_itm & and_dcpl_109);
  assign COMP_LOOP_or_38_nl = (COMP_LOOP_COMP_LOOP_and_100_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_36_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_288_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_286_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_285_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_284_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_30_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_39_nl = (COMP_LOOP_COMP_LOOP_and_101_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_37_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_36_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_288_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_34_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_286_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_285_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_284_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_40_nl = (COMP_LOOP_COMP_LOOP_and_102_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_38_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_37_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_36_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_288_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_286_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_285_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_41_nl = (COMP_LOOP_COMP_LOOP_and_103_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_39_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_38_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_37_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_36_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_288_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_34_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_286_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_42_nl = (COMP_LOOP_COMP_LOOP_and_104_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_40_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_39_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_38_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_37_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_36_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_288_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_34_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_43_nl = (COMP_LOOP_COMP_LOOP_and_105_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_41_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_40_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_39_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_38_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_37_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_36_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_288_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_44_nl = (COMP_LOOP_COMP_LOOP_and_106_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_42_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_41_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_40_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_39_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_38_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_37_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_36_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_45_nl = (COMP_LOOP_COMP_LOOP_and_107_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_43_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_42_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_41_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_40_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_39_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_38_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_37_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_46_nl = (COMP_LOOP_COMP_LOOP_and_108_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_44_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_43_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_42_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_41_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_40_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_39_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_38_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_47_nl = (COMP_LOOP_COMP_LOOP_and_109_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_45_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_44_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_43_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_42_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_41_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_40_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_39_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_48_nl = (COMP_LOOP_COMP_LOOP_and_110_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_46_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_45_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_44_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_43_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_42_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_41_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_40_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_49_nl = (COMP_LOOP_COMP_LOOP_and_1104_itm & and_dcpl_77) |
      (COMP_LOOP_COMP_LOOP_and_47_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_46_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_45_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_44_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_43_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_42_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_41_itm & and_dcpl_109);
  assign COMP_LOOP_or_50_nl = (COMP_LOOP_COMP_LOOP_and_1106_itm & and_dcpl_77) |
      (COMP_LOOP_COMP_LOOP_and_48_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_47_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_46_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_45_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_44_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_43_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_42_itm & and_dcpl_109);
  assign COMP_LOOP_or_51_nl = (COMP_LOOP_COMP_LOOP_and_1110_itm & and_dcpl_77) |
      (COMP_LOOP_COMP_LOOP_and_49_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_48_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_47_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_46_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_45_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_44_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_43_itm & and_dcpl_109);
  assign COMP_LOOP_or_52_nl = (COMP_LOOP_COMP_LOOP_and_1118_itm & and_dcpl_77) |
      (COMP_LOOP_COMP_LOOP_and_50_itm & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_49_itm
      & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_48_itm & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_47_itm
      & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_46_itm & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_45_itm
      & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_44_itm & and_dcpl_109);
  assign COMP_LOOP_or_53_nl = (COMP_LOOP_COMP_LOOP_and_115_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_51_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_50_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_49_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_48_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_47_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_46_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_45_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_54_nl = (COMP_LOOP_COMP_LOOP_and_116_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_52_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_51_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_50_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_49_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_48_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_47_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_46_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_55_nl = (COMP_LOOP_COMP_LOOP_and_117_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_53_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_52_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_51_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_50_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_49_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_48_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_47_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_56_nl = (COMP_LOOP_COMP_LOOP_and_118_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_54_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_53_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_52_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_51_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_50_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_49_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_48_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_57_nl = (COMP_LOOP_COMP_LOOP_and_119_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_55_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_54_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_53_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_52_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_51_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_50_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_49_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_58_nl = (COMP_LOOP_COMP_LOOP_and_120_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_56_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_55_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_54_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_53_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_52_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_51_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_50_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_59_nl = (COMP_LOOP_COMP_LOOP_and_121_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_57_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_56_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_55_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_54_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_53_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_52_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_51_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_60_nl = (COMP_LOOP_COMP_LOOP_and_122_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_58_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_57_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_56_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_55_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_54_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_53_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_52_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_61_nl = (COMP_LOOP_COMP_LOOP_and_123_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_59_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_58_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_57_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_56_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_55_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_54_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_53_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_62_nl = (COMP_LOOP_COMP_LOOP_and_124_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_60_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_59_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_58_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_57_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_56_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_55_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_54_itm
      & and_dcpl_109);
  assign COMP_LOOP_or_63_nl = (COMP_LOOP_COMP_LOOP_and_125_itm & and_dcpl_77) | (COMP_LOOP_COMP_LOOP_and_61_itm
      & and_dcpl_86) | (COMP_LOOP_COMP_LOOP_and_60_itm & and_dcpl_90) | (COMP_LOOP_COMP_LOOP_and_59_itm
      & and_dcpl_95) | (COMP_LOOP_COMP_LOOP_and_58_itm & and_dcpl_99) | (COMP_LOOP_COMP_LOOP_and_57_itm
      & and_dcpl_104) | (COMP_LOOP_COMP_LOOP_and_56_itm & and_dcpl_106) | (COMP_LOOP_COMP_LOOP_and_55_itm
      & and_dcpl_109);
  assign COMP_LOOP_tmp_and_249_nl = COMP_LOOP_COMP_LOOP_and_119_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_7_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_153_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_8_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[1])
      & COMP_LOOP_tmp_nor_165_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_250_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_10_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[2])
      & COMP_LOOP_tmp_nor_180_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_251_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_252_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_253_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_14_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_10_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_254_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_255_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_256_nl = COMP_LOOP_COMP_LOOP_and_102_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_257_nl = COMP_LOOP_COMP_LOOP_and_106_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_258_nl = COMP_LOOP_COMP_LOOP_and_107_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_259_nl = COMP_LOOP_COMP_LOOP_and_108_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_260_nl = COMP_LOOP_COMP_LOOP_and_109_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_22_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[4])
      & COMP_LOOP_tmp_nor_151_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_261_nl = COMP_LOOP_COMP_LOOP_and_110_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_262_nl = COMP_LOOP_COMP_LOOP_and_1104_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_263_nl = COMP_LOOP_COMP_LOOP_and_1106_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_264_nl = COMP_LOOP_COMP_LOOP_and_1118_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_265_nl = COMP_LOOP_COMP_LOOP_and_115_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_266_nl = COMP_LOOP_COMP_LOOP_and_116_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_267_nl = COMP_LOOP_COMP_LOOP_and_117_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_268_nl = COMP_LOOP_COMP_LOOP_and_118_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_269_nl = COMP_LOOP_COMP_LOOP_and_120_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_270_nl = COMP_LOOP_COMP_LOOP_and_121_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_271_nl = COMP_LOOP_COMP_LOOP_and_122_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_272_nl = COMP_LOOP_COMP_LOOP_and_123_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_273_nl = COMP_LOOP_COMP_LOOP_and_124_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_274_nl = COMP_LOOP_COMP_LOOP_and_125_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_275_nl = COMP_LOOP_COMP_LOOP_and_1370_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_38_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[5])
      & COMP_LOOP_tmp_nor_157_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_276_nl = COMP_LOOP_COMP_LOOP_and_1831_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_277_nl = COMP_LOOP_COMP_LOOP_and_1874_itm & (~ and_474_tmp);
  assign COMP_LOOP_tmp_and_278_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_279_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_280_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_281_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_282_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_283_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_284_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_285_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_286_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_287_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_288_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_289_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_290_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_291_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_292_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_293_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_294_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_295_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_296_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_297_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_298_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_299_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_300_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_301_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_302_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_303_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_304_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_305_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_306_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm & (~
      and_474_tmp);
  assign COMP_LOOP_tmp_and_222_nl = COMP_LOOP_COMP_LOOP_and_1874_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_70_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_4_0[0])
      & COMP_LOOP_tmp_nor_206_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_71_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_4_0[1])
      & COMP_LOOP_tmp_nor_207_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_223_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~
      nor_1579_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_73_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_4_0[2])
      & COMP_LOOP_tmp_nor_209_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_224_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & (~
      nor_1579_tmp);
  assign COMP_LOOP_tmp_and_225_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~
      nor_1579_tmp);
  assign COMP_LOOP_tmp_and_226_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~
      nor_1579_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_77_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_4_0[3])
      & COMP_LOOP_tmp_nor_213_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_227_nl = COMP_LOOP_COMP_LOOP_and_102_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_228_nl = COMP_LOOP_COMP_LOOP_and_106_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_229_nl = COMP_LOOP_COMP_LOOP_and_107_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_230_nl = COMP_LOOP_COMP_LOOP_and_108_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_231_nl = COMP_LOOP_COMP_LOOP_and_109_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_232_nl = COMP_LOOP_COMP_LOOP_and_110_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_233_nl = COMP_LOOP_COMP_LOOP_and_1104_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_85_nl = (COMP_LOOP_3_tmp_mul_idiv_sva_4_0[4])
      & COMP_LOOP_tmp_nor_220_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_234_nl = COMP_LOOP_COMP_LOOP_and_1106_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_235_nl = COMP_LOOP_COMP_LOOP_and_1118_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_236_nl = COMP_LOOP_COMP_LOOP_and_115_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_237_nl = COMP_LOOP_COMP_LOOP_and_116_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_238_nl = COMP_LOOP_COMP_LOOP_and_117_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_239_nl = COMP_LOOP_COMP_LOOP_and_118_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_240_nl = COMP_LOOP_COMP_LOOP_and_120_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_241_nl = COMP_LOOP_COMP_LOOP_and_121_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_242_nl = COMP_LOOP_COMP_LOOP_and_122_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_243_nl = COMP_LOOP_COMP_LOOP_and_123_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_244_nl = COMP_LOOP_COMP_LOOP_and_124_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_245_nl = COMP_LOOP_COMP_LOOP_and_125_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_246_nl = COMP_LOOP_COMP_LOOP_and_1370_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_247_nl = COMP_LOOP_COMP_LOOP_and_1831_itm & (~ nor_1579_tmp);
  assign COMP_LOOP_tmp_and_248_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & (~
      nor_1579_tmp);
  assign COMP_LOOP_tmp_and_164_nl = COMP_LOOP_COMP_LOOP_and_119_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_101_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_151_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_102_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[1])
      & COMP_LOOP_tmp_nor_153_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_165_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_104_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[2])
      & COMP_LOOP_tmp_nor_157_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_166_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_167_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_168_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_108_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_165_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_169_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_170_nl = COMP_LOOP_COMP_LOOP_and_102_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_171_nl = COMP_LOOP_COMP_LOOP_and_106_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_172_nl = COMP_LOOP_COMP_LOOP_and_107_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_173_nl = COMP_LOOP_COMP_LOOP_and_108_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_174_nl = COMP_LOOP_COMP_LOOP_and_109_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_175_nl = COMP_LOOP_COMP_LOOP_and_110_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_116_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[4])
      & COMP_LOOP_tmp_nor_180_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_176_nl = COMP_LOOP_COMP_LOOP_and_1104_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_177_nl = COMP_LOOP_COMP_LOOP_and_1106_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_178_nl = COMP_LOOP_COMP_LOOP_and_1118_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_179_nl = COMP_LOOP_COMP_LOOP_and_115_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_180_nl = COMP_LOOP_COMP_LOOP_and_116_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_181_nl = COMP_LOOP_COMP_LOOP_and_117_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_182_nl = COMP_LOOP_COMP_LOOP_and_118_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_183_nl = COMP_LOOP_COMP_LOOP_and_120_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_184_nl = COMP_LOOP_COMP_LOOP_and_121_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_185_nl = COMP_LOOP_COMP_LOOP_and_122_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_186_nl = COMP_LOOP_COMP_LOOP_and_123_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_187_nl = COMP_LOOP_COMP_LOOP_and_124_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_188_nl = COMP_LOOP_COMP_LOOP_and_125_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_189_nl = COMP_LOOP_COMP_LOOP_and_1370_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_190_nl = COMP_LOOP_COMP_LOOP_and_1831_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_132_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[5])
      & COMP_LOOP_tmp_nor_10_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_191_nl = COMP_LOOP_COMP_LOOP_and_1874_itm & (~ and_476_tmp);
  assign COMP_LOOP_tmp_and_192_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_193_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_194_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_195_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_196_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_197_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_198_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_199_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_200_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_201_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_202_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_203_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_204_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_205_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_206_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_207_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_208_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_209_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_210_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_211_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_212_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_213_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_214_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_215_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_216_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_217_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_218_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_219_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_220_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_221_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm & (~
      and_476_tmp);
  assign COMP_LOOP_tmp_and_152_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_4_itm & (~ nor_tmp_396);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_164_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_140_itm & (~ nor_tmp_396);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_165_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[1])
      & COMP_LOOP_tmp_nor_141_itm & (~ nor_tmp_396);
  assign COMP_LOOP_tmp_and_153_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_166_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_167_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[2])
      & COMP_LOOP_tmp_nor_143_itm & (~ nor_tmp_396);
  assign COMP_LOOP_tmp_and_154_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_168_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_155_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_169_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_156_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_170_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_171_nl = (COMP_LOOP_5_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_146_itm & (~ nor_tmp_396);
  assign COMP_LOOP_tmp_and_157_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_172_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_158_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_173_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_159_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_174_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_160_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_175_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_161_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_176_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_162_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_177_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_163_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_178_itm & (~
      nor_tmp_396);
  assign COMP_LOOP_tmp_and_89_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_90_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_274_rgt & and_478_m1c;
  assign COMP_LOOP_tmp_and_91_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_92_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_276_rgt & and_478_m1c;
  assign COMP_LOOP_tmp_and_93_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_94_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_95_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_96_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_280_rgt & and_478_m1c;
  assign COMP_LOOP_tmp_and_97_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_98_nl = COMP_LOOP_COMP_LOOP_and_102_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_99_nl = COMP_LOOP_COMP_LOOP_and_106_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_100_nl = COMP_LOOP_COMP_LOOP_and_107_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_101_nl = COMP_LOOP_COMP_LOOP_and_108_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_102_nl = COMP_LOOP_COMP_LOOP_and_109_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_103_nl = COMP_LOOP_COMP_LOOP_and_110_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_104_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_288_rgt & and_478_m1c;
  assign COMP_LOOP_tmp_and_105_nl = COMP_LOOP_COMP_LOOP_and_1104_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_106_nl = COMP_LOOP_COMP_LOOP_and_1106_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_107_nl = COMP_LOOP_COMP_LOOP_and_1118_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_108_nl = COMP_LOOP_COMP_LOOP_and_115_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_109_nl = COMP_LOOP_COMP_LOOP_and_116_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_110_nl = COMP_LOOP_COMP_LOOP_and_117_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_111_nl = COMP_LOOP_COMP_LOOP_and_118_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_112_nl = COMP_LOOP_COMP_LOOP_and_120_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_113_nl = COMP_LOOP_COMP_LOOP_and_121_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_114_nl = COMP_LOOP_COMP_LOOP_and_122_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_115_nl = COMP_LOOP_COMP_LOOP_and_123_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_116_nl = COMP_LOOP_COMP_LOOP_and_124_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_117_nl = COMP_LOOP_COMP_LOOP_and_125_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_118_nl = COMP_LOOP_COMP_LOOP_and_1370_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_119_nl = COMP_LOOP_COMP_LOOP_and_1831_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_120_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_304_rgt & and_478_m1c;
  assign COMP_LOOP_tmp_and_121_nl = COMP_LOOP_COMP_LOOP_and_1874_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_122_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_123_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_124_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_125_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_126_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_127_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_128_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_129_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_130_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_131_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_132_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_133_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_134_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_135_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_136_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_137_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_138_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_139_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_140_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_141_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_142_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_143_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_144_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_145_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_146_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_147_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_148_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_149_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_150_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm & and_478_m1c;
  assign COMP_LOOP_tmp_and_151_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm & and_478_m1c;
  assign mux_3350_nl = MUX_s_1_2_2(not_tmp_88, nor_tmp_391, fsm_output[6]);
  assign mux_3351_nl = MUX_s_1_2_2(mux_3350_nl, mux_tmp_3280, fsm_output[2]);
  assign mux_3348_nl = MUX_s_1_2_2(not_tmp_868, nor_tmp_391, fsm_output[6]);
  assign mux_3349_nl = MUX_s_1_2_2(mux_3348_nl, mux_tmp_3280, fsm_output[2]);
  assign mux_3352_nl = MUX_s_1_2_2(mux_3351_nl, mux_3349_nl, fsm_output[1]);
  assign mux_3353_nl = MUX_s_1_2_2(mux_3352_nl, and_705_cse, fsm_output[5]);
  assign COMP_LOOP_tmp_and_31_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_5_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_179_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[0])
      & COMP_LOOP_tmp_nor_10_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_180_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[1])
      & COMP_LOOP_tmp_nor_151_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_32_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_100_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_182_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[2])
      & COMP_LOOP_tmp_nor_153_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_33_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_105_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_34_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_106_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_35_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_107_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_186_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[3])
      & COMP_LOOP_tmp_nor_157_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_36_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_109_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_37_nl = COMP_LOOP_COMP_LOOP_and_102_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_38_nl = COMP_LOOP_COMP_LOOP_and_106_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_39_nl = COMP_LOOP_COMP_LOOP_and_107_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_40_nl = COMP_LOOP_COMP_LOOP_and_108_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_41_nl = COMP_LOOP_COMP_LOOP_and_109_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_42_nl = COMP_LOOP_COMP_LOOP_and_110_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_194_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[4])
      & COMP_LOOP_tmp_nor_165_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_43_nl = COMP_LOOP_COMP_LOOP_and_1104_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_44_nl = COMP_LOOP_COMP_LOOP_and_1106_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_45_nl = COMP_LOOP_COMP_LOOP_and_1118_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_46_nl = COMP_LOOP_COMP_LOOP_and_115_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_47_nl = COMP_LOOP_COMP_LOOP_and_116_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_48_nl = COMP_LOOP_COMP_LOOP_and_117_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_49_nl = COMP_LOOP_COMP_LOOP_and_118_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_50_nl = COMP_LOOP_COMP_LOOP_and_120_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_51_nl = COMP_LOOP_COMP_LOOP_and_121_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_52_nl = COMP_LOOP_COMP_LOOP_and_122_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_53_nl = COMP_LOOP_COMP_LOOP_and_123_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_54_nl = COMP_LOOP_COMP_LOOP_and_124_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_55_nl = COMP_LOOP_COMP_LOOP_and_125_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_56_nl = COMP_LOOP_COMP_LOOP_and_1370_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_57_nl = COMP_LOOP_COMP_LOOP_and_1831_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_210_nl = (COMP_LOOP_2_tmp_mul_idiv_sva[5])
      & COMP_LOOP_tmp_nor_180_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_58_nl = COMP_LOOP_COMP_LOOP_and_1874_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_59_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_134_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_60_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_135_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_61_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_136_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_62_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_137_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_63_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_138_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_64_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_139_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_65_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_140_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_66_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_141_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_67_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_142_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_68_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_143_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_69_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_144_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_70_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_145_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_71_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_146_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_72_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_147_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_73_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_148_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_74_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_149_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_75_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_150_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_76_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_151_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_77_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_152_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_78_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_153_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_79_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_154_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_80_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_155_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_81_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_156_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_82_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_157_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_83_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_158_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_84_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_159_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_85_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_160_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_86_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_161_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_87_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_162_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_88_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_163_itm & mux_3360_tmp;
  assign COMP_LOOP_tmp_and_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_nor_6_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_1_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_243_rgt & and_dcpl_265;
  assign COMP_LOOP_tmp_and_2_nl = COMP_LOOP_COMP_LOOP_and_119_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_3_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_245_rgt & and_dcpl_265;
  assign COMP_LOOP_tmp_and_4_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_246_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_5_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_247_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_6_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_248_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_7_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_249_rgt & and_dcpl_265;
  assign COMP_LOOP_tmp_and_8_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_250_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_9_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_251_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_10_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_252_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_11_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_253_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_12_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_254_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_13_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_255_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_14_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_256_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_15_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_257_rgt & and_dcpl_265;
  assign COMP_LOOP_tmp_and_16_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_258_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_17_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_259_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_18_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_260_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_19_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_261_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_20_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_262_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_21_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_263_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_22_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_264_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_23_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_265_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_24_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_266_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_25_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_267_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_26_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_268_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_27_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_269_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_28_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_270_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_29_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_271_itm & and_dcpl_265;
  assign COMP_LOOP_tmp_and_30_nl = COMP_LOOP_tmp_COMP_LOOP_tmp_and_272_itm & and_dcpl_265;
  assign mux_3362_nl = MUX_s_1_2_2(not_tmp_88, (fsm_output[7]), fsm_output[6]);
  assign mux_3363_nl = MUX_s_1_2_2(mux_3362_nl, mux_tmp_3100, or_359_cse);
  assign mux_3361_nl = MUX_s_1_2_2(nor_tmp_391, (fsm_output[7]), fsm_output[6]);
  assign mux_3364_nl = MUX_s_1_2_2(mux_3363_nl, mux_3361_nl, fsm_output[5]);
  assign and_1047_nl = and_dcpl_58 & (~ (fsm_output[3])) & (fsm_output[6]) & (fsm_output[2])
      & (~ (fsm_output[1])) & (fsm_output[7]) & (fsm_output[5]);
  assign COMP_LOOP_mux_721_nl = MUX_v_7_2_2(COMP_LOOP_k_10_3_sva_6_0, ({3'b001 ,
      (~ z_out_4)}), and_1047_nl);
  assign nl_z_out_2 = conv_u2u_7_8(COMP_LOOP_mux_721_nl) + 8'b00000001;
  assign z_out_2 = nl_z_out_2[7:0];
  assign COMP_LOOP_mux_722_nl = MUX_v_11_2_2(({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[10:1]))}),
      STAGE_LOOP_lshift_psp_sva, and_dcpl_488);
  assign COMP_LOOP_COMP_LOOP_nand_1_nl = ~(and_dcpl_488 & (~(and_dcpl_58 & nor_1715_cse
      & and_dcpl_477 & nor_1716_cse)));
  assign COMP_LOOP_mux_723_nl = MUX_v_10_2_2(({COMP_LOOP_k_10_3_sva_6_0 , 3'b001}),
      VEC_LOOP_j_10_0_sva_9_0, and_dcpl_488);
  assign nl_acc_1_nl = ({COMP_LOOP_mux_722_nl , COMP_LOOP_COMP_LOOP_nand_1_nl}) +
      conv_u2u_11_12({COMP_LOOP_mux_723_nl , 1'b1});
  assign acc_1_nl = nl_acc_1_nl[11:0];
  assign z_out_3 = readslicef_12_11_1(acc_1_nl);
  assign STAGE_LOOP_mux_4_nl = MUX_v_4_2_2(STAGE_LOOP_i_3_0_sva, (~ STAGE_LOOP_i_3_0_sva),
      and_dcpl_501);
  assign nl_z_out_4 = STAGE_LOOP_mux_4_nl + ({1'b1 , (~ and_dcpl_501) , 2'b11});
  assign z_out_4 = nl_z_out_4[3:0];
  assign COMP_LOOP_mux_724_cse = MUX_v_64_2_2(z_out_9, COMP_LOOP_1_acc_8_itm, COMP_LOOP_or_65_itm);
  assign COMP_LOOP_tmp_nor_300_cse = ~(and_dcpl_574 | and_dcpl_589 | and_dcpl_590);
  assign COMP_LOOP_tmp_mux_64_nl = MUX_s_1_2_2((z_out_1[9]), (COMP_LOOP_2_tmp_lshift_ncse_sva[9]),
      COMP_LOOP_tmp_or_54_ssc);
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_and_337_nl = COMP_LOOP_tmp_mux_64_nl & COMP_LOOP_tmp_nor_300_cse;
  assign COMP_LOOP_tmp_or_88_nl = and_dcpl_577 | and_dcpl_589;
  assign COMP_LOOP_tmp_mux1h_146_nl = MUX1HOT_v_9_4_2(({1'b0 , (z_out[7:0])}), (z_out_1[8:0]),
      (COMP_LOOP_2_tmp_lshift_ncse_sva[8:0]), COMP_LOOP_3_tmp_lshift_ncse_sva, {and_dcpl_574
      , COMP_LOOP_tmp_or_88_nl , COMP_LOOP_tmp_or_54_ssc , and_dcpl_590});
  assign COMP_LOOP_tmp_and_312_nl = (COMP_LOOP_k_10_3_sva_6_0[6]) & COMP_LOOP_tmp_nor_300_cse;
  assign COMP_LOOP_tmp_or_89_nl = and_dcpl_577 | and_dcpl_580 | and_dcpl_583 | and_dcpl_588;
  assign COMP_LOOP_tmp_mux1h_147_nl = MUX1HOT_v_6_3_2(({1'b0 , (COMP_LOOP_k_10_3_sva_6_0[6:2])}),
      (COMP_LOOP_k_10_3_sva_6_0[5:0]), (COMP_LOOP_k_10_3_sva_6_0[6:1]), {and_dcpl_574
      , COMP_LOOP_tmp_or_89_nl , COMP_LOOP_tmp_or_83_itm});
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_mux_17_nl = MUX_s_1_2_2((COMP_LOOP_k_10_3_sva_6_0[1]),
      (COMP_LOOP_k_10_3_sva_6_0[0]), COMP_LOOP_tmp_or_83_itm);
  assign COMP_LOOP_tmp_or_90_nl = (COMP_LOOP_tmp_COMP_LOOP_tmp_mux_17_nl & (~(and_dcpl_577
      | and_dcpl_580))) | and_dcpl_583 | and_dcpl_588;
  assign COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl = ((COMP_LOOP_k_10_3_sva_6_0[0]) & (~(and_dcpl_577
      | and_dcpl_583 | and_dcpl_589))) | and_dcpl_580 | and_dcpl_588 | and_dcpl_590;
  assign nl_z_out_7 = ({COMP_LOOP_tmp_COMP_LOOP_tmp_and_337_nl , COMP_LOOP_tmp_mux1h_146_nl})
      * ({COMP_LOOP_tmp_and_312_nl , COMP_LOOP_tmp_mux1h_147_nl , COMP_LOOP_tmp_or_90_nl
      , COMP_LOOP_tmp_COMP_LOOP_tmp_or_1_nl , 1'b1});
  assign z_out_7 = nl_z_out_7[9:0];
  assign and_1048_nl = and_dcpl_573 & (fsm_output[2:1]==2'b01) & nor_1716_cse;
  assign COMP_LOOP_tmp_mux1h_148_nl = MUX1HOT_v_64_9_2(({57'b000000000000000000000000000000000000000000000000000000000
      , (z_out_1[6:0])}), COMP_LOOP_tmp_mux1h_itm, COMP_LOOP_tmp_mux1h_1_itm, COMP_LOOP_tmp_mux1h_2_itm,
      COMP_LOOP_tmp_mux1h_3_itm, COMP_LOOP_tmp_mux1h_4_itm, COMP_LOOP_tmp_mux1h_5_itm,
      COMP_LOOP_tmp_mux1h_6_itm, tmp_21_sva_1, {and_1048_nl , and_dcpl_602 , and_dcpl_608
      , and_dcpl_611 , and_dcpl_614 , and_dcpl_617 , and_dcpl_620 , and_dcpl_623
      , and_dcpl_625});
  assign COMP_LOOP_tmp_or_91_nl = and_dcpl_602 | and_dcpl_608 | and_dcpl_611 | and_dcpl_614
      | and_dcpl_617 | and_dcpl_620 | and_dcpl_623 | and_dcpl_625;
  assign COMP_LOOP_tmp_mux_65_nl = MUX_v_64_2_2(({57'b000000000000000000000000000000000000000000000000000000000
      , COMP_LOOP_k_10_3_sva_6_0}), COMP_LOOP_1_modulo_dev_cmp_return_rsc_z, COMP_LOOP_tmp_or_91_nl);
  assign nl_z_out_8 = COMP_LOOP_tmp_mux1h_148_nl * COMP_LOOP_tmp_mux_65_nl;
  assign z_out_8 = nl_z_out_8[63:0];
  assign COMP_LOOP_mux1h_1267_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_nor_itm, COMP_LOOP_COMP_LOOP_nor_5_itm,
      COMP_LOOP_COMP_LOOP_nor_9_itm, COMP_LOOP_COMP_LOOP_nor_13_itm, COMP_LOOP_COMP_LOOP_nor_17_itm,
      COMP_LOOP_COMP_LOOP_nor_21_itm, COMP_LOOP_COMP_LOOP_nor_25_itm, COMP_LOOP_COMP_LOOP_nor_29_itm,
      {and_dcpl_632 , and_dcpl_636 , and_903_cse , and_907_cse , and_910_cse , and_914_cse
      , and_918_cse , and_920_cse});
  assign COMP_LOOP_COMP_LOOP_and_1890_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[0]) &
      COMP_LOOP_nor_281_itm;
  assign COMP_LOOP_COMP_LOOP_and_1891_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[0]) &
      COMP_LOOP_nor_505_itm;
  assign COMP_LOOP_COMP_LOOP_and_1892_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[0]) &
      COMP_LOOP_nor_729_itm;
  assign COMP_LOOP_COMP_LOOP_and_1893_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[0]) &
      COMP_LOOP_nor_953_itm;
  assign COMP_LOOP_COMP_LOOP_and_1894_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[0]) &
      COMP_LOOP_nor_1177_itm;
  assign COMP_LOOP_COMP_LOOP_and_1895_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[0]) &
      COMP_LOOP_nor_1401_itm;
  assign COMP_LOOP_COMP_LOOP_and_1896_nl = (COMP_LOOP_acc_10_cse_10_1_sva[0]) & COMP_LOOP_nor_1625_itm;
  assign COMP_LOOP_mux1h_1268_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_1518_itm,
      COMP_LOOP_COMP_LOOP_and_1890_nl, COMP_LOOP_COMP_LOOP_and_1891_nl, COMP_LOOP_COMP_LOOP_and_1892_nl,
      COMP_LOOP_COMP_LOOP_and_1893_nl, COMP_LOOP_COMP_LOOP_and_1894_nl, COMP_LOOP_COMP_LOOP_and_1895_nl,
      COMP_LOOP_COMP_LOOP_and_1896_nl, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_COMP_LOOP_and_1897_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[1]) &
      COMP_LOOP_nor_282_itm;
  assign COMP_LOOP_COMP_LOOP_and_1898_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[1]) &
      COMP_LOOP_nor_506_itm;
  assign COMP_LOOP_COMP_LOOP_and_1899_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[1]) &
      COMP_LOOP_nor_730_itm;
  assign COMP_LOOP_COMP_LOOP_and_1900_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[1]) &
      COMP_LOOP_nor_954_itm;
  assign COMP_LOOP_COMP_LOOP_and_1901_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[1]) &
      COMP_LOOP_nor_1178_itm;
  assign COMP_LOOP_COMP_LOOP_and_1902_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[1]) &
      COMP_LOOP_nor_1402_itm;
  assign COMP_LOOP_COMP_LOOP_and_1903_nl = (COMP_LOOP_acc_10_cse_10_1_sva[1]) & COMP_LOOP_nor_1626_itm;
  assign COMP_LOOP_mux1h_1269_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_760_itm,
      COMP_LOOP_COMP_LOOP_and_1897_nl, COMP_LOOP_COMP_LOOP_and_1898_nl, COMP_LOOP_COMP_LOOP_and_1899_nl,
      COMP_LOOP_COMP_LOOP_and_1900_nl, COMP_LOOP_COMP_LOOP_and_1901_nl, COMP_LOOP_COMP_LOOP_and_1902_nl,
      COMP_LOOP_COMP_LOOP_and_1903_nl, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1270_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_761_itm,
      COMP_LOOP_COMP_LOOP_and_1594_itm, COMP_LOOP_COMP_LOOP_and_569_itm, COMP_LOOP_COMP_LOOP_and_821_itm,
      COMP_LOOP_COMP_LOOP_and_100_itm, COMP_LOOP_COMP_LOOP_and_1325_itm, COMP_LOOP_COMP_LOOP_and_1577_itm,
      COMP_LOOP_COMP_LOOP_and_1829_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_COMP_LOOP_and_1904_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[2]) &
      COMP_LOOP_nor_284_itm;
  assign COMP_LOOP_COMP_LOOP_and_1905_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[2]) &
      COMP_LOOP_nor_508_itm;
  assign COMP_LOOP_COMP_LOOP_and_1906_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[2]) &
      COMP_LOOP_nor_732_itm;
  assign COMP_LOOP_COMP_LOOP_and_1907_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[2]) &
      COMP_LOOP_nor_956_itm;
  assign COMP_LOOP_COMP_LOOP_and_1908_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[2]) &
      COMP_LOOP_nor_1180_itm;
  assign COMP_LOOP_COMP_LOOP_and_1909_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[2]) &
      COMP_LOOP_nor_1404_itm;
  assign COMP_LOOP_COMP_LOOP_and_1910_nl = (COMP_LOOP_acc_10_cse_10_1_sva[2]) & COMP_LOOP_nor_1628_itm;
  assign COMP_LOOP_mux1h_1271_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_509_itm,
      COMP_LOOP_COMP_LOOP_and_1904_nl, COMP_LOOP_COMP_LOOP_and_1905_nl, COMP_LOOP_COMP_LOOP_and_1906_nl,
      COMP_LOOP_COMP_LOOP_and_1907_nl, COMP_LOOP_COMP_LOOP_and_1908_nl, COMP_LOOP_COMP_LOOP_and_1909_nl,
      COMP_LOOP_COMP_LOOP_and_1910_nl, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1272_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_510_itm,
      COMP_LOOP_COMP_LOOP_and_1598_itm, COMP_LOOP_COMP_LOOP_and_571_itm, COMP_LOOP_COMP_LOOP_and_823_itm,
      COMP_LOOP_COMP_LOOP_and_101_itm, COMP_LOOP_COMP_LOOP_and_1327_itm, COMP_LOOP_COMP_LOOP_and_1579_itm,
      COMP_LOOP_COMP_LOOP_and_1831_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1273_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_258_itm,
      COMP_LOOP_COMP_LOOP_and_1607_itm, COMP_LOOP_COMP_LOOP_and_572_itm, COMP_LOOP_COMP_LOOP_and_73_itm,
      COMP_LOOP_COMP_LOOP_and_102_itm, COMP_LOOP_COMP_LOOP_and_115_itm, COMP_LOOP_COMP_LOOP_and_1580_itm,
      COMP_LOOP_COMP_LOOP_and_1832_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1274_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_6_itm,
      COMP_LOOP_COMP_LOOP_and_1610_itm, COMP_LOOP_COMP_LOOP_and_573_itm, COMP_LOOP_COMP_LOOP_and_825_itm,
      COMP_LOOP_COMP_LOOP_and_1077_itm, COMP_LOOP_COMP_LOOP_and_1329_itm, COMP_LOOP_COMP_LOOP_and_1581_itm,
      COMP_LOOP_COMP_LOOP_and_1833_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_COMP_LOOP_and_1911_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[3]) &
      COMP_LOOP_nor_288_itm;
  assign COMP_LOOP_COMP_LOOP_and_1912_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[3]) &
      COMP_LOOP_nor_512_itm;
  assign COMP_LOOP_COMP_LOOP_and_1913_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[3]) &
      COMP_LOOP_nor_736_itm;
  assign COMP_LOOP_COMP_LOOP_and_1914_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[3]) &
      COMP_LOOP_nor_960_itm;
  assign COMP_LOOP_COMP_LOOP_and_1915_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[3]) &
      COMP_LOOP_nor_1184_itm;
  assign COMP_LOOP_COMP_LOOP_and_1916_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[3]) &
      COMP_LOOP_nor_1408_itm;
  assign COMP_LOOP_COMP_LOOP_and_1917_nl = (COMP_LOOP_acc_10_cse_10_1_sva[3]) & COMP_LOOP_nor_1632_itm;
  assign COMP_LOOP_mux1h_1275_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_260_itm,
      COMP_LOOP_COMP_LOOP_and_1911_nl, COMP_LOOP_COMP_LOOP_and_1912_nl, COMP_LOOP_COMP_LOOP_and_1913_nl,
      COMP_LOOP_COMP_LOOP_and_1914_nl, COMP_LOOP_COMP_LOOP_and_1915_nl, COMP_LOOP_COMP_LOOP_and_1916_nl,
      COMP_LOOP_COMP_LOOP_and_1917_nl, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1276_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_261_itm,
      COMP_LOOP_COMP_LOOP_and_100_itm, COMP_LOOP_COMP_LOOP_and_575_itm, COMP_LOOP_COMP_LOOP_and_827_itm,
      COMP_LOOP_COMP_LOOP_and_103_itm, COMP_LOOP_COMP_LOOP_and_116_itm, COMP_LOOP_COMP_LOOP_and_1583_itm,
      COMP_LOOP_COMP_LOOP_and_1835_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1277_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_262_itm,
      COMP_LOOP_COMP_LOOP_and_1614_itm, COMP_LOOP_COMP_LOOP_and_576_itm, COMP_LOOP_COMP_LOOP_and_828_itm,
      COMP_LOOP_COMP_LOOP_and_104_itm, COMP_LOOP_COMP_LOOP_and_117_itm, COMP_LOOP_COMP_LOOP_and_1584_itm,
      COMP_LOOP_COMP_LOOP_and_1836_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1278_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_10_itm,
      COMP_LOOP_COMP_LOOP_and_1622_itm, COMP_LOOP_COMP_LOOP_and_577_itm, COMP_LOOP_COMP_LOOP_and_829_itm,
      COMP_LOOP_COMP_LOOP_and_1081_itm, COMP_LOOP_COMP_LOOP_and_1333_itm, COMP_LOOP_COMP_LOOP_and_1585_itm,
      COMP_LOOP_COMP_LOOP_and_1837_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1279_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_264_itm,
      COMP_LOOP_COMP_LOOP_and_1832_itm, COMP_LOOP_COMP_LOOP_and_578_itm, COMP_LOOP_COMP_LOOP_and_830_itm,
      COMP_LOOP_COMP_LOOP_and_105_itm, COMP_LOOP_COMP_LOOP_and_118_itm, COMP_LOOP_COMP_LOOP_and_1586_itm,
      COMP_LOOP_COMP_LOOP_and_1838_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1280_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_12_itm,
      COMP_LOOP_COMP_LOOP_and_1835_itm, COMP_LOOP_COMP_LOOP_and_579_itm, COMP_LOOP_COMP_LOOP_and_831_itm,
      COMP_LOOP_COMP_LOOP_and_1083_itm, COMP_LOOP_COMP_LOOP_and_1335_itm, COMP_LOOP_COMP_LOOP_and_1587_itm,
      COMP_LOOP_COMP_LOOP_and_1839_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1281_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_13_itm,
      COMP_LOOP_COMP_LOOP_and_1844_itm, COMP_LOOP_COMP_LOOP_and_580_itm, COMP_LOOP_COMP_LOOP_and_832_itm,
      COMP_LOOP_COMP_LOOP_and_1084_itm, COMP_LOOP_COMP_LOOP_and_1336_itm, COMP_LOOP_COMP_LOOP_and_1588_itm,
      COMP_LOOP_COMP_LOOP_and_1840_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1282_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_14_itm,
      COMP_LOOP_COMP_LOOP_and_1850_itm, COMP_LOOP_COMP_LOOP_and_581_itm, COMP_LOOP_COMP_LOOP_and_833_itm,
      COMP_LOOP_COMP_LOOP_and_1085_itm, COMP_LOOP_COMP_LOOP_and_1337_itm, COMP_LOOP_COMP_LOOP_and_1589_itm,
      COMP_LOOP_COMP_LOOP_and_1841_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_COMP_LOOP_and_1918_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[4]) &
      COMP_LOOP_nor_296_itm;
  assign COMP_LOOP_COMP_LOOP_and_1919_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[4]) &
      COMP_LOOP_nor_520_itm;
  assign COMP_LOOP_COMP_LOOP_and_1920_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[4]) &
      COMP_LOOP_nor_744_itm;
  assign COMP_LOOP_COMP_LOOP_and_1921_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[4]) &
      COMP_LOOP_nor_968_itm;
  assign COMP_LOOP_COMP_LOOP_and_1922_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[4]) &
      COMP_LOOP_nor_1192_itm;
  assign COMP_LOOP_COMP_LOOP_and_1923_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[4]) &
      COMP_LOOP_nor_1416_itm;
  assign COMP_LOOP_COMP_LOOP_and_1924_nl = (COMP_LOOP_acc_10_cse_10_1_sva[4]) & COMP_LOOP_nor_1640_itm;
  assign COMP_LOOP_mux1h_1283_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_268_itm,
      COMP_LOOP_COMP_LOOP_and_1918_nl, COMP_LOOP_COMP_LOOP_and_1919_nl, COMP_LOOP_COMP_LOOP_and_1920_nl,
      COMP_LOOP_COMP_LOOP_and_1921_nl, COMP_LOOP_COMP_LOOP_and_1922_nl, COMP_LOOP_COMP_LOOP_and_1923_nl,
      COMP_LOOP_COMP_LOOP_and_1924_nl, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1284_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_522_itm,
      COMP_LOOP_COMP_LOOP_and_1862_itm, COMP_LOOP_COMP_LOOP_and_583_itm, COMP_LOOP_COMP_LOOP_and_835_itm,
      COMP_LOOP_COMP_LOOP_and_106_itm, COMP_LOOP_COMP_LOOP_and_119_itm, COMP_LOOP_COMP_LOOP_and_1591_itm,
      COMP_LOOP_COMP_LOOP_and_1843_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1285_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_270_itm,
      COMP_LOOP_COMP_LOOP_and_1866_itm, COMP_LOOP_COMP_LOOP_and_584_itm, COMP_LOOP_COMP_LOOP_and_836_itm,
      COMP_LOOP_COMP_LOOP_and_107_itm, COMP_LOOP_COMP_LOOP_and_120_itm, COMP_LOOP_COMP_LOOP_and_1592_itm,
      COMP_LOOP_COMP_LOOP_and_1844_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1286_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_18_itm,
      COMP_LOOP_COMP_LOOP_and_333_itm, COMP_LOOP_COMP_LOOP_and_585_itm, COMP_LOOP_COMP_LOOP_and_837_itm,
      COMP_LOOP_COMP_LOOP_and_1089_itm, COMP_LOOP_COMP_LOOP_and_1341_itm, COMP_LOOP_COMP_LOOP_and_1593_itm,
      COMP_LOOP_COMP_LOOP_and_1845_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1287_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_272_itm,
      COMP_LOOP_COMP_LOOP_and_334_itm, COMP_LOOP_COMP_LOOP_and_586_itm, COMP_LOOP_COMP_LOOP_and_838_itm,
      COMP_LOOP_COMP_LOOP_and_108_itm, COMP_LOOP_COMP_LOOP_and_121_itm, COMP_LOOP_COMP_LOOP_and_1594_itm,
      COMP_LOOP_COMP_LOOP_and_1846_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1288_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_20_itm,
      COMP_LOOP_COMP_LOOP_and_335_itm, COMP_LOOP_COMP_LOOP_and_587_itm, COMP_LOOP_COMP_LOOP_and_839_itm,
      COMP_LOOP_COMP_LOOP_and_1091_itm, COMP_LOOP_COMP_LOOP_and_1343_itm, COMP_LOOP_COMP_LOOP_and_1595_itm,
      COMP_LOOP_COMP_LOOP_and_1847_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1289_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_21_itm,
      COMP_LOOP_COMP_LOOP_and_336_itm, COMP_LOOP_COMP_LOOP_and_588_itm, COMP_LOOP_COMP_LOOP_and_840_itm,
      COMP_LOOP_COMP_LOOP_and_1092_itm, COMP_LOOP_COMP_LOOP_and_1344_itm, COMP_LOOP_COMP_LOOP_and_1596_itm,
      COMP_LOOP_COMP_LOOP_and_1848_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1290_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_22_itm,
      COMP_LOOP_COMP_LOOP_and_337_itm, COMP_LOOP_COMP_LOOP_and_589_itm, COMP_LOOP_COMP_LOOP_and_841_itm,
      COMP_LOOP_COMP_LOOP_and_1093_itm, COMP_LOOP_COMP_LOOP_and_1345_itm, COMP_LOOP_COMP_LOOP_and_1597_itm,
      COMP_LOOP_COMP_LOOP_and_1849_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1291_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_23_itm,
      COMP_LOOP_COMP_LOOP_and_338_itm, COMP_LOOP_COMP_LOOP_and_590_itm, COMP_LOOP_COMP_LOOP_and_842_itm,
      COMP_LOOP_COMP_LOOP_and_109_itm, COMP_LOOP_COMP_LOOP_and_1346_itm, COMP_LOOP_COMP_LOOP_and_1598_itm,
      COMP_LOOP_COMP_LOOP_and_1850_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1292_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_24_itm,
      COMP_LOOP_COMP_LOOP_and_339_itm, COMP_LOOP_COMP_LOOP_and_591_itm, COMP_LOOP_COMP_LOOP_and_843_itm,
      COMP_LOOP_COMP_LOOP_and_1095_itm, COMP_LOOP_COMP_LOOP_and_1347_itm, COMP_LOOP_COMP_LOOP_and_1599_itm,
      COMP_LOOP_COMP_LOOP_and_1851_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1293_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_25_itm,
      COMP_LOOP_COMP_LOOP_and_340_itm, COMP_LOOP_COMP_LOOP_and_592_itm, COMP_LOOP_COMP_LOOP_and_844_itm,
      COMP_LOOP_COMP_LOOP_and_1096_itm, COMP_LOOP_COMP_LOOP_and_1348_itm, COMP_LOOP_COMP_LOOP_and_1600_itm,
      COMP_LOOP_COMP_LOOP_and_1852_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1294_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_26_itm,
      COMP_LOOP_COMP_LOOP_and_341_itm, COMP_LOOP_COMP_LOOP_and_593_itm, COMP_LOOP_COMP_LOOP_and_845_itm,
      COMP_LOOP_COMP_LOOP_and_1097_itm, COMP_LOOP_COMP_LOOP_and_1349_itm, COMP_LOOP_COMP_LOOP_and_1601_itm,
      COMP_LOOP_COMP_LOOP_and_1853_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1295_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_27_itm,
      COMP_LOOP_COMP_LOOP_and_342_itm, COMP_LOOP_COMP_LOOP_and_594_itm, COMP_LOOP_COMP_LOOP_and_846_itm,
      COMP_LOOP_COMP_LOOP_and_1098_itm, COMP_LOOP_COMP_LOOP_and_1350_itm, COMP_LOOP_COMP_LOOP_and_1602_itm,
      COMP_LOOP_COMP_LOOP_and_1854_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1296_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_28_itm,
      COMP_LOOP_COMP_LOOP_and_343_itm, COMP_LOOP_COMP_LOOP_and_595_itm, COMP_LOOP_COMP_LOOP_and_847_itm,
      COMP_LOOP_COMP_LOOP_and_1099_itm, COMP_LOOP_COMP_LOOP_and_1351_itm, COMP_LOOP_COMP_LOOP_and_1603_itm,
      COMP_LOOP_COMP_LOOP_and_1855_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1297_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_29_itm,
      COMP_LOOP_COMP_LOOP_and_344_itm, COMP_LOOP_COMP_LOOP_and_596_itm, COMP_LOOP_COMP_LOOP_and_848_itm,
      COMP_LOOP_COMP_LOOP_and_1100_itm, COMP_LOOP_COMP_LOOP_and_1352_itm, COMP_LOOP_COMP_LOOP_and_1604_itm,
      COMP_LOOP_COMP_LOOP_and_1856_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1298_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_30_itm,
      COMP_LOOP_COMP_LOOP_and_345_itm, COMP_LOOP_COMP_LOOP_and_597_itm, COMP_LOOP_COMP_LOOP_and_849_itm,
      COMP_LOOP_COMP_LOOP_and_1101_itm, COMP_LOOP_COMP_LOOP_and_1353_itm, COMP_LOOP_COMP_LOOP_and_1605_itm,
      COMP_LOOP_COMP_LOOP_and_1857_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_COMP_LOOP_and_1925_nl = (COMP_LOOP_acc_10_cse_10_1_2_sva[5]) &
      COMP_LOOP_nor_311_itm;
  assign COMP_LOOP_COMP_LOOP_and_1926_nl = (COMP_LOOP_acc_10_cse_10_1_3_sva[5]) &
      COMP_LOOP_nor_535_itm;
  assign COMP_LOOP_COMP_LOOP_and_1927_nl = (COMP_LOOP_acc_10_cse_10_1_4_sva[5]) &
      COMP_LOOP_nor_759_itm;
  assign COMP_LOOP_COMP_LOOP_and_1928_nl = (COMP_LOOP_acc_10_cse_10_1_5_sva[5]) &
      COMP_LOOP_nor_983_itm;
  assign COMP_LOOP_COMP_LOOP_and_1929_nl = (COMP_LOOP_acc_10_cse_10_1_6_sva[5]) &
      COMP_LOOP_nor_1207_itm;
  assign COMP_LOOP_COMP_LOOP_and_1930_nl = (COMP_LOOP_acc_10_cse_10_1_7_sva[5]) &
      COMP_LOOP_nor_1431_itm;
  assign COMP_LOOP_COMP_LOOP_and_1931_nl = (COMP_LOOP_acc_10_cse_10_1_sva[5]) & COMP_LOOP_nor_1655_itm;
  assign COMP_LOOP_mux1h_1299_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_284_itm,
      COMP_LOOP_COMP_LOOP_and_1925_nl, COMP_LOOP_COMP_LOOP_and_1926_nl, COMP_LOOP_COMP_LOOP_and_1927_nl,
      COMP_LOOP_COMP_LOOP_and_1928_nl, COMP_LOOP_COMP_LOOP_and_1929_nl, COMP_LOOP_COMP_LOOP_and_1930_nl,
      COMP_LOOP_COMP_LOOP_and_1931_nl, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1300_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_285_itm,
      COMP_LOOP_COMP_LOOP_and_347_itm, COMP_LOOP_COMP_LOOP_and_599_itm, COMP_LOOP_COMP_LOOP_and_74_itm,
      COMP_LOOP_COMP_LOOP_and_110_itm, COMP_LOOP_COMP_LOOP_and_122_itm, COMP_LOOP_COMP_LOOP_and_1607_itm,
      COMP_LOOP_COMP_LOOP_and_1859_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1301_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_286_itm,
      COMP_LOOP_COMP_LOOP_and_101_itm, COMP_LOOP_COMP_LOOP_and_600_itm, COMP_LOOP_COMP_LOOP_and_852_itm,
      COMP_LOOP_COMP_LOOP_and_1104_itm, COMP_LOOP_COMP_LOOP_and_123_itm, COMP_LOOP_COMP_LOOP_and_1608_itm,
      COMP_LOOP_COMP_LOOP_and_1860_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1302_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_34_itm,
      COMP_LOOP_COMP_LOOP_and_349_itm, COMP_LOOP_COMP_LOOP_and_601_itm, COMP_LOOP_COMP_LOOP_and_853_itm,
      COMP_LOOP_COMP_LOOP_and_1105_itm, COMP_LOOP_COMP_LOOP_and_1357_itm, COMP_LOOP_COMP_LOOP_and_1609_itm,
      COMP_LOOP_COMP_LOOP_and_1861_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1303_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_288_itm,
      COMP_LOOP_COMP_LOOP_and_103_itm, COMP_LOOP_COMP_LOOP_and_602_itm, COMP_LOOP_COMP_LOOP_and_854_itm,
      COMP_LOOP_COMP_LOOP_and_1106_itm, COMP_LOOP_COMP_LOOP_and_124_itm, COMP_LOOP_COMP_LOOP_and_1610_itm,
      COMP_LOOP_COMP_LOOP_and_1862_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1304_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_36_itm,
      COMP_LOOP_COMP_LOOP_and_351_itm, COMP_LOOP_COMP_LOOP_and_603_itm, COMP_LOOP_COMP_LOOP_and_855_itm,
      COMP_LOOP_COMP_LOOP_and_1107_itm, COMP_LOOP_COMP_LOOP_and_1359_itm, COMP_LOOP_COMP_LOOP_and_1611_itm,
      COMP_LOOP_COMP_LOOP_and_1863_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1305_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_37_itm,
      COMP_LOOP_COMP_LOOP_and_352_itm, COMP_LOOP_COMP_LOOP_and_604_itm, COMP_LOOP_COMP_LOOP_and_856_itm,
      COMP_LOOP_COMP_LOOP_and_1108_itm, COMP_LOOP_COMP_LOOP_and_1360_itm, COMP_LOOP_COMP_LOOP_and_1612_itm,
      COMP_LOOP_COMP_LOOP_and_1864_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1306_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_38_itm,
      COMP_LOOP_COMP_LOOP_and_353_itm, COMP_LOOP_COMP_LOOP_and_605_itm, COMP_LOOP_COMP_LOOP_and_857_itm,
      COMP_LOOP_COMP_LOOP_and_1109_itm, COMP_LOOP_COMP_LOOP_and_1361_itm, COMP_LOOP_COMP_LOOP_and_1613_itm,
      COMP_LOOP_COMP_LOOP_and_1865_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1307_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_39_itm,
      COMP_LOOP_COMP_LOOP_and_104_itm, COMP_LOOP_COMP_LOOP_and_606_itm, COMP_LOOP_COMP_LOOP_and_75_itm,
      COMP_LOOP_COMP_LOOP_and_1110_itm, COMP_LOOP_COMP_LOOP_and_125_itm, COMP_LOOP_COMP_LOOP_and_1614_itm,
      COMP_LOOP_COMP_LOOP_and_1866_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1308_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_40_itm,
      COMP_LOOP_COMP_LOOP_and_355_itm, COMP_LOOP_COMP_LOOP_and_607_itm, COMP_LOOP_COMP_LOOP_and_859_itm,
      COMP_LOOP_COMP_LOOP_and_1111_itm, COMP_LOOP_COMP_LOOP_and_1363_itm, COMP_LOOP_COMP_LOOP_and_1615_itm,
      COMP_LOOP_COMP_LOOP_and_1867_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1309_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_41_itm,
      COMP_LOOP_COMP_LOOP_and_356_itm, COMP_LOOP_COMP_LOOP_and_608_itm, COMP_LOOP_COMP_LOOP_and_860_itm,
      COMP_LOOP_COMP_LOOP_and_1112_itm, COMP_LOOP_COMP_LOOP_and_1364_itm, COMP_LOOP_COMP_LOOP_and_1616_itm,
      COMP_LOOP_COMP_LOOP_and_1868_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1310_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_42_itm,
      COMP_LOOP_COMP_LOOP_and_357_itm, COMP_LOOP_COMP_LOOP_and_609_itm, COMP_LOOP_COMP_LOOP_and_861_itm,
      COMP_LOOP_COMP_LOOP_and_1113_itm, COMP_LOOP_COMP_LOOP_and_1365_itm, COMP_LOOP_COMP_LOOP_and_1617_itm,
      COMP_LOOP_COMP_LOOP_and_1869_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1311_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_43_itm,
      COMP_LOOP_COMP_LOOP_and_358_itm, COMP_LOOP_COMP_LOOP_and_610_itm, COMP_LOOP_COMP_LOOP_and_862_itm,
      COMP_LOOP_COMP_LOOP_and_1114_itm, COMP_LOOP_COMP_LOOP_and_1366_itm, COMP_LOOP_COMP_LOOP_and_1618_itm,
      COMP_LOOP_COMP_LOOP_and_1870_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1312_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_44_itm,
      COMP_LOOP_COMP_LOOP_and_359_itm, COMP_LOOP_COMP_LOOP_and_611_itm, COMP_LOOP_COMP_LOOP_and_863_itm,
      COMP_LOOP_COMP_LOOP_and_1115_itm, COMP_LOOP_COMP_LOOP_and_1367_itm, COMP_LOOP_COMP_LOOP_and_1619_itm,
      COMP_LOOP_COMP_LOOP_and_1871_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1313_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_45_itm,
      COMP_LOOP_COMP_LOOP_and_360_itm, COMP_LOOP_COMP_LOOP_and_612_itm, COMP_LOOP_COMP_LOOP_and_864_itm,
      COMP_LOOP_COMP_LOOP_and_1116_itm, COMP_LOOP_COMP_LOOP_and_1368_itm, COMP_LOOP_COMP_LOOP_and_1620_itm,
      COMP_LOOP_COMP_LOOP_and_1872_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1314_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_46_itm,
      COMP_LOOP_COMP_LOOP_and_361_itm, COMP_LOOP_COMP_LOOP_and_613_itm, COMP_LOOP_COMP_LOOP_and_865_itm,
      COMP_LOOP_COMP_LOOP_and_1117_itm, COMP_LOOP_COMP_LOOP_and_1369_itm, COMP_LOOP_COMP_LOOP_and_1621_itm,
      COMP_LOOP_COMP_LOOP_and_1873_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1315_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_47_itm,
      COMP_LOOP_COMP_LOOP_and_105_itm, COMP_LOOP_COMP_LOOP_and_614_itm, COMP_LOOP_COMP_LOOP_and_866_itm,
      COMP_LOOP_COMP_LOOP_and_1118_itm, COMP_LOOP_COMP_LOOP_and_1370_itm, COMP_LOOP_COMP_LOOP_and_1622_itm,
      COMP_LOOP_COMP_LOOP_and_1874_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1316_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_48_itm,
      COMP_LOOP_COMP_LOOP_and_363_itm, COMP_LOOP_COMP_LOOP_and_615_itm, COMP_LOOP_COMP_LOOP_and_867_itm,
      COMP_LOOP_COMP_LOOP_and_1119_itm, COMP_LOOP_COMP_LOOP_and_1371_itm, COMP_LOOP_COMP_LOOP_and_1623_itm,
      COMP_LOOP_COMP_LOOP_and_1875_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1317_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_49_itm,
      COMP_LOOP_COMP_LOOP_and_364_itm, COMP_LOOP_COMP_LOOP_and_616_itm, COMP_LOOP_COMP_LOOP_and_868_itm,
      COMP_LOOP_COMP_LOOP_and_1120_itm, COMP_LOOP_COMP_LOOP_and_1372_itm, COMP_LOOP_COMP_LOOP_and_1624_itm,
      COMP_LOOP_COMP_LOOP_and_1876_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1318_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_50_itm,
      COMP_LOOP_COMP_LOOP_and_365_itm, COMP_LOOP_COMP_LOOP_and_617_itm, COMP_LOOP_COMP_LOOP_and_869_itm,
      COMP_LOOP_COMP_LOOP_and_1121_itm, COMP_LOOP_COMP_LOOP_and_1373_itm, COMP_LOOP_COMP_LOOP_and_1625_itm,
      COMP_LOOP_COMP_LOOP_and_1877_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1319_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_51_itm,
      COMP_LOOP_COMP_LOOP_and_366_itm, COMP_LOOP_COMP_LOOP_and_618_itm, COMP_LOOP_COMP_LOOP_and_870_itm,
      COMP_LOOP_COMP_LOOP_and_1122_itm, COMP_LOOP_COMP_LOOP_and_1374_itm, COMP_LOOP_COMP_LOOP_and_1626_itm,
      COMP_LOOP_COMP_LOOP_and_1878_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1320_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_52_itm,
      COMP_LOOP_COMP_LOOP_and_367_itm, COMP_LOOP_COMP_LOOP_and_619_itm, COMP_LOOP_COMP_LOOP_and_871_itm,
      COMP_LOOP_COMP_LOOP_and_1123_itm, COMP_LOOP_COMP_LOOP_and_1375_itm, COMP_LOOP_COMP_LOOP_and_1627_itm,
      COMP_LOOP_COMP_LOOP_and_1879_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1321_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_53_itm,
      COMP_LOOP_COMP_LOOP_and_368_itm, COMP_LOOP_COMP_LOOP_and_620_itm, COMP_LOOP_COMP_LOOP_and_872_itm,
      COMP_LOOP_COMP_LOOP_and_1124_itm, COMP_LOOP_COMP_LOOP_and_1376_itm, COMP_LOOP_COMP_LOOP_and_1628_itm,
      COMP_LOOP_COMP_LOOP_and_1880_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1322_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_54_itm,
      COMP_LOOP_COMP_LOOP_and_369_itm, COMP_LOOP_COMP_LOOP_and_621_itm, COMP_LOOP_COMP_LOOP_and_873_itm,
      COMP_LOOP_COMP_LOOP_and_1125_itm, COMP_LOOP_COMP_LOOP_and_1377_itm, COMP_LOOP_COMP_LOOP_and_1629_itm,
      COMP_LOOP_COMP_LOOP_and_1881_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1323_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_55_itm,
      COMP_LOOP_COMP_LOOP_and_370_itm, COMP_LOOP_COMP_LOOP_and_622_itm, COMP_LOOP_COMP_LOOP_and_874_itm,
      COMP_LOOP_COMP_LOOP_and_1126_itm, COMP_LOOP_COMP_LOOP_and_1378_itm, COMP_LOOP_COMP_LOOP_and_1630_itm,
      COMP_LOOP_COMP_LOOP_and_1882_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1324_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_56_itm,
      COMP_LOOP_COMP_LOOP_and_371_itm, COMP_LOOP_COMP_LOOP_and_623_itm, COMP_LOOP_COMP_LOOP_and_875_itm,
      COMP_LOOP_COMP_LOOP_and_1127_itm, COMP_LOOP_COMP_LOOP_and_1379_itm, COMP_LOOP_COMP_LOOP_and_1631_itm,
      COMP_LOOP_COMP_LOOP_and_1883_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1325_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_57_itm,
      COMP_LOOP_COMP_LOOP_and_372_itm, COMP_LOOP_COMP_LOOP_and_624_itm, COMP_LOOP_COMP_LOOP_and_876_itm,
      COMP_LOOP_COMP_LOOP_and_1128_itm, COMP_LOOP_COMP_LOOP_and_1380_itm, COMP_LOOP_COMP_LOOP_and_1632_itm,
      COMP_LOOP_COMP_LOOP_and_1884_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1326_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_58_itm,
      COMP_LOOP_COMP_LOOP_and_373_itm, COMP_LOOP_COMP_LOOP_and_625_itm, COMP_LOOP_COMP_LOOP_and_877_itm,
      COMP_LOOP_COMP_LOOP_and_1129_itm, COMP_LOOP_COMP_LOOP_and_1381_itm, COMP_LOOP_COMP_LOOP_and_1633_itm,
      COMP_LOOP_COMP_LOOP_and_1885_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1327_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_59_itm,
      COMP_LOOP_COMP_LOOP_and_374_itm, COMP_LOOP_COMP_LOOP_and_626_itm, COMP_LOOP_COMP_LOOP_and_878_itm,
      COMP_LOOP_COMP_LOOP_and_1130_itm, COMP_LOOP_COMP_LOOP_and_1382_itm, COMP_LOOP_COMP_LOOP_and_1634_itm,
      COMP_LOOP_COMP_LOOP_and_1886_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1328_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_60_itm,
      COMP_LOOP_COMP_LOOP_and_375_itm, COMP_LOOP_COMP_LOOP_and_627_itm, COMP_LOOP_COMP_LOOP_and_879_itm,
      COMP_LOOP_COMP_LOOP_and_1131_itm, COMP_LOOP_COMP_LOOP_and_1383_itm, COMP_LOOP_COMP_LOOP_and_1635_itm,
      COMP_LOOP_COMP_LOOP_and_1887_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1329_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_61_itm,
      COMP_LOOP_COMP_LOOP_and_376_itm, COMP_LOOP_COMP_LOOP_and_628_itm, COMP_LOOP_COMP_LOOP_and_880_itm,
      COMP_LOOP_COMP_LOOP_and_1132_itm, COMP_LOOP_COMP_LOOP_and_1384_itm, COMP_LOOP_COMP_LOOP_and_1636_itm,
      COMP_LOOP_COMP_LOOP_and_1888_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign COMP_LOOP_mux1h_1330_nl = MUX1HOT_s_1_8_2(COMP_LOOP_COMP_LOOP_and_62_itm,
      COMP_LOOP_COMP_LOOP_and_377_itm, COMP_LOOP_COMP_LOOP_and_629_itm, COMP_LOOP_COMP_LOOP_and_881_itm,
      COMP_LOOP_COMP_LOOP_and_1133_itm, COMP_LOOP_COMP_LOOP_and_1385_itm, COMP_LOOP_COMP_LOOP_and_1637_itm,
      COMP_LOOP_COMP_LOOP_and_1889_itm, {and_dcpl_632 , and_dcpl_636 , and_903_cse
      , and_907_cse , and_910_cse , and_914_cse , and_918_cse , and_920_cse});
  assign z_out_9 = MUX1HOT_v_64_64_2(vec_rsc_0_0_i_q_d, vec_rsc_0_1_i_q_d, vec_rsc_0_2_i_q_d,
      vec_rsc_0_3_i_q_d, vec_rsc_0_4_i_q_d, vec_rsc_0_5_i_q_d, vec_rsc_0_6_i_q_d,
      vec_rsc_0_7_i_q_d, vec_rsc_0_8_i_q_d, vec_rsc_0_9_i_q_d, vec_rsc_0_10_i_q_d,
      vec_rsc_0_11_i_q_d, vec_rsc_0_12_i_q_d, vec_rsc_0_13_i_q_d, vec_rsc_0_14_i_q_d,
      vec_rsc_0_15_i_q_d, vec_rsc_0_16_i_q_d, vec_rsc_0_17_i_q_d, vec_rsc_0_18_i_q_d,
      vec_rsc_0_19_i_q_d, vec_rsc_0_20_i_q_d, vec_rsc_0_21_i_q_d, vec_rsc_0_22_i_q_d,
      vec_rsc_0_23_i_q_d, vec_rsc_0_24_i_q_d, vec_rsc_0_25_i_q_d, vec_rsc_0_26_i_q_d,
      vec_rsc_0_27_i_q_d, vec_rsc_0_28_i_q_d, vec_rsc_0_29_i_q_d, vec_rsc_0_30_i_q_d,
      vec_rsc_0_31_i_q_d, vec_rsc_0_32_i_q_d, vec_rsc_0_33_i_q_d, vec_rsc_0_34_i_q_d,
      vec_rsc_0_35_i_q_d, vec_rsc_0_36_i_q_d, vec_rsc_0_37_i_q_d, vec_rsc_0_38_i_q_d,
      vec_rsc_0_39_i_q_d, vec_rsc_0_40_i_q_d, vec_rsc_0_41_i_q_d, vec_rsc_0_42_i_q_d,
      vec_rsc_0_43_i_q_d, vec_rsc_0_44_i_q_d, vec_rsc_0_45_i_q_d, vec_rsc_0_46_i_q_d,
      vec_rsc_0_47_i_q_d, vec_rsc_0_48_i_q_d, vec_rsc_0_49_i_q_d, vec_rsc_0_50_i_q_d,
      vec_rsc_0_51_i_q_d, vec_rsc_0_52_i_q_d, vec_rsc_0_53_i_q_d, vec_rsc_0_54_i_q_d,
      vec_rsc_0_55_i_q_d, vec_rsc_0_56_i_q_d, vec_rsc_0_57_i_q_d, vec_rsc_0_58_i_q_d,
      vec_rsc_0_59_i_q_d, vec_rsc_0_60_i_q_d, vec_rsc_0_61_i_q_d, vec_rsc_0_62_i_q_d,
      vec_rsc_0_63_i_q_d, {COMP_LOOP_mux1h_1267_nl , COMP_LOOP_mux1h_1268_nl , COMP_LOOP_mux1h_1269_nl
      , COMP_LOOP_mux1h_1270_nl , COMP_LOOP_mux1h_1271_nl , COMP_LOOP_mux1h_1272_nl
      , COMP_LOOP_mux1h_1273_nl , COMP_LOOP_mux1h_1274_nl , COMP_LOOP_mux1h_1275_nl
      , COMP_LOOP_mux1h_1276_nl , COMP_LOOP_mux1h_1277_nl , COMP_LOOP_mux1h_1278_nl
      , COMP_LOOP_mux1h_1279_nl , COMP_LOOP_mux1h_1280_nl , COMP_LOOP_mux1h_1281_nl
      , COMP_LOOP_mux1h_1282_nl , COMP_LOOP_mux1h_1283_nl , COMP_LOOP_mux1h_1284_nl
      , COMP_LOOP_mux1h_1285_nl , COMP_LOOP_mux1h_1286_nl , COMP_LOOP_mux1h_1287_nl
      , COMP_LOOP_mux1h_1288_nl , COMP_LOOP_mux1h_1289_nl , COMP_LOOP_mux1h_1290_nl
      , COMP_LOOP_mux1h_1291_nl , COMP_LOOP_mux1h_1292_nl , COMP_LOOP_mux1h_1293_nl
      , COMP_LOOP_mux1h_1294_nl , COMP_LOOP_mux1h_1295_nl , COMP_LOOP_mux1h_1296_nl
      , COMP_LOOP_mux1h_1297_nl , COMP_LOOP_mux1h_1298_nl , COMP_LOOP_mux1h_1299_nl
      , COMP_LOOP_mux1h_1300_nl , COMP_LOOP_mux1h_1301_nl , COMP_LOOP_mux1h_1302_nl
      , COMP_LOOP_mux1h_1303_nl , COMP_LOOP_mux1h_1304_nl , COMP_LOOP_mux1h_1305_nl
      , COMP_LOOP_mux1h_1306_nl , COMP_LOOP_mux1h_1307_nl , COMP_LOOP_mux1h_1308_nl
      , COMP_LOOP_mux1h_1309_nl , COMP_LOOP_mux1h_1310_nl , COMP_LOOP_mux1h_1311_nl
      , COMP_LOOP_mux1h_1312_nl , COMP_LOOP_mux1h_1313_nl , COMP_LOOP_mux1h_1314_nl
      , COMP_LOOP_mux1h_1315_nl , COMP_LOOP_mux1h_1316_nl , COMP_LOOP_mux1h_1317_nl
      , COMP_LOOP_mux1h_1318_nl , COMP_LOOP_mux1h_1319_nl , COMP_LOOP_mux1h_1320_nl
      , COMP_LOOP_mux1h_1321_nl , COMP_LOOP_mux1h_1322_nl , COMP_LOOP_mux1h_1323_nl
      , COMP_LOOP_mux1h_1324_nl , COMP_LOOP_mux1h_1325_nl , COMP_LOOP_mux1h_1326_nl
      , COMP_LOOP_mux1h_1327_nl , COMP_LOOP_mux1h_1328_nl , COMP_LOOP_mux1h_1329_nl
      , COMP_LOOP_mux1h_1330_nl});

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_5_2;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [4:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_8_2;
    input [0:0] input_7;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [7:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    result = result | ( input_7 & {1{sel[7]}});
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_16_2;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [15:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    result = result | ( input_7 & {4{sel[7]}});
    result = result | ( input_8 & {4{sel[8]}});
    result = result | ( input_9 & {4{sel[9]}});
    result = result | ( input_10 & {4{sel[10]}});
    result = result | ( input_11 & {4{sel[11]}});
    result = result | ( input_12 & {4{sel[12]}});
    result = result | ( input_13 & {4{sel[13]}});
    result = result | ( input_14 & {4{sel[14]}});
    result = result | ( input_15 & {4{sel[15]}});
    MUX1HOT_v_4_16_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_16_2;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [15:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    MUX1HOT_v_64_16_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_32_2;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [31:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    MUX1HOT_v_64_32_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_64_2;
    input [63:0] input_63;
    input [63:0] input_62;
    input [63:0] input_61;
    input [63:0] input_60;
    input [63:0] input_59;
    input [63:0] input_58;
    input [63:0] input_57;
    input [63:0] input_56;
    input [63:0] input_55;
    input [63:0] input_54;
    input [63:0] input_53;
    input [63:0] input_52;
    input [63:0] input_51;
    input [63:0] input_50;
    input [63:0] input_49;
    input [63:0] input_48;
    input [63:0] input_47;
    input [63:0] input_46;
    input [63:0] input_45;
    input [63:0] input_44;
    input [63:0] input_43;
    input [63:0] input_42;
    input [63:0] input_41;
    input [63:0] input_40;
    input [63:0] input_39;
    input [63:0] input_38;
    input [63:0] input_37;
    input [63:0] input_36;
    input [63:0] input_35;
    input [63:0] input_34;
    input [63:0] input_33;
    input [63:0] input_32;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [63:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    result = result | ( input_32 & {64{sel[32]}});
    result = result | ( input_33 & {64{sel[33]}});
    result = result | ( input_34 & {64{sel[34]}});
    result = result | ( input_35 & {64{sel[35]}});
    result = result | ( input_36 & {64{sel[36]}});
    result = result | ( input_37 & {64{sel[37]}});
    result = result | ( input_38 & {64{sel[38]}});
    result = result | ( input_39 & {64{sel[39]}});
    result = result | ( input_40 & {64{sel[40]}});
    result = result | ( input_41 & {64{sel[41]}});
    result = result | ( input_42 & {64{sel[42]}});
    result = result | ( input_43 & {64{sel[43]}});
    result = result | ( input_44 & {64{sel[44]}});
    result = result | ( input_45 & {64{sel[45]}});
    result = result | ( input_46 & {64{sel[46]}});
    result = result | ( input_47 & {64{sel[47]}});
    result = result | ( input_48 & {64{sel[48]}});
    result = result | ( input_49 & {64{sel[49]}});
    result = result | ( input_50 & {64{sel[50]}});
    result = result | ( input_51 & {64{sel[51]}});
    result = result | ( input_52 & {64{sel[52]}});
    result = result | ( input_53 & {64{sel[53]}});
    result = result | ( input_54 & {64{sel[54]}});
    result = result | ( input_55 & {64{sel[55]}});
    result = result | ( input_56 & {64{sel[56]}});
    result = result | ( input_57 & {64{sel[57]}});
    result = result | ( input_58 & {64{sel[58]}});
    result = result | ( input_59 & {64{sel[59]}});
    result = result | ( input_60 & {64{sel[60]}});
    result = result | ( input_61 & {64{sel[61]}});
    result = result | ( input_62 & {64{sel[62]}});
    result = result | ( input_63 & {64{sel[63]}});
    MUX1HOT_v_64_64_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_65_2;
    input [63:0] input_64;
    input [63:0] input_63;
    input [63:0] input_62;
    input [63:0] input_61;
    input [63:0] input_60;
    input [63:0] input_59;
    input [63:0] input_58;
    input [63:0] input_57;
    input [63:0] input_56;
    input [63:0] input_55;
    input [63:0] input_54;
    input [63:0] input_53;
    input [63:0] input_52;
    input [63:0] input_51;
    input [63:0] input_50;
    input [63:0] input_49;
    input [63:0] input_48;
    input [63:0] input_47;
    input [63:0] input_46;
    input [63:0] input_45;
    input [63:0] input_44;
    input [63:0] input_43;
    input [63:0] input_42;
    input [63:0] input_41;
    input [63:0] input_40;
    input [63:0] input_39;
    input [63:0] input_38;
    input [63:0] input_37;
    input [63:0] input_36;
    input [63:0] input_35;
    input [63:0] input_34;
    input [63:0] input_33;
    input [63:0] input_32;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [64:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    result = result | ( input_32 & {64{sel[32]}});
    result = result | ( input_33 & {64{sel[33]}});
    result = result | ( input_34 & {64{sel[34]}});
    result = result | ( input_35 & {64{sel[35]}});
    result = result | ( input_36 & {64{sel[36]}});
    result = result | ( input_37 & {64{sel[37]}});
    result = result | ( input_38 & {64{sel[38]}});
    result = result | ( input_39 & {64{sel[39]}});
    result = result | ( input_40 & {64{sel[40]}});
    result = result | ( input_41 & {64{sel[41]}});
    result = result | ( input_42 & {64{sel[42]}});
    result = result | ( input_43 & {64{sel[43]}});
    result = result | ( input_44 & {64{sel[44]}});
    result = result | ( input_45 & {64{sel[45]}});
    result = result | ( input_46 & {64{sel[46]}});
    result = result | ( input_47 & {64{sel[47]}});
    result = result | ( input_48 & {64{sel[48]}});
    result = result | ( input_49 & {64{sel[49]}});
    result = result | ( input_50 & {64{sel[50]}});
    result = result | ( input_51 & {64{sel[51]}});
    result = result | ( input_52 & {64{sel[52]}});
    result = result | ( input_53 & {64{sel[53]}});
    result = result | ( input_54 & {64{sel[54]}});
    result = result | ( input_55 & {64{sel[55]}});
    result = result | ( input_56 & {64{sel[56]}});
    result = result | ( input_57 & {64{sel[57]}});
    result = result | ( input_58 & {64{sel[58]}});
    result = result | ( input_59 & {64{sel[59]}});
    result = result | ( input_60 & {64{sel[60]}});
    result = result | ( input_61 & {64{sel[61]}});
    result = result | ( input_62 & {64{sel[62]}});
    result = result | ( input_63 & {64{sel[63]}});
    result = result | ( input_64 & {64{sel[64]}});
    MUX1HOT_v_64_65_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_68_2;
    input [63:0] input_67;
    input [63:0] input_66;
    input [63:0] input_65;
    input [63:0] input_64;
    input [63:0] input_63;
    input [63:0] input_62;
    input [63:0] input_61;
    input [63:0] input_60;
    input [63:0] input_59;
    input [63:0] input_58;
    input [63:0] input_57;
    input [63:0] input_56;
    input [63:0] input_55;
    input [63:0] input_54;
    input [63:0] input_53;
    input [63:0] input_52;
    input [63:0] input_51;
    input [63:0] input_50;
    input [63:0] input_49;
    input [63:0] input_48;
    input [63:0] input_47;
    input [63:0] input_46;
    input [63:0] input_45;
    input [63:0] input_44;
    input [63:0] input_43;
    input [63:0] input_42;
    input [63:0] input_41;
    input [63:0] input_40;
    input [63:0] input_39;
    input [63:0] input_38;
    input [63:0] input_37;
    input [63:0] input_36;
    input [63:0] input_35;
    input [63:0] input_34;
    input [63:0] input_33;
    input [63:0] input_32;
    input [63:0] input_31;
    input [63:0] input_30;
    input [63:0] input_29;
    input [63:0] input_28;
    input [63:0] input_27;
    input [63:0] input_26;
    input [63:0] input_25;
    input [63:0] input_24;
    input [63:0] input_23;
    input [63:0] input_22;
    input [63:0] input_21;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [67:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    result = result | ( input_21 & {64{sel[21]}});
    result = result | ( input_22 & {64{sel[22]}});
    result = result | ( input_23 & {64{sel[23]}});
    result = result | ( input_24 & {64{sel[24]}});
    result = result | ( input_25 & {64{sel[25]}});
    result = result | ( input_26 & {64{sel[26]}});
    result = result | ( input_27 & {64{sel[27]}});
    result = result | ( input_28 & {64{sel[28]}});
    result = result | ( input_29 & {64{sel[29]}});
    result = result | ( input_30 & {64{sel[30]}});
    result = result | ( input_31 & {64{sel[31]}});
    result = result | ( input_32 & {64{sel[32]}});
    result = result | ( input_33 & {64{sel[33]}});
    result = result | ( input_34 & {64{sel[34]}});
    result = result | ( input_35 & {64{sel[35]}});
    result = result | ( input_36 & {64{sel[36]}});
    result = result | ( input_37 & {64{sel[37]}});
    result = result | ( input_38 & {64{sel[38]}});
    result = result | ( input_39 & {64{sel[39]}});
    result = result | ( input_40 & {64{sel[40]}});
    result = result | ( input_41 & {64{sel[41]}});
    result = result | ( input_42 & {64{sel[42]}});
    result = result | ( input_43 & {64{sel[43]}});
    result = result | ( input_44 & {64{sel[44]}});
    result = result | ( input_45 & {64{sel[45]}});
    result = result | ( input_46 & {64{sel[46]}});
    result = result | ( input_47 & {64{sel[47]}});
    result = result | ( input_48 & {64{sel[48]}});
    result = result | ( input_49 & {64{sel[49]}});
    result = result | ( input_50 & {64{sel[50]}});
    result = result | ( input_51 & {64{sel[51]}});
    result = result | ( input_52 & {64{sel[52]}});
    result = result | ( input_53 & {64{sel[53]}});
    result = result | ( input_54 & {64{sel[54]}});
    result = result | ( input_55 & {64{sel[55]}});
    result = result | ( input_56 & {64{sel[56]}});
    result = result | ( input_57 & {64{sel[57]}});
    result = result | ( input_58 & {64{sel[58]}});
    result = result | ( input_59 & {64{sel[59]}});
    result = result | ( input_60 & {64{sel[60]}});
    result = result | ( input_61 & {64{sel[61]}});
    result = result | ( input_62 & {64{sel[62]}});
    result = result | ( input_63 & {64{sel[63]}});
    result = result | ( input_64 & {64{sel[64]}});
    result = result | ( input_65 & {64{sel[65]}});
    result = result | ( input_66 & {64{sel[66]}});
    result = result | ( input_67 & {64{sel[67]}});
    MUX1HOT_v_64_68_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_8_2;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [7:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    MUX1HOT_v_64_8_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_9_2;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [8:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    MUX1HOT_v_64_9_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [8:0] MUX1HOT_v_9_4_2;
    input [8:0] input_3;
    input [8:0] input_2;
    input [8:0] input_1;
    input [8:0] input_0;
    input [3:0] sel;
    reg [8:0] result;
  begin
    result = input_0 & {9{sel[0]}};
    result = result | ( input_1 & {9{sel[1]}});
    result = result | ( input_2 & {9{sel[2]}});
    result = result | ( input_3 & {9{sel[3]}});
    MUX1HOT_v_9_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input [0:0] sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [0:0] readslicef_11_1_10;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 10;
    readslicef_11_1_10 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] readslicef_12_11_1;
    input [11:0] vector;
    reg [11:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_12_11_1 = tmp[10:0];
  end
  endfunction


  function automatic [63:0] readslicef_65_64_1;
    input [64:0] vector;
    reg [64:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_65_64_1 = tmp[63:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [10:0] conv_u2s_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2s_10_11 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_u2u_11_12 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIF
// ------------------------------------------------------------------


module inPlaceNTT_DIF (
  clk, rst, vec_rsc_0_0_wadr, vec_rsc_0_0_d, vec_rsc_0_0_we, vec_rsc_0_0_radr, vec_rsc_0_0_q,
      vec_rsc_triosy_0_0_lz, vec_rsc_0_1_wadr, vec_rsc_0_1_d, vec_rsc_0_1_we, vec_rsc_0_1_radr,
      vec_rsc_0_1_q, vec_rsc_triosy_0_1_lz, vec_rsc_0_2_wadr, vec_rsc_0_2_d, vec_rsc_0_2_we,
      vec_rsc_0_2_radr, vec_rsc_0_2_q, vec_rsc_triosy_0_2_lz, vec_rsc_0_3_wadr, vec_rsc_0_3_d,
      vec_rsc_0_3_we, vec_rsc_0_3_radr, vec_rsc_0_3_q, vec_rsc_triosy_0_3_lz, vec_rsc_0_4_wadr,
      vec_rsc_0_4_d, vec_rsc_0_4_we, vec_rsc_0_4_radr, vec_rsc_0_4_q, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_wadr, vec_rsc_0_5_d, vec_rsc_0_5_we, vec_rsc_0_5_radr, vec_rsc_0_5_q,
      vec_rsc_triosy_0_5_lz, vec_rsc_0_6_wadr, vec_rsc_0_6_d, vec_rsc_0_6_we, vec_rsc_0_6_radr,
      vec_rsc_0_6_q, vec_rsc_triosy_0_6_lz, vec_rsc_0_7_wadr, vec_rsc_0_7_d, vec_rsc_0_7_we,
      vec_rsc_0_7_radr, vec_rsc_0_7_q, vec_rsc_triosy_0_7_lz, vec_rsc_0_8_wadr, vec_rsc_0_8_d,
      vec_rsc_0_8_we, vec_rsc_0_8_radr, vec_rsc_0_8_q, vec_rsc_triosy_0_8_lz, vec_rsc_0_9_wadr,
      vec_rsc_0_9_d, vec_rsc_0_9_we, vec_rsc_0_9_radr, vec_rsc_0_9_q, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_wadr, vec_rsc_0_10_d, vec_rsc_0_10_we, vec_rsc_0_10_radr, vec_rsc_0_10_q,
      vec_rsc_triosy_0_10_lz, vec_rsc_0_11_wadr, vec_rsc_0_11_d, vec_rsc_0_11_we,
      vec_rsc_0_11_radr, vec_rsc_0_11_q, vec_rsc_triosy_0_11_lz, vec_rsc_0_12_wadr,
      vec_rsc_0_12_d, vec_rsc_0_12_we, vec_rsc_0_12_radr, vec_rsc_0_12_q, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_wadr, vec_rsc_0_13_d, vec_rsc_0_13_we, vec_rsc_0_13_radr, vec_rsc_0_13_q,
      vec_rsc_triosy_0_13_lz, vec_rsc_0_14_wadr, vec_rsc_0_14_d, vec_rsc_0_14_we,
      vec_rsc_0_14_radr, vec_rsc_0_14_q, vec_rsc_triosy_0_14_lz, vec_rsc_0_15_wadr,
      vec_rsc_0_15_d, vec_rsc_0_15_we, vec_rsc_0_15_radr, vec_rsc_0_15_q, vec_rsc_triosy_0_15_lz,
      vec_rsc_0_16_wadr, vec_rsc_0_16_d, vec_rsc_0_16_we, vec_rsc_0_16_radr, vec_rsc_0_16_q,
      vec_rsc_triosy_0_16_lz, vec_rsc_0_17_wadr, vec_rsc_0_17_d, vec_rsc_0_17_we,
      vec_rsc_0_17_radr, vec_rsc_0_17_q, vec_rsc_triosy_0_17_lz, vec_rsc_0_18_wadr,
      vec_rsc_0_18_d, vec_rsc_0_18_we, vec_rsc_0_18_radr, vec_rsc_0_18_q, vec_rsc_triosy_0_18_lz,
      vec_rsc_0_19_wadr, vec_rsc_0_19_d, vec_rsc_0_19_we, vec_rsc_0_19_radr, vec_rsc_0_19_q,
      vec_rsc_triosy_0_19_lz, vec_rsc_0_20_wadr, vec_rsc_0_20_d, vec_rsc_0_20_we,
      vec_rsc_0_20_radr, vec_rsc_0_20_q, vec_rsc_triosy_0_20_lz, vec_rsc_0_21_wadr,
      vec_rsc_0_21_d, vec_rsc_0_21_we, vec_rsc_0_21_radr, vec_rsc_0_21_q, vec_rsc_triosy_0_21_lz,
      vec_rsc_0_22_wadr, vec_rsc_0_22_d, vec_rsc_0_22_we, vec_rsc_0_22_radr, vec_rsc_0_22_q,
      vec_rsc_triosy_0_22_lz, vec_rsc_0_23_wadr, vec_rsc_0_23_d, vec_rsc_0_23_we,
      vec_rsc_0_23_radr, vec_rsc_0_23_q, vec_rsc_triosy_0_23_lz, vec_rsc_0_24_wadr,
      vec_rsc_0_24_d, vec_rsc_0_24_we, vec_rsc_0_24_radr, vec_rsc_0_24_q, vec_rsc_triosy_0_24_lz,
      vec_rsc_0_25_wadr, vec_rsc_0_25_d, vec_rsc_0_25_we, vec_rsc_0_25_radr, vec_rsc_0_25_q,
      vec_rsc_triosy_0_25_lz, vec_rsc_0_26_wadr, vec_rsc_0_26_d, vec_rsc_0_26_we,
      vec_rsc_0_26_radr, vec_rsc_0_26_q, vec_rsc_triosy_0_26_lz, vec_rsc_0_27_wadr,
      vec_rsc_0_27_d, vec_rsc_0_27_we, vec_rsc_0_27_radr, vec_rsc_0_27_q, vec_rsc_triosy_0_27_lz,
      vec_rsc_0_28_wadr, vec_rsc_0_28_d, vec_rsc_0_28_we, vec_rsc_0_28_radr, vec_rsc_0_28_q,
      vec_rsc_triosy_0_28_lz, vec_rsc_0_29_wadr, vec_rsc_0_29_d, vec_rsc_0_29_we,
      vec_rsc_0_29_radr, vec_rsc_0_29_q, vec_rsc_triosy_0_29_lz, vec_rsc_0_30_wadr,
      vec_rsc_0_30_d, vec_rsc_0_30_we, vec_rsc_0_30_radr, vec_rsc_0_30_q, vec_rsc_triosy_0_30_lz,
      vec_rsc_0_31_wadr, vec_rsc_0_31_d, vec_rsc_0_31_we, vec_rsc_0_31_radr, vec_rsc_0_31_q,
      vec_rsc_triosy_0_31_lz, vec_rsc_0_32_wadr, vec_rsc_0_32_d, vec_rsc_0_32_we,
      vec_rsc_0_32_radr, vec_rsc_0_32_q, vec_rsc_triosy_0_32_lz, vec_rsc_0_33_wadr,
      vec_rsc_0_33_d, vec_rsc_0_33_we, vec_rsc_0_33_radr, vec_rsc_0_33_q, vec_rsc_triosy_0_33_lz,
      vec_rsc_0_34_wadr, vec_rsc_0_34_d, vec_rsc_0_34_we, vec_rsc_0_34_radr, vec_rsc_0_34_q,
      vec_rsc_triosy_0_34_lz, vec_rsc_0_35_wadr, vec_rsc_0_35_d, vec_rsc_0_35_we,
      vec_rsc_0_35_radr, vec_rsc_0_35_q, vec_rsc_triosy_0_35_lz, vec_rsc_0_36_wadr,
      vec_rsc_0_36_d, vec_rsc_0_36_we, vec_rsc_0_36_radr, vec_rsc_0_36_q, vec_rsc_triosy_0_36_lz,
      vec_rsc_0_37_wadr, vec_rsc_0_37_d, vec_rsc_0_37_we, vec_rsc_0_37_radr, vec_rsc_0_37_q,
      vec_rsc_triosy_0_37_lz, vec_rsc_0_38_wadr, vec_rsc_0_38_d, vec_rsc_0_38_we,
      vec_rsc_0_38_radr, vec_rsc_0_38_q, vec_rsc_triosy_0_38_lz, vec_rsc_0_39_wadr,
      vec_rsc_0_39_d, vec_rsc_0_39_we, vec_rsc_0_39_radr, vec_rsc_0_39_q, vec_rsc_triosy_0_39_lz,
      vec_rsc_0_40_wadr, vec_rsc_0_40_d, vec_rsc_0_40_we, vec_rsc_0_40_radr, vec_rsc_0_40_q,
      vec_rsc_triosy_0_40_lz, vec_rsc_0_41_wadr, vec_rsc_0_41_d, vec_rsc_0_41_we,
      vec_rsc_0_41_radr, vec_rsc_0_41_q, vec_rsc_triosy_0_41_lz, vec_rsc_0_42_wadr,
      vec_rsc_0_42_d, vec_rsc_0_42_we, vec_rsc_0_42_radr, vec_rsc_0_42_q, vec_rsc_triosy_0_42_lz,
      vec_rsc_0_43_wadr, vec_rsc_0_43_d, vec_rsc_0_43_we, vec_rsc_0_43_radr, vec_rsc_0_43_q,
      vec_rsc_triosy_0_43_lz, vec_rsc_0_44_wadr, vec_rsc_0_44_d, vec_rsc_0_44_we,
      vec_rsc_0_44_radr, vec_rsc_0_44_q, vec_rsc_triosy_0_44_lz, vec_rsc_0_45_wadr,
      vec_rsc_0_45_d, vec_rsc_0_45_we, vec_rsc_0_45_radr, vec_rsc_0_45_q, vec_rsc_triosy_0_45_lz,
      vec_rsc_0_46_wadr, vec_rsc_0_46_d, vec_rsc_0_46_we, vec_rsc_0_46_radr, vec_rsc_0_46_q,
      vec_rsc_triosy_0_46_lz, vec_rsc_0_47_wadr, vec_rsc_0_47_d, vec_rsc_0_47_we,
      vec_rsc_0_47_radr, vec_rsc_0_47_q, vec_rsc_triosy_0_47_lz, vec_rsc_0_48_wadr,
      vec_rsc_0_48_d, vec_rsc_0_48_we, vec_rsc_0_48_radr, vec_rsc_0_48_q, vec_rsc_triosy_0_48_lz,
      vec_rsc_0_49_wadr, vec_rsc_0_49_d, vec_rsc_0_49_we, vec_rsc_0_49_radr, vec_rsc_0_49_q,
      vec_rsc_triosy_0_49_lz, vec_rsc_0_50_wadr, vec_rsc_0_50_d, vec_rsc_0_50_we,
      vec_rsc_0_50_radr, vec_rsc_0_50_q, vec_rsc_triosy_0_50_lz, vec_rsc_0_51_wadr,
      vec_rsc_0_51_d, vec_rsc_0_51_we, vec_rsc_0_51_radr, vec_rsc_0_51_q, vec_rsc_triosy_0_51_lz,
      vec_rsc_0_52_wadr, vec_rsc_0_52_d, vec_rsc_0_52_we, vec_rsc_0_52_radr, vec_rsc_0_52_q,
      vec_rsc_triosy_0_52_lz, vec_rsc_0_53_wadr, vec_rsc_0_53_d, vec_rsc_0_53_we,
      vec_rsc_0_53_radr, vec_rsc_0_53_q, vec_rsc_triosy_0_53_lz, vec_rsc_0_54_wadr,
      vec_rsc_0_54_d, vec_rsc_0_54_we, vec_rsc_0_54_radr, vec_rsc_0_54_q, vec_rsc_triosy_0_54_lz,
      vec_rsc_0_55_wadr, vec_rsc_0_55_d, vec_rsc_0_55_we, vec_rsc_0_55_radr, vec_rsc_0_55_q,
      vec_rsc_triosy_0_55_lz, vec_rsc_0_56_wadr, vec_rsc_0_56_d, vec_rsc_0_56_we,
      vec_rsc_0_56_radr, vec_rsc_0_56_q, vec_rsc_triosy_0_56_lz, vec_rsc_0_57_wadr,
      vec_rsc_0_57_d, vec_rsc_0_57_we, vec_rsc_0_57_radr, vec_rsc_0_57_q, vec_rsc_triosy_0_57_lz,
      vec_rsc_0_58_wadr, vec_rsc_0_58_d, vec_rsc_0_58_we, vec_rsc_0_58_radr, vec_rsc_0_58_q,
      vec_rsc_triosy_0_58_lz, vec_rsc_0_59_wadr, vec_rsc_0_59_d, vec_rsc_0_59_we,
      vec_rsc_0_59_radr, vec_rsc_0_59_q, vec_rsc_triosy_0_59_lz, vec_rsc_0_60_wadr,
      vec_rsc_0_60_d, vec_rsc_0_60_we, vec_rsc_0_60_radr, vec_rsc_0_60_q, vec_rsc_triosy_0_60_lz,
      vec_rsc_0_61_wadr, vec_rsc_0_61_d, vec_rsc_0_61_we, vec_rsc_0_61_radr, vec_rsc_0_61_q,
      vec_rsc_triosy_0_61_lz, vec_rsc_0_62_wadr, vec_rsc_0_62_d, vec_rsc_0_62_we,
      vec_rsc_0_62_radr, vec_rsc_0_62_q, vec_rsc_triosy_0_62_lz, vec_rsc_0_63_wadr,
      vec_rsc_0_63_d, vec_rsc_0_63_we, vec_rsc_0_63_radr, vec_rsc_0_63_q, vec_rsc_triosy_0_63_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz, twiddle_rsc_0_0_radr,
      twiddle_rsc_0_0_q, twiddle_rsc_triosy_0_0_lz, twiddle_rsc_0_1_radr, twiddle_rsc_0_1_q,
      twiddle_rsc_triosy_0_1_lz, twiddle_rsc_0_2_radr, twiddle_rsc_0_2_q, twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_0_3_radr, twiddle_rsc_0_3_q, twiddle_rsc_triosy_0_3_lz, twiddle_rsc_0_4_radr,
      twiddle_rsc_0_4_q, twiddle_rsc_triosy_0_4_lz, twiddle_rsc_0_5_radr, twiddle_rsc_0_5_q,
      twiddle_rsc_triosy_0_5_lz, twiddle_rsc_0_6_radr, twiddle_rsc_0_6_q, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_0_7_radr, twiddle_rsc_0_7_q, twiddle_rsc_triosy_0_7_lz, twiddle_rsc_0_8_radr,
      twiddle_rsc_0_8_q, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_0_9_radr, twiddle_rsc_0_9_q,
      twiddle_rsc_triosy_0_9_lz, twiddle_rsc_0_10_radr, twiddle_rsc_0_10_q, twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_0_11_radr, twiddle_rsc_0_11_q, twiddle_rsc_triosy_0_11_lz, twiddle_rsc_0_12_radr,
      twiddle_rsc_0_12_q, twiddle_rsc_triosy_0_12_lz, twiddle_rsc_0_13_radr, twiddle_rsc_0_13_q,
      twiddle_rsc_triosy_0_13_lz, twiddle_rsc_0_14_radr, twiddle_rsc_0_14_q, twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_0_15_radr, twiddle_rsc_0_15_q, twiddle_rsc_triosy_0_15_lz, twiddle_rsc_0_16_radr,
      twiddle_rsc_0_16_q, twiddle_rsc_triosy_0_16_lz, twiddle_rsc_0_17_radr, twiddle_rsc_0_17_q,
      twiddle_rsc_triosy_0_17_lz, twiddle_rsc_0_18_radr, twiddle_rsc_0_18_q, twiddle_rsc_triosy_0_18_lz,
      twiddle_rsc_0_19_radr, twiddle_rsc_0_19_q, twiddle_rsc_triosy_0_19_lz, twiddle_rsc_0_20_radr,
      twiddle_rsc_0_20_q, twiddle_rsc_triosy_0_20_lz, twiddle_rsc_0_21_radr, twiddle_rsc_0_21_q,
      twiddle_rsc_triosy_0_21_lz, twiddle_rsc_0_22_radr, twiddle_rsc_0_22_q, twiddle_rsc_triosy_0_22_lz,
      twiddle_rsc_0_23_radr, twiddle_rsc_0_23_q, twiddle_rsc_triosy_0_23_lz, twiddle_rsc_0_24_radr,
      twiddle_rsc_0_24_q, twiddle_rsc_triosy_0_24_lz, twiddle_rsc_0_25_radr, twiddle_rsc_0_25_q,
      twiddle_rsc_triosy_0_25_lz, twiddle_rsc_0_26_radr, twiddle_rsc_0_26_q, twiddle_rsc_triosy_0_26_lz,
      twiddle_rsc_0_27_radr, twiddle_rsc_0_27_q, twiddle_rsc_triosy_0_27_lz, twiddle_rsc_0_28_radr,
      twiddle_rsc_0_28_q, twiddle_rsc_triosy_0_28_lz, twiddle_rsc_0_29_radr, twiddle_rsc_0_29_q,
      twiddle_rsc_triosy_0_29_lz, twiddle_rsc_0_30_radr, twiddle_rsc_0_30_q, twiddle_rsc_triosy_0_30_lz,
      twiddle_rsc_0_31_radr, twiddle_rsc_0_31_q, twiddle_rsc_triosy_0_31_lz, twiddle_rsc_0_32_radr,
      twiddle_rsc_0_32_q, twiddle_rsc_triosy_0_32_lz, twiddle_rsc_0_33_radr, twiddle_rsc_0_33_q,
      twiddle_rsc_triosy_0_33_lz, twiddle_rsc_0_34_radr, twiddle_rsc_0_34_q, twiddle_rsc_triosy_0_34_lz,
      twiddle_rsc_0_35_radr, twiddle_rsc_0_35_q, twiddle_rsc_triosy_0_35_lz, twiddle_rsc_0_36_radr,
      twiddle_rsc_0_36_q, twiddle_rsc_triosy_0_36_lz, twiddle_rsc_0_37_radr, twiddle_rsc_0_37_q,
      twiddle_rsc_triosy_0_37_lz, twiddle_rsc_0_38_radr, twiddle_rsc_0_38_q, twiddle_rsc_triosy_0_38_lz,
      twiddle_rsc_0_39_radr, twiddle_rsc_0_39_q, twiddle_rsc_triosy_0_39_lz, twiddle_rsc_0_40_radr,
      twiddle_rsc_0_40_q, twiddle_rsc_triosy_0_40_lz, twiddle_rsc_0_41_radr, twiddle_rsc_0_41_q,
      twiddle_rsc_triosy_0_41_lz, twiddle_rsc_0_42_radr, twiddle_rsc_0_42_q, twiddle_rsc_triosy_0_42_lz,
      twiddle_rsc_0_43_radr, twiddle_rsc_0_43_q, twiddle_rsc_triosy_0_43_lz, twiddle_rsc_0_44_radr,
      twiddle_rsc_0_44_q, twiddle_rsc_triosy_0_44_lz, twiddle_rsc_0_45_radr, twiddle_rsc_0_45_q,
      twiddle_rsc_triosy_0_45_lz, twiddle_rsc_0_46_radr, twiddle_rsc_0_46_q, twiddle_rsc_triosy_0_46_lz,
      twiddle_rsc_0_47_radr, twiddle_rsc_0_47_q, twiddle_rsc_triosy_0_47_lz, twiddle_rsc_0_48_radr,
      twiddle_rsc_0_48_q, twiddle_rsc_triosy_0_48_lz, twiddle_rsc_0_49_radr, twiddle_rsc_0_49_q,
      twiddle_rsc_triosy_0_49_lz, twiddle_rsc_0_50_radr, twiddle_rsc_0_50_q, twiddle_rsc_triosy_0_50_lz,
      twiddle_rsc_0_51_radr, twiddle_rsc_0_51_q, twiddle_rsc_triosy_0_51_lz, twiddle_rsc_0_52_radr,
      twiddle_rsc_0_52_q, twiddle_rsc_triosy_0_52_lz, twiddle_rsc_0_53_radr, twiddle_rsc_0_53_q,
      twiddle_rsc_triosy_0_53_lz, twiddle_rsc_0_54_radr, twiddle_rsc_0_54_q, twiddle_rsc_triosy_0_54_lz,
      twiddle_rsc_0_55_radr, twiddle_rsc_0_55_q, twiddle_rsc_triosy_0_55_lz, twiddle_rsc_0_56_radr,
      twiddle_rsc_0_56_q, twiddle_rsc_triosy_0_56_lz, twiddle_rsc_0_57_radr, twiddle_rsc_0_57_q,
      twiddle_rsc_triosy_0_57_lz, twiddle_rsc_0_58_radr, twiddle_rsc_0_58_q, twiddle_rsc_triosy_0_58_lz,
      twiddle_rsc_0_59_radr, twiddle_rsc_0_59_q, twiddle_rsc_triosy_0_59_lz, twiddle_rsc_0_60_radr,
      twiddle_rsc_0_60_q, twiddle_rsc_triosy_0_60_lz, twiddle_rsc_0_61_radr, twiddle_rsc_0_61_q,
      twiddle_rsc_triosy_0_61_lz, twiddle_rsc_0_62_radr, twiddle_rsc_0_62_q, twiddle_rsc_triosy_0_62_lz,
      twiddle_rsc_0_63_radr, twiddle_rsc_0_63_q, twiddle_rsc_triosy_0_63_lz
);
  input clk;
  input rst;
  output [3:0] vec_rsc_0_0_wadr;
  output [63:0] vec_rsc_0_0_d;
  output vec_rsc_0_0_we;
  output [3:0] vec_rsc_0_0_radr;
  input [63:0] vec_rsc_0_0_q;
  output vec_rsc_triosy_0_0_lz;
  output [3:0] vec_rsc_0_1_wadr;
  output [63:0] vec_rsc_0_1_d;
  output vec_rsc_0_1_we;
  output [3:0] vec_rsc_0_1_radr;
  input [63:0] vec_rsc_0_1_q;
  output vec_rsc_triosy_0_1_lz;
  output [3:0] vec_rsc_0_2_wadr;
  output [63:0] vec_rsc_0_2_d;
  output vec_rsc_0_2_we;
  output [3:0] vec_rsc_0_2_radr;
  input [63:0] vec_rsc_0_2_q;
  output vec_rsc_triosy_0_2_lz;
  output [3:0] vec_rsc_0_3_wadr;
  output [63:0] vec_rsc_0_3_d;
  output vec_rsc_0_3_we;
  output [3:0] vec_rsc_0_3_radr;
  input [63:0] vec_rsc_0_3_q;
  output vec_rsc_triosy_0_3_lz;
  output [3:0] vec_rsc_0_4_wadr;
  output [63:0] vec_rsc_0_4_d;
  output vec_rsc_0_4_we;
  output [3:0] vec_rsc_0_4_radr;
  input [63:0] vec_rsc_0_4_q;
  output vec_rsc_triosy_0_4_lz;
  output [3:0] vec_rsc_0_5_wadr;
  output [63:0] vec_rsc_0_5_d;
  output vec_rsc_0_5_we;
  output [3:0] vec_rsc_0_5_radr;
  input [63:0] vec_rsc_0_5_q;
  output vec_rsc_triosy_0_5_lz;
  output [3:0] vec_rsc_0_6_wadr;
  output [63:0] vec_rsc_0_6_d;
  output vec_rsc_0_6_we;
  output [3:0] vec_rsc_0_6_radr;
  input [63:0] vec_rsc_0_6_q;
  output vec_rsc_triosy_0_6_lz;
  output [3:0] vec_rsc_0_7_wadr;
  output [63:0] vec_rsc_0_7_d;
  output vec_rsc_0_7_we;
  output [3:0] vec_rsc_0_7_radr;
  input [63:0] vec_rsc_0_7_q;
  output vec_rsc_triosy_0_7_lz;
  output [3:0] vec_rsc_0_8_wadr;
  output [63:0] vec_rsc_0_8_d;
  output vec_rsc_0_8_we;
  output [3:0] vec_rsc_0_8_radr;
  input [63:0] vec_rsc_0_8_q;
  output vec_rsc_triosy_0_8_lz;
  output [3:0] vec_rsc_0_9_wadr;
  output [63:0] vec_rsc_0_9_d;
  output vec_rsc_0_9_we;
  output [3:0] vec_rsc_0_9_radr;
  input [63:0] vec_rsc_0_9_q;
  output vec_rsc_triosy_0_9_lz;
  output [3:0] vec_rsc_0_10_wadr;
  output [63:0] vec_rsc_0_10_d;
  output vec_rsc_0_10_we;
  output [3:0] vec_rsc_0_10_radr;
  input [63:0] vec_rsc_0_10_q;
  output vec_rsc_triosy_0_10_lz;
  output [3:0] vec_rsc_0_11_wadr;
  output [63:0] vec_rsc_0_11_d;
  output vec_rsc_0_11_we;
  output [3:0] vec_rsc_0_11_radr;
  input [63:0] vec_rsc_0_11_q;
  output vec_rsc_triosy_0_11_lz;
  output [3:0] vec_rsc_0_12_wadr;
  output [63:0] vec_rsc_0_12_d;
  output vec_rsc_0_12_we;
  output [3:0] vec_rsc_0_12_radr;
  input [63:0] vec_rsc_0_12_q;
  output vec_rsc_triosy_0_12_lz;
  output [3:0] vec_rsc_0_13_wadr;
  output [63:0] vec_rsc_0_13_d;
  output vec_rsc_0_13_we;
  output [3:0] vec_rsc_0_13_radr;
  input [63:0] vec_rsc_0_13_q;
  output vec_rsc_triosy_0_13_lz;
  output [3:0] vec_rsc_0_14_wadr;
  output [63:0] vec_rsc_0_14_d;
  output vec_rsc_0_14_we;
  output [3:0] vec_rsc_0_14_radr;
  input [63:0] vec_rsc_0_14_q;
  output vec_rsc_triosy_0_14_lz;
  output [3:0] vec_rsc_0_15_wadr;
  output [63:0] vec_rsc_0_15_d;
  output vec_rsc_0_15_we;
  output [3:0] vec_rsc_0_15_radr;
  input [63:0] vec_rsc_0_15_q;
  output vec_rsc_triosy_0_15_lz;
  output [3:0] vec_rsc_0_16_wadr;
  output [63:0] vec_rsc_0_16_d;
  output vec_rsc_0_16_we;
  output [3:0] vec_rsc_0_16_radr;
  input [63:0] vec_rsc_0_16_q;
  output vec_rsc_triosy_0_16_lz;
  output [3:0] vec_rsc_0_17_wadr;
  output [63:0] vec_rsc_0_17_d;
  output vec_rsc_0_17_we;
  output [3:0] vec_rsc_0_17_radr;
  input [63:0] vec_rsc_0_17_q;
  output vec_rsc_triosy_0_17_lz;
  output [3:0] vec_rsc_0_18_wadr;
  output [63:0] vec_rsc_0_18_d;
  output vec_rsc_0_18_we;
  output [3:0] vec_rsc_0_18_radr;
  input [63:0] vec_rsc_0_18_q;
  output vec_rsc_triosy_0_18_lz;
  output [3:0] vec_rsc_0_19_wadr;
  output [63:0] vec_rsc_0_19_d;
  output vec_rsc_0_19_we;
  output [3:0] vec_rsc_0_19_radr;
  input [63:0] vec_rsc_0_19_q;
  output vec_rsc_triosy_0_19_lz;
  output [3:0] vec_rsc_0_20_wadr;
  output [63:0] vec_rsc_0_20_d;
  output vec_rsc_0_20_we;
  output [3:0] vec_rsc_0_20_radr;
  input [63:0] vec_rsc_0_20_q;
  output vec_rsc_triosy_0_20_lz;
  output [3:0] vec_rsc_0_21_wadr;
  output [63:0] vec_rsc_0_21_d;
  output vec_rsc_0_21_we;
  output [3:0] vec_rsc_0_21_radr;
  input [63:0] vec_rsc_0_21_q;
  output vec_rsc_triosy_0_21_lz;
  output [3:0] vec_rsc_0_22_wadr;
  output [63:0] vec_rsc_0_22_d;
  output vec_rsc_0_22_we;
  output [3:0] vec_rsc_0_22_radr;
  input [63:0] vec_rsc_0_22_q;
  output vec_rsc_triosy_0_22_lz;
  output [3:0] vec_rsc_0_23_wadr;
  output [63:0] vec_rsc_0_23_d;
  output vec_rsc_0_23_we;
  output [3:0] vec_rsc_0_23_radr;
  input [63:0] vec_rsc_0_23_q;
  output vec_rsc_triosy_0_23_lz;
  output [3:0] vec_rsc_0_24_wadr;
  output [63:0] vec_rsc_0_24_d;
  output vec_rsc_0_24_we;
  output [3:0] vec_rsc_0_24_radr;
  input [63:0] vec_rsc_0_24_q;
  output vec_rsc_triosy_0_24_lz;
  output [3:0] vec_rsc_0_25_wadr;
  output [63:0] vec_rsc_0_25_d;
  output vec_rsc_0_25_we;
  output [3:0] vec_rsc_0_25_radr;
  input [63:0] vec_rsc_0_25_q;
  output vec_rsc_triosy_0_25_lz;
  output [3:0] vec_rsc_0_26_wadr;
  output [63:0] vec_rsc_0_26_d;
  output vec_rsc_0_26_we;
  output [3:0] vec_rsc_0_26_radr;
  input [63:0] vec_rsc_0_26_q;
  output vec_rsc_triosy_0_26_lz;
  output [3:0] vec_rsc_0_27_wadr;
  output [63:0] vec_rsc_0_27_d;
  output vec_rsc_0_27_we;
  output [3:0] vec_rsc_0_27_radr;
  input [63:0] vec_rsc_0_27_q;
  output vec_rsc_triosy_0_27_lz;
  output [3:0] vec_rsc_0_28_wadr;
  output [63:0] vec_rsc_0_28_d;
  output vec_rsc_0_28_we;
  output [3:0] vec_rsc_0_28_radr;
  input [63:0] vec_rsc_0_28_q;
  output vec_rsc_triosy_0_28_lz;
  output [3:0] vec_rsc_0_29_wadr;
  output [63:0] vec_rsc_0_29_d;
  output vec_rsc_0_29_we;
  output [3:0] vec_rsc_0_29_radr;
  input [63:0] vec_rsc_0_29_q;
  output vec_rsc_triosy_0_29_lz;
  output [3:0] vec_rsc_0_30_wadr;
  output [63:0] vec_rsc_0_30_d;
  output vec_rsc_0_30_we;
  output [3:0] vec_rsc_0_30_radr;
  input [63:0] vec_rsc_0_30_q;
  output vec_rsc_triosy_0_30_lz;
  output [3:0] vec_rsc_0_31_wadr;
  output [63:0] vec_rsc_0_31_d;
  output vec_rsc_0_31_we;
  output [3:0] vec_rsc_0_31_radr;
  input [63:0] vec_rsc_0_31_q;
  output vec_rsc_triosy_0_31_lz;
  output [3:0] vec_rsc_0_32_wadr;
  output [63:0] vec_rsc_0_32_d;
  output vec_rsc_0_32_we;
  output [3:0] vec_rsc_0_32_radr;
  input [63:0] vec_rsc_0_32_q;
  output vec_rsc_triosy_0_32_lz;
  output [3:0] vec_rsc_0_33_wadr;
  output [63:0] vec_rsc_0_33_d;
  output vec_rsc_0_33_we;
  output [3:0] vec_rsc_0_33_radr;
  input [63:0] vec_rsc_0_33_q;
  output vec_rsc_triosy_0_33_lz;
  output [3:0] vec_rsc_0_34_wadr;
  output [63:0] vec_rsc_0_34_d;
  output vec_rsc_0_34_we;
  output [3:0] vec_rsc_0_34_radr;
  input [63:0] vec_rsc_0_34_q;
  output vec_rsc_triosy_0_34_lz;
  output [3:0] vec_rsc_0_35_wadr;
  output [63:0] vec_rsc_0_35_d;
  output vec_rsc_0_35_we;
  output [3:0] vec_rsc_0_35_radr;
  input [63:0] vec_rsc_0_35_q;
  output vec_rsc_triosy_0_35_lz;
  output [3:0] vec_rsc_0_36_wadr;
  output [63:0] vec_rsc_0_36_d;
  output vec_rsc_0_36_we;
  output [3:0] vec_rsc_0_36_radr;
  input [63:0] vec_rsc_0_36_q;
  output vec_rsc_triosy_0_36_lz;
  output [3:0] vec_rsc_0_37_wadr;
  output [63:0] vec_rsc_0_37_d;
  output vec_rsc_0_37_we;
  output [3:0] vec_rsc_0_37_radr;
  input [63:0] vec_rsc_0_37_q;
  output vec_rsc_triosy_0_37_lz;
  output [3:0] vec_rsc_0_38_wadr;
  output [63:0] vec_rsc_0_38_d;
  output vec_rsc_0_38_we;
  output [3:0] vec_rsc_0_38_radr;
  input [63:0] vec_rsc_0_38_q;
  output vec_rsc_triosy_0_38_lz;
  output [3:0] vec_rsc_0_39_wadr;
  output [63:0] vec_rsc_0_39_d;
  output vec_rsc_0_39_we;
  output [3:0] vec_rsc_0_39_radr;
  input [63:0] vec_rsc_0_39_q;
  output vec_rsc_triosy_0_39_lz;
  output [3:0] vec_rsc_0_40_wadr;
  output [63:0] vec_rsc_0_40_d;
  output vec_rsc_0_40_we;
  output [3:0] vec_rsc_0_40_radr;
  input [63:0] vec_rsc_0_40_q;
  output vec_rsc_triosy_0_40_lz;
  output [3:0] vec_rsc_0_41_wadr;
  output [63:0] vec_rsc_0_41_d;
  output vec_rsc_0_41_we;
  output [3:0] vec_rsc_0_41_radr;
  input [63:0] vec_rsc_0_41_q;
  output vec_rsc_triosy_0_41_lz;
  output [3:0] vec_rsc_0_42_wadr;
  output [63:0] vec_rsc_0_42_d;
  output vec_rsc_0_42_we;
  output [3:0] vec_rsc_0_42_radr;
  input [63:0] vec_rsc_0_42_q;
  output vec_rsc_triosy_0_42_lz;
  output [3:0] vec_rsc_0_43_wadr;
  output [63:0] vec_rsc_0_43_d;
  output vec_rsc_0_43_we;
  output [3:0] vec_rsc_0_43_radr;
  input [63:0] vec_rsc_0_43_q;
  output vec_rsc_triosy_0_43_lz;
  output [3:0] vec_rsc_0_44_wadr;
  output [63:0] vec_rsc_0_44_d;
  output vec_rsc_0_44_we;
  output [3:0] vec_rsc_0_44_radr;
  input [63:0] vec_rsc_0_44_q;
  output vec_rsc_triosy_0_44_lz;
  output [3:0] vec_rsc_0_45_wadr;
  output [63:0] vec_rsc_0_45_d;
  output vec_rsc_0_45_we;
  output [3:0] vec_rsc_0_45_radr;
  input [63:0] vec_rsc_0_45_q;
  output vec_rsc_triosy_0_45_lz;
  output [3:0] vec_rsc_0_46_wadr;
  output [63:0] vec_rsc_0_46_d;
  output vec_rsc_0_46_we;
  output [3:0] vec_rsc_0_46_radr;
  input [63:0] vec_rsc_0_46_q;
  output vec_rsc_triosy_0_46_lz;
  output [3:0] vec_rsc_0_47_wadr;
  output [63:0] vec_rsc_0_47_d;
  output vec_rsc_0_47_we;
  output [3:0] vec_rsc_0_47_radr;
  input [63:0] vec_rsc_0_47_q;
  output vec_rsc_triosy_0_47_lz;
  output [3:0] vec_rsc_0_48_wadr;
  output [63:0] vec_rsc_0_48_d;
  output vec_rsc_0_48_we;
  output [3:0] vec_rsc_0_48_radr;
  input [63:0] vec_rsc_0_48_q;
  output vec_rsc_triosy_0_48_lz;
  output [3:0] vec_rsc_0_49_wadr;
  output [63:0] vec_rsc_0_49_d;
  output vec_rsc_0_49_we;
  output [3:0] vec_rsc_0_49_radr;
  input [63:0] vec_rsc_0_49_q;
  output vec_rsc_triosy_0_49_lz;
  output [3:0] vec_rsc_0_50_wadr;
  output [63:0] vec_rsc_0_50_d;
  output vec_rsc_0_50_we;
  output [3:0] vec_rsc_0_50_radr;
  input [63:0] vec_rsc_0_50_q;
  output vec_rsc_triosy_0_50_lz;
  output [3:0] vec_rsc_0_51_wadr;
  output [63:0] vec_rsc_0_51_d;
  output vec_rsc_0_51_we;
  output [3:0] vec_rsc_0_51_radr;
  input [63:0] vec_rsc_0_51_q;
  output vec_rsc_triosy_0_51_lz;
  output [3:0] vec_rsc_0_52_wadr;
  output [63:0] vec_rsc_0_52_d;
  output vec_rsc_0_52_we;
  output [3:0] vec_rsc_0_52_radr;
  input [63:0] vec_rsc_0_52_q;
  output vec_rsc_triosy_0_52_lz;
  output [3:0] vec_rsc_0_53_wadr;
  output [63:0] vec_rsc_0_53_d;
  output vec_rsc_0_53_we;
  output [3:0] vec_rsc_0_53_radr;
  input [63:0] vec_rsc_0_53_q;
  output vec_rsc_triosy_0_53_lz;
  output [3:0] vec_rsc_0_54_wadr;
  output [63:0] vec_rsc_0_54_d;
  output vec_rsc_0_54_we;
  output [3:0] vec_rsc_0_54_radr;
  input [63:0] vec_rsc_0_54_q;
  output vec_rsc_triosy_0_54_lz;
  output [3:0] vec_rsc_0_55_wadr;
  output [63:0] vec_rsc_0_55_d;
  output vec_rsc_0_55_we;
  output [3:0] vec_rsc_0_55_radr;
  input [63:0] vec_rsc_0_55_q;
  output vec_rsc_triosy_0_55_lz;
  output [3:0] vec_rsc_0_56_wadr;
  output [63:0] vec_rsc_0_56_d;
  output vec_rsc_0_56_we;
  output [3:0] vec_rsc_0_56_radr;
  input [63:0] vec_rsc_0_56_q;
  output vec_rsc_triosy_0_56_lz;
  output [3:0] vec_rsc_0_57_wadr;
  output [63:0] vec_rsc_0_57_d;
  output vec_rsc_0_57_we;
  output [3:0] vec_rsc_0_57_radr;
  input [63:0] vec_rsc_0_57_q;
  output vec_rsc_triosy_0_57_lz;
  output [3:0] vec_rsc_0_58_wadr;
  output [63:0] vec_rsc_0_58_d;
  output vec_rsc_0_58_we;
  output [3:0] vec_rsc_0_58_radr;
  input [63:0] vec_rsc_0_58_q;
  output vec_rsc_triosy_0_58_lz;
  output [3:0] vec_rsc_0_59_wadr;
  output [63:0] vec_rsc_0_59_d;
  output vec_rsc_0_59_we;
  output [3:0] vec_rsc_0_59_radr;
  input [63:0] vec_rsc_0_59_q;
  output vec_rsc_triosy_0_59_lz;
  output [3:0] vec_rsc_0_60_wadr;
  output [63:0] vec_rsc_0_60_d;
  output vec_rsc_0_60_we;
  output [3:0] vec_rsc_0_60_radr;
  input [63:0] vec_rsc_0_60_q;
  output vec_rsc_triosy_0_60_lz;
  output [3:0] vec_rsc_0_61_wadr;
  output [63:0] vec_rsc_0_61_d;
  output vec_rsc_0_61_we;
  output [3:0] vec_rsc_0_61_radr;
  input [63:0] vec_rsc_0_61_q;
  output vec_rsc_triosy_0_61_lz;
  output [3:0] vec_rsc_0_62_wadr;
  output [63:0] vec_rsc_0_62_d;
  output vec_rsc_0_62_we;
  output [3:0] vec_rsc_0_62_radr;
  input [63:0] vec_rsc_0_62_q;
  output vec_rsc_triosy_0_62_lz;
  output [3:0] vec_rsc_0_63_wadr;
  output [63:0] vec_rsc_0_63_d;
  output vec_rsc_0_63_we;
  output [3:0] vec_rsc_0_63_radr;
  input [63:0] vec_rsc_0_63_q;
  output vec_rsc_triosy_0_63_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [3:0] twiddle_rsc_0_0_radr;
  input [63:0] twiddle_rsc_0_0_q;
  output twiddle_rsc_triosy_0_0_lz;
  output [3:0] twiddle_rsc_0_1_radr;
  input [63:0] twiddle_rsc_0_1_q;
  output twiddle_rsc_triosy_0_1_lz;
  output [3:0] twiddle_rsc_0_2_radr;
  input [63:0] twiddle_rsc_0_2_q;
  output twiddle_rsc_triosy_0_2_lz;
  output [3:0] twiddle_rsc_0_3_radr;
  input [63:0] twiddle_rsc_0_3_q;
  output twiddle_rsc_triosy_0_3_lz;
  output [3:0] twiddle_rsc_0_4_radr;
  input [63:0] twiddle_rsc_0_4_q;
  output twiddle_rsc_triosy_0_4_lz;
  output [3:0] twiddle_rsc_0_5_radr;
  input [63:0] twiddle_rsc_0_5_q;
  output twiddle_rsc_triosy_0_5_lz;
  output [3:0] twiddle_rsc_0_6_radr;
  input [63:0] twiddle_rsc_0_6_q;
  output twiddle_rsc_triosy_0_6_lz;
  output [3:0] twiddle_rsc_0_7_radr;
  input [63:0] twiddle_rsc_0_7_q;
  output twiddle_rsc_triosy_0_7_lz;
  output [3:0] twiddle_rsc_0_8_radr;
  input [63:0] twiddle_rsc_0_8_q;
  output twiddle_rsc_triosy_0_8_lz;
  output [3:0] twiddle_rsc_0_9_radr;
  input [63:0] twiddle_rsc_0_9_q;
  output twiddle_rsc_triosy_0_9_lz;
  output [3:0] twiddle_rsc_0_10_radr;
  input [63:0] twiddle_rsc_0_10_q;
  output twiddle_rsc_triosy_0_10_lz;
  output [3:0] twiddle_rsc_0_11_radr;
  input [63:0] twiddle_rsc_0_11_q;
  output twiddle_rsc_triosy_0_11_lz;
  output [3:0] twiddle_rsc_0_12_radr;
  input [63:0] twiddle_rsc_0_12_q;
  output twiddle_rsc_triosy_0_12_lz;
  output [3:0] twiddle_rsc_0_13_radr;
  input [63:0] twiddle_rsc_0_13_q;
  output twiddle_rsc_triosy_0_13_lz;
  output [3:0] twiddle_rsc_0_14_radr;
  input [63:0] twiddle_rsc_0_14_q;
  output twiddle_rsc_triosy_0_14_lz;
  output [3:0] twiddle_rsc_0_15_radr;
  input [63:0] twiddle_rsc_0_15_q;
  output twiddle_rsc_triosy_0_15_lz;
  output [3:0] twiddle_rsc_0_16_radr;
  input [63:0] twiddle_rsc_0_16_q;
  output twiddle_rsc_triosy_0_16_lz;
  output [3:0] twiddle_rsc_0_17_radr;
  input [63:0] twiddle_rsc_0_17_q;
  output twiddle_rsc_triosy_0_17_lz;
  output [3:0] twiddle_rsc_0_18_radr;
  input [63:0] twiddle_rsc_0_18_q;
  output twiddle_rsc_triosy_0_18_lz;
  output [3:0] twiddle_rsc_0_19_radr;
  input [63:0] twiddle_rsc_0_19_q;
  output twiddle_rsc_triosy_0_19_lz;
  output [3:0] twiddle_rsc_0_20_radr;
  input [63:0] twiddle_rsc_0_20_q;
  output twiddle_rsc_triosy_0_20_lz;
  output [3:0] twiddle_rsc_0_21_radr;
  input [63:0] twiddle_rsc_0_21_q;
  output twiddle_rsc_triosy_0_21_lz;
  output [3:0] twiddle_rsc_0_22_radr;
  input [63:0] twiddle_rsc_0_22_q;
  output twiddle_rsc_triosy_0_22_lz;
  output [3:0] twiddle_rsc_0_23_radr;
  input [63:0] twiddle_rsc_0_23_q;
  output twiddle_rsc_triosy_0_23_lz;
  output [3:0] twiddle_rsc_0_24_radr;
  input [63:0] twiddle_rsc_0_24_q;
  output twiddle_rsc_triosy_0_24_lz;
  output [3:0] twiddle_rsc_0_25_radr;
  input [63:0] twiddle_rsc_0_25_q;
  output twiddle_rsc_triosy_0_25_lz;
  output [3:0] twiddle_rsc_0_26_radr;
  input [63:0] twiddle_rsc_0_26_q;
  output twiddle_rsc_triosy_0_26_lz;
  output [3:0] twiddle_rsc_0_27_radr;
  input [63:0] twiddle_rsc_0_27_q;
  output twiddle_rsc_triosy_0_27_lz;
  output [3:0] twiddle_rsc_0_28_radr;
  input [63:0] twiddle_rsc_0_28_q;
  output twiddle_rsc_triosy_0_28_lz;
  output [3:0] twiddle_rsc_0_29_radr;
  input [63:0] twiddle_rsc_0_29_q;
  output twiddle_rsc_triosy_0_29_lz;
  output [3:0] twiddle_rsc_0_30_radr;
  input [63:0] twiddle_rsc_0_30_q;
  output twiddle_rsc_triosy_0_30_lz;
  output [3:0] twiddle_rsc_0_31_radr;
  input [63:0] twiddle_rsc_0_31_q;
  output twiddle_rsc_triosy_0_31_lz;
  output [3:0] twiddle_rsc_0_32_radr;
  input [63:0] twiddle_rsc_0_32_q;
  output twiddle_rsc_triosy_0_32_lz;
  output [3:0] twiddle_rsc_0_33_radr;
  input [63:0] twiddle_rsc_0_33_q;
  output twiddle_rsc_triosy_0_33_lz;
  output [3:0] twiddle_rsc_0_34_radr;
  input [63:0] twiddle_rsc_0_34_q;
  output twiddle_rsc_triosy_0_34_lz;
  output [3:0] twiddle_rsc_0_35_radr;
  input [63:0] twiddle_rsc_0_35_q;
  output twiddle_rsc_triosy_0_35_lz;
  output [3:0] twiddle_rsc_0_36_radr;
  input [63:0] twiddle_rsc_0_36_q;
  output twiddle_rsc_triosy_0_36_lz;
  output [3:0] twiddle_rsc_0_37_radr;
  input [63:0] twiddle_rsc_0_37_q;
  output twiddle_rsc_triosy_0_37_lz;
  output [3:0] twiddle_rsc_0_38_radr;
  input [63:0] twiddle_rsc_0_38_q;
  output twiddle_rsc_triosy_0_38_lz;
  output [3:0] twiddle_rsc_0_39_radr;
  input [63:0] twiddle_rsc_0_39_q;
  output twiddle_rsc_triosy_0_39_lz;
  output [3:0] twiddle_rsc_0_40_radr;
  input [63:0] twiddle_rsc_0_40_q;
  output twiddle_rsc_triosy_0_40_lz;
  output [3:0] twiddle_rsc_0_41_radr;
  input [63:0] twiddle_rsc_0_41_q;
  output twiddle_rsc_triosy_0_41_lz;
  output [3:0] twiddle_rsc_0_42_radr;
  input [63:0] twiddle_rsc_0_42_q;
  output twiddle_rsc_triosy_0_42_lz;
  output [3:0] twiddle_rsc_0_43_radr;
  input [63:0] twiddle_rsc_0_43_q;
  output twiddle_rsc_triosy_0_43_lz;
  output [3:0] twiddle_rsc_0_44_radr;
  input [63:0] twiddle_rsc_0_44_q;
  output twiddle_rsc_triosy_0_44_lz;
  output [3:0] twiddle_rsc_0_45_radr;
  input [63:0] twiddle_rsc_0_45_q;
  output twiddle_rsc_triosy_0_45_lz;
  output [3:0] twiddle_rsc_0_46_radr;
  input [63:0] twiddle_rsc_0_46_q;
  output twiddle_rsc_triosy_0_46_lz;
  output [3:0] twiddle_rsc_0_47_radr;
  input [63:0] twiddle_rsc_0_47_q;
  output twiddle_rsc_triosy_0_47_lz;
  output [3:0] twiddle_rsc_0_48_radr;
  input [63:0] twiddle_rsc_0_48_q;
  output twiddle_rsc_triosy_0_48_lz;
  output [3:0] twiddle_rsc_0_49_radr;
  input [63:0] twiddle_rsc_0_49_q;
  output twiddle_rsc_triosy_0_49_lz;
  output [3:0] twiddle_rsc_0_50_radr;
  input [63:0] twiddle_rsc_0_50_q;
  output twiddle_rsc_triosy_0_50_lz;
  output [3:0] twiddle_rsc_0_51_radr;
  input [63:0] twiddle_rsc_0_51_q;
  output twiddle_rsc_triosy_0_51_lz;
  output [3:0] twiddle_rsc_0_52_radr;
  input [63:0] twiddle_rsc_0_52_q;
  output twiddle_rsc_triosy_0_52_lz;
  output [3:0] twiddle_rsc_0_53_radr;
  input [63:0] twiddle_rsc_0_53_q;
  output twiddle_rsc_triosy_0_53_lz;
  output [3:0] twiddle_rsc_0_54_radr;
  input [63:0] twiddle_rsc_0_54_q;
  output twiddle_rsc_triosy_0_54_lz;
  output [3:0] twiddle_rsc_0_55_radr;
  input [63:0] twiddle_rsc_0_55_q;
  output twiddle_rsc_triosy_0_55_lz;
  output [3:0] twiddle_rsc_0_56_radr;
  input [63:0] twiddle_rsc_0_56_q;
  output twiddle_rsc_triosy_0_56_lz;
  output [3:0] twiddle_rsc_0_57_radr;
  input [63:0] twiddle_rsc_0_57_q;
  output twiddle_rsc_triosy_0_57_lz;
  output [3:0] twiddle_rsc_0_58_radr;
  input [63:0] twiddle_rsc_0_58_q;
  output twiddle_rsc_triosy_0_58_lz;
  output [3:0] twiddle_rsc_0_59_radr;
  input [63:0] twiddle_rsc_0_59_q;
  output twiddle_rsc_triosy_0_59_lz;
  output [3:0] twiddle_rsc_0_60_radr;
  input [63:0] twiddle_rsc_0_60_q;
  output twiddle_rsc_triosy_0_60_lz;
  output [3:0] twiddle_rsc_0_61_radr;
  input [63:0] twiddle_rsc_0_61_q;
  output twiddle_rsc_triosy_0_61_lz;
  output [3:0] twiddle_rsc_0_62_radr;
  input [63:0] twiddle_rsc_0_62_q;
  output twiddle_rsc_triosy_0_62_lz;
  output [3:0] twiddle_rsc_0_63_radr;
  input [63:0] twiddle_rsc_0_63_q;
  output twiddle_rsc_triosy_0_63_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_q_d;
  wire vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_q_d;
  wire vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_q_d;
  wire vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_q_d;
  wire vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_q_d;
  wire vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_q_d;
  wire vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_q_d;
  wire vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_q_d;
  wire vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_q_d;
  wire vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_q_d;
  wire vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_q_d;
  wire vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_q_d;
  wire vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_q_d;
  wire vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_q_d;
  wire vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_q_d;
  wire vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_q_d;
  wire vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_16_i_q_d;
  wire vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_17_i_q_d;
  wire vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_18_i_q_d;
  wire vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_19_i_q_d;
  wire vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_20_i_q_d;
  wire vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_21_i_q_d;
  wire vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_22_i_q_d;
  wire vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_23_i_q_d;
  wire vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_24_i_q_d;
  wire vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_25_i_q_d;
  wire vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_26_i_q_d;
  wire vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_27_i_q_d;
  wire vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_28_i_q_d;
  wire vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_29_i_q_d;
  wire vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_30_i_q_d;
  wire vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_31_i_q_d;
  wire vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_32_i_q_d;
  wire vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_33_i_q_d;
  wire vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_34_i_q_d;
  wire vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_35_i_q_d;
  wire vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_36_i_q_d;
  wire vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_37_i_q_d;
  wire vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_38_i_q_d;
  wire vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_39_i_q_d;
  wire vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_40_i_q_d;
  wire vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_41_i_q_d;
  wire vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_42_i_q_d;
  wire vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_43_i_q_d;
  wire vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_44_i_q_d;
  wire vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_45_i_q_d;
  wire vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_46_i_q_d;
  wire vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_47_i_q_d;
  wire vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_48_i_q_d;
  wire vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_49_i_q_d;
  wire vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_50_i_q_d;
  wire vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_51_i_q_d;
  wire vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_52_i_q_d;
  wire vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_53_i_q_d;
  wire vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_54_i_q_d;
  wire vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_55_i_q_d;
  wire vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_56_i_q_d;
  wire vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_57_i_q_d;
  wire vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_58_i_q_d;
  wire vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_59_i_q_d;
  wire vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_60_i_q_d;
  wire vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_61_i_q_d;
  wire vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_62_i_q_d;
  wire vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_63_i_q_d;
  wire vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_0_i_q_d;
  wire twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_1_i_q_d;
  wire twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_2_i_q_d;
  wire twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_3_i_q_d;
  wire twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_4_i_q_d;
  wire twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_5_i_q_d;
  wire twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_6_i_q_d;
  wire twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_7_i_q_d;
  wire twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_8_i_q_d;
  wire twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_9_i_q_d;
  wire twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_10_i_q_d;
  wire twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_11_i_q_d;
  wire twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_12_i_q_d;
  wire twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_13_i_q_d;
  wire twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_14_i_q_d;
  wire twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_15_i_q_d;
  wire twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_16_i_q_d;
  wire twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_17_i_q_d;
  wire twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_18_i_q_d;
  wire twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_19_i_q_d;
  wire twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_20_i_q_d;
  wire twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_21_i_q_d;
  wire twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_22_i_q_d;
  wire twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_23_i_q_d;
  wire twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_24_i_q_d;
  wire twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_25_i_q_d;
  wire twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_26_i_q_d;
  wire twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_27_i_q_d;
  wire twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_28_i_q_d;
  wire twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_29_i_q_d;
  wire twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_30_i_q_d;
  wire twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_31_i_q_d;
  wire twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_32_i_q_d;
  wire twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_33_i_q_d;
  wire twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_34_i_q_d;
  wire twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_35_i_q_d;
  wire twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_36_i_q_d;
  wire twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_37_i_q_d;
  wire twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_38_i_q_d;
  wire twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_39_i_q_d;
  wire twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_40_i_q_d;
  wire twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_41_i_q_d;
  wire twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_42_i_q_d;
  wire twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_43_i_q_d;
  wire twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_44_i_q_d;
  wire twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_45_i_q_d;
  wire twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_46_i_q_d;
  wire twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_47_i_q_d;
  wire twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_48_i_q_d;
  wire twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_49_i_q_d;
  wire twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_50_i_q_d;
  wire twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_51_i_q_d;
  wire twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_52_i_q_d;
  wire twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_53_i_q_d;
  wire twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_54_i_q_d;
  wire twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_55_i_q_d;
  wire twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_56_i_q_d;
  wire twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_57_i_q_d;
  wire twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_58_i_q_d;
  wire twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_59_i_q_d;
  wire twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_60_i_q_d;
  wire twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_61_i_q_d;
  wire twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_62_i_q_d;
  wire twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] twiddle_rsc_0_63_i_q_d;
  wire twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_0_i_d_d_iff;
  wire [3:0] vec_rsc_0_0_i_radr_d_iff;
  wire [3:0] vec_rsc_0_0_i_wadr_d_iff;
  wire vec_rsc_0_0_i_we_d_iff;
  wire vec_rsc_0_1_i_we_d_iff;
  wire vec_rsc_0_2_i_we_d_iff;
  wire vec_rsc_0_3_i_we_d_iff;
  wire vec_rsc_0_4_i_we_d_iff;
  wire vec_rsc_0_5_i_we_d_iff;
  wire vec_rsc_0_6_i_we_d_iff;
  wire vec_rsc_0_7_i_we_d_iff;
  wire vec_rsc_0_8_i_we_d_iff;
  wire vec_rsc_0_9_i_we_d_iff;
  wire vec_rsc_0_10_i_we_d_iff;
  wire vec_rsc_0_11_i_we_d_iff;
  wire vec_rsc_0_12_i_we_d_iff;
  wire vec_rsc_0_13_i_we_d_iff;
  wire vec_rsc_0_14_i_we_d_iff;
  wire vec_rsc_0_15_i_we_d_iff;
  wire vec_rsc_0_16_i_we_d_iff;
  wire vec_rsc_0_17_i_we_d_iff;
  wire vec_rsc_0_18_i_we_d_iff;
  wire vec_rsc_0_19_i_we_d_iff;
  wire vec_rsc_0_20_i_we_d_iff;
  wire vec_rsc_0_21_i_we_d_iff;
  wire vec_rsc_0_22_i_we_d_iff;
  wire vec_rsc_0_23_i_we_d_iff;
  wire vec_rsc_0_24_i_we_d_iff;
  wire vec_rsc_0_25_i_we_d_iff;
  wire vec_rsc_0_26_i_we_d_iff;
  wire vec_rsc_0_27_i_we_d_iff;
  wire vec_rsc_0_28_i_we_d_iff;
  wire vec_rsc_0_29_i_we_d_iff;
  wire vec_rsc_0_30_i_we_d_iff;
  wire vec_rsc_0_31_i_we_d_iff;
  wire vec_rsc_0_32_i_we_d_iff;
  wire vec_rsc_0_33_i_we_d_iff;
  wire vec_rsc_0_34_i_we_d_iff;
  wire vec_rsc_0_35_i_we_d_iff;
  wire vec_rsc_0_36_i_we_d_iff;
  wire vec_rsc_0_37_i_we_d_iff;
  wire vec_rsc_0_38_i_we_d_iff;
  wire vec_rsc_0_39_i_we_d_iff;
  wire vec_rsc_0_40_i_we_d_iff;
  wire vec_rsc_0_41_i_we_d_iff;
  wire vec_rsc_0_42_i_we_d_iff;
  wire vec_rsc_0_43_i_we_d_iff;
  wire vec_rsc_0_44_i_we_d_iff;
  wire vec_rsc_0_45_i_we_d_iff;
  wire vec_rsc_0_46_i_we_d_iff;
  wire vec_rsc_0_47_i_we_d_iff;
  wire vec_rsc_0_48_i_we_d_iff;
  wire vec_rsc_0_49_i_we_d_iff;
  wire vec_rsc_0_50_i_we_d_iff;
  wire vec_rsc_0_51_i_we_d_iff;
  wire vec_rsc_0_52_i_we_d_iff;
  wire vec_rsc_0_53_i_we_d_iff;
  wire vec_rsc_0_54_i_we_d_iff;
  wire vec_rsc_0_55_i_we_d_iff;
  wire vec_rsc_0_56_i_we_d_iff;
  wire vec_rsc_0_57_i_we_d_iff;
  wire vec_rsc_0_58_i_we_d_iff;
  wire vec_rsc_0_59_i_we_d_iff;
  wire vec_rsc_0_60_i_we_d_iff;
  wire vec_rsc_0_61_i_we_d_iff;
  wire vec_rsc_0_62_i_we_d_iff;
  wire vec_rsc_0_63_i_we_d_iff;
  wire [3:0] twiddle_rsc_0_0_i_radr_d_iff;
  wire [3:0] twiddle_rsc_0_1_i_radr_d_iff;
  wire [3:0] twiddle_rsc_0_2_i_radr_d_iff;
  wire [3:0] twiddle_rsc_0_4_i_radr_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_9_4_64_16_16_64_1_gen vec_rsc_0_0_i
      (
      .q(vec_rsc_0_0_q),
      .radr(vec_rsc_0_0_radr),
      .we(vec_rsc_0_0_we),
      .d(vec_rsc_0_0_d),
      .wadr(vec_rsc_0_0_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_0_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_0_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_10_4_64_16_16_64_1_gen vec_rsc_0_1_i
      (
      .q(vec_rsc_0_1_q),
      .radr(vec_rsc_0_1_radr),
      .we(vec_rsc_0_1_we),
      .d(vec_rsc_0_1_d),
      .wadr(vec_rsc_0_1_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_1_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_1_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_11_4_64_16_16_64_1_gen vec_rsc_0_2_i
      (
      .q(vec_rsc_0_2_q),
      .radr(vec_rsc_0_2_radr),
      .we(vec_rsc_0_2_we),
      .d(vec_rsc_0_2_d),
      .wadr(vec_rsc_0_2_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_2_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_2_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_12_4_64_16_16_64_1_gen vec_rsc_0_3_i
      (
      .q(vec_rsc_0_3_q),
      .radr(vec_rsc_0_3_radr),
      .we(vec_rsc_0_3_we),
      .d(vec_rsc_0_3_d),
      .wadr(vec_rsc_0_3_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_3_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_3_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_13_4_64_16_16_64_1_gen vec_rsc_0_4_i
      (
      .q(vec_rsc_0_4_q),
      .radr(vec_rsc_0_4_radr),
      .we(vec_rsc_0_4_we),
      .d(vec_rsc_0_4_d),
      .wadr(vec_rsc_0_4_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_4_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_4_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_14_4_64_16_16_64_1_gen vec_rsc_0_5_i
      (
      .q(vec_rsc_0_5_q),
      .radr(vec_rsc_0_5_radr),
      .we(vec_rsc_0_5_we),
      .d(vec_rsc_0_5_d),
      .wadr(vec_rsc_0_5_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_5_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_5_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_15_4_64_16_16_64_1_gen vec_rsc_0_6_i
      (
      .q(vec_rsc_0_6_q),
      .radr(vec_rsc_0_6_radr),
      .we(vec_rsc_0_6_we),
      .d(vec_rsc_0_6_d),
      .wadr(vec_rsc_0_6_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_6_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_6_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_16_4_64_16_16_64_1_gen vec_rsc_0_7_i
      (
      .q(vec_rsc_0_7_q),
      .radr(vec_rsc_0_7_radr),
      .we(vec_rsc_0_7_we),
      .d(vec_rsc_0_7_d),
      .wadr(vec_rsc_0_7_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_7_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_7_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_17_4_64_16_16_64_1_gen vec_rsc_0_8_i
      (
      .q(vec_rsc_0_8_q),
      .radr(vec_rsc_0_8_radr),
      .we(vec_rsc_0_8_we),
      .d(vec_rsc_0_8_d),
      .wadr(vec_rsc_0_8_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_8_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_8_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_18_4_64_16_16_64_1_gen vec_rsc_0_9_i
      (
      .q(vec_rsc_0_9_q),
      .radr(vec_rsc_0_9_radr),
      .we(vec_rsc_0_9_we),
      .d(vec_rsc_0_9_d),
      .wadr(vec_rsc_0_9_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_9_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_9_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_19_4_64_16_16_64_1_gen vec_rsc_0_10_i
      (
      .q(vec_rsc_0_10_q),
      .radr(vec_rsc_0_10_radr),
      .we(vec_rsc_0_10_we),
      .d(vec_rsc_0_10_d),
      .wadr(vec_rsc_0_10_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_10_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_10_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_20_4_64_16_16_64_1_gen vec_rsc_0_11_i
      (
      .q(vec_rsc_0_11_q),
      .radr(vec_rsc_0_11_radr),
      .we(vec_rsc_0_11_we),
      .d(vec_rsc_0_11_d),
      .wadr(vec_rsc_0_11_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_11_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_11_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_21_4_64_16_16_64_1_gen vec_rsc_0_12_i
      (
      .q(vec_rsc_0_12_q),
      .radr(vec_rsc_0_12_radr),
      .we(vec_rsc_0_12_we),
      .d(vec_rsc_0_12_d),
      .wadr(vec_rsc_0_12_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_12_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_12_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_22_4_64_16_16_64_1_gen vec_rsc_0_13_i
      (
      .q(vec_rsc_0_13_q),
      .radr(vec_rsc_0_13_radr),
      .we(vec_rsc_0_13_we),
      .d(vec_rsc_0_13_d),
      .wadr(vec_rsc_0_13_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_13_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_13_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_23_4_64_16_16_64_1_gen vec_rsc_0_14_i
      (
      .q(vec_rsc_0_14_q),
      .radr(vec_rsc_0_14_radr),
      .we(vec_rsc_0_14_we),
      .d(vec_rsc_0_14_d),
      .wadr(vec_rsc_0_14_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_14_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_14_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_24_4_64_16_16_64_1_gen vec_rsc_0_15_i
      (
      .q(vec_rsc_0_15_q),
      .radr(vec_rsc_0_15_radr),
      .we(vec_rsc_0_15_we),
      .d(vec_rsc_0_15_d),
      .wadr(vec_rsc_0_15_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_15_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_15_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_25_4_64_16_16_64_1_gen vec_rsc_0_16_i
      (
      .q(vec_rsc_0_16_q),
      .radr(vec_rsc_0_16_radr),
      .we(vec_rsc_0_16_we),
      .d(vec_rsc_0_16_d),
      .wadr(vec_rsc_0_16_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_16_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_16_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_16_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_26_4_64_16_16_64_1_gen vec_rsc_0_17_i
      (
      .q(vec_rsc_0_17_q),
      .radr(vec_rsc_0_17_radr),
      .we(vec_rsc_0_17_we),
      .d(vec_rsc_0_17_d),
      .wadr(vec_rsc_0_17_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_17_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_17_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_17_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_27_4_64_16_16_64_1_gen vec_rsc_0_18_i
      (
      .q(vec_rsc_0_18_q),
      .radr(vec_rsc_0_18_radr),
      .we(vec_rsc_0_18_we),
      .d(vec_rsc_0_18_d),
      .wadr(vec_rsc_0_18_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_18_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_18_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_18_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_28_4_64_16_16_64_1_gen vec_rsc_0_19_i
      (
      .q(vec_rsc_0_19_q),
      .radr(vec_rsc_0_19_radr),
      .we(vec_rsc_0_19_we),
      .d(vec_rsc_0_19_d),
      .wadr(vec_rsc_0_19_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_19_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_19_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_19_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_29_4_64_16_16_64_1_gen vec_rsc_0_20_i
      (
      .q(vec_rsc_0_20_q),
      .radr(vec_rsc_0_20_radr),
      .we(vec_rsc_0_20_we),
      .d(vec_rsc_0_20_d),
      .wadr(vec_rsc_0_20_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_20_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_20_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_20_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_30_4_64_16_16_64_1_gen vec_rsc_0_21_i
      (
      .q(vec_rsc_0_21_q),
      .radr(vec_rsc_0_21_radr),
      .we(vec_rsc_0_21_we),
      .d(vec_rsc_0_21_d),
      .wadr(vec_rsc_0_21_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_21_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_21_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_21_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_31_4_64_16_16_64_1_gen vec_rsc_0_22_i
      (
      .q(vec_rsc_0_22_q),
      .radr(vec_rsc_0_22_radr),
      .we(vec_rsc_0_22_we),
      .d(vec_rsc_0_22_d),
      .wadr(vec_rsc_0_22_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_22_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_22_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_22_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_32_4_64_16_16_64_1_gen vec_rsc_0_23_i
      (
      .q(vec_rsc_0_23_q),
      .radr(vec_rsc_0_23_radr),
      .we(vec_rsc_0_23_we),
      .d(vec_rsc_0_23_d),
      .wadr(vec_rsc_0_23_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_23_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_23_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_23_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_33_4_64_16_16_64_1_gen vec_rsc_0_24_i
      (
      .q(vec_rsc_0_24_q),
      .radr(vec_rsc_0_24_radr),
      .we(vec_rsc_0_24_we),
      .d(vec_rsc_0_24_d),
      .wadr(vec_rsc_0_24_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_24_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_24_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_24_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_34_4_64_16_16_64_1_gen vec_rsc_0_25_i
      (
      .q(vec_rsc_0_25_q),
      .radr(vec_rsc_0_25_radr),
      .we(vec_rsc_0_25_we),
      .d(vec_rsc_0_25_d),
      .wadr(vec_rsc_0_25_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_25_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_25_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_25_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_35_4_64_16_16_64_1_gen vec_rsc_0_26_i
      (
      .q(vec_rsc_0_26_q),
      .radr(vec_rsc_0_26_radr),
      .we(vec_rsc_0_26_we),
      .d(vec_rsc_0_26_d),
      .wadr(vec_rsc_0_26_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_26_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_26_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_26_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_36_4_64_16_16_64_1_gen vec_rsc_0_27_i
      (
      .q(vec_rsc_0_27_q),
      .radr(vec_rsc_0_27_radr),
      .we(vec_rsc_0_27_we),
      .d(vec_rsc_0_27_d),
      .wadr(vec_rsc_0_27_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_27_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_27_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_27_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_37_4_64_16_16_64_1_gen vec_rsc_0_28_i
      (
      .q(vec_rsc_0_28_q),
      .radr(vec_rsc_0_28_radr),
      .we(vec_rsc_0_28_we),
      .d(vec_rsc_0_28_d),
      .wadr(vec_rsc_0_28_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_28_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_28_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_28_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_38_4_64_16_16_64_1_gen vec_rsc_0_29_i
      (
      .q(vec_rsc_0_29_q),
      .radr(vec_rsc_0_29_radr),
      .we(vec_rsc_0_29_we),
      .d(vec_rsc_0_29_d),
      .wadr(vec_rsc_0_29_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_29_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_29_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_29_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_39_4_64_16_16_64_1_gen vec_rsc_0_30_i
      (
      .q(vec_rsc_0_30_q),
      .radr(vec_rsc_0_30_radr),
      .we(vec_rsc_0_30_we),
      .d(vec_rsc_0_30_d),
      .wadr(vec_rsc_0_30_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_30_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_30_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_30_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_40_4_64_16_16_64_1_gen vec_rsc_0_31_i
      (
      .q(vec_rsc_0_31_q),
      .radr(vec_rsc_0_31_radr),
      .we(vec_rsc_0_31_we),
      .d(vec_rsc_0_31_d),
      .wadr(vec_rsc_0_31_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_31_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_31_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_31_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_41_4_64_16_16_64_1_gen vec_rsc_0_32_i
      (
      .q(vec_rsc_0_32_q),
      .radr(vec_rsc_0_32_radr),
      .we(vec_rsc_0_32_we),
      .d(vec_rsc_0_32_d),
      .wadr(vec_rsc_0_32_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_32_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_32_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_32_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_42_4_64_16_16_64_1_gen vec_rsc_0_33_i
      (
      .q(vec_rsc_0_33_q),
      .radr(vec_rsc_0_33_radr),
      .we(vec_rsc_0_33_we),
      .d(vec_rsc_0_33_d),
      .wadr(vec_rsc_0_33_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_33_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_33_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_33_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_43_4_64_16_16_64_1_gen vec_rsc_0_34_i
      (
      .q(vec_rsc_0_34_q),
      .radr(vec_rsc_0_34_radr),
      .we(vec_rsc_0_34_we),
      .d(vec_rsc_0_34_d),
      .wadr(vec_rsc_0_34_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_34_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_34_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_34_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_44_4_64_16_16_64_1_gen vec_rsc_0_35_i
      (
      .q(vec_rsc_0_35_q),
      .radr(vec_rsc_0_35_radr),
      .we(vec_rsc_0_35_we),
      .d(vec_rsc_0_35_d),
      .wadr(vec_rsc_0_35_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_35_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_35_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_35_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_45_4_64_16_16_64_1_gen vec_rsc_0_36_i
      (
      .q(vec_rsc_0_36_q),
      .radr(vec_rsc_0_36_radr),
      .we(vec_rsc_0_36_we),
      .d(vec_rsc_0_36_d),
      .wadr(vec_rsc_0_36_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_36_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_36_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_36_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_46_4_64_16_16_64_1_gen vec_rsc_0_37_i
      (
      .q(vec_rsc_0_37_q),
      .radr(vec_rsc_0_37_radr),
      .we(vec_rsc_0_37_we),
      .d(vec_rsc_0_37_d),
      .wadr(vec_rsc_0_37_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_37_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_37_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_37_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_47_4_64_16_16_64_1_gen vec_rsc_0_38_i
      (
      .q(vec_rsc_0_38_q),
      .radr(vec_rsc_0_38_radr),
      .we(vec_rsc_0_38_we),
      .d(vec_rsc_0_38_d),
      .wadr(vec_rsc_0_38_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_38_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_38_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_38_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_48_4_64_16_16_64_1_gen vec_rsc_0_39_i
      (
      .q(vec_rsc_0_39_q),
      .radr(vec_rsc_0_39_radr),
      .we(vec_rsc_0_39_we),
      .d(vec_rsc_0_39_d),
      .wadr(vec_rsc_0_39_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_39_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_39_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_39_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_49_4_64_16_16_64_1_gen vec_rsc_0_40_i
      (
      .q(vec_rsc_0_40_q),
      .radr(vec_rsc_0_40_radr),
      .we(vec_rsc_0_40_we),
      .d(vec_rsc_0_40_d),
      .wadr(vec_rsc_0_40_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_40_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_40_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_40_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_50_4_64_16_16_64_1_gen vec_rsc_0_41_i
      (
      .q(vec_rsc_0_41_q),
      .radr(vec_rsc_0_41_radr),
      .we(vec_rsc_0_41_we),
      .d(vec_rsc_0_41_d),
      .wadr(vec_rsc_0_41_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_41_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_41_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_41_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_51_4_64_16_16_64_1_gen vec_rsc_0_42_i
      (
      .q(vec_rsc_0_42_q),
      .radr(vec_rsc_0_42_radr),
      .we(vec_rsc_0_42_we),
      .d(vec_rsc_0_42_d),
      .wadr(vec_rsc_0_42_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_42_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_42_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_42_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_52_4_64_16_16_64_1_gen vec_rsc_0_43_i
      (
      .q(vec_rsc_0_43_q),
      .radr(vec_rsc_0_43_radr),
      .we(vec_rsc_0_43_we),
      .d(vec_rsc_0_43_d),
      .wadr(vec_rsc_0_43_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_43_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_43_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_43_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_53_4_64_16_16_64_1_gen vec_rsc_0_44_i
      (
      .q(vec_rsc_0_44_q),
      .radr(vec_rsc_0_44_radr),
      .we(vec_rsc_0_44_we),
      .d(vec_rsc_0_44_d),
      .wadr(vec_rsc_0_44_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_44_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_44_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_44_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_54_4_64_16_16_64_1_gen vec_rsc_0_45_i
      (
      .q(vec_rsc_0_45_q),
      .radr(vec_rsc_0_45_radr),
      .we(vec_rsc_0_45_we),
      .d(vec_rsc_0_45_d),
      .wadr(vec_rsc_0_45_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_45_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_45_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_45_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_55_4_64_16_16_64_1_gen vec_rsc_0_46_i
      (
      .q(vec_rsc_0_46_q),
      .radr(vec_rsc_0_46_radr),
      .we(vec_rsc_0_46_we),
      .d(vec_rsc_0_46_d),
      .wadr(vec_rsc_0_46_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_46_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_46_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_46_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_56_4_64_16_16_64_1_gen vec_rsc_0_47_i
      (
      .q(vec_rsc_0_47_q),
      .radr(vec_rsc_0_47_radr),
      .we(vec_rsc_0_47_we),
      .d(vec_rsc_0_47_d),
      .wadr(vec_rsc_0_47_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_47_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_47_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_47_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_57_4_64_16_16_64_1_gen vec_rsc_0_48_i
      (
      .q(vec_rsc_0_48_q),
      .radr(vec_rsc_0_48_radr),
      .we(vec_rsc_0_48_we),
      .d(vec_rsc_0_48_d),
      .wadr(vec_rsc_0_48_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_48_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_48_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_48_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_58_4_64_16_16_64_1_gen vec_rsc_0_49_i
      (
      .q(vec_rsc_0_49_q),
      .radr(vec_rsc_0_49_radr),
      .we(vec_rsc_0_49_we),
      .d(vec_rsc_0_49_d),
      .wadr(vec_rsc_0_49_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_49_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_49_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_49_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_59_4_64_16_16_64_1_gen vec_rsc_0_50_i
      (
      .q(vec_rsc_0_50_q),
      .radr(vec_rsc_0_50_radr),
      .we(vec_rsc_0_50_we),
      .d(vec_rsc_0_50_d),
      .wadr(vec_rsc_0_50_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_50_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_50_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_50_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_60_4_64_16_16_64_1_gen vec_rsc_0_51_i
      (
      .q(vec_rsc_0_51_q),
      .radr(vec_rsc_0_51_radr),
      .we(vec_rsc_0_51_we),
      .d(vec_rsc_0_51_d),
      .wadr(vec_rsc_0_51_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_51_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_51_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_51_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_61_4_64_16_16_64_1_gen vec_rsc_0_52_i
      (
      .q(vec_rsc_0_52_q),
      .radr(vec_rsc_0_52_radr),
      .we(vec_rsc_0_52_we),
      .d(vec_rsc_0_52_d),
      .wadr(vec_rsc_0_52_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_52_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_52_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_52_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_62_4_64_16_16_64_1_gen vec_rsc_0_53_i
      (
      .q(vec_rsc_0_53_q),
      .radr(vec_rsc_0_53_radr),
      .we(vec_rsc_0_53_we),
      .d(vec_rsc_0_53_d),
      .wadr(vec_rsc_0_53_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_53_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_53_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_53_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_63_4_64_16_16_64_1_gen vec_rsc_0_54_i
      (
      .q(vec_rsc_0_54_q),
      .radr(vec_rsc_0_54_radr),
      .we(vec_rsc_0_54_we),
      .d(vec_rsc_0_54_d),
      .wadr(vec_rsc_0_54_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_54_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_54_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_54_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_64_4_64_16_16_64_1_gen vec_rsc_0_55_i
      (
      .q(vec_rsc_0_55_q),
      .radr(vec_rsc_0_55_radr),
      .we(vec_rsc_0_55_we),
      .d(vec_rsc_0_55_d),
      .wadr(vec_rsc_0_55_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_55_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_55_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_55_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_65_4_64_16_16_64_1_gen vec_rsc_0_56_i
      (
      .q(vec_rsc_0_56_q),
      .radr(vec_rsc_0_56_radr),
      .we(vec_rsc_0_56_we),
      .d(vec_rsc_0_56_d),
      .wadr(vec_rsc_0_56_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_56_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_56_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_56_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_66_4_64_16_16_64_1_gen vec_rsc_0_57_i
      (
      .q(vec_rsc_0_57_q),
      .radr(vec_rsc_0_57_radr),
      .we(vec_rsc_0_57_we),
      .d(vec_rsc_0_57_d),
      .wadr(vec_rsc_0_57_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_57_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_57_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_57_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_67_4_64_16_16_64_1_gen vec_rsc_0_58_i
      (
      .q(vec_rsc_0_58_q),
      .radr(vec_rsc_0_58_radr),
      .we(vec_rsc_0_58_we),
      .d(vec_rsc_0_58_d),
      .wadr(vec_rsc_0_58_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_58_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_58_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_58_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_68_4_64_16_16_64_1_gen vec_rsc_0_59_i
      (
      .q(vec_rsc_0_59_q),
      .radr(vec_rsc_0_59_radr),
      .we(vec_rsc_0_59_we),
      .d(vec_rsc_0_59_d),
      .wadr(vec_rsc_0_59_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_59_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_59_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_59_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_69_4_64_16_16_64_1_gen vec_rsc_0_60_i
      (
      .q(vec_rsc_0_60_q),
      .radr(vec_rsc_0_60_radr),
      .we(vec_rsc_0_60_we),
      .d(vec_rsc_0_60_d),
      .wadr(vec_rsc_0_60_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_60_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_60_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_60_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_70_4_64_16_16_64_1_gen vec_rsc_0_61_i
      (
      .q(vec_rsc_0_61_q),
      .radr(vec_rsc_0_61_radr),
      .we(vec_rsc_0_61_we),
      .d(vec_rsc_0_61_d),
      .wadr(vec_rsc_0_61_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_61_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_61_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_61_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_71_4_64_16_16_64_1_gen vec_rsc_0_62_i
      (
      .q(vec_rsc_0_62_q),
      .radr(vec_rsc_0_62_radr),
      .we(vec_rsc_0_62_we),
      .d(vec_rsc_0_62_d),
      .wadr(vec_rsc_0_62_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_62_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_62_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_62_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rwport_72_4_64_16_16_64_1_gen vec_rsc_0_63_i
      (
      .q(vec_rsc_0_63_q),
      .radr(vec_rsc_0_63_radr),
      .we(vec_rsc_0_63_we),
      .d(vec_rsc_0_63_d),
      .wadr(vec_rsc_0_63_wadr),
      .d_d(vec_rsc_0_0_i_d_d_iff),
      .q_d(vec_rsc_0_63_i_q_d),
      .radr_d(vec_rsc_0_0_i_radr_d_iff),
      .wadr_d(vec_rsc_0_0_i_wadr_d_iff),
      .we_d(vec_rsc_0_63_i_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(vec_rsc_0_63_i_we_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_73_4_64_16_16_64_1_gen twiddle_rsc_0_0_i
      (
      .q(twiddle_rsc_0_0_q),
      .radr(twiddle_rsc_0_0_radr),
      .q_d(twiddle_rsc_0_0_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_74_4_64_16_16_64_1_gen twiddle_rsc_0_1_i
      (
      .q(twiddle_rsc_0_1_q),
      .radr(twiddle_rsc_0_1_radr),
      .q_d(twiddle_rsc_0_1_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_75_4_64_16_16_64_1_gen twiddle_rsc_0_2_i
      (
      .q(twiddle_rsc_0_2_q),
      .radr(twiddle_rsc_0_2_radr),
      .q_d(twiddle_rsc_0_2_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_76_4_64_16_16_64_1_gen twiddle_rsc_0_3_i
      (
      .q(twiddle_rsc_0_3_q),
      .radr(twiddle_rsc_0_3_radr),
      .q_d(twiddle_rsc_0_3_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_77_4_64_16_16_64_1_gen twiddle_rsc_0_4_i
      (
      .q(twiddle_rsc_0_4_q),
      .radr(twiddle_rsc_0_4_radr),
      .q_d(twiddle_rsc_0_4_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_78_4_64_16_16_64_1_gen twiddle_rsc_0_5_i
      (
      .q(twiddle_rsc_0_5_q),
      .radr(twiddle_rsc_0_5_radr),
      .q_d(twiddle_rsc_0_5_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_79_4_64_16_16_64_1_gen twiddle_rsc_0_6_i
      (
      .q(twiddle_rsc_0_6_q),
      .radr(twiddle_rsc_0_6_radr),
      .q_d(twiddle_rsc_0_6_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_80_4_64_16_16_64_1_gen twiddle_rsc_0_7_i
      (
      .q(twiddle_rsc_0_7_q),
      .radr(twiddle_rsc_0_7_radr),
      .q_d(twiddle_rsc_0_7_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_81_4_64_16_16_64_1_gen twiddle_rsc_0_8_i
      (
      .q(twiddle_rsc_0_8_q),
      .radr(twiddle_rsc_0_8_radr),
      .q_d(twiddle_rsc_0_8_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_82_4_64_16_16_64_1_gen twiddle_rsc_0_9_i
      (
      .q(twiddle_rsc_0_9_q),
      .radr(twiddle_rsc_0_9_radr),
      .q_d(twiddle_rsc_0_9_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_83_4_64_16_16_64_1_gen twiddle_rsc_0_10_i
      (
      .q(twiddle_rsc_0_10_q),
      .radr(twiddle_rsc_0_10_radr),
      .q_d(twiddle_rsc_0_10_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_84_4_64_16_16_64_1_gen twiddle_rsc_0_11_i
      (
      .q(twiddle_rsc_0_11_q),
      .radr(twiddle_rsc_0_11_radr),
      .q_d(twiddle_rsc_0_11_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_85_4_64_16_16_64_1_gen twiddle_rsc_0_12_i
      (
      .q(twiddle_rsc_0_12_q),
      .radr(twiddle_rsc_0_12_radr),
      .q_d(twiddle_rsc_0_12_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_86_4_64_16_16_64_1_gen twiddle_rsc_0_13_i
      (
      .q(twiddle_rsc_0_13_q),
      .radr(twiddle_rsc_0_13_radr),
      .q_d(twiddle_rsc_0_13_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_87_4_64_16_16_64_1_gen twiddle_rsc_0_14_i
      (
      .q(twiddle_rsc_0_14_q),
      .radr(twiddle_rsc_0_14_radr),
      .q_d(twiddle_rsc_0_14_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_88_4_64_16_16_64_1_gen twiddle_rsc_0_15_i
      (
      .q(twiddle_rsc_0_15_q),
      .radr(twiddle_rsc_0_15_radr),
      .q_d(twiddle_rsc_0_15_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_89_4_64_16_16_64_1_gen twiddle_rsc_0_16_i
      (
      .q(twiddle_rsc_0_16_q),
      .radr(twiddle_rsc_0_16_radr),
      .q_d(twiddle_rsc_0_16_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_90_4_64_16_16_64_1_gen twiddle_rsc_0_17_i
      (
      .q(twiddle_rsc_0_17_q),
      .radr(twiddle_rsc_0_17_radr),
      .q_d(twiddle_rsc_0_17_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_91_4_64_16_16_64_1_gen twiddle_rsc_0_18_i
      (
      .q(twiddle_rsc_0_18_q),
      .radr(twiddle_rsc_0_18_radr),
      .q_d(twiddle_rsc_0_18_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_92_4_64_16_16_64_1_gen twiddle_rsc_0_19_i
      (
      .q(twiddle_rsc_0_19_q),
      .radr(twiddle_rsc_0_19_radr),
      .q_d(twiddle_rsc_0_19_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_93_4_64_16_16_64_1_gen twiddle_rsc_0_20_i
      (
      .q(twiddle_rsc_0_20_q),
      .radr(twiddle_rsc_0_20_radr),
      .q_d(twiddle_rsc_0_20_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_94_4_64_16_16_64_1_gen twiddle_rsc_0_21_i
      (
      .q(twiddle_rsc_0_21_q),
      .radr(twiddle_rsc_0_21_radr),
      .q_d(twiddle_rsc_0_21_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_95_4_64_16_16_64_1_gen twiddle_rsc_0_22_i
      (
      .q(twiddle_rsc_0_22_q),
      .radr(twiddle_rsc_0_22_radr),
      .q_d(twiddle_rsc_0_22_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_96_4_64_16_16_64_1_gen twiddle_rsc_0_23_i
      (
      .q(twiddle_rsc_0_23_q),
      .radr(twiddle_rsc_0_23_radr),
      .q_d(twiddle_rsc_0_23_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_97_4_64_16_16_64_1_gen twiddle_rsc_0_24_i
      (
      .q(twiddle_rsc_0_24_q),
      .radr(twiddle_rsc_0_24_radr),
      .q_d(twiddle_rsc_0_24_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_98_4_64_16_16_64_1_gen twiddle_rsc_0_25_i
      (
      .q(twiddle_rsc_0_25_q),
      .radr(twiddle_rsc_0_25_radr),
      .q_d(twiddle_rsc_0_25_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_99_4_64_16_16_64_1_gen twiddle_rsc_0_26_i
      (
      .q(twiddle_rsc_0_26_q),
      .radr(twiddle_rsc_0_26_radr),
      .q_d(twiddle_rsc_0_26_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_100_4_64_16_16_64_1_gen twiddle_rsc_0_27_i
      (
      .q(twiddle_rsc_0_27_q),
      .radr(twiddle_rsc_0_27_radr),
      .q_d(twiddle_rsc_0_27_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_101_4_64_16_16_64_1_gen twiddle_rsc_0_28_i
      (
      .q(twiddle_rsc_0_28_q),
      .radr(twiddle_rsc_0_28_radr),
      .q_d(twiddle_rsc_0_28_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_102_4_64_16_16_64_1_gen twiddle_rsc_0_29_i
      (
      .q(twiddle_rsc_0_29_q),
      .radr(twiddle_rsc_0_29_radr),
      .q_d(twiddle_rsc_0_29_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_103_4_64_16_16_64_1_gen twiddle_rsc_0_30_i
      (
      .q(twiddle_rsc_0_30_q),
      .radr(twiddle_rsc_0_30_radr),
      .q_d(twiddle_rsc_0_30_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_104_4_64_16_16_64_1_gen twiddle_rsc_0_31_i
      (
      .q(twiddle_rsc_0_31_q),
      .radr(twiddle_rsc_0_31_radr),
      .q_d(twiddle_rsc_0_31_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_105_4_64_16_16_64_1_gen twiddle_rsc_0_32_i
      (
      .q(twiddle_rsc_0_32_q),
      .radr(twiddle_rsc_0_32_radr),
      .q_d(twiddle_rsc_0_32_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_106_4_64_16_16_64_1_gen twiddle_rsc_0_33_i
      (
      .q(twiddle_rsc_0_33_q),
      .radr(twiddle_rsc_0_33_radr),
      .q_d(twiddle_rsc_0_33_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_107_4_64_16_16_64_1_gen twiddle_rsc_0_34_i
      (
      .q(twiddle_rsc_0_34_q),
      .radr(twiddle_rsc_0_34_radr),
      .q_d(twiddle_rsc_0_34_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_108_4_64_16_16_64_1_gen twiddle_rsc_0_35_i
      (
      .q(twiddle_rsc_0_35_q),
      .radr(twiddle_rsc_0_35_radr),
      .q_d(twiddle_rsc_0_35_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_109_4_64_16_16_64_1_gen twiddle_rsc_0_36_i
      (
      .q(twiddle_rsc_0_36_q),
      .radr(twiddle_rsc_0_36_radr),
      .q_d(twiddle_rsc_0_36_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_110_4_64_16_16_64_1_gen twiddle_rsc_0_37_i
      (
      .q(twiddle_rsc_0_37_q),
      .radr(twiddle_rsc_0_37_radr),
      .q_d(twiddle_rsc_0_37_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_111_4_64_16_16_64_1_gen twiddle_rsc_0_38_i
      (
      .q(twiddle_rsc_0_38_q),
      .radr(twiddle_rsc_0_38_radr),
      .q_d(twiddle_rsc_0_38_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_112_4_64_16_16_64_1_gen twiddle_rsc_0_39_i
      (
      .q(twiddle_rsc_0_39_q),
      .radr(twiddle_rsc_0_39_radr),
      .q_d(twiddle_rsc_0_39_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_113_4_64_16_16_64_1_gen twiddle_rsc_0_40_i
      (
      .q(twiddle_rsc_0_40_q),
      .radr(twiddle_rsc_0_40_radr),
      .q_d(twiddle_rsc_0_40_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_114_4_64_16_16_64_1_gen twiddle_rsc_0_41_i
      (
      .q(twiddle_rsc_0_41_q),
      .radr(twiddle_rsc_0_41_radr),
      .q_d(twiddle_rsc_0_41_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_115_4_64_16_16_64_1_gen twiddle_rsc_0_42_i
      (
      .q(twiddle_rsc_0_42_q),
      .radr(twiddle_rsc_0_42_radr),
      .q_d(twiddle_rsc_0_42_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_116_4_64_16_16_64_1_gen twiddle_rsc_0_43_i
      (
      .q(twiddle_rsc_0_43_q),
      .radr(twiddle_rsc_0_43_radr),
      .q_d(twiddle_rsc_0_43_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_117_4_64_16_16_64_1_gen twiddle_rsc_0_44_i
      (
      .q(twiddle_rsc_0_44_q),
      .radr(twiddle_rsc_0_44_radr),
      .q_d(twiddle_rsc_0_44_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_118_4_64_16_16_64_1_gen twiddle_rsc_0_45_i
      (
      .q(twiddle_rsc_0_45_q),
      .radr(twiddle_rsc_0_45_radr),
      .q_d(twiddle_rsc_0_45_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_119_4_64_16_16_64_1_gen twiddle_rsc_0_46_i
      (
      .q(twiddle_rsc_0_46_q),
      .radr(twiddle_rsc_0_46_radr),
      .q_d(twiddle_rsc_0_46_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_120_4_64_16_16_64_1_gen twiddle_rsc_0_47_i
      (
      .q(twiddle_rsc_0_47_q),
      .radr(twiddle_rsc_0_47_radr),
      .q_d(twiddle_rsc_0_47_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_121_4_64_16_16_64_1_gen twiddle_rsc_0_48_i
      (
      .q(twiddle_rsc_0_48_q),
      .radr(twiddle_rsc_0_48_radr),
      .q_d(twiddle_rsc_0_48_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_122_4_64_16_16_64_1_gen twiddle_rsc_0_49_i
      (
      .q(twiddle_rsc_0_49_q),
      .radr(twiddle_rsc_0_49_radr),
      .q_d(twiddle_rsc_0_49_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_123_4_64_16_16_64_1_gen twiddle_rsc_0_50_i
      (
      .q(twiddle_rsc_0_50_q),
      .radr(twiddle_rsc_0_50_radr),
      .q_d(twiddle_rsc_0_50_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_124_4_64_16_16_64_1_gen twiddle_rsc_0_51_i
      (
      .q(twiddle_rsc_0_51_q),
      .radr(twiddle_rsc_0_51_radr),
      .q_d(twiddle_rsc_0_51_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_125_4_64_16_16_64_1_gen twiddle_rsc_0_52_i
      (
      .q(twiddle_rsc_0_52_q),
      .radr(twiddle_rsc_0_52_radr),
      .q_d(twiddle_rsc_0_52_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_126_4_64_16_16_64_1_gen twiddle_rsc_0_53_i
      (
      .q(twiddle_rsc_0_53_q),
      .radr(twiddle_rsc_0_53_radr),
      .q_d(twiddle_rsc_0_53_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_127_4_64_16_16_64_1_gen twiddle_rsc_0_54_i
      (
      .q(twiddle_rsc_0_54_q),
      .radr(twiddle_rsc_0_54_radr),
      .q_d(twiddle_rsc_0_54_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_128_4_64_16_16_64_1_gen twiddle_rsc_0_55_i
      (
      .q(twiddle_rsc_0_55_q),
      .radr(twiddle_rsc_0_55_radr),
      .q_d(twiddle_rsc_0_55_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_129_4_64_16_16_64_1_gen twiddle_rsc_0_56_i
      (
      .q(twiddle_rsc_0_56_q),
      .radr(twiddle_rsc_0_56_radr),
      .q_d(twiddle_rsc_0_56_i_q_d),
      .radr_d(twiddle_rsc_0_0_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_130_4_64_16_16_64_1_gen twiddle_rsc_0_57_i
      (
      .q(twiddle_rsc_0_57_q),
      .radr(twiddle_rsc_0_57_radr),
      .q_d(twiddle_rsc_0_57_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_131_4_64_16_16_64_1_gen twiddle_rsc_0_58_i
      (
      .q(twiddle_rsc_0_58_q),
      .radr(twiddle_rsc_0_58_radr),
      .q_d(twiddle_rsc_0_58_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_132_4_64_16_16_64_1_gen twiddle_rsc_0_59_i
      (
      .q(twiddle_rsc_0_59_q),
      .radr(twiddle_rsc_0_59_radr),
      .q_d(twiddle_rsc_0_59_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_133_4_64_16_16_64_1_gen twiddle_rsc_0_60_i
      (
      .q(twiddle_rsc_0_60_q),
      .radr(twiddle_rsc_0_60_radr),
      .q_d(twiddle_rsc_0_60_i_q_d),
      .radr_d(twiddle_rsc_0_4_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_134_4_64_16_16_64_1_gen twiddle_rsc_0_61_i
      (
      .q(twiddle_rsc_0_61_q),
      .radr(twiddle_rsc_0_61_radr),
      .q_d(twiddle_rsc_0_61_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_135_4_64_16_16_64_1_gen twiddle_rsc_0_62_i
      (
      .q(twiddle_rsc_0_62_q),
      .radr(twiddle_rsc_0_62_radr),
      .q_d(twiddle_rsc_0_62_i_q_d),
      .radr_d(twiddle_rsc_0_2_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_136_4_64_16_16_64_1_gen twiddle_rsc_0_63_i
      (
      .q(twiddle_rsc_0_63_q),
      .radr(twiddle_rsc_0_63_radr),
      .q_d(twiddle_rsc_0_63_i_q_d),
      .radr_d(twiddle_rsc_0_1_i_radr_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d)
    );
  inPlaceNTT_DIF_core inPlaceNTT_DIF_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .vec_rsc_triosy_0_16_lz(vec_rsc_triosy_0_16_lz),
      .vec_rsc_triosy_0_17_lz(vec_rsc_triosy_0_17_lz),
      .vec_rsc_triosy_0_18_lz(vec_rsc_triosy_0_18_lz),
      .vec_rsc_triosy_0_19_lz(vec_rsc_triosy_0_19_lz),
      .vec_rsc_triosy_0_20_lz(vec_rsc_triosy_0_20_lz),
      .vec_rsc_triosy_0_21_lz(vec_rsc_triosy_0_21_lz),
      .vec_rsc_triosy_0_22_lz(vec_rsc_triosy_0_22_lz),
      .vec_rsc_triosy_0_23_lz(vec_rsc_triosy_0_23_lz),
      .vec_rsc_triosy_0_24_lz(vec_rsc_triosy_0_24_lz),
      .vec_rsc_triosy_0_25_lz(vec_rsc_triosy_0_25_lz),
      .vec_rsc_triosy_0_26_lz(vec_rsc_triosy_0_26_lz),
      .vec_rsc_triosy_0_27_lz(vec_rsc_triosy_0_27_lz),
      .vec_rsc_triosy_0_28_lz(vec_rsc_triosy_0_28_lz),
      .vec_rsc_triosy_0_29_lz(vec_rsc_triosy_0_29_lz),
      .vec_rsc_triosy_0_30_lz(vec_rsc_triosy_0_30_lz),
      .vec_rsc_triosy_0_31_lz(vec_rsc_triosy_0_31_lz),
      .vec_rsc_triosy_0_32_lz(vec_rsc_triosy_0_32_lz),
      .vec_rsc_triosy_0_33_lz(vec_rsc_triosy_0_33_lz),
      .vec_rsc_triosy_0_34_lz(vec_rsc_triosy_0_34_lz),
      .vec_rsc_triosy_0_35_lz(vec_rsc_triosy_0_35_lz),
      .vec_rsc_triosy_0_36_lz(vec_rsc_triosy_0_36_lz),
      .vec_rsc_triosy_0_37_lz(vec_rsc_triosy_0_37_lz),
      .vec_rsc_triosy_0_38_lz(vec_rsc_triosy_0_38_lz),
      .vec_rsc_triosy_0_39_lz(vec_rsc_triosy_0_39_lz),
      .vec_rsc_triosy_0_40_lz(vec_rsc_triosy_0_40_lz),
      .vec_rsc_triosy_0_41_lz(vec_rsc_triosy_0_41_lz),
      .vec_rsc_triosy_0_42_lz(vec_rsc_triosy_0_42_lz),
      .vec_rsc_triosy_0_43_lz(vec_rsc_triosy_0_43_lz),
      .vec_rsc_triosy_0_44_lz(vec_rsc_triosy_0_44_lz),
      .vec_rsc_triosy_0_45_lz(vec_rsc_triosy_0_45_lz),
      .vec_rsc_triosy_0_46_lz(vec_rsc_triosy_0_46_lz),
      .vec_rsc_triosy_0_47_lz(vec_rsc_triosy_0_47_lz),
      .vec_rsc_triosy_0_48_lz(vec_rsc_triosy_0_48_lz),
      .vec_rsc_triosy_0_49_lz(vec_rsc_triosy_0_49_lz),
      .vec_rsc_triosy_0_50_lz(vec_rsc_triosy_0_50_lz),
      .vec_rsc_triosy_0_51_lz(vec_rsc_triosy_0_51_lz),
      .vec_rsc_triosy_0_52_lz(vec_rsc_triosy_0_52_lz),
      .vec_rsc_triosy_0_53_lz(vec_rsc_triosy_0_53_lz),
      .vec_rsc_triosy_0_54_lz(vec_rsc_triosy_0_54_lz),
      .vec_rsc_triosy_0_55_lz(vec_rsc_triosy_0_55_lz),
      .vec_rsc_triosy_0_56_lz(vec_rsc_triosy_0_56_lz),
      .vec_rsc_triosy_0_57_lz(vec_rsc_triosy_0_57_lz),
      .vec_rsc_triosy_0_58_lz(vec_rsc_triosy_0_58_lz),
      .vec_rsc_triosy_0_59_lz(vec_rsc_triosy_0_59_lz),
      .vec_rsc_triosy_0_60_lz(vec_rsc_triosy_0_60_lz),
      .vec_rsc_triosy_0_61_lz(vec_rsc_triosy_0_61_lz),
      .vec_rsc_triosy_0_62_lz(vec_rsc_triosy_0_62_lz),
      .vec_rsc_triosy_0_63_lz(vec_rsc_triosy_0_63_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_0_0_lz(twiddle_rsc_triosy_0_0_lz),
      .twiddle_rsc_triosy_0_1_lz(twiddle_rsc_triosy_0_1_lz),
      .twiddle_rsc_triosy_0_2_lz(twiddle_rsc_triosy_0_2_lz),
      .twiddle_rsc_triosy_0_3_lz(twiddle_rsc_triosy_0_3_lz),
      .twiddle_rsc_triosy_0_4_lz(twiddle_rsc_triosy_0_4_lz),
      .twiddle_rsc_triosy_0_5_lz(twiddle_rsc_triosy_0_5_lz),
      .twiddle_rsc_triosy_0_6_lz(twiddle_rsc_triosy_0_6_lz),
      .twiddle_rsc_triosy_0_7_lz(twiddle_rsc_triosy_0_7_lz),
      .twiddle_rsc_triosy_0_8_lz(twiddle_rsc_triosy_0_8_lz),
      .twiddle_rsc_triosy_0_9_lz(twiddle_rsc_triosy_0_9_lz),
      .twiddle_rsc_triosy_0_10_lz(twiddle_rsc_triosy_0_10_lz),
      .twiddle_rsc_triosy_0_11_lz(twiddle_rsc_triosy_0_11_lz),
      .twiddle_rsc_triosy_0_12_lz(twiddle_rsc_triosy_0_12_lz),
      .twiddle_rsc_triosy_0_13_lz(twiddle_rsc_triosy_0_13_lz),
      .twiddle_rsc_triosy_0_14_lz(twiddle_rsc_triosy_0_14_lz),
      .twiddle_rsc_triosy_0_15_lz(twiddle_rsc_triosy_0_15_lz),
      .twiddle_rsc_triosy_0_16_lz(twiddle_rsc_triosy_0_16_lz),
      .twiddle_rsc_triosy_0_17_lz(twiddle_rsc_triosy_0_17_lz),
      .twiddle_rsc_triosy_0_18_lz(twiddle_rsc_triosy_0_18_lz),
      .twiddle_rsc_triosy_0_19_lz(twiddle_rsc_triosy_0_19_lz),
      .twiddle_rsc_triosy_0_20_lz(twiddle_rsc_triosy_0_20_lz),
      .twiddle_rsc_triosy_0_21_lz(twiddle_rsc_triosy_0_21_lz),
      .twiddle_rsc_triosy_0_22_lz(twiddle_rsc_triosy_0_22_lz),
      .twiddle_rsc_triosy_0_23_lz(twiddle_rsc_triosy_0_23_lz),
      .twiddle_rsc_triosy_0_24_lz(twiddle_rsc_triosy_0_24_lz),
      .twiddle_rsc_triosy_0_25_lz(twiddle_rsc_triosy_0_25_lz),
      .twiddle_rsc_triosy_0_26_lz(twiddle_rsc_triosy_0_26_lz),
      .twiddle_rsc_triosy_0_27_lz(twiddle_rsc_triosy_0_27_lz),
      .twiddle_rsc_triosy_0_28_lz(twiddle_rsc_triosy_0_28_lz),
      .twiddle_rsc_triosy_0_29_lz(twiddle_rsc_triosy_0_29_lz),
      .twiddle_rsc_triosy_0_30_lz(twiddle_rsc_triosy_0_30_lz),
      .twiddle_rsc_triosy_0_31_lz(twiddle_rsc_triosy_0_31_lz),
      .twiddle_rsc_triosy_0_32_lz(twiddle_rsc_triosy_0_32_lz),
      .twiddle_rsc_triosy_0_33_lz(twiddle_rsc_triosy_0_33_lz),
      .twiddle_rsc_triosy_0_34_lz(twiddle_rsc_triosy_0_34_lz),
      .twiddle_rsc_triosy_0_35_lz(twiddle_rsc_triosy_0_35_lz),
      .twiddle_rsc_triosy_0_36_lz(twiddle_rsc_triosy_0_36_lz),
      .twiddle_rsc_triosy_0_37_lz(twiddle_rsc_triosy_0_37_lz),
      .twiddle_rsc_triosy_0_38_lz(twiddle_rsc_triosy_0_38_lz),
      .twiddle_rsc_triosy_0_39_lz(twiddle_rsc_triosy_0_39_lz),
      .twiddle_rsc_triosy_0_40_lz(twiddle_rsc_triosy_0_40_lz),
      .twiddle_rsc_triosy_0_41_lz(twiddle_rsc_triosy_0_41_lz),
      .twiddle_rsc_triosy_0_42_lz(twiddle_rsc_triosy_0_42_lz),
      .twiddle_rsc_triosy_0_43_lz(twiddle_rsc_triosy_0_43_lz),
      .twiddle_rsc_triosy_0_44_lz(twiddle_rsc_triosy_0_44_lz),
      .twiddle_rsc_triosy_0_45_lz(twiddle_rsc_triosy_0_45_lz),
      .twiddle_rsc_triosy_0_46_lz(twiddle_rsc_triosy_0_46_lz),
      .twiddle_rsc_triosy_0_47_lz(twiddle_rsc_triosy_0_47_lz),
      .twiddle_rsc_triosy_0_48_lz(twiddle_rsc_triosy_0_48_lz),
      .twiddle_rsc_triosy_0_49_lz(twiddle_rsc_triosy_0_49_lz),
      .twiddle_rsc_triosy_0_50_lz(twiddle_rsc_triosy_0_50_lz),
      .twiddle_rsc_triosy_0_51_lz(twiddle_rsc_triosy_0_51_lz),
      .twiddle_rsc_triosy_0_52_lz(twiddle_rsc_triosy_0_52_lz),
      .twiddle_rsc_triosy_0_53_lz(twiddle_rsc_triosy_0_53_lz),
      .twiddle_rsc_triosy_0_54_lz(twiddle_rsc_triosy_0_54_lz),
      .twiddle_rsc_triosy_0_55_lz(twiddle_rsc_triosy_0_55_lz),
      .twiddle_rsc_triosy_0_56_lz(twiddle_rsc_triosy_0_56_lz),
      .twiddle_rsc_triosy_0_57_lz(twiddle_rsc_triosy_0_57_lz),
      .twiddle_rsc_triosy_0_58_lz(twiddle_rsc_triosy_0_58_lz),
      .twiddle_rsc_triosy_0_59_lz(twiddle_rsc_triosy_0_59_lz),
      .twiddle_rsc_triosy_0_60_lz(twiddle_rsc_triosy_0_60_lz),
      .twiddle_rsc_triosy_0_61_lz(twiddle_rsc_triosy_0_61_lz),
      .twiddle_rsc_triosy_0_62_lz(twiddle_rsc_triosy_0_62_lz),
      .twiddle_rsc_triosy_0_63_lz(twiddle_rsc_triosy_0_63_lz),
      .vec_rsc_0_0_i_q_d(vec_rsc_0_0_i_q_d),
      .vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_q_d(vec_rsc_0_1_i_q_d),
      .vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_q_d(vec_rsc_0_2_i_q_d),
      .vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_q_d(vec_rsc_0_3_i_q_d),
      .vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_q_d(vec_rsc_0_4_i_q_d),
      .vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_q_d(vec_rsc_0_5_i_q_d),
      .vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_q_d(vec_rsc_0_6_i_q_d),
      .vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_q_d(vec_rsc_0_7_i_q_d),
      .vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_q_d(vec_rsc_0_8_i_q_d),
      .vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_q_d(vec_rsc_0_9_i_q_d),
      .vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_q_d(vec_rsc_0_10_i_q_d),
      .vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_q_d(vec_rsc_0_11_i_q_d),
      .vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_q_d(vec_rsc_0_12_i_q_d),
      .vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_q_d(vec_rsc_0_13_i_q_d),
      .vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_q_d(vec_rsc_0_14_i_q_d),
      .vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_q_d(vec_rsc_0_15_i_q_d),
      .vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_16_i_q_d(vec_rsc_0_16_i_q_d),
      .vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_17_i_q_d(vec_rsc_0_17_i_q_d),
      .vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_18_i_q_d(vec_rsc_0_18_i_q_d),
      .vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_19_i_q_d(vec_rsc_0_19_i_q_d),
      .vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_20_i_q_d(vec_rsc_0_20_i_q_d),
      .vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_21_i_q_d(vec_rsc_0_21_i_q_d),
      .vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_22_i_q_d(vec_rsc_0_22_i_q_d),
      .vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_23_i_q_d(vec_rsc_0_23_i_q_d),
      .vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_24_i_q_d(vec_rsc_0_24_i_q_d),
      .vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_25_i_q_d(vec_rsc_0_25_i_q_d),
      .vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_26_i_q_d(vec_rsc_0_26_i_q_d),
      .vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_27_i_q_d(vec_rsc_0_27_i_q_d),
      .vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_28_i_q_d(vec_rsc_0_28_i_q_d),
      .vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_29_i_q_d(vec_rsc_0_29_i_q_d),
      .vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_30_i_q_d(vec_rsc_0_30_i_q_d),
      .vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_31_i_q_d(vec_rsc_0_31_i_q_d),
      .vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_32_i_q_d(vec_rsc_0_32_i_q_d),
      .vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_33_i_q_d(vec_rsc_0_33_i_q_d),
      .vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_34_i_q_d(vec_rsc_0_34_i_q_d),
      .vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_35_i_q_d(vec_rsc_0_35_i_q_d),
      .vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_36_i_q_d(vec_rsc_0_36_i_q_d),
      .vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_37_i_q_d(vec_rsc_0_37_i_q_d),
      .vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_38_i_q_d(vec_rsc_0_38_i_q_d),
      .vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_39_i_q_d(vec_rsc_0_39_i_q_d),
      .vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_40_i_q_d(vec_rsc_0_40_i_q_d),
      .vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_41_i_q_d(vec_rsc_0_41_i_q_d),
      .vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_42_i_q_d(vec_rsc_0_42_i_q_d),
      .vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_43_i_q_d(vec_rsc_0_43_i_q_d),
      .vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_44_i_q_d(vec_rsc_0_44_i_q_d),
      .vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_45_i_q_d(vec_rsc_0_45_i_q_d),
      .vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_46_i_q_d(vec_rsc_0_46_i_q_d),
      .vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_47_i_q_d(vec_rsc_0_47_i_q_d),
      .vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_48_i_q_d(vec_rsc_0_48_i_q_d),
      .vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_49_i_q_d(vec_rsc_0_49_i_q_d),
      .vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_50_i_q_d(vec_rsc_0_50_i_q_d),
      .vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_51_i_q_d(vec_rsc_0_51_i_q_d),
      .vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_52_i_q_d(vec_rsc_0_52_i_q_d),
      .vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_53_i_q_d(vec_rsc_0_53_i_q_d),
      .vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_54_i_q_d(vec_rsc_0_54_i_q_d),
      .vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_55_i_q_d(vec_rsc_0_55_i_q_d),
      .vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_56_i_q_d(vec_rsc_0_56_i_q_d),
      .vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_57_i_q_d(vec_rsc_0_57_i_q_d),
      .vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_58_i_q_d(vec_rsc_0_58_i_q_d),
      .vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_59_i_q_d(vec_rsc_0_59_i_q_d),
      .vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_60_i_q_d(vec_rsc_0_60_i_q_d),
      .vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_61_i_q_d(vec_rsc_0_61_i_q_d),
      .vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_62_i_q_d(vec_rsc_0_62_i_q_d),
      .vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_63_i_q_d(vec_rsc_0_63_i_q_d),
      .vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d(vec_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_0_i_q_d(twiddle_rsc_0_0_i_q_d),
      .twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_1_i_q_d(twiddle_rsc_0_1_i_q_d),
      .twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_2_i_q_d(twiddle_rsc_0_2_i_q_d),
      .twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_3_i_q_d(twiddle_rsc_0_3_i_q_d),
      .twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_4_i_q_d(twiddle_rsc_0_4_i_q_d),
      .twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_5_i_q_d(twiddle_rsc_0_5_i_q_d),
      .twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_6_i_q_d(twiddle_rsc_0_6_i_q_d),
      .twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_7_i_q_d(twiddle_rsc_0_7_i_q_d),
      .twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_8_i_q_d(twiddle_rsc_0_8_i_q_d),
      .twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_9_i_q_d(twiddle_rsc_0_9_i_q_d),
      .twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_10_i_q_d(twiddle_rsc_0_10_i_q_d),
      .twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_11_i_q_d(twiddle_rsc_0_11_i_q_d),
      .twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_12_i_q_d(twiddle_rsc_0_12_i_q_d),
      .twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_13_i_q_d(twiddle_rsc_0_13_i_q_d),
      .twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_14_i_q_d(twiddle_rsc_0_14_i_q_d),
      .twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_15_i_q_d(twiddle_rsc_0_15_i_q_d),
      .twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_16_i_q_d(twiddle_rsc_0_16_i_q_d),
      .twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_16_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_17_i_q_d(twiddle_rsc_0_17_i_q_d),
      .twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_17_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_18_i_q_d(twiddle_rsc_0_18_i_q_d),
      .twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_18_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_19_i_q_d(twiddle_rsc_0_19_i_q_d),
      .twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_19_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_20_i_q_d(twiddle_rsc_0_20_i_q_d),
      .twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_20_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_21_i_q_d(twiddle_rsc_0_21_i_q_d),
      .twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_21_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_22_i_q_d(twiddle_rsc_0_22_i_q_d),
      .twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_22_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_23_i_q_d(twiddle_rsc_0_23_i_q_d),
      .twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_23_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_24_i_q_d(twiddle_rsc_0_24_i_q_d),
      .twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_24_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_25_i_q_d(twiddle_rsc_0_25_i_q_d),
      .twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_25_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_26_i_q_d(twiddle_rsc_0_26_i_q_d),
      .twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_26_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_27_i_q_d(twiddle_rsc_0_27_i_q_d),
      .twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_27_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_28_i_q_d(twiddle_rsc_0_28_i_q_d),
      .twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_28_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_29_i_q_d(twiddle_rsc_0_29_i_q_d),
      .twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_29_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_30_i_q_d(twiddle_rsc_0_30_i_q_d),
      .twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_30_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_31_i_q_d(twiddle_rsc_0_31_i_q_d),
      .twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_31_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_32_i_q_d(twiddle_rsc_0_32_i_q_d),
      .twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_32_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_33_i_q_d(twiddle_rsc_0_33_i_q_d),
      .twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_33_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_34_i_q_d(twiddle_rsc_0_34_i_q_d),
      .twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_34_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_35_i_q_d(twiddle_rsc_0_35_i_q_d),
      .twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_35_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_36_i_q_d(twiddle_rsc_0_36_i_q_d),
      .twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_36_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_37_i_q_d(twiddle_rsc_0_37_i_q_d),
      .twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_37_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_38_i_q_d(twiddle_rsc_0_38_i_q_d),
      .twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_38_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_39_i_q_d(twiddle_rsc_0_39_i_q_d),
      .twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_39_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_40_i_q_d(twiddle_rsc_0_40_i_q_d),
      .twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_40_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_41_i_q_d(twiddle_rsc_0_41_i_q_d),
      .twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_41_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_42_i_q_d(twiddle_rsc_0_42_i_q_d),
      .twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_42_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_43_i_q_d(twiddle_rsc_0_43_i_q_d),
      .twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_43_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_44_i_q_d(twiddle_rsc_0_44_i_q_d),
      .twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_44_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_45_i_q_d(twiddle_rsc_0_45_i_q_d),
      .twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_45_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_46_i_q_d(twiddle_rsc_0_46_i_q_d),
      .twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_46_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_47_i_q_d(twiddle_rsc_0_47_i_q_d),
      .twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_47_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_48_i_q_d(twiddle_rsc_0_48_i_q_d),
      .twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_48_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_49_i_q_d(twiddle_rsc_0_49_i_q_d),
      .twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_49_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_50_i_q_d(twiddle_rsc_0_50_i_q_d),
      .twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_50_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_51_i_q_d(twiddle_rsc_0_51_i_q_d),
      .twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_51_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_52_i_q_d(twiddle_rsc_0_52_i_q_d),
      .twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_52_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_53_i_q_d(twiddle_rsc_0_53_i_q_d),
      .twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_53_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_54_i_q_d(twiddle_rsc_0_54_i_q_d),
      .twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_54_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_55_i_q_d(twiddle_rsc_0_55_i_q_d),
      .twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_55_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_56_i_q_d(twiddle_rsc_0_56_i_q_d),
      .twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_56_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_57_i_q_d(twiddle_rsc_0_57_i_q_d),
      .twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_57_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_58_i_q_d(twiddle_rsc_0_58_i_q_d),
      .twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_58_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_59_i_q_d(twiddle_rsc_0_59_i_q_d),
      .twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_59_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_60_i_q_d(twiddle_rsc_0_60_i_q_d),
      .twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_60_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_61_i_q_d(twiddle_rsc_0_61_i_q_d),
      .twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_61_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_62_i_q_d(twiddle_rsc_0_62_i_q_d),
      .twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_62_i_readA_r_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_63_i_q_d(twiddle_rsc_0_63_i_q_d),
      .twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_63_i_readA_r_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_d_d_pff(vec_rsc_0_0_i_d_d_iff),
      .vec_rsc_0_0_i_radr_d_pff(vec_rsc_0_0_i_radr_d_iff),
      .vec_rsc_0_0_i_wadr_d_pff(vec_rsc_0_0_i_wadr_d_iff),
      .vec_rsc_0_0_i_we_d_pff(vec_rsc_0_0_i_we_d_iff),
      .vec_rsc_0_1_i_we_d_pff(vec_rsc_0_1_i_we_d_iff),
      .vec_rsc_0_2_i_we_d_pff(vec_rsc_0_2_i_we_d_iff),
      .vec_rsc_0_3_i_we_d_pff(vec_rsc_0_3_i_we_d_iff),
      .vec_rsc_0_4_i_we_d_pff(vec_rsc_0_4_i_we_d_iff),
      .vec_rsc_0_5_i_we_d_pff(vec_rsc_0_5_i_we_d_iff),
      .vec_rsc_0_6_i_we_d_pff(vec_rsc_0_6_i_we_d_iff),
      .vec_rsc_0_7_i_we_d_pff(vec_rsc_0_7_i_we_d_iff),
      .vec_rsc_0_8_i_we_d_pff(vec_rsc_0_8_i_we_d_iff),
      .vec_rsc_0_9_i_we_d_pff(vec_rsc_0_9_i_we_d_iff),
      .vec_rsc_0_10_i_we_d_pff(vec_rsc_0_10_i_we_d_iff),
      .vec_rsc_0_11_i_we_d_pff(vec_rsc_0_11_i_we_d_iff),
      .vec_rsc_0_12_i_we_d_pff(vec_rsc_0_12_i_we_d_iff),
      .vec_rsc_0_13_i_we_d_pff(vec_rsc_0_13_i_we_d_iff),
      .vec_rsc_0_14_i_we_d_pff(vec_rsc_0_14_i_we_d_iff),
      .vec_rsc_0_15_i_we_d_pff(vec_rsc_0_15_i_we_d_iff),
      .vec_rsc_0_16_i_we_d_pff(vec_rsc_0_16_i_we_d_iff),
      .vec_rsc_0_17_i_we_d_pff(vec_rsc_0_17_i_we_d_iff),
      .vec_rsc_0_18_i_we_d_pff(vec_rsc_0_18_i_we_d_iff),
      .vec_rsc_0_19_i_we_d_pff(vec_rsc_0_19_i_we_d_iff),
      .vec_rsc_0_20_i_we_d_pff(vec_rsc_0_20_i_we_d_iff),
      .vec_rsc_0_21_i_we_d_pff(vec_rsc_0_21_i_we_d_iff),
      .vec_rsc_0_22_i_we_d_pff(vec_rsc_0_22_i_we_d_iff),
      .vec_rsc_0_23_i_we_d_pff(vec_rsc_0_23_i_we_d_iff),
      .vec_rsc_0_24_i_we_d_pff(vec_rsc_0_24_i_we_d_iff),
      .vec_rsc_0_25_i_we_d_pff(vec_rsc_0_25_i_we_d_iff),
      .vec_rsc_0_26_i_we_d_pff(vec_rsc_0_26_i_we_d_iff),
      .vec_rsc_0_27_i_we_d_pff(vec_rsc_0_27_i_we_d_iff),
      .vec_rsc_0_28_i_we_d_pff(vec_rsc_0_28_i_we_d_iff),
      .vec_rsc_0_29_i_we_d_pff(vec_rsc_0_29_i_we_d_iff),
      .vec_rsc_0_30_i_we_d_pff(vec_rsc_0_30_i_we_d_iff),
      .vec_rsc_0_31_i_we_d_pff(vec_rsc_0_31_i_we_d_iff),
      .vec_rsc_0_32_i_we_d_pff(vec_rsc_0_32_i_we_d_iff),
      .vec_rsc_0_33_i_we_d_pff(vec_rsc_0_33_i_we_d_iff),
      .vec_rsc_0_34_i_we_d_pff(vec_rsc_0_34_i_we_d_iff),
      .vec_rsc_0_35_i_we_d_pff(vec_rsc_0_35_i_we_d_iff),
      .vec_rsc_0_36_i_we_d_pff(vec_rsc_0_36_i_we_d_iff),
      .vec_rsc_0_37_i_we_d_pff(vec_rsc_0_37_i_we_d_iff),
      .vec_rsc_0_38_i_we_d_pff(vec_rsc_0_38_i_we_d_iff),
      .vec_rsc_0_39_i_we_d_pff(vec_rsc_0_39_i_we_d_iff),
      .vec_rsc_0_40_i_we_d_pff(vec_rsc_0_40_i_we_d_iff),
      .vec_rsc_0_41_i_we_d_pff(vec_rsc_0_41_i_we_d_iff),
      .vec_rsc_0_42_i_we_d_pff(vec_rsc_0_42_i_we_d_iff),
      .vec_rsc_0_43_i_we_d_pff(vec_rsc_0_43_i_we_d_iff),
      .vec_rsc_0_44_i_we_d_pff(vec_rsc_0_44_i_we_d_iff),
      .vec_rsc_0_45_i_we_d_pff(vec_rsc_0_45_i_we_d_iff),
      .vec_rsc_0_46_i_we_d_pff(vec_rsc_0_46_i_we_d_iff),
      .vec_rsc_0_47_i_we_d_pff(vec_rsc_0_47_i_we_d_iff),
      .vec_rsc_0_48_i_we_d_pff(vec_rsc_0_48_i_we_d_iff),
      .vec_rsc_0_49_i_we_d_pff(vec_rsc_0_49_i_we_d_iff),
      .vec_rsc_0_50_i_we_d_pff(vec_rsc_0_50_i_we_d_iff),
      .vec_rsc_0_51_i_we_d_pff(vec_rsc_0_51_i_we_d_iff),
      .vec_rsc_0_52_i_we_d_pff(vec_rsc_0_52_i_we_d_iff),
      .vec_rsc_0_53_i_we_d_pff(vec_rsc_0_53_i_we_d_iff),
      .vec_rsc_0_54_i_we_d_pff(vec_rsc_0_54_i_we_d_iff),
      .vec_rsc_0_55_i_we_d_pff(vec_rsc_0_55_i_we_d_iff),
      .vec_rsc_0_56_i_we_d_pff(vec_rsc_0_56_i_we_d_iff),
      .vec_rsc_0_57_i_we_d_pff(vec_rsc_0_57_i_we_d_iff),
      .vec_rsc_0_58_i_we_d_pff(vec_rsc_0_58_i_we_d_iff),
      .vec_rsc_0_59_i_we_d_pff(vec_rsc_0_59_i_we_d_iff),
      .vec_rsc_0_60_i_we_d_pff(vec_rsc_0_60_i_we_d_iff),
      .vec_rsc_0_61_i_we_d_pff(vec_rsc_0_61_i_we_d_iff),
      .vec_rsc_0_62_i_we_d_pff(vec_rsc_0_62_i_we_d_iff),
      .vec_rsc_0_63_i_we_d_pff(vec_rsc_0_63_i_we_d_iff),
      .twiddle_rsc_0_0_i_radr_d_pff(twiddle_rsc_0_0_i_radr_d_iff),
      .twiddle_rsc_0_1_i_radr_d_pff(twiddle_rsc_0_1_i_radr_d_iff),
      .twiddle_rsc_0_2_i_radr_d_pff(twiddle_rsc_0_2_i_radr_d_iff),
      .twiddle_rsc_0_4_i_radr_d_pff(twiddle_rsc_0_4_i_radr_d_iff)
    );
endmodule



