
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_rem_beh.v 
module mgc_rem(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_b-1:0] z;  
   reg  [width_b-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  rem_s(a,b,z);
	else
          rem_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_div_beh.v 
module mgc_div(a,b,z);
   parameter width_a = 8;
   parameter width_b = 8;
   parameter signd = 1;
   input [width_a-1:0] a;
   input [width_b-1:0] b; 
   output [width_a-1:0] z;  
   reg  [width_a-1:0] z;

   always@(a or b)
     begin
	if(signd)
	  div_s(a,b,z);
	else
          div_u(a,b,z);
     end


//-----------------------------------------------------------------
//     -- Vectorized Overloaded Arithmetic Operators
//-----------------------------------------------------------------
   
   function [width_a-1:0] fabs_l; 
      input [width_a-1:0] arg1;
      begin
         case(arg1[width_a-1])
            1'b1:
               fabs_l = {(width_a){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_l = arg1;
         endcase
      end
   endfunction
   
   function [width_b-1:0] fabs_r; 
      input [width_b-1:0] arg1;
      begin
         case (arg1[width_b-1])
            1'b1:
               fabs_r =  {(width_b){1'b0}} - arg1;
            default: // was: 1'b0:
               fabs_r = arg1;
         endcase
      end
   endfunction

   function [width_b:0] minus;
     input [width_b:0] in1;
     input [width_b:0] in2;
     reg [width_b+1:0] tmp;
     begin
       tmp = in1 - in2;
       minus = tmp[width_b:0];
     end
   endfunction

   
   task divmod;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      output [width_b-1:0] rmod;
      
      parameter llen = width_a;
      parameter rlen = width_b;
      reg [(llen+rlen)-1:0] lbuf;
      reg [rlen:0] diff;
	  integer i;
      begin
	 lbuf = {(llen+rlen){1'b0}};
//64'b0;
	 lbuf[llen-1:0] = l;
	 for(i=width_a-1;i>=0;i=i-1)
	   begin
              diff = minus(lbuf[(llen+rlen)-1:llen-1], {1'b0,r});
	      rdiv[i] = ~diff[rlen];
	      if(diff[rlen] == 0)
		lbuf[(llen+rlen)-1:llen-1] = diff;
	      lbuf[(llen+rlen)-1:1] = lbuf[(llen+rlen)-2:0];
	   end
	 rmod = lbuf[(llen+rlen)-1:llen];
      end
   endtask
      

   task div_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask
   
   task mod_u;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(l, r, rdiv, rmod);
      end
   endtask

   task rem_u; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;
      begin
	 mod_u(l,r,rmod);
      end
   endtask // rem_u

   task div_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_a-1:0] rdiv;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l), fabs_r(r),rdiv,rmod);
	 if(l[width_a-1] != r[width_b-1])
	   rdiv = {(width_a){1'b0}} - rdiv;
      end
   endtask

   task mod_s;
      input [width_a-1:0] l;
      input [width_b-1:0] r;
      output [width_b-1:0] rmod;
      
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      reg [width_b-1:0] rnul;
      reg [width_b:0] rmod_t;
      begin
         rnul = {width_b{1'b0}};
	 divmod(fabs_l(l), fabs_r(r), rdiv, rmod);
         if (l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
	 if((rmod != rnul) && (l[width_a-1] != r[width_b-1]))
            begin
               rmod_t = r + rmod;
               rmod = rmod_t[width_b-1:0];
            end
      end
   endtask // mod_s
   
   task rem_s; 
      input [width_a-1:0] l;
      input [width_b-1:0] r;    
      output [width_b-1:0] rmod;   
      reg [width_a-01:0] rdiv;
      reg [width_b-1:0] rmod;
      begin
	 divmod(fabs_l(l),fabs_r(r),rdiv,rmod);
	 if(l[width_a-1])
	   rmod = {(width_b){1'b0}} - rmod;
      end
   endtask

  endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Thu Jul  1 13:33:43 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
// ------------------------------------------------------------------


module inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen
    (
  qa, wea, da, adra, adra_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [63:0] qa;
  output wea;
  output [63:0] da;
  output [7:0] adra;
  input [7:0] adra_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input wea_d;
  input rwA_rw_ram_ir_internal_RMASK_B_d;
  input rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d);
  assign da = (da_d);
  assign adra = (adra_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core_core_fsm (
  clk, rst, fsm_output, STAGE_LOOP_C_8_tr0, modExp_while_C_38_tr0, COMP_LOOP_C_1_tr0,
      COMP_LOOP_1_modExp_1_while_C_38_tr0, COMP_LOOP_C_64_tr0, COMP_LOOP_2_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_128_tr0, COMP_LOOP_3_modExp_1_while_C_38_tr0, COMP_LOOP_C_192_tr0,
      COMP_LOOP_4_modExp_1_while_C_38_tr0, COMP_LOOP_C_256_tr0, COMP_LOOP_5_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_320_tr0, COMP_LOOP_6_modExp_1_while_C_38_tr0, COMP_LOOP_C_384_tr0,
      COMP_LOOP_7_modExp_1_while_C_38_tr0, COMP_LOOP_C_448_tr0, COMP_LOOP_8_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_512_tr0, COMP_LOOP_9_modExp_1_while_C_38_tr0, COMP_LOOP_C_576_tr0,
      COMP_LOOP_10_modExp_1_while_C_38_tr0, COMP_LOOP_C_640_tr0, COMP_LOOP_11_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_704_tr0, COMP_LOOP_12_modExp_1_while_C_38_tr0, COMP_LOOP_C_768_tr0,
      COMP_LOOP_13_modExp_1_while_C_38_tr0, COMP_LOOP_C_832_tr0, COMP_LOOP_14_modExp_1_while_C_38_tr0,
      COMP_LOOP_C_896_tr0, COMP_LOOP_15_modExp_1_while_C_38_tr0, COMP_LOOP_C_960_tr0,
      COMP_LOOP_16_modExp_1_while_C_38_tr0, COMP_LOOP_C_1024_tr0, VEC_LOOP_C_0_tr0,
      STAGE_LOOP_C_9_tr0
);
  input clk;
  input rst;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input STAGE_LOOP_C_8_tr0;
  input modExp_while_C_38_tr0;
  input COMP_LOOP_C_1_tr0;
  input COMP_LOOP_1_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_64_tr0;
  input COMP_LOOP_2_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_128_tr0;
  input COMP_LOOP_3_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_192_tr0;
  input COMP_LOOP_4_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_256_tr0;
  input COMP_LOOP_5_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_320_tr0;
  input COMP_LOOP_6_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_384_tr0;
  input COMP_LOOP_7_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_448_tr0;
  input COMP_LOOP_8_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_512_tr0;
  input COMP_LOOP_9_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_576_tr0;
  input COMP_LOOP_10_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_640_tr0;
  input COMP_LOOP_11_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_704_tr0;
  input COMP_LOOP_12_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_768_tr0;
  input COMP_LOOP_13_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_832_tr0;
  input COMP_LOOP_14_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_896_tr0;
  input COMP_LOOP_15_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_960_tr0;
  input COMP_LOOP_16_modExp_1_while_C_38_tr0;
  input COMP_LOOP_C_1024_tr0;
  input VEC_LOOP_C_0_tr0;
  input STAGE_LOOP_C_9_tr0;


  // FSM State Type Declaration for inPlaceNTT_DIT_core_core_fsm_1
  parameter
    main_C_0 = 11'd0,
    STAGE_LOOP_C_0 = 11'd1,
    STAGE_LOOP_C_1 = 11'd2,
    STAGE_LOOP_C_2 = 11'd3,
    STAGE_LOOP_C_3 = 11'd4,
    STAGE_LOOP_C_4 = 11'd5,
    STAGE_LOOP_C_5 = 11'd6,
    STAGE_LOOP_C_6 = 11'd7,
    STAGE_LOOP_C_7 = 11'd8,
    STAGE_LOOP_C_8 = 11'd9,
    modExp_while_C_0 = 11'd10,
    modExp_while_C_1 = 11'd11,
    modExp_while_C_2 = 11'd12,
    modExp_while_C_3 = 11'd13,
    modExp_while_C_4 = 11'd14,
    modExp_while_C_5 = 11'd15,
    modExp_while_C_6 = 11'd16,
    modExp_while_C_7 = 11'd17,
    modExp_while_C_8 = 11'd18,
    modExp_while_C_9 = 11'd19,
    modExp_while_C_10 = 11'd20,
    modExp_while_C_11 = 11'd21,
    modExp_while_C_12 = 11'd22,
    modExp_while_C_13 = 11'd23,
    modExp_while_C_14 = 11'd24,
    modExp_while_C_15 = 11'd25,
    modExp_while_C_16 = 11'd26,
    modExp_while_C_17 = 11'd27,
    modExp_while_C_18 = 11'd28,
    modExp_while_C_19 = 11'd29,
    modExp_while_C_20 = 11'd30,
    modExp_while_C_21 = 11'd31,
    modExp_while_C_22 = 11'd32,
    modExp_while_C_23 = 11'd33,
    modExp_while_C_24 = 11'd34,
    modExp_while_C_25 = 11'd35,
    modExp_while_C_26 = 11'd36,
    modExp_while_C_27 = 11'd37,
    modExp_while_C_28 = 11'd38,
    modExp_while_C_29 = 11'd39,
    modExp_while_C_30 = 11'd40,
    modExp_while_C_31 = 11'd41,
    modExp_while_C_32 = 11'd42,
    modExp_while_C_33 = 11'd43,
    modExp_while_C_34 = 11'd44,
    modExp_while_C_35 = 11'd45,
    modExp_while_C_36 = 11'd46,
    modExp_while_C_37 = 11'd47,
    modExp_while_C_38 = 11'd48,
    COMP_LOOP_C_0 = 11'd49,
    COMP_LOOP_C_1 = 11'd50,
    COMP_LOOP_1_modExp_1_while_C_0 = 11'd51,
    COMP_LOOP_1_modExp_1_while_C_1 = 11'd52,
    COMP_LOOP_1_modExp_1_while_C_2 = 11'd53,
    COMP_LOOP_1_modExp_1_while_C_3 = 11'd54,
    COMP_LOOP_1_modExp_1_while_C_4 = 11'd55,
    COMP_LOOP_1_modExp_1_while_C_5 = 11'd56,
    COMP_LOOP_1_modExp_1_while_C_6 = 11'd57,
    COMP_LOOP_1_modExp_1_while_C_7 = 11'd58,
    COMP_LOOP_1_modExp_1_while_C_8 = 11'd59,
    COMP_LOOP_1_modExp_1_while_C_9 = 11'd60,
    COMP_LOOP_1_modExp_1_while_C_10 = 11'd61,
    COMP_LOOP_1_modExp_1_while_C_11 = 11'd62,
    COMP_LOOP_1_modExp_1_while_C_12 = 11'd63,
    COMP_LOOP_1_modExp_1_while_C_13 = 11'd64,
    COMP_LOOP_1_modExp_1_while_C_14 = 11'd65,
    COMP_LOOP_1_modExp_1_while_C_15 = 11'd66,
    COMP_LOOP_1_modExp_1_while_C_16 = 11'd67,
    COMP_LOOP_1_modExp_1_while_C_17 = 11'd68,
    COMP_LOOP_1_modExp_1_while_C_18 = 11'd69,
    COMP_LOOP_1_modExp_1_while_C_19 = 11'd70,
    COMP_LOOP_1_modExp_1_while_C_20 = 11'd71,
    COMP_LOOP_1_modExp_1_while_C_21 = 11'd72,
    COMP_LOOP_1_modExp_1_while_C_22 = 11'd73,
    COMP_LOOP_1_modExp_1_while_C_23 = 11'd74,
    COMP_LOOP_1_modExp_1_while_C_24 = 11'd75,
    COMP_LOOP_1_modExp_1_while_C_25 = 11'd76,
    COMP_LOOP_1_modExp_1_while_C_26 = 11'd77,
    COMP_LOOP_1_modExp_1_while_C_27 = 11'd78,
    COMP_LOOP_1_modExp_1_while_C_28 = 11'd79,
    COMP_LOOP_1_modExp_1_while_C_29 = 11'd80,
    COMP_LOOP_1_modExp_1_while_C_30 = 11'd81,
    COMP_LOOP_1_modExp_1_while_C_31 = 11'd82,
    COMP_LOOP_1_modExp_1_while_C_32 = 11'd83,
    COMP_LOOP_1_modExp_1_while_C_33 = 11'd84,
    COMP_LOOP_1_modExp_1_while_C_34 = 11'd85,
    COMP_LOOP_1_modExp_1_while_C_35 = 11'd86,
    COMP_LOOP_1_modExp_1_while_C_36 = 11'd87,
    COMP_LOOP_1_modExp_1_while_C_37 = 11'd88,
    COMP_LOOP_1_modExp_1_while_C_38 = 11'd89,
    COMP_LOOP_C_2 = 11'd90,
    COMP_LOOP_C_3 = 11'd91,
    COMP_LOOP_C_4 = 11'd92,
    COMP_LOOP_C_5 = 11'd93,
    COMP_LOOP_C_6 = 11'd94,
    COMP_LOOP_C_7 = 11'd95,
    COMP_LOOP_C_8 = 11'd96,
    COMP_LOOP_C_9 = 11'd97,
    COMP_LOOP_C_10 = 11'd98,
    COMP_LOOP_C_11 = 11'd99,
    COMP_LOOP_C_12 = 11'd100,
    COMP_LOOP_C_13 = 11'd101,
    COMP_LOOP_C_14 = 11'd102,
    COMP_LOOP_C_15 = 11'd103,
    COMP_LOOP_C_16 = 11'd104,
    COMP_LOOP_C_17 = 11'd105,
    COMP_LOOP_C_18 = 11'd106,
    COMP_LOOP_C_19 = 11'd107,
    COMP_LOOP_C_20 = 11'd108,
    COMP_LOOP_C_21 = 11'd109,
    COMP_LOOP_C_22 = 11'd110,
    COMP_LOOP_C_23 = 11'd111,
    COMP_LOOP_C_24 = 11'd112,
    COMP_LOOP_C_25 = 11'd113,
    COMP_LOOP_C_26 = 11'd114,
    COMP_LOOP_C_27 = 11'd115,
    COMP_LOOP_C_28 = 11'd116,
    COMP_LOOP_C_29 = 11'd117,
    COMP_LOOP_C_30 = 11'd118,
    COMP_LOOP_C_31 = 11'd119,
    COMP_LOOP_C_32 = 11'd120,
    COMP_LOOP_C_33 = 11'd121,
    COMP_LOOP_C_34 = 11'd122,
    COMP_LOOP_C_35 = 11'd123,
    COMP_LOOP_C_36 = 11'd124,
    COMP_LOOP_C_37 = 11'd125,
    COMP_LOOP_C_38 = 11'd126,
    COMP_LOOP_C_39 = 11'd127,
    COMP_LOOP_C_40 = 11'd128,
    COMP_LOOP_C_41 = 11'd129,
    COMP_LOOP_C_42 = 11'd130,
    COMP_LOOP_C_43 = 11'd131,
    COMP_LOOP_C_44 = 11'd132,
    COMP_LOOP_C_45 = 11'd133,
    COMP_LOOP_C_46 = 11'd134,
    COMP_LOOP_C_47 = 11'd135,
    COMP_LOOP_C_48 = 11'd136,
    COMP_LOOP_C_49 = 11'd137,
    COMP_LOOP_C_50 = 11'd138,
    COMP_LOOP_C_51 = 11'd139,
    COMP_LOOP_C_52 = 11'd140,
    COMP_LOOP_C_53 = 11'd141,
    COMP_LOOP_C_54 = 11'd142,
    COMP_LOOP_C_55 = 11'd143,
    COMP_LOOP_C_56 = 11'd144,
    COMP_LOOP_C_57 = 11'd145,
    COMP_LOOP_C_58 = 11'd146,
    COMP_LOOP_C_59 = 11'd147,
    COMP_LOOP_C_60 = 11'd148,
    COMP_LOOP_C_61 = 11'd149,
    COMP_LOOP_C_62 = 11'd150,
    COMP_LOOP_C_63 = 11'd151,
    COMP_LOOP_C_64 = 11'd152,
    COMP_LOOP_C_65 = 11'd153,
    COMP_LOOP_2_modExp_1_while_C_0 = 11'd154,
    COMP_LOOP_2_modExp_1_while_C_1 = 11'd155,
    COMP_LOOP_2_modExp_1_while_C_2 = 11'd156,
    COMP_LOOP_2_modExp_1_while_C_3 = 11'd157,
    COMP_LOOP_2_modExp_1_while_C_4 = 11'd158,
    COMP_LOOP_2_modExp_1_while_C_5 = 11'd159,
    COMP_LOOP_2_modExp_1_while_C_6 = 11'd160,
    COMP_LOOP_2_modExp_1_while_C_7 = 11'd161,
    COMP_LOOP_2_modExp_1_while_C_8 = 11'd162,
    COMP_LOOP_2_modExp_1_while_C_9 = 11'd163,
    COMP_LOOP_2_modExp_1_while_C_10 = 11'd164,
    COMP_LOOP_2_modExp_1_while_C_11 = 11'd165,
    COMP_LOOP_2_modExp_1_while_C_12 = 11'd166,
    COMP_LOOP_2_modExp_1_while_C_13 = 11'd167,
    COMP_LOOP_2_modExp_1_while_C_14 = 11'd168,
    COMP_LOOP_2_modExp_1_while_C_15 = 11'd169,
    COMP_LOOP_2_modExp_1_while_C_16 = 11'd170,
    COMP_LOOP_2_modExp_1_while_C_17 = 11'd171,
    COMP_LOOP_2_modExp_1_while_C_18 = 11'd172,
    COMP_LOOP_2_modExp_1_while_C_19 = 11'd173,
    COMP_LOOP_2_modExp_1_while_C_20 = 11'd174,
    COMP_LOOP_2_modExp_1_while_C_21 = 11'd175,
    COMP_LOOP_2_modExp_1_while_C_22 = 11'd176,
    COMP_LOOP_2_modExp_1_while_C_23 = 11'd177,
    COMP_LOOP_2_modExp_1_while_C_24 = 11'd178,
    COMP_LOOP_2_modExp_1_while_C_25 = 11'd179,
    COMP_LOOP_2_modExp_1_while_C_26 = 11'd180,
    COMP_LOOP_2_modExp_1_while_C_27 = 11'd181,
    COMP_LOOP_2_modExp_1_while_C_28 = 11'd182,
    COMP_LOOP_2_modExp_1_while_C_29 = 11'd183,
    COMP_LOOP_2_modExp_1_while_C_30 = 11'd184,
    COMP_LOOP_2_modExp_1_while_C_31 = 11'd185,
    COMP_LOOP_2_modExp_1_while_C_32 = 11'd186,
    COMP_LOOP_2_modExp_1_while_C_33 = 11'd187,
    COMP_LOOP_2_modExp_1_while_C_34 = 11'd188,
    COMP_LOOP_2_modExp_1_while_C_35 = 11'd189,
    COMP_LOOP_2_modExp_1_while_C_36 = 11'd190,
    COMP_LOOP_2_modExp_1_while_C_37 = 11'd191,
    COMP_LOOP_2_modExp_1_while_C_38 = 11'd192,
    COMP_LOOP_C_66 = 11'd193,
    COMP_LOOP_C_67 = 11'd194,
    COMP_LOOP_C_68 = 11'd195,
    COMP_LOOP_C_69 = 11'd196,
    COMP_LOOP_C_70 = 11'd197,
    COMP_LOOP_C_71 = 11'd198,
    COMP_LOOP_C_72 = 11'd199,
    COMP_LOOP_C_73 = 11'd200,
    COMP_LOOP_C_74 = 11'd201,
    COMP_LOOP_C_75 = 11'd202,
    COMP_LOOP_C_76 = 11'd203,
    COMP_LOOP_C_77 = 11'd204,
    COMP_LOOP_C_78 = 11'd205,
    COMP_LOOP_C_79 = 11'd206,
    COMP_LOOP_C_80 = 11'd207,
    COMP_LOOP_C_81 = 11'd208,
    COMP_LOOP_C_82 = 11'd209,
    COMP_LOOP_C_83 = 11'd210,
    COMP_LOOP_C_84 = 11'd211,
    COMP_LOOP_C_85 = 11'd212,
    COMP_LOOP_C_86 = 11'd213,
    COMP_LOOP_C_87 = 11'd214,
    COMP_LOOP_C_88 = 11'd215,
    COMP_LOOP_C_89 = 11'd216,
    COMP_LOOP_C_90 = 11'd217,
    COMP_LOOP_C_91 = 11'd218,
    COMP_LOOP_C_92 = 11'd219,
    COMP_LOOP_C_93 = 11'd220,
    COMP_LOOP_C_94 = 11'd221,
    COMP_LOOP_C_95 = 11'd222,
    COMP_LOOP_C_96 = 11'd223,
    COMP_LOOP_C_97 = 11'd224,
    COMP_LOOP_C_98 = 11'd225,
    COMP_LOOP_C_99 = 11'd226,
    COMP_LOOP_C_100 = 11'd227,
    COMP_LOOP_C_101 = 11'd228,
    COMP_LOOP_C_102 = 11'd229,
    COMP_LOOP_C_103 = 11'd230,
    COMP_LOOP_C_104 = 11'd231,
    COMP_LOOP_C_105 = 11'd232,
    COMP_LOOP_C_106 = 11'd233,
    COMP_LOOP_C_107 = 11'd234,
    COMP_LOOP_C_108 = 11'd235,
    COMP_LOOP_C_109 = 11'd236,
    COMP_LOOP_C_110 = 11'd237,
    COMP_LOOP_C_111 = 11'd238,
    COMP_LOOP_C_112 = 11'd239,
    COMP_LOOP_C_113 = 11'd240,
    COMP_LOOP_C_114 = 11'd241,
    COMP_LOOP_C_115 = 11'd242,
    COMP_LOOP_C_116 = 11'd243,
    COMP_LOOP_C_117 = 11'd244,
    COMP_LOOP_C_118 = 11'd245,
    COMP_LOOP_C_119 = 11'd246,
    COMP_LOOP_C_120 = 11'd247,
    COMP_LOOP_C_121 = 11'd248,
    COMP_LOOP_C_122 = 11'd249,
    COMP_LOOP_C_123 = 11'd250,
    COMP_LOOP_C_124 = 11'd251,
    COMP_LOOP_C_125 = 11'd252,
    COMP_LOOP_C_126 = 11'd253,
    COMP_LOOP_C_127 = 11'd254,
    COMP_LOOP_C_128 = 11'd255,
    COMP_LOOP_C_129 = 11'd256,
    COMP_LOOP_3_modExp_1_while_C_0 = 11'd257,
    COMP_LOOP_3_modExp_1_while_C_1 = 11'd258,
    COMP_LOOP_3_modExp_1_while_C_2 = 11'd259,
    COMP_LOOP_3_modExp_1_while_C_3 = 11'd260,
    COMP_LOOP_3_modExp_1_while_C_4 = 11'd261,
    COMP_LOOP_3_modExp_1_while_C_5 = 11'd262,
    COMP_LOOP_3_modExp_1_while_C_6 = 11'd263,
    COMP_LOOP_3_modExp_1_while_C_7 = 11'd264,
    COMP_LOOP_3_modExp_1_while_C_8 = 11'd265,
    COMP_LOOP_3_modExp_1_while_C_9 = 11'd266,
    COMP_LOOP_3_modExp_1_while_C_10 = 11'd267,
    COMP_LOOP_3_modExp_1_while_C_11 = 11'd268,
    COMP_LOOP_3_modExp_1_while_C_12 = 11'd269,
    COMP_LOOP_3_modExp_1_while_C_13 = 11'd270,
    COMP_LOOP_3_modExp_1_while_C_14 = 11'd271,
    COMP_LOOP_3_modExp_1_while_C_15 = 11'd272,
    COMP_LOOP_3_modExp_1_while_C_16 = 11'd273,
    COMP_LOOP_3_modExp_1_while_C_17 = 11'd274,
    COMP_LOOP_3_modExp_1_while_C_18 = 11'd275,
    COMP_LOOP_3_modExp_1_while_C_19 = 11'd276,
    COMP_LOOP_3_modExp_1_while_C_20 = 11'd277,
    COMP_LOOP_3_modExp_1_while_C_21 = 11'd278,
    COMP_LOOP_3_modExp_1_while_C_22 = 11'd279,
    COMP_LOOP_3_modExp_1_while_C_23 = 11'd280,
    COMP_LOOP_3_modExp_1_while_C_24 = 11'd281,
    COMP_LOOP_3_modExp_1_while_C_25 = 11'd282,
    COMP_LOOP_3_modExp_1_while_C_26 = 11'd283,
    COMP_LOOP_3_modExp_1_while_C_27 = 11'd284,
    COMP_LOOP_3_modExp_1_while_C_28 = 11'd285,
    COMP_LOOP_3_modExp_1_while_C_29 = 11'd286,
    COMP_LOOP_3_modExp_1_while_C_30 = 11'd287,
    COMP_LOOP_3_modExp_1_while_C_31 = 11'd288,
    COMP_LOOP_3_modExp_1_while_C_32 = 11'd289,
    COMP_LOOP_3_modExp_1_while_C_33 = 11'd290,
    COMP_LOOP_3_modExp_1_while_C_34 = 11'd291,
    COMP_LOOP_3_modExp_1_while_C_35 = 11'd292,
    COMP_LOOP_3_modExp_1_while_C_36 = 11'd293,
    COMP_LOOP_3_modExp_1_while_C_37 = 11'd294,
    COMP_LOOP_3_modExp_1_while_C_38 = 11'd295,
    COMP_LOOP_C_130 = 11'd296,
    COMP_LOOP_C_131 = 11'd297,
    COMP_LOOP_C_132 = 11'd298,
    COMP_LOOP_C_133 = 11'd299,
    COMP_LOOP_C_134 = 11'd300,
    COMP_LOOP_C_135 = 11'd301,
    COMP_LOOP_C_136 = 11'd302,
    COMP_LOOP_C_137 = 11'd303,
    COMP_LOOP_C_138 = 11'd304,
    COMP_LOOP_C_139 = 11'd305,
    COMP_LOOP_C_140 = 11'd306,
    COMP_LOOP_C_141 = 11'd307,
    COMP_LOOP_C_142 = 11'd308,
    COMP_LOOP_C_143 = 11'd309,
    COMP_LOOP_C_144 = 11'd310,
    COMP_LOOP_C_145 = 11'd311,
    COMP_LOOP_C_146 = 11'd312,
    COMP_LOOP_C_147 = 11'd313,
    COMP_LOOP_C_148 = 11'd314,
    COMP_LOOP_C_149 = 11'd315,
    COMP_LOOP_C_150 = 11'd316,
    COMP_LOOP_C_151 = 11'd317,
    COMP_LOOP_C_152 = 11'd318,
    COMP_LOOP_C_153 = 11'd319,
    COMP_LOOP_C_154 = 11'd320,
    COMP_LOOP_C_155 = 11'd321,
    COMP_LOOP_C_156 = 11'd322,
    COMP_LOOP_C_157 = 11'd323,
    COMP_LOOP_C_158 = 11'd324,
    COMP_LOOP_C_159 = 11'd325,
    COMP_LOOP_C_160 = 11'd326,
    COMP_LOOP_C_161 = 11'd327,
    COMP_LOOP_C_162 = 11'd328,
    COMP_LOOP_C_163 = 11'd329,
    COMP_LOOP_C_164 = 11'd330,
    COMP_LOOP_C_165 = 11'd331,
    COMP_LOOP_C_166 = 11'd332,
    COMP_LOOP_C_167 = 11'd333,
    COMP_LOOP_C_168 = 11'd334,
    COMP_LOOP_C_169 = 11'd335,
    COMP_LOOP_C_170 = 11'd336,
    COMP_LOOP_C_171 = 11'd337,
    COMP_LOOP_C_172 = 11'd338,
    COMP_LOOP_C_173 = 11'd339,
    COMP_LOOP_C_174 = 11'd340,
    COMP_LOOP_C_175 = 11'd341,
    COMP_LOOP_C_176 = 11'd342,
    COMP_LOOP_C_177 = 11'd343,
    COMP_LOOP_C_178 = 11'd344,
    COMP_LOOP_C_179 = 11'd345,
    COMP_LOOP_C_180 = 11'd346,
    COMP_LOOP_C_181 = 11'd347,
    COMP_LOOP_C_182 = 11'd348,
    COMP_LOOP_C_183 = 11'd349,
    COMP_LOOP_C_184 = 11'd350,
    COMP_LOOP_C_185 = 11'd351,
    COMP_LOOP_C_186 = 11'd352,
    COMP_LOOP_C_187 = 11'd353,
    COMP_LOOP_C_188 = 11'd354,
    COMP_LOOP_C_189 = 11'd355,
    COMP_LOOP_C_190 = 11'd356,
    COMP_LOOP_C_191 = 11'd357,
    COMP_LOOP_C_192 = 11'd358,
    COMP_LOOP_C_193 = 11'd359,
    COMP_LOOP_4_modExp_1_while_C_0 = 11'd360,
    COMP_LOOP_4_modExp_1_while_C_1 = 11'd361,
    COMP_LOOP_4_modExp_1_while_C_2 = 11'd362,
    COMP_LOOP_4_modExp_1_while_C_3 = 11'd363,
    COMP_LOOP_4_modExp_1_while_C_4 = 11'd364,
    COMP_LOOP_4_modExp_1_while_C_5 = 11'd365,
    COMP_LOOP_4_modExp_1_while_C_6 = 11'd366,
    COMP_LOOP_4_modExp_1_while_C_7 = 11'd367,
    COMP_LOOP_4_modExp_1_while_C_8 = 11'd368,
    COMP_LOOP_4_modExp_1_while_C_9 = 11'd369,
    COMP_LOOP_4_modExp_1_while_C_10 = 11'd370,
    COMP_LOOP_4_modExp_1_while_C_11 = 11'd371,
    COMP_LOOP_4_modExp_1_while_C_12 = 11'd372,
    COMP_LOOP_4_modExp_1_while_C_13 = 11'd373,
    COMP_LOOP_4_modExp_1_while_C_14 = 11'd374,
    COMP_LOOP_4_modExp_1_while_C_15 = 11'd375,
    COMP_LOOP_4_modExp_1_while_C_16 = 11'd376,
    COMP_LOOP_4_modExp_1_while_C_17 = 11'd377,
    COMP_LOOP_4_modExp_1_while_C_18 = 11'd378,
    COMP_LOOP_4_modExp_1_while_C_19 = 11'd379,
    COMP_LOOP_4_modExp_1_while_C_20 = 11'd380,
    COMP_LOOP_4_modExp_1_while_C_21 = 11'd381,
    COMP_LOOP_4_modExp_1_while_C_22 = 11'd382,
    COMP_LOOP_4_modExp_1_while_C_23 = 11'd383,
    COMP_LOOP_4_modExp_1_while_C_24 = 11'd384,
    COMP_LOOP_4_modExp_1_while_C_25 = 11'd385,
    COMP_LOOP_4_modExp_1_while_C_26 = 11'd386,
    COMP_LOOP_4_modExp_1_while_C_27 = 11'd387,
    COMP_LOOP_4_modExp_1_while_C_28 = 11'd388,
    COMP_LOOP_4_modExp_1_while_C_29 = 11'd389,
    COMP_LOOP_4_modExp_1_while_C_30 = 11'd390,
    COMP_LOOP_4_modExp_1_while_C_31 = 11'd391,
    COMP_LOOP_4_modExp_1_while_C_32 = 11'd392,
    COMP_LOOP_4_modExp_1_while_C_33 = 11'd393,
    COMP_LOOP_4_modExp_1_while_C_34 = 11'd394,
    COMP_LOOP_4_modExp_1_while_C_35 = 11'd395,
    COMP_LOOP_4_modExp_1_while_C_36 = 11'd396,
    COMP_LOOP_4_modExp_1_while_C_37 = 11'd397,
    COMP_LOOP_4_modExp_1_while_C_38 = 11'd398,
    COMP_LOOP_C_194 = 11'd399,
    COMP_LOOP_C_195 = 11'd400,
    COMP_LOOP_C_196 = 11'd401,
    COMP_LOOP_C_197 = 11'd402,
    COMP_LOOP_C_198 = 11'd403,
    COMP_LOOP_C_199 = 11'd404,
    COMP_LOOP_C_200 = 11'd405,
    COMP_LOOP_C_201 = 11'd406,
    COMP_LOOP_C_202 = 11'd407,
    COMP_LOOP_C_203 = 11'd408,
    COMP_LOOP_C_204 = 11'd409,
    COMP_LOOP_C_205 = 11'd410,
    COMP_LOOP_C_206 = 11'd411,
    COMP_LOOP_C_207 = 11'd412,
    COMP_LOOP_C_208 = 11'd413,
    COMP_LOOP_C_209 = 11'd414,
    COMP_LOOP_C_210 = 11'd415,
    COMP_LOOP_C_211 = 11'd416,
    COMP_LOOP_C_212 = 11'd417,
    COMP_LOOP_C_213 = 11'd418,
    COMP_LOOP_C_214 = 11'd419,
    COMP_LOOP_C_215 = 11'd420,
    COMP_LOOP_C_216 = 11'd421,
    COMP_LOOP_C_217 = 11'd422,
    COMP_LOOP_C_218 = 11'd423,
    COMP_LOOP_C_219 = 11'd424,
    COMP_LOOP_C_220 = 11'd425,
    COMP_LOOP_C_221 = 11'd426,
    COMP_LOOP_C_222 = 11'd427,
    COMP_LOOP_C_223 = 11'd428,
    COMP_LOOP_C_224 = 11'd429,
    COMP_LOOP_C_225 = 11'd430,
    COMP_LOOP_C_226 = 11'd431,
    COMP_LOOP_C_227 = 11'd432,
    COMP_LOOP_C_228 = 11'd433,
    COMP_LOOP_C_229 = 11'd434,
    COMP_LOOP_C_230 = 11'd435,
    COMP_LOOP_C_231 = 11'd436,
    COMP_LOOP_C_232 = 11'd437,
    COMP_LOOP_C_233 = 11'd438,
    COMP_LOOP_C_234 = 11'd439,
    COMP_LOOP_C_235 = 11'd440,
    COMP_LOOP_C_236 = 11'd441,
    COMP_LOOP_C_237 = 11'd442,
    COMP_LOOP_C_238 = 11'd443,
    COMP_LOOP_C_239 = 11'd444,
    COMP_LOOP_C_240 = 11'd445,
    COMP_LOOP_C_241 = 11'd446,
    COMP_LOOP_C_242 = 11'd447,
    COMP_LOOP_C_243 = 11'd448,
    COMP_LOOP_C_244 = 11'd449,
    COMP_LOOP_C_245 = 11'd450,
    COMP_LOOP_C_246 = 11'd451,
    COMP_LOOP_C_247 = 11'd452,
    COMP_LOOP_C_248 = 11'd453,
    COMP_LOOP_C_249 = 11'd454,
    COMP_LOOP_C_250 = 11'd455,
    COMP_LOOP_C_251 = 11'd456,
    COMP_LOOP_C_252 = 11'd457,
    COMP_LOOP_C_253 = 11'd458,
    COMP_LOOP_C_254 = 11'd459,
    COMP_LOOP_C_255 = 11'd460,
    COMP_LOOP_C_256 = 11'd461,
    COMP_LOOP_C_257 = 11'd462,
    COMP_LOOP_5_modExp_1_while_C_0 = 11'd463,
    COMP_LOOP_5_modExp_1_while_C_1 = 11'd464,
    COMP_LOOP_5_modExp_1_while_C_2 = 11'd465,
    COMP_LOOP_5_modExp_1_while_C_3 = 11'd466,
    COMP_LOOP_5_modExp_1_while_C_4 = 11'd467,
    COMP_LOOP_5_modExp_1_while_C_5 = 11'd468,
    COMP_LOOP_5_modExp_1_while_C_6 = 11'd469,
    COMP_LOOP_5_modExp_1_while_C_7 = 11'd470,
    COMP_LOOP_5_modExp_1_while_C_8 = 11'd471,
    COMP_LOOP_5_modExp_1_while_C_9 = 11'd472,
    COMP_LOOP_5_modExp_1_while_C_10 = 11'd473,
    COMP_LOOP_5_modExp_1_while_C_11 = 11'd474,
    COMP_LOOP_5_modExp_1_while_C_12 = 11'd475,
    COMP_LOOP_5_modExp_1_while_C_13 = 11'd476,
    COMP_LOOP_5_modExp_1_while_C_14 = 11'd477,
    COMP_LOOP_5_modExp_1_while_C_15 = 11'd478,
    COMP_LOOP_5_modExp_1_while_C_16 = 11'd479,
    COMP_LOOP_5_modExp_1_while_C_17 = 11'd480,
    COMP_LOOP_5_modExp_1_while_C_18 = 11'd481,
    COMP_LOOP_5_modExp_1_while_C_19 = 11'd482,
    COMP_LOOP_5_modExp_1_while_C_20 = 11'd483,
    COMP_LOOP_5_modExp_1_while_C_21 = 11'd484,
    COMP_LOOP_5_modExp_1_while_C_22 = 11'd485,
    COMP_LOOP_5_modExp_1_while_C_23 = 11'd486,
    COMP_LOOP_5_modExp_1_while_C_24 = 11'd487,
    COMP_LOOP_5_modExp_1_while_C_25 = 11'd488,
    COMP_LOOP_5_modExp_1_while_C_26 = 11'd489,
    COMP_LOOP_5_modExp_1_while_C_27 = 11'd490,
    COMP_LOOP_5_modExp_1_while_C_28 = 11'd491,
    COMP_LOOP_5_modExp_1_while_C_29 = 11'd492,
    COMP_LOOP_5_modExp_1_while_C_30 = 11'd493,
    COMP_LOOP_5_modExp_1_while_C_31 = 11'd494,
    COMP_LOOP_5_modExp_1_while_C_32 = 11'd495,
    COMP_LOOP_5_modExp_1_while_C_33 = 11'd496,
    COMP_LOOP_5_modExp_1_while_C_34 = 11'd497,
    COMP_LOOP_5_modExp_1_while_C_35 = 11'd498,
    COMP_LOOP_5_modExp_1_while_C_36 = 11'd499,
    COMP_LOOP_5_modExp_1_while_C_37 = 11'd500,
    COMP_LOOP_5_modExp_1_while_C_38 = 11'd501,
    COMP_LOOP_C_258 = 11'd502,
    COMP_LOOP_C_259 = 11'd503,
    COMP_LOOP_C_260 = 11'd504,
    COMP_LOOP_C_261 = 11'd505,
    COMP_LOOP_C_262 = 11'd506,
    COMP_LOOP_C_263 = 11'd507,
    COMP_LOOP_C_264 = 11'd508,
    COMP_LOOP_C_265 = 11'd509,
    COMP_LOOP_C_266 = 11'd510,
    COMP_LOOP_C_267 = 11'd511,
    COMP_LOOP_C_268 = 11'd512,
    COMP_LOOP_C_269 = 11'd513,
    COMP_LOOP_C_270 = 11'd514,
    COMP_LOOP_C_271 = 11'd515,
    COMP_LOOP_C_272 = 11'd516,
    COMP_LOOP_C_273 = 11'd517,
    COMP_LOOP_C_274 = 11'd518,
    COMP_LOOP_C_275 = 11'd519,
    COMP_LOOP_C_276 = 11'd520,
    COMP_LOOP_C_277 = 11'd521,
    COMP_LOOP_C_278 = 11'd522,
    COMP_LOOP_C_279 = 11'd523,
    COMP_LOOP_C_280 = 11'd524,
    COMP_LOOP_C_281 = 11'd525,
    COMP_LOOP_C_282 = 11'd526,
    COMP_LOOP_C_283 = 11'd527,
    COMP_LOOP_C_284 = 11'd528,
    COMP_LOOP_C_285 = 11'd529,
    COMP_LOOP_C_286 = 11'd530,
    COMP_LOOP_C_287 = 11'd531,
    COMP_LOOP_C_288 = 11'd532,
    COMP_LOOP_C_289 = 11'd533,
    COMP_LOOP_C_290 = 11'd534,
    COMP_LOOP_C_291 = 11'd535,
    COMP_LOOP_C_292 = 11'd536,
    COMP_LOOP_C_293 = 11'd537,
    COMP_LOOP_C_294 = 11'd538,
    COMP_LOOP_C_295 = 11'd539,
    COMP_LOOP_C_296 = 11'd540,
    COMP_LOOP_C_297 = 11'd541,
    COMP_LOOP_C_298 = 11'd542,
    COMP_LOOP_C_299 = 11'd543,
    COMP_LOOP_C_300 = 11'd544,
    COMP_LOOP_C_301 = 11'd545,
    COMP_LOOP_C_302 = 11'd546,
    COMP_LOOP_C_303 = 11'd547,
    COMP_LOOP_C_304 = 11'd548,
    COMP_LOOP_C_305 = 11'd549,
    COMP_LOOP_C_306 = 11'd550,
    COMP_LOOP_C_307 = 11'd551,
    COMP_LOOP_C_308 = 11'd552,
    COMP_LOOP_C_309 = 11'd553,
    COMP_LOOP_C_310 = 11'd554,
    COMP_LOOP_C_311 = 11'd555,
    COMP_LOOP_C_312 = 11'd556,
    COMP_LOOP_C_313 = 11'd557,
    COMP_LOOP_C_314 = 11'd558,
    COMP_LOOP_C_315 = 11'd559,
    COMP_LOOP_C_316 = 11'd560,
    COMP_LOOP_C_317 = 11'd561,
    COMP_LOOP_C_318 = 11'd562,
    COMP_LOOP_C_319 = 11'd563,
    COMP_LOOP_C_320 = 11'd564,
    COMP_LOOP_C_321 = 11'd565,
    COMP_LOOP_6_modExp_1_while_C_0 = 11'd566,
    COMP_LOOP_6_modExp_1_while_C_1 = 11'd567,
    COMP_LOOP_6_modExp_1_while_C_2 = 11'd568,
    COMP_LOOP_6_modExp_1_while_C_3 = 11'd569,
    COMP_LOOP_6_modExp_1_while_C_4 = 11'd570,
    COMP_LOOP_6_modExp_1_while_C_5 = 11'd571,
    COMP_LOOP_6_modExp_1_while_C_6 = 11'd572,
    COMP_LOOP_6_modExp_1_while_C_7 = 11'd573,
    COMP_LOOP_6_modExp_1_while_C_8 = 11'd574,
    COMP_LOOP_6_modExp_1_while_C_9 = 11'd575,
    COMP_LOOP_6_modExp_1_while_C_10 = 11'd576,
    COMP_LOOP_6_modExp_1_while_C_11 = 11'd577,
    COMP_LOOP_6_modExp_1_while_C_12 = 11'd578,
    COMP_LOOP_6_modExp_1_while_C_13 = 11'd579,
    COMP_LOOP_6_modExp_1_while_C_14 = 11'd580,
    COMP_LOOP_6_modExp_1_while_C_15 = 11'd581,
    COMP_LOOP_6_modExp_1_while_C_16 = 11'd582,
    COMP_LOOP_6_modExp_1_while_C_17 = 11'd583,
    COMP_LOOP_6_modExp_1_while_C_18 = 11'd584,
    COMP_LOOP_6_modExp_1_while_C_19 = 11'd585,
    COMP_LOOP_6_modExp_1_while_C_20 = 11'd586,
    COMP_LOOP_6_modExp_1_while_C_21 = 11'd587,
    COMP_LOOP_6_modExp_1_while_C_22 = 11'd588,
    COMP_LOOP_6_modExp_1_while_C_23 = 11'd589,
    COMP_LOOP_6_modExp_1_while_C_24 = 11'd590,
    COMP_LOOP_6_modExp_1_while_C_25 = 11'd591,
    COMP_LOOP_6_modExp_1_while_C_26 = 11'd592,
    COMP_LOOP_6_modExp_1_while_C_27 = 11'd593,
    COMP_LOOP_6_modExp_1_while_C_28 = 11'd594,
    COMP_LOOP_6_modExp_1_while_C_29 = 11'd595,
    COMP_LOOP_6_modExp_1_while_C_30 = 11'd596,
    COMP_LOOP_6_modExp_1_while_C_31 = 11'd597,
    COMP_LOOP_6_modExp_1_while_C_32 = 11'd598,
    COMP_LOOP_6_modExp_1_while_C_33 = 11'd599,
    COMP_LOOP_6_modExp_1_while_C_34 = 11'd600,
    COMP_LOOP_6_modExp_1_while_C_35 = 11'd601,
    COMP_LOOP_6_modExp_1_while_C_36 = 11'd602,
    COMP_LOOP_6_modExp_1_while_C_37 = 11'd603,
    COMP_LOOP_6_modExp_1_while_C_38 = 11'd604,
    COMP_LOOP_C_322 = 11'd605,
    COMP_LOOP_C_323 = 11'd606,
    COMP_LOOP_C_324 = 11'd607,
    COMP_LOOP_C_325 = 11'd608,
    COMP_LOOP_C_326 = 11'd609,
    COMP_LOOP_C_327 = 11'd610,
    COMP_LOOP_C_328 = 11'd611,
    COMP_LOOP_C_329 = 11'd612,
    COMP_LOOP_C_330 = 11'd613,
    COMP_LOOP_C_331 = 11'd614,
    COMP_LOOP_C_332 = 11'd615,
    COMP_LOOP_C_333 = 11'd616,
    COMP_LOOP_C_334 = 11'd617,
    COMP_LOOP_C_335 = 11'd618,
    COMP_LOOP_C_336 = 11'd619,
    COMP_LOOP_C_337 = 11'd620,
    COMP_LOOP_C_338 = 11'd621,
    COMP_LOOP_C_339 = 11'd622,
    COMP_LOOP_C_340 = 11'd623,
    COMP_LOOP_C_341 = 11'd624,
    COMP_LOOP_C_342 = 11'd625,
    COMP_LOOP_C_343 = 11'd626,
    COMP_LOOP_C_344 = 11'd627,
    COMP_LOOP_C_345 = 11'd628,
    COMP_LOOP_C_346 = 11'd629,
    COMP_LOOP_C_347 = 11'd630,
    COMP_LOOP_C_348 = 11'd631,
    COMP_LOOP_C_349 = 11'd632,
    COMP_LOOP_C_350 = 11'd633,
    COMP_LOOP_C_351 = 11'd634,
    COMP_LOOP_C_352 = 11'd635,
    COMP_LOOP_C_353 = 11'd636,
    COMP_LOOP_C_354 = 11'd637,
    COMP_LOOP_C_355 = 11'd638,
    COMP_LOOP_C_356 = 11'd639,
    COMP_LOOP_C_357 = 11'd640,
    COMP_LOOP_C_358 = 11'd641,
    COMP_LOOP_C_359 = 11'd642,
    COMP_LOOP_C_360 = 11'd643,
    COMP_LOOP_C_361 = 11'd644,
    COMP_LOOP_C_362 = 11'd645,
    COMP_LOOP_C_363 = 11'd646,
    COMP_LOOP_C_364 = 11'd647,
    COMP_LOOP_C_365 = 11'd648,
    COMP_LOOP_C_366 = 11'd649,
    COMP_LOOP_C_367 = 11'd650,
    COMP_LOOP_C_368 = 11'd651,
    COMP_LOOP_C_369 = 11'd652,
    COMP_LOOP_C_370 = 11'd653,
    COMP_LOOP_C_371 = 11'd654,
    COMP_LOOP_C_372 = 11'd655,
    COMP_LOOP_C_373 = 11'd656,
    COMP_LOOP_C_374 = 11'd657,
    COMP_LOOP_C_375 = 11'd658,
    COMP_LOOP_C_376 = 11'd659,
    COMP_LOOP_C_377 = 11'd660,
    COMP_LOOP_C_378 = 11'd661,
    COMP_LOOP_C_379 = 11'd662,
    COMP_LOOP_C_380 = 11'd663,
    COMP_LOOP_C_381 = 11'd664,
    COMP_LOOP_C_382 = 11'd665,
    COMP_LOOP_C_383 = 11'd666,
    COMP_LOOP_C_384 = 11'd667,
    COMP_LOOP_C_385 = 11'd668,
    COMP_LOOP_7_modExp_1_while_C_0 = 11'd669,
    COMP_LOOP_7_modExp_1_while_C_1 = 11'd670,
    COMP_LOOP_7_modExp_1_while_C_2 = 11'd671,
    COMP_LOOP_7_modExp_1_while_C_3 = 11'd672,
    COMP_LOOP_7_modExp_1_while_C_4 = 11'd673,
    COMP_LOOP_7_modExp_1_while_C_5 = 11'd674,
    COMP_LOOP_7_modExp_1_while_C_6 = 11'd675,
    COMP_LOOP_7_modExp_1_while_C_7 = 11'd676,
    COMP_LOOP_7_modExp_1_while_C_8 = 11'd677,
    COMP_LOOP_7_modExp_1_while_C_9 = 11'd678,
    COMP_LOOP_7_modExp_1_while_C_10 = 11'd679,
    COMP_LOOP_7_modExp_1_while_C_11 = 11'd680,
    COMP_LOOP_7_modExp_1_while_C_12 = 11'd681,
    COMP_LOOP_7_modExp_1_while_C_13 = 11'd682,
    COMP_LOOP_7_modExp_1_while_C_14 = 11'd683,
    COMP_LOOP_7_modExp_1_while_C_15 = 11'd684,
    COMP_LOOP_7_modExp_1_while_C_16 = 11'd685,
    COMP_LOOP_7_modExp_1_while_C_17 = 11'd686,
    COMP_LOOP_7_modExp_1_while_C_18 = 11'd687,
    COMP_LOOP_7_modExp_1_while_C_19 = 11'd688,
    COMP_LOOP_7_modExp_1_while_C_20 = 11'd689,
    COMP_LOOP_7_modExp_1_while_C_21 = 11'd690,
    COMP_LOOP_7_modExp_1_while_C_22 = 11'd691,
    COMP_LOOP_7_modExp_1_while_C_23 = 11'd692,
    COMP_LOOP_7_modExp_1_while_C_24 = 11'd693,
    COMP_LOOP_7_modExp_1_while_C_25 = 11'd694,
    COMP_LOOP_7_modExp_1_while_C_26 = 11'd695,
    COMP_LOOP_7_modExp_1_while_C_27 = 11'd696,
    COMP_LOOP_7_modExp_1_while_C_28 = 11'd697,
    COMP_LOOP_7_modExp_1_while_C_29 = 11'd698,
    COMP_LOOP_7_modExp_1_while_C_30 = 11'd699,
    COMP_LOOP_7_modExp_1_while_C_31 = 11'd700,
    COMP_LOOP_7_modExp_1_while_C_32 = 11'd701,
    COMP_LOOP_7_modExp_1_while_C_33 = 11'd702,
    COMP_LOOP_7_modExp_1_while_C_34 = 11'd703,
    COMP_LOOP_7_modExp_1_while_C_35 = 11'd704,
    COMP_LOOP_7_modExp_1_while_C_36 = 11'd705,
    COMP_LOOP_7_modExp_1_while_C_37 = 11'd706,
    COMP_LOOP_7_modExp_1_while_C_38 = 11'd707,
    COMP_LOOP_C_386 = 11'd708,
    COMP_LOOP_C_387 = 11'd709,
    COMP_LOOP_C_388 = 11'd710,
    COMP_LOOP_C_389 = 11'd711,
    COMP_LOOP_C_390 = 11'd712,
    COMP_LOOP_C_391 = 11'd713,
    COMP_LOOP_C_392 = 11'd714,
    COMP_LOOP_C_393 = 11'd715,
    COMP_LOOP_C_394 = 11'd716,
    COMP_LOOP_C_395 = 11'd717,
    COMP_LOOP_C_396 = 11'd718,
    COMP_LOOP_C_397 = 11'd719,
    COMP_LOOP_C_398 = 11'd720,
    COMP_LOOP_C_399 = 11'd721,
    COMP_LOOP_C_400 = 11'd722,
    COMP_LOOP_C_401 = 11'd723,
    COMP_LOOP_C_402 = 11'd724,
    COMP_LOOP_C_403 = 11'd725,
    COMP_LOOP_C_404 = 11'd726,
    COMP_LOOP_C_405 = 11'd727,
    COMP_LOOP_C_406 = 11'd728,
    COMP_LOOP_C_407 = 11'd729,
    COMP_LOOP_C_408 = 11'd730,
    COMP_LOOP_C_409 = 11'd731,
    COMP_LOOP_C_410 = 11'd732,
    COMP_LOOP_C_411 = 11'd733,
    COMP_LOOP_C_412 = 11'd734,
    COMP_LOOP_C_413 = 11'd735,
    COMP_LOOP_C_414 = 11'd736,
    COMP_LOOP_C_415 = 11'd737,
    COMP_LOOP_C_416 = 11'd738,
    COMP_LOOP_C_417 = 11'd739,
    COMP_LOOP_C_418 = 11'd740,
    COMP_LOOP_C_419 = 11'd741,
    COMP_LOOP_C_420 = 11'd742,
    COMP_LOOP_C_421 = 11'd743,
    COMP_LOOP_C_422 = 11'd744,
    COMP_LOOP_C_423 = 11'd745,
    COMP_LOOP_C_424 = 11'd746,
    COMP_LOOP_C_425 = 11'd747,
    COMP_LOOP_C_426 = 11'd748,
    COMP_LOOP_C_427 = 11'd749,
    COMP_LOOP_C_428 = 11'd750,
    COMP_LOOP_C_429 = 11'd751,
    COMP_LOOP_C_430 = 11'd752,
    COMP_LOOP_C_431 = 11'd753,
    COMP_LOOP_C_432 = 11'd754,
    COMP_LOOP_C_433 = 11'd755,
    COMP_LOOP_C_434 = 11'd756,
    COMP_LOOP_C_435 = 11'd757,
    COMP_LOOP_C_436 = 11'd758,
    COMP_LOOP_C_437 = 11'd759,
    COMP_LOOP_C_438 = 11'd760,
    COMP_LOOP_C_439 = 11'd761,
    COMP_LOOP_C_440 = 11'd762,
    COMP_LOOP_C_441 = 11'd763,
    COMP_LOOP_C_442 = 11'd764,
    COMP_LOOP_C_443 = 11'd765,
    COMP_LOOP_C_444 = 11'd766,
    COMP_LOOP_C_445 = 11'd767,
    COMP_LOOP_C_446 = 11'd768,
    COMP_LOOP_C_447 = 11'd769,
    COMP_LOOP_C_448 = 11'd770,
    COMP_LOOP_C_449 = 11'd771,
    COMP_LOOP_8_modExp_1_while_C_0 = 11'd772,
    COMP_LOOP_8_modExp_1_while_C_1 = 11'd773,
    COMP_LOOP_8_modExp_1_while_C_2 = 11'd774,
    COMP_LOOP_8_modExp_1_while_C_3 = 11'd775,
    COMP_LOOP_8_modExp_1_while_C_4 = 11'd776,
    COMP_LOOP_8_modExp_1_while_C_5 = 11'd777,
    COMP_LOOP_8_modExp_1_while_C_6 = 11'd778,
    COMP_LOOP_8_modExp_1_while_C_7 = 11'd779,
    COMP_LOOP_8_modExp_1_while_C_8 = 11'd780,
    COMP_LOOP_8_modExp_1_while_C_9 = 11'd781,
    COMP_LOOP_8_modExp_1_while_C_10 = 11'd782,
    COMP_LOOP_8_modExp_1_while_C_11 = 11'd783,
    COMP_LOOP_8_modExp_1_while_C_12 = 11'd784,
    COMP_LOOP_8_modExp_1_while_C_13 = 11'd785,
    COMP_LOOP_8_modExp_1_while_C_14 = 11'd786,
    COMP_LOOP_8_modExp_1_while_C_15 = 11'd787,
    COMP_LOOP_8_modExp_1_while_C_16 = 11'd788,
    COMP_LOOP_8_modExp_1_while_C_17 = 11'd789,
    COMP_LOOP_8_modExp_1_while_C_18 = 11'd790,
    COMP_LOOP_8_modExp_1_while_C_19 = 11'd791,
    COMP_LOOP_8_modExp_1_while_C_20 = 11'd792,
    COMP_LOOP_8_modExp_1_while_C_21 = 11'd793,
    COMP_LOOP_8_modExp_1_while_C_22 = 11'd794,
    COMP_LOOP_8_modExp_1_while_C_23 = 11'd795,
    COMP_LOOP_8_modExp_1_while_C_24 = 11'd796,
    COMP_LOOP_8_modExp_1_while_C_25 = 11'd797,
    COMP_LOOP_8_modExp_1_while_C_26 = 11'd798,
    COMP_LOOP_8_modExp_1_while_C_27 = 11'd799,
    COMP_LOOP_8_modExp_1_while_C_28 = 11'd800,
    COMP_LOOP_8_modExp_1_while_C_29 = 11'd801,
    COMP_LOOP_8_modExp_1_while_C_30 = 11'd802,
    COMP_LOOP_8_modExp_1_while_C_31 = 11'd803,
    COMP_LOOP_8_modExp_1_while_C_32 = 11'd804,
    COMP_LOOP_8_modExp_1_while_C_33 = 11'd805,
    COMP_LOOP_8_modExp_1_while_C_34 = 11'd806,
    COMP_LOOP_8_modExp_1_while_C_35 = 11'd807,
    COMP_LOOP_8_modExp_1_while_C_36 = 11'd808,
    COMP_LOOP_8_modExp_1_while_C_37 = 11'd809,
    COMP_LOOP_8_modExp_1_while_C_38 = 11'd810,
    COMP_LOOP_C_450 = 11'd811,
    COMP_LOOP_C_451 = 11'd812,
    COMP_LOOP_C_452 = 11'd813,
    COMP_LOOP_C_453 = 11'd814,
    COMP_LOOP_C_454 = 11'd815,
    COMP_LOOP_C_455 = 11'd816,
    COMP_LOOP_C_456 = 11'd817,
    COMP_LOOP_C_457 = 11'd818,
    COMP_LOOP_C_458 = 11'd819,
    COMP_LOOP_C_459 = 11'd820,
    COMP_LOOP_C_460 = 11'd821,
    COMP_LOOP_C_461 = 11'd822,
    COMP_LOOP_C_462 = 11'd823,
    COMP_LOOP_C_463 = 11'd824,
    COMP_LOOP_C_464 = 11'd825,
    COMP_LOOP_C_465 = 11'd826,
    COMP_LOOP_C_466 = 11'd827,
    COMP_LOOP_C_467 = 11'd828,
    COMP_LOOP_C_468 = 11'd829,
    COMP_LOOP_C_469 = 11'd830,
    COMP_LOOP_C_470 = 11'd831,
    COMP_LOOP_C_471 = 11'd832,
    COMP_LOOP_C_472 = 11'd833,
    COMP_LOOP_C_473 = 11'd834,
    COMP_LOOP_C_474 = 11'd835,
    COMP_LOOP_C_475 = 11'd836,
    COMP_LOOP_C_476 = 11'd837,
    COMP_LOOP_C_477 = 11'd838,
    COMP_LOOP_C_478 = 11'd839,
    COMP_LOOP_C_479 = 11'd840,
    COMP_LOOP_C_480 = 11'd841,
    COMP_LOOP_C_481 = 11'd842,
    COMP_LOOP_C_482 = 11'd843,
    COMP_LOOP_C_483 = 11'd844,
    COMP_LOOP_C_484 = 11'd845,
    COMP_LOOP_C_485 = 11'd846,
    COMP_LOOP_C_486 = 11'd847,
    COMP_LOOP_C_487 = 11'd848,
    COMP_LOOP_C_488 = 11'd849,
    COMP_LOOP_C_489 = 11'd850,
    COMP_LOOP_C_490 = 11'd851,
    COMP_LOOP_C_491 = 11'd852,
    COMP_LOOP_C_492 = 11'd853,
    COMP_LOOP_C_493 = 11'd854,
    COMP_LOOP_C_494 = 11'd855,
    COMP_LOOP_C_495 = 11'd856,
    COMP_LOOP_C_496 = 11'd857,
    COMP_LOOP_C_497 = 11'd858,
    COMP_LOOP_C_498 = 11'd859,
    COMP_LOOP_C_499 = 11'd860,
    COMP_LOOP_C_500 = 11'd861,
    COMP_LOOP_C_501 = 11'd862,
    COMP_LOOP_C_502 = 11'd863,
    COMP_LOOP_C_503 = 11'd864,
    COMP_LOOP_C_504 = 11'd865,
    COMP_LOOP_C_505 = 11'd866,
    COMP_LOOP_C_506 = 11'd867,
    COMP_LOOP_C_507 = 11'd868,
    COMP_LOOP_C_508 = 11'd869,
    COMP_LOOP_C_509 = 11'd870,
    COMP_LOOP_C_510 = 11'd871,
    COMP_LOOP_C_511 = 11'd872,
    COMP_LOOP_C_512 = 11'd873,
    COMP_LOOP_C_513 = 11'd874,
    COMP_LOOP_9_modExp_1_while_C_0 = 11'd875,
    COMP_LOOP_9_modExp_1_while_C_1 = 11'd876,
    COMP_LOOP_9_modExp_1_while_C_2 = 11'd877,
    COMP_LOOP_9_modExp_1_while_C_3 = 11'd878,
    COMP_LOOP_9_modExp_1_while_C_4 = 11'd879,
    COMP_LOOP_9_modExp_1_while_C_5 = 11'd880,
    COMP_LOOP_9_modExp_1_while_C_6 = 11'd881,
    COMP_LOOP_9_modExp_1_while_C_7 = 11'd882,
    COMP_LOOP_9_modExp_1_while_C_8 = 11'd883,
    COMP_LOOP_9_modExp_1_while_C_9 = 11'd884,
    COMP_LOOP_9_modExp_1_while_C_10 = 11'd885,
    COMP_LOOP_9_modExp_1_while_C_11 = 11'd886,
    COMP_LOOP_9_modExp_1_while_C_12 = 11'd887,
    COMP_LOOP_9_modExp_1_while_C_13 = 11'd888,
    COMP_LOOP_9_modExp_1_while_C_14 = 11'd889,
    COMP_LOOP_9_modExp_1_while_C_15 = 11'd890,
    COMP_LOOP_9_modExp_1_while_C_16 = 11'd891,
    COMP_LOOP_9_modExp_1_while_C_17 = 11'd892,
    COMP_LOOP_9_modExp_1_while_C_18 = 11'd893,
    COMP_LOOP_9_modExp_1_while_C_19 = 11'd894,
    COMP_LOOP_9_modExp_1_while_C_20 = 11'd895,
    COMP_LOOP_9_modExp_1_while_C_21 = 11'd896,
    COMP_LOOP_9_modExp_1_while_C_22 = 11'd897,
    COMP_LOOP_9_modExp_1_while_C_23 = 11'd898,
    COMP_LOOP_9_modExp_1_while_C_24 = 11'd899,
    COMP_LOOP_9_modExp_1_while_C_25 = 11'd900,
    COMP_LOOP_9_modExp_1_while_C_26 = 11'd901,
    COMP_LOOP_9_modExp_1_while_C_27 = 11'd902,
    COMP_LOOP_9_modExp_1_while_C_28 = 11'd903,
    COMP_LOOP_9_modExp_1_while_C_29 = 11'd904,
    COMP_LOOP_9_modExp_1_while_C_30 = 11'd905,
    COMP_LOOP_9_modExp_1_while_C_31 = 11'd906,
    COMP_LOOP_9_modExp_1_while_C_32 = 11'd907,
    COMP_LOOP_9_modExp_1_while_C_33 = 11'd908,
    COMP_LOOP_9_modExp_1_while_C_34 = 11'd909,
    COMP_LOOP_9_modExp_1_while_C_35 = 11'd910,
    COMP_LOOP_9_modExp_1_while_C_36 = 11'd911,
    COMP_LOOP_9_modExp_1_while_C_37 = 11'd912,
    COMP_LOOP_9_modExp_1_while_C_38 = 11'd913,
    COMP_LOOP_C_514 = 11'd914,
    COMP_LOOP_C_515 = 11'd915,
    COMP_LOOP_C_516 = 11'd916,
    COMP_LOOP_C_517 = 11'd917,
    COMP_LOOP_C_518 = 11'd918,
    COMP_LOOP_C_519 = 11'd919,
    COMP_LOOP_C_520 = 11'd920,
    COMP_LOOP_C_521 = 11'd921,
    COMP_LOOP_C_522 = 11'd922,
    COMP_LOOP_C_523 = 11'd923,
    COMP_LOOP_C_524 = 11'd924,
    COMP_LOOP_C_525 = 11'd925,
    COMP_LOOP_C_526 = 11'd926,
    COMP_LOOP_C_527 = 11'd927,
    COMP_LOOP_C_528 = 11'd928,
    COMP_LOOP_C_529 = 11'd929,
    COMP_LOOP_C_530 = 11'd930,
    COMP_LOOP_C_531 = 11'd931,
    COMP_LOOP_C_532 = 11'd932,
    COMP_LOOP_C_533 = 11'd933,
    COMP_LOOP_C_534 = 11'd934,
    COMP_LOOP_C_535 = 11'd935,
    COMP_LOOP_C_536 = 11'd936,
    COMP_LOOP_C_537 = 11'd937,
    COMP_LOOP_C_538 = 11'd938,
    COMP_LOOP_C_539 = 11'd939,
    COMP_LOOP_C_540 = 11'd940,
    COMP_LOOP_C_541 = 11'd941,
    COMP_LOOP_C_542 = 11'd942,
    COMP_LOOP_C_543 = 11'd943,
    COMP_LOOP_C_544 = 11'd944,
    COMP_LOOP_C_545 = 11'd945,
    COMP_LOOP_C_546 = 11'd946,
    COMP_LOOP_C_547 = 11'd947,
    COMP_LOOP_C_548 = 11'd948,
    COMP_LOOP_C_549 = 11'd949,
    COMP_LOOP_C_550 = 11'd950,
    COMP_LOOP_C_551 = 11'd951,
    COMP_LOOP_C_552 = 11'd952,
    COMP_LOOP_C_553 = 11'd953,
    COMP_LOOP_C_554 = 11'd954,
    COMP_LOOP_C_555 = 11'd955,
    COMP_LOOP_C_556 = 11'd956,
    COMP_LOOP_C_557 = 11'd957,
    COMP_LOOP_C_558 = 11'd958,
    COMP_LOOP_C_559 = 11'd959,
    COMP_LOOP_C_560 = 11'd960,
    COMP_LOOP_C_561 = 11'd961,
    COMP_LOOP_C_562 = 11'd962,
    COMP_LOOP_C_563 = 11'd963,
    COMP_LOOP_C_564 = 11'd964,
    COMP_LOOP_C_565 = 11'd965,
    COMP_LOOP_C_566 = 11'd966,
    COMP_LOOP_C_567 = 11'd967,
    COMP_LOOP_C_568 = 11'd968,
    COMP_LOOP_C_569 = 11'd969,
    COMP_LOOP_C_570 = 11'd970,
    COMP_LOOP_C_571 = 11'd971,
    COMP_LOOP_C_572 = 11'd972,
    COMP_LOOP_C_573 = 11'd973,
    COMP_LOOP_C_574 = 11'd974,
    COMP_LOOP_C_575 = 11'd975,
    COMP_LOOP_C_576 = 11'd976,
    COMP_LOOP_C_577 = 11'd977,
    COMP_LOOP_10_modExp_1_while_C_0 = 11'd978,
    COMP_LOOP_10_modExp_1_while_C_1 = 11'd979,
    COMP_LOOP_10_modExp_1_while_C_2 = 11'd980,
    COMP_LOOP_10_modExp_1_while_C_3 = 11'd981,
    COMP_LOOP_10_modExp_1_while_C_4 = 11'd982,
    COMP_LOOP_10_modExp_1_while_C_5 = 11'd983,
    COMP_LOOP_10_modExp_1_while_C_6 = 11'd984,
    COMP_LOOP_10_modExp_1_while_C_7 = 11'd985,
    COMP_LOOP_10_modExp_1_while_C_8 = 11'd986,
    COMP_LOOP_10_modExp_1_while_C_9 = 11'd987,
    COMP_LOOP_10_modExp_1_while_C_10 = 11'd988,
    COMP_LOOP_10_modExp_1_while_C_11 = 11'd989,
    COMP_LOOP_10_modExp_1_while_C_12 = 11'd990,
    COMP_LOOP_10_modExp_1_while_C_13 = 11'd991,
    COMP_LOOP_10_modExp_1_while_C_14 = 11'd992,
    COMP_LOOP_10_modExp_1_while_C_15 = 11'd993,
    COMP_LOOP_10_modExp_1_while_C_16 = 11'd994,
    COMP_LOOP_10_modExp_1_while_C_17 = 11'd995,
    COMP_LOOP_10_modExp_1_while_C_18 = 11'd996,
    COMP_LOOP_10_modExp_1_while_C_19 = 11'd997,
    COMP_LOOP_10_modExp_1_while_C_20 = 11'd998,
    COMP_LOOP_10_modExp_1_while_C_21 = 11'd999,
    COMP_LOOP_10_modExp_1_while_C_22 = 11'd1000,
    COMP_LOOP_10_modExp_1_while_C_23 = 11'd1001,
    COMP_LOOP_10_modExp_1_while_C_24 = 11'd1002,
    COMP_LOOP_10_modExp_1_while_C_25 = 11'd1003,
    COMP_LOOP_10_modExp_1_while_C_26 = 11'd1004,
    COMP_LOOP_10_modExp_1_while_C_27 = 11'd1005,
    COMP_LOOP_10_modExp_1_while_C_28 = 11'd1006,
    COMP_LOOP_10_modExp_1_while_C_29 = 11'd1007,
    COMP_LOOP_10_modExp_1_while_C_30 = 11'd1008,
    COMP_LOOP_10_modExp_1_while_C_31 = 11'd1009,
    COMP_LOOP_10_modExp_1_while_C_32 = 11'd1010,
    COMP_LOOP_10_modExp_1_while_C_33 = 11'd1011,
    COMP_LOOP_10_modExp_1_while_C_34 = 11'd1012,
    COMP_LOOP_10_modExp_1_while_C_35 = 11'd1013,
    COMP_LOOP_10_modExp_1_while_C_36 = 11'd1014,
    COMP_LOOP_10_modExp_1_while_C_37 = 11'd1015,
    COMP_LOOP_10_modExp_1_while_C_38 = 11'd1016,
    COMP_LOOP_C_578 = 11'd1017,
    COMP_LOOP_C_579 = 11'd1018,
    COMP_LOOP_C_580 = 11'd1019,
    COMP_LOOP_C_581 = 11'd1020,
    COMP_LOOP_C_582 = 11'd1021,
    COMP_LOOP_C_583 = 11'd1022,
    COMP_LOOP_C_584 = 11'd1023,
    COMP_LOOP_C_585 = 11'd1024,
    COMP_LOOP_C_586 = 11'd1025,
    COMP_LOOP_C_587 = 11'd1026,
    COMP_LOOP_C_588 = 11'd1027,
    COMP_LOOP_C_589 = 11'd1028,
    COMP_LOOP_C_590 = 11'd1029,
    COMP_LOOP_C_591 = 11'd1030,
    COMP_LOOP_C_592 = 11'd1031,
    COMP_LOOP_C_593 = 11'd1032,
    COMP_LOOP_C_594 = 11'd1033,
    COMP_LOOP_C_595 = 11'd1034,
    COMP_LOOP_C_596 = 11'd1035,
    COMP_LOOP_C_597 = 11'd1036,
    COMP_LOOP_C_598 = 11'd1037,
    COMP_LOOP_C_599 = 11'd1038,
    COMP_LOOP_C_600 = 11'd1039,
    COMP_LOOP_C_601 = 11'd1040,
    COMP_LOOP_C_602 = 11'd1041,
    COMP_LOOP_C_603 = 11'd1042,
    COMP_LOOP_C_604 = 11'd1043,
    COMP_LOOP_C_605 = 11'd1044,
    COMP_LOOP_C_606 = 11'd1045,
    COMP_LOOP_C_607 = 11'd1046,
    COMP_LOOP_C_608 = 11'd1047,
    COMP_LOOP_C_609 = 11'd1048,
    COMP_LOOP_C_610 = 11'd1049,
    COMP_LOOP_C_611 = 11'd1050,
    COMP_LOOP_C_612 = 11'd1051,
    COMP_LOOP_C_613 = 11'd1052,
    COMP_LOOP_C_614 = 11'd1053,
    COMP_LOOP_C_615 = 11'd1054,
    COMP_LOOP_C_616 = 11'd1055,
    COMP_LOOP_C_617 = 11'd1056,
    COMP_LOOP_C_618 = 11'd1057,
    COMP_LOOP_C_619 = 11'd1058,
    COMP_LOOP_C_620 = 11'd1059,
    COMP_LOOP_C_621 = 11'd1060,
    COMP_LOOP_C_622 = 11'd1061,
    COMP_LOOP_C_623 = 11'd1062,
    COMP_LOOP_C_624 = 11'd1063,
    COMP_LOOP_C_625 = 11'd1064,
    COMP_LOOP_C_626 = 11'd1065,
    COMP_LOOP_C_627 = 11'd1066,
    COMP_LOOP_C_628 = 11'd1067,
    COMP_LOOP_C_629 = 11'd1068,
    COMP_LOOP_C_630 = 11'd1069,
    COMP_LOOP_C_631 = 11'd1070,
    COMP_LOOP_C_632 = 11'd1071,
    COMP_LOOP_C_633 = 11'd1072,
    COMP_LOOP_C_634 = 11'd1073,
    COMP_LOOP_C_635 = 11'd1074,
    COMP_LOOP_C_636 = 11'd1075,
    COMP_LOOP_C_637 = 11'd1076,
    COMP_LOOP_C_638 = 11'd1077,
    COMP_LOOP_C_639 = 11'd1078,
    COMP_LOOP_C_640 = 11'd1079,
    COMP_LOOP_C_641 = 11'd1080,
    COMP_LOOP_11_modExp_1_while_C_0 = 11'd1081,
    COMP_LOOP_11_modExp_1_while_C_1 = 11'd1082,
    COMP_LOOP_11_modExp_1_while_C_2 = 11'd1083,
    COMP_LOOP_11_modExp_1_while_C_3 = 11'd1084,
    COMP_LOOP_11_modExp_1_while_C_4 = 11'd1085,
    COMP_LOOP_11_modExp_1_while_C_5 = 11'd1086,
    COMP_LOOP_11_modExp_1_while_C_6 = 11'd1087,
    COMP_LOOP_11_modExp_1_while_C_7 = 11'd1088,
    COMP_LOOP_11_modExp_1_while_C_8 = 11'd1089,
    COMP_LOOP_11_modExp_1_while_C_9 = 11'd1090,
    COMP_LOOP_11_modExp_1_while_C_10 = 11'd1091,
    COMP_LOOP_11_modExp_1_while_C_11 = 11'd1092,
    COMP_LOOP_11_modExp_1_while_C_12 = 11'd1093,
    COMP_LOOP_11_modExp_1_while_C_13 = 11'd1094,
    COMP_LOOP_11_modExp_1_while_C_14 = 11'd1095,
    COMP_LOOP_11_modExp_1_while_C_15 = 11'd1096,
    COMP_LOOP_11_modExp_1_while_C_16 = 11'd1097,
    COMP_LOOP_11_modExp_1_while_C_17 = 11'd1098,
    COMP_LOOP_11_modExp_1_while_C_18 = 11'd1099,
    COMP_LOOP_11_modExp_1_while_C_19 = 11'd1100,
    COMP_LOOP_11_modExp_1_while_C_20 = 11'd1101,
    COMP_LOOP_11_modExp_1_while_C_21 = 11'd1102,
    COMP_LOOP_11_modExp_1_while_C_22 = 11'd1103,
    COMP_LOOP_11_modExp_1_while_C_23 = 11'd1104,
    COMP_LOOP_11_modExp_1_while_C_24 = 11'd1105,
    COMP_LOOP_11_modExp_1_while_C_25 = 11'd1106,
    COMP_LOOP_11_modExp_1_while_C_26 = 11'd1107,
    COMP_LOOP_11_modExp_1_while_C_27 = 11'd1108,
    COMP_LOOP_11_modExp_1_while_C_28 = 11'd1109,
    COMP_LOOP_11_modExp_1_while_C_29 = 11'd1110,
    COMP_LOOP_11_modExp_1_while_C_30 = 11'd1111,
    COMP_LOOP_11_modExp_1_while_C_31 = 11'd1112,
    COMP_LOOP_11_modExp_1_while_C_32 = 11'd1113,
    COMP_LOOP_11_modExp_1_while_C_33 = 11'd1114,
    COMP_LOOP_11_modExp_1_while_C_34 = 11'd1115,
    COMP_LOOP_11_modExp_1_while_C_35 = 11'd1116,
    COMP_LOOP_11_modExp_1_while_C_36 = 11'd1117,
    COMP_LOOP_11_modExp_1_while_C_37 = 11'd1118,
    COMP_LOOP_11_modExp_1_while_C_38 = 11'd1119,
    COMP_LOOP_C_642 = 11'd1120,
    COMP_LOOP_C_643 = 11'd1121,
    COMP_LOOP_C_644 = 11'd1122,
    COMP_LOOP_C_645 = 11'd1123,
    COMP_LOOP_C_646 = 11'd1124,
    COMP_LOOP_C_647 = 11'd1125,
    COMP_LOOP_C_648 = 11'd1126,
    COMP_LOOP_C_649 = 11'd1127,
    COMP_LOOP_C_650 = 11'd1128,
    COMP_LOOP_C_651 = 11'd1129,
    COMP_LOOP_C_652 = 11'd1130,
    COMP_LOOP_C_653 = 11'd1131,
    COMP_LOOP_C_654 = 11'd1132,
    COMP_LOOP_C_655 = 11'd1133,
    COMP_LOOP_C_656 = 11'd1134,
    COMP_LOOP_C_657 = 11'd1135,
    COMP_LOOP_C_658 = 11'd1136,
    COMP_LOOP_C_659 = 11'd1137,
    COMP_LOOP_C_660 = 11'd1138,
    COMP_LOOP_C_661 = 11'd1139,
    COMP_LOOP_C_662 = 11'd1140,
    COMP_LOOP_C_663 = 11'd1141,
    COMP_LOOP_C_664 = 11'd1142,
    COMP_LOOP_C_665 = 11'd1143,
    COMP_LOOP_C_666 = 11'd1144,
    COMP_LOOP_C_667 = 11'd1145,
    COMP_LOOP_C_668 = 11'd1146,
    COMP_LOOP_C_669 = 11'd1147,
    COMP_LOOP_C_670 = 11'd1148,
    COMP_LOOP_C_671 = 11'd1149,
    COMP_LOOP_C_672 = 11'd1150,
    COMP_LOOP_C_673 = 11'd1151,
    COMP_LOOP_C_674 = 11'd1152,
    COMP_LOOP_C_675 = 11'd1153,
    COMP_LOOP_C_676 = 11'd1154,
    COMP_LOOP_C_677 = 11'd1155,
    COMP_LOOP_C_678 = 11'd1156,
    COMP_LOOP_C_679 = 11'd1157,
    COMP_LOOP_C_680 = 11'd1158,
    COMP_LOOP_C_681 = 11'd1159,
    COMP_LOOP_C_682 = 11'd1160,
    COMP_LOOP_C_683 = 11'd1161,
    COMP_LOOP_C_684 = 11'd1162,
    COMP_LOOP_C_685 = 11'd1163,
    COMP_LOOP_C_686 = 11'd1164,
    COMP_LOOP_C_687 = 11'd1165,
    COMP_LOOP_C_688 = 11'd1166,
    COMP_LOOP_C_689 = 11'd1167,
    COMP_LOOP_C_690 = 11'd1168,
    COMP_LOOP_C_691 = 11'd1169,
    COMP_LOOP_C_692 = 11'd1170,
    COMP_LOOP_C_693 = 11'd1171,
    COMP_LOOP_C_694 = 11'd1172,
    COMP_LOOP_C_695 = 11'd1173,
    COMP_LOOP_C_696 = 11'd1174,
    COMP_LOOP_C_697 = 11'd1175,
    COMP_LOOP_C_698 = 11'd1176,
    COMP_LOOP_C_699 = 11'd1177,
    COMP_LOOP_C_700 = 11'd1178,
    COMP_LOOP_C_701 = 11'd1179,
    COMP_LOOP_C_702 = 11'd1180,
    COMP_LOOP_C_703 = 11'd1181,
    COMP_LOOP_C_704 = 11'd1182,
    COMP_LOOP_C_705 = 11'd1183,
    COMP_LOOP_12_modExp_1_while_C_0 = 11'd1184,
    COMP_LOOP_12_modExp_1_while_C_1 = 11'd1185,
    COMP_LOOP_12_modExp_1_while_C_2 = 11'd1186,
    COMP_LOOP_12_modExp_1_while_C_3 = 11'd1187,
    COMP_LOOP_12_modExp_1_while_C_4 = 11'd1188,
    COMP_LOOP_12_modExp_1_while_C_5 = 11'd1189,
    COMP_LOOP_12_modExp_1_while_C_6 = 11'd1190,
    COMP_LOOP_12_modExp_1_while_C_7 = 11'd1191,
    COMP_LOOP_12_modExp_1_while_C_8 = 11'd1192,
    COMP_LOOP_12_modExp_1_while_C_9 = 11'd1193,
    COMP_LOOP_12_modExp_1_while_C_10 = 11'd1194,
    COMP_LOOP_12_modExp_1_while_C_11 = 11'd1195,
    COMP_LOOP_12_modExp_1_while_C_12 = 11'd1196,
    COMP_LOOP_12_modExp_1_while_C_13 = 11'd1197,
    COMP_LOOP_12_modExp_1_while_C_14 = 11'd1198,
    COMP_LOOP_12_modExp_1_while_C_15 = 11'd1199,
    COMP_LOOP_12_modExp_1_while_C_16 = 11'd1200,
    COMP_LOOP_12_modExp_1_while_C_17 = 11'd1201,
    COMP_LOOP_12_modExp_1_while_C_18 = 11'd1202,
    COMP_LOOP_12_modExp_1_while_C_19 = 11'd1203,
    COMP_LOOP_12_modExp_1_while_C_20 = 11'd1204,
    COMP_LOOP_12_modExp_1_while_C_21 = 11'd1205,
    COMP_LOOP_12_modExp_1_while_C_22 = 11'd1206,
    COMP_LOOP_12_modExp_1_while_C_23 = 11'd1207,
    COMP_LOOP_12_modExp_1_while_C_24 = 11'd1208,
    COMP_LOOP_12_modExp_1_while_C_25 = 11'd1209,
    COMP_LOOP_12_modExp_1_while_C_26 = 11'd1210,
    COMP_LOOP_12_modExp_1_while_C_27 = 11'd1211,
    COMP_LOOP_12_modExp_1_while_C_28 = 11'd1212,
    COMP_LOOP_12_modExp_1_while_C_29 = 11'd1213,
    COMP_LOOP_12_modExp_1_while_C_30 = 11'd1214,
    COMP_LOOP_12_modExp_1_while_C_31 = 11'd1215,
    COMP_LOOP_12_modExp_1_while_C_32 = 11'd1216,
    COMP_LOOP_12_modExp_1_while_C_33 = 11'd1217,
    COMP_LOOP_12_modExp_1_while_C_34 = 11'd1218,
    COMP_LOOP_12_modExp_1_while_C_35 = 11'd1219,
    COMP_LOOP_12_modExp_1_while_C_36 = 11'd1220,
    COMP_LOOP_12_modExp_1_while_C_37 = 11'd1221,
    COMP_LOOP_12_modExp_1_while_C_38 = 11'd1222,
    COMP_LOOP_C_706 = 11'd1223,
    COMP_LOOP_C_707 = 11'd1224,
    COMP_LOOP_C_708 = 11'd1225,
    COMP_LOOP_C_709 = 11'd1226,
    COMP_LOOP_C_710 = 11'd1227,
    COMP_LOOP_C_711 = 11'd1228,
    COMP_LOOP_C_712 = 11'd1229,
    COMP_LOOP_C_713 = 11'd1230,
    COMP_LOOP_C_714 = 11'd1231,
    COMP_LOOP_C_715 = 11'd1232,
    COMP_LOOP_C_716 = 11'd1233,
    COMP_LOOP_C_717 = 11'd1234,
    COMP_LOOP_C_718 = 11'd1235,
    COMP_LOOP_C_719 = 11'd1236,
    COMP_LOOP_C_720 = 11'd1237,
    COMP_LOOP_C_721 = 11'd1238,
    COMP_LOOP_C_722 = 11'd1239,
    COMP_LOOP_C_723 = 11'd1240,
    COMP_LOOP_C_724 = 11'd1241,
    COMP_LOOP_C_725 = 11'd1242,
    COMP_LOOP_C_726 = 11'd1243,
    COMP_LOOP_C_727 = 11'd1244,
    COMP_LOOP_C_728 = 11'd1245,
    COMP_LOOP_C_729 = 11'd1246,
    COMP_LOOP_C_730 = 11'd1247,
    COMP_LOOP_C_731 = 11'd1248,
    COMP_LOOP_C_732 = 11'd1249,
    COMP_LOOP_C_733 = 11'd1250,
    COMP_LOOP_C_734 = 11'd1251,
    COMP_LOOP_C_735 = 11'd1252,
    COMP_LOOP_C_736 = 11'd1253,
    COMP_LOOP_C_737 = 11'd1254,
    COMP_LOOP_C_738 = 11'd1255,
    COMP_LOOP_C_739 = 11'd1256,
    COMP_LOOP_C_740 = 11'd1257,
    COMP_LOOP_C_741 = 11'd1258,
    COMP_LOOP_C_742 = 11'd1259,
    COMP_LOOP_C_743 = 11'd1260,
    COMP_LOOP_C_744 = 11'd1261,
    COMP_LOOP_C_745 = 11'd1262,
    COMP_LOOP_C_746 = 11'd1263,
    COMP_LOOP_C_747 = 11'd1264,
    COMP_LOOP_C_748 = 11'd1265,
    COMP_LOOP_C_749 = 11'd1266,
    COMP_LOOP_C_750 = 11'd1267,
    COMP_LOOP_C_751 = 11'd1268,
    COMP_LOOP_C_752 = 11'd1269,
    COMP_LOOP_C_753 = 11'd1270,
    COMP_LOOP_C_754 = 11'd1271,
    COMP_LOOP_C_755 = 11'd1272,
    COMP_LOOP_C_756 = 11'd1273,
    COMP_LOOP_C_757 = 11'd1274,
    COMP_LOOP_C_758 = 11'd1275,
    COMP_LOOP_C_759 = 11'd1276,
    COMP_LOOP_C_760 = 11'd1277,
    COMP_LOOP_C_761 = 11'd1278,
    COMP_LOOP_C_762 = 11'd1279,
    COMP_LOOP_C_763 = 11'd1280,
    COMP_LOOP_C_764 = 11'd1281,
    COMP_LOOP_C_765 = 11'd1282,
    COMP_LOOP_C_766 = 11'd1283,
    COMP_LOOP_C_767 = 11'd1284,
    COMP_LOOP_C_768 = 11'd1285,
    COMP_LOOP_C_769 = 11'd1286,
    COMP_LOOP_13_modExp_1_while_C_0 = 11'd1287,
    COMP_LOOP_13_modExp_1_while_C_1 = 11'd1288,
    COMP_LOOP_13_modExp_1_while_C_2 = 11'd1289,
    COMP_LOOP_13_modExp_1_while_C_3 = 11'd1290,
    COMP_LOOP_13_modExp_1_while_C_4 = 11'd1291,
    COMP_LOOP_13_modExp_1_while_C_5 = 11'd1292,
    COMP_LOOP_13_modExp_1_while_C_6 = 11'd1293,
    COMP_LOOP_13_modExp_1_while_C_7 = 11'd1294,
    COMP_LOOP_13_modExp_1_while_C_8 = 11'd1295,
    COMP_LOOP_13_modExp_1_while_C_9 = 11'd1296,
    COMP_LOOP_13_modExp_1_while_C_10 = 11'd1297,
    COMP_LOOP_13_modExp_1_while_C_11 = 11'd1298,
    COMP_LOOP_13_modExp_1_while_C_12 = 11'd1299,
    COMP_LOOP_13_modExp_1_while_C_13 = 11'd1300,
    COMP_LOOP_13_modExp_1_while_C_14 = 11'd1301,
    COMP_LOOP_13_modExp_1_while_C_15 = 11'd1302,
    COMP_LOOP_13_modExp_1_while_C_16 = 11'd1303,
    COMP_LOOP_13_modExp_1_while_C_17 = 11'd1304,
    COMP_LOOP_13_modExp_1_while_C_18 = 11'd1305,
    COMP_LOOP_13_modExp_1_while_C_19 = 11'd1306,
    COMP_LOOP_13_modExp_1_while_C_20 = 11'd1307,
    COMP_LOOP_13_modExp_1_while_C_21 = 11'd1308,
    COMP_LOOP_13_modExp_1_while_C_22 = 11'd1309,
    COMP_LOOP_13_modExp_1_while_C_23 = 11'd1310,
    COMP_LOOP_13_modExp_1_while_C_24 = 11'd1311,
    COMP_LOOP_13_modExp_1_while_C_25 = 11'd1312,
    COMP_LOOP_13_modExp_1_while_C_26 = 11'd1313,
    COMP_LOOP_13_modExp_1_while_C_27 = 11'd1314,
    COMP_LOOP_13_modExp_1_while_C_28 = 11'd1315,
    COMP_LOOP_13_modExp_1_while_C_29 = 11'd1316,
    COMP_LOOP_13_modExp_1_while_C_30 = 11'd1317,
    COMP_LOOP_13_modExp_1_while_C_31 = 11'd1318,
    COMP_LOOP_13_modExp_1_while_C_32 = 11'd1319,
    COMP_LOOP_13_modExp_1_while_C_33 = 11'd1320,
    COMP_LOOP_13_modExp_1_while_C_34 = 11'd1321,
    COMP_LOOP_13_modExp_1_while_C_35 = 11'd1322,
    COMP_LOOP_13_modExp_1_while_C_36 = 11'd1323,
    COMP_LOOP_13_modExp_1_while_C_37 = 11'd1324,
    COMP_LOOP_13_modExp_1_while_C_38 = 11'd1325,
    COMP_LOOP_C_770 = 11'd1326,
    COMP_LOOP_C_771 = 11'd1327,
    COMP_LOOP_C_772 = 11'd1328,
    COMP_LOOP_C_773 = 11'd1329,
    COMP_LOOP_C_774 = 11'd1330,
    COMP_LOOP_C_775 = 11'd1331,
    COMP_LOOP_C_776 = 11'd1332,
    COMP_LOOP_C_777 = 11'd1333,
    COMP_LOOP_C_778 = 11'd1334,
    COMP_LOOP_C_779 = 11'd1335,
    COMP_LOOP_C_780 = 11'd1336,
    COMP_LOOP_C_781 = 11'd1337,
    COMP_LOOP_C_782 = 11'd1338,
    COMP_LOOP_C_783 = 11'd1339,
    COMP_LOOP_C_784 = 11'd1340,
    COMP_LOOP_C_785 = 11'd1341,
    COMP_LOOP_C_786 = 11'd1342,
    COMP_LOOP_C_787 = 11'd1343,
    COMP_LOOP_C_788 = 11'd1344,
    COMP_LOOP_C_789 = 11'd1345,
    COMP_LOOP_C_790 = 11'd1346,
    COMP_LOOP_C_791 = 11'd1347,
    COMP_LOOP_C_792 = 11'd1348,
    COMP_LOOP_C_793 = 11'd1349,
    COMP_LOOP_C_794 = 11'd1350,
    COMP_LOOP_C_795 = 11'd1351,
    COMP_LOOP_C_796 = 11'd1352,
    COMP_LOOP_C_797 = 11'd1353,
    COMP_LOOP_C_798 = 11'd1354,
    COMP_LOOP_C_799 = 11'd1355,
    COMP_LOOP_C_800 = 11'd1356,
    COMP_LOOP_C_801 = 11'd1357,
    COMP_LOOP_C_802 = 11'd1358,
    COMP_LOOP_C_803 = 11'd1359,
    COMP_LOOP_C_804 = 11'd1360,
    COMP_LOOP_C_805 = 11'd1361,
    COMP_LOOP_C_806 = 11'd1362,
    COMP_LOOP_C_807 = 11'd1363,
    COMP_LOOP_C_808 = 11'd1364,
    COMP_LOOP_C_809 = 11'd1365,
    COMP_LOOP_C_810 = 11'd1366,
    COMP_LOOP_C_811 = 11'd1367,
    COMP_LOOP_C_812 = 11'd1368,
    COMP_LOOP_C_813 = 11'd1369,
    COMP_LOOP_C_814 = 11'd1370,
    COMP_LOOP_C_815 = 11'd1371,
    COMP_LOOP_C_816 = 11'd1372,
    COMP_LOOP_C_817 = 11'd1373,
    COMP_LOOP_C_818 = 11'd1374,
    COMP_LOOP_C_819 = 11'd1375,
    COMP_LOOP_C_820 = 11'd1376,
    COMP_LOOP_C_821 = 11'd1377,
    COMP_LOOP_C_822 = 11'd1378,
    COMP_LOOP_C_823 = 11'd1379,
    COMP_LOOP_C_824 = 11'd1380,
    COMP_LOOP_C_825 = 11'd1381,
    COMP_LOOP_C_826 = 11'd1382,
    COMP_LOOP_C_827 = 11'd1383,
    COMP_LOOP_C_828 = 11'd1384,
    COMP_LOOP_C_829 = 11'd1385,
    COMP_LOOP_C_830 = 11'd1386,
    COMP_LOOP_C_831 = 11'd1387,
    COMP_LOOP_C_832 = 11'd1388,
    COMP_LOOP_C_833 = 11'd1389,
    COMP_LOOP_14_modExp_1_while_C_0 = 11'd1390,
    COMP_LOOP_14_modExp_1_while_C_1 = 11'd1391,
    COMP_LOOP_14_modExp_1_while_C_2 = 11'd1392,
    COMP_LOOP_14_modExp_1_while_C_3 = 11'd1393,
    COMP_LOOP_14_modExp_1_while_C_4 = 11'd1394,
    COMP_LOOP_14_modExp_1_while_C_5 = 11'd1395,
    COMP_LOOP_14_modExp_1_while_C_6 = 11'd1396,
    COMP_LOOP_14_modExp_1_while_C_7 = 11'd1397,
    COMP_LOOP_14_modExp_1_while_C_8 = 11'd1398,
    COMP_LOOP_14_modExp_1_while_C_9 = 11'd1399,
    COMP_LOOP_14_modExp_1_while_C_10 = 11'd1400,
    COMP_LOOP_14_modExp_1_while_C_11 = 11'd1401,
    COMP_LOOP_14_modExp_1_while_C_12 = 11'd1402,
    COMP_LOOP_14_modExp_1_while_C_13 = 11'd1403,
    COMP_LOOP_14_modExp_1_while_C_14 = 11'd1404,
    COMP_LOOP_14_modExp_1_while_C_15 = 11'd1405,
    COMP_LOOP_14_modExp_1_while_C_16 = 11'd1406,
    COMP_LOOP_14_modExp_1_while_C_17 = 11'd1407,
    COMP_LOOP_14_modExp_1_while_C_18 = 11'd1408,
    COMP_LOOP_14_modExp_1_while_C_19 = 11'd1409,
    COMP_LOOP_14_modExp_1_while_C_20 = 11'd1410,
    COMP_LOOP_14_modExp_1_while_C_21 = 11'd1411,
    COMP_LOOP_14_modExp_1_while_C_22 = 11'd1412,
    COMP_LOOP_14_modExp_1_while_C_23 = 11'd1413,
    COMP_LOOP_14_modExp_1_while_C_24 = 11'd1414,
    COMP_LOOP_14_modExp_1_while_C_25 = 11'd1415,
    COMP_LOOP_14_modExp_1_while_C_26 = 11'd1416,
    COMP_LOOP_14_modExp_1_while_C_27 = 11'd1417,
    COMP_LOOP_14_modExp_1_while_C_28 = 11'd1418,
    COMP_LOOP_14_modExp_1_while_C_29 = 11'd1419,
    COMP_LOOP_14_modExp_1_while_C_30 = 11'd1420,
    COMP_LOOP_14_modExp_1_while_C_31 = 11'd1421,
    COMP_LOOP_14_modExp_1_while_C_32 = 11'd1422,
    COMP_LOOP_14_modExp_1_while_C_33 = 11'd1423,
    COMP_LOOP_14_modExp_1_while_C_34 = 11'd1424,
    COMP_LOOP_14_modExp_1_while_C_35 = 11'd1425,
    COMP_LOOP_14_modExp_1_while_C_36 = 11'd1426,
    COMP_LOOP_14_modExp_1_while_C_37 = 11'd1427,
    COMP_LOOP_14_modExp_1_while_C_38 = 11'd1428,
    COMP_LOOP_C_834 = 11'd1429,
    COMP_LOOP_C_835 = 11'd1430,
    COMP_LOOP_C_836 = 11'd1431,
    COMP_LOOP_C_837 = 11'd1432,
    COMP_LOOP_C_838 = 11'd1433,
    COMP_LOOP_C_839 = 11'd1434,
    COMP_LOOP_C_840 = 11'd1435,
    COMP_LOOP_C_841 = 11'd1436,
    COMP_LOOP_C_842 = 11'd1437,
    COMP_LOOP_C_843 = 11'd1438,
    COMP_LOOP_C_844 = 11'd1439,
    COMP_LOOP_C_845 = 11'd1440,
    COMP_LOOP_C_846 = 11'd1441,
    COMP_LOOP_C_847 = 11'd1442,
    COMP_LOOP_C_848 = 11'd1443,
    COMP_LOOP_C_849 = 11'd1444,
    COMP_LOOP_C_850 = 11'd1445,
    COMP_LOOP_C_851 = 11'd1446,
    COMP_LOOP_C_852 = 11'd1447,
    COMP_LOOP_C_853 = 11'd1448,
    COMP_LOOP_C_854 = 11'd1449,
    COMP_LOOP_C_855 = 11'd1450,
    COMP_LOOP_C_856 = 11'd1451,
    COMP_LOOP_C_857 = 11'd1452,
    COMP_LOOP_C_858 = 11'd1453,
    COMP_LOOP_C_859 = 11'd1454,
    COMP_LOOP_C_860 = 11'd1455,
    COMP_LOOP_C_861 = 11'd1456,
    COMP_LOOP_C_862 = 11'd1457,
    COMP_LOOP_C_863 = 11'd1458,
    COMP_LOOP_C_864 = 11'd1459,
    COMP_LOOP_C_865 = 11'd1460,
    COMP_LOOP_C_866 = 11'd1461,
    COMP_LOOP_C_867 = 11'd1462,
    COMP_LOOP_C_868 = 11'd1463,
    COMP_LOOP_C_869 = 11'd1464,
    COMP_LOOP_C_870 = 11'd1465,
    COMP_LOOP_C_871 = 11'd1466,
    COMP_LOOP_C_872 = 11'd1467,
    COMP_LOOP_C_873 = 11'd1468,
    COMP_LOOP_C_874 = 11'd1469,
    COMP_LOOP_C_875 = 11'd1470,
    COMP_LOOP_C_876 = 11'd1471,
    COMP_LOOP_C_877 = 11'd1472,
    COMP_LOOP_C_878 = 11'd1473,
    COMP_LOOP_C_879 = 11'd1474,
    COMP_LOOP_C_880 = 11'd1475,
    COMP_LOOP_C_881 = 11'd1476,
    COMP_LOOP_C_882 = 11'd1477,
    COMP_LOOP_C_883 = 11'd1478,
    COMP_LOOP_C_884 = 11'd1479,
    COMP_LOOP_C_885 = 11'd1480,
    COMP_LOOP_C_886 = 11'd1481,
    COMP_LOOP_C_887 = 11'd1482,
    COMP_LOOP_C_888 = 11'd1483,
    COMP_LOOP_C_889 = 11'd1484,
    COMP_LOOP_C_890 = 11'd1485,
    COMP_LOOP_C_891 = 11'd1486,
    COMP_LOOP_C_892 = 11'd1487,
    COMP_LOOP_C_893 = 11'd1488,
    COMP_LOOP_C_894 = 11'd1489,
    COMP_LOOP_C_895 = 11'd1490,
    COMP_LOOP_C_896 = 11'd1491,
    COMP_LOOP_C_897 = 11'd1492,
    COMP_LOOP_15_modExp_1_while_C_0 = 11'd1493,
    COMP_LOOP_15_modExp_1_while_C_1 = 11'd1494,
    COMP_LOOP_15_modExp_1_while_C_2 = 11'd1495,
    COMP_LOOP_15_modExp_1_while_C_3 = 11'd1496,
    COMP_LOOP_15_modExp_1_while_C_4 = 11'd1497,
    COMP_LOOP_15_modExp_1_while_C_5 = 11'd1498,
    COMP_LOOP_15_modExp_1_while_C_6 = 11'd1499,
    COMP_LOOP_15_modExp_1_while_C_7 = 11'd1500,
    COMP_LOOP_15_modExp_1_while_C_8 = 11'd1501,
    COMP_LOOP_15_modExp_1_while_C_9 = 11'd1502,
    COMP_LOOP_15_modExp_1_while_C_10 = 11'd1503,
    COMP_LOOP_15_modExp_1_while_C_11 = 11'd1504,
    COMP_LOOP_15_modExp_1_while_C_12 = 11'd1505,
    COMP_LOOP_15_modExp_1_while_C_13 = 11'd1506,
    COMP_LOOP_15_modExp_1_while_C_14 = 11'd1507,
    COMP_LOOP_15_modExp_1_while_C_15 = 11'd1508,
    COMP_LOOP_15_modExp_1_while_C_16 = 11'd1509,
    COMP_LOOP_15_modExp_1_while_C_17 = 11'd1510,
    COMP_LOOP_15_modExp_1_while_C_18 = 11'd1511,
    COMP_LOOP_15_modExp_1_while_C_19 = 11'd1512,
    COMP_LOOP_15_modExp_1_while_C_20 = 11'd1513,
    COMP_LOOP_15_modExp_1_while_C_21 = 11'd1514,
    COMP_LOOP_15_modExp_1_while_C_22 = 11'd1515,
    COMP_LOOP_15_modExp_1_while_C_23 = 11'd1516,
    COMP_LOOP_15_modExp_1_while_C_24 = 11'd1517,
    COMP_LOOP_15_modExp_1_while_C_25 = 11'd1518,
    COMP_LOOP_15_modExp_1_while_C_26 = 11'd1519,
    COMP_LOOP_15_modExp_1_while_C_27 = 11'd1520,
    COMP_LOOP_15_modExp_1_while_C_28 = 11'd1521,
    COMP_LOOP_15_modExp_1_while_C_29 = 11'd1522,
    COMP_LOOP_15_modExp_1_while_C_30 = 11'd1523,
    COMP_LOOP_15_modExp_1_while_C_31 = 11'd1524,
    COMP_LOOP_15_modExp_1_while_C_32 = 11'd1525,
    COMP_LOOP_15_modExp_1_while_C_33 = 11'd1526,
    COMP_LOOP_15_modExp_1_while_C_34 = 11'd1527,
    COMP_LOOP_15_modExp_1_while_C_35 = 11'd1528,
    COMP_LOOP_15_modExp_1_while_C_36 = 11'd1529,
    COMP_LOOP_15_modExp_1_while_C_37 = 11'd1530,
    COMP_LOOP_15_modExp_1_while_C_38 = 11'd1531,
    COMP_LOOP_C_898 = 11'd1532,
    COMP_LOOP_C_899 = 11'd1533,
    COMP_LOOP_C_900 = 11'd1534,
    COMP_LOOP_C_901 = 11'd1535,
    COMP_LOOP_C_902 = 11'd1536,
    COMP_LOOP_C_903 = 11'd1537,
    COMP_LOOP_C_904 = 11'd1538,
    COMP_LOOP_C_905 = 11'd1539,
    COMP_LOOP_C_906 = 11'd1540,
    COMP_LOOP_C_907 = 11'd1541,
    COMP_LOOP_C_908 = 11'd1542,
    COMP_LOOP_C_909 = 11'd1543,
    COMP_LOOP_C_910 = 11'd1544,
    COMP_LOOP_C_911 = 11'd1545,
    COMP_LOOP_C_912 = 11'd1546,
    COMP_LOOP_C_913 = 11'd1547,
    COMP_LOOP_C_914 = 11'd1548,
    COMP_LOOP_C_915 = 11'd1549,
    COMP_LOOP_C_916 = 11'd1550,
    COMP_LOOP_C_917 = 11'd1551,
    COMP_LOOP_C_918 = 11'd1552,
    COMP_LOOP_C_919 = 11'd1553,
    COMP_LOOP_C_920 = 11'd1554,
    COMP_LOOP_C_921 = 11'd1555,
    COMP_LOOP_C_922 = 11'd1556,
    COMP_LOOP_C_923 = 11'd1557,
    COMP_LOOP_C_924 = 11'd1558,
    COMP_LOOP_C_925 = 11'd1559,
    COMP_LOOP_C_926 = 11'd1560,
    COMP_LOOP_C_927 = 11'd1561,
    COMP_LOOP_C_928 = 11'd1562,
    COMP_LOOP_C_929 = 11'd1563,
    COMP_LOOP_C_930 = 11'd1564,
    COMP_LOOP_C_931 = 11'd1565,
    COMP_LOOP_C_932 = 11'd1566,
    COMP_LOOP_C_933 = 11'd1567,
    COMP_LOOP_C_934 = 11'd1568,
    COMP_LOOP_C_935 = 11'd1569,
    COMP_LOOP_C_936 = 11'd1570,
    COMP_LOOP_C_937 = 11'd1571,
    COMP_LOOP_C_938 = 11'd1572,
    COMP_LOOP_C_939 = 11'd1573,
    COMP_LOOP_C_940 = 11'd1574,
    COMP_LOOP_C_941 = 11'd1575,
    COMP_LOOP_C_942 = 11'd1576,
    COMP_LOOP_C_943 = 11'd1577,
    COMP_LOOP_C_944 = 11'd1578,
    COMP_LOOP_C_945 = 11'd1579,
    COMP_LOOP_C_946 = 11'd1580,
    COMP_LOOP_C_947 = 11'd1581,
    COMP_LOOP_C_948 = 11'd1582,
    COMP_LOOP_C_949 = 11'd1583,
    COMP_LOOP_C_950 = 11'd1584,
    COMP_LOOP_C_951 = 11'd1585,
    COMP_LOOP_C_952 = 11'd1586,
    COMP_LOOP_C_953 = 11'd1587,
    COMP_LOOP_C_954 = 11'd1588,
    COMP_LOOP_C_955 = 11'd1589,
    COMP_LOOP_C_956 = 11'd1590,
    COMP_LOOP_C_957 = 11'd1591,
    COMP_LOOP_C_958 = 11'd1592,
    COMP_LOOP_C_959 = 11'd1593,
    COMP_LOOP_C_960 = 11'd1594,
    COMP_LOOP_C_961 = 11'd1595,
    COMP_LOOP_16_modExp_1_while_C_0 = 11'd1596,
    COMP_LOOP_16_modExp_1_while_C_1 = 11'd1597,
    COMP_LOOP_16_modExp_1_while_C_2 = 11'd1598,
    COMP_LOOP_16_modExp_1_while_C_3 = 11'd1599,
    COMP_LOOP_16_modExp_1_while_C_4 = 11'd1600,
    COMP_LOOP_16_modExp_1_while_C_5 = 11'd1601,
    COMP_LOOP_16_modExp_1_while_C_6 = 11'd1602,
    COMP_LOOP_16_modExp_1_while_C_7 = 11'd1603,
    COMP_LOOP_16_modExp_1_while_C_8 = 11'd1604,
    COMP_LOOP_16_modExp_1_while_C_9 = 11'd1605,
    COMP_LOOP_16_modExp_1_while_C_10 = 11'd1606,
    COMP_LOOP_16_modExp_1_while_C_11 = 11'd1607,
    COMP_LOOP_16_modExp_1_while_C_12 = 11'd1608,
    COMP_LOOP_16_modExp_1_while_C_13 = 11'd1609,
    COMP_LOOP_16_modExp_1_while_C_14 = 11'd1610,
    COMP_LOOP_16_modExp_1_while_C_15 = 11'd1611,
    COMP_LOOP_16_modExp_1_while_C_16 = 11'd1612,
    COMP_LOOP_16_modExp_1_while_C_17 = 11'd1613,
    COMP_LOOP_16_modExp_1_while_C_18 = 11'd1614,
    COMP_LOOP_16_modExp_1_while_C_19 = 11'd1615,
    COMP_LOOP_16_modExp_1_while_C_20 = 11'd1616,
    COMP_LOOP_16_modExp_1_while_C_21 = 11'd1617,
    COMP_LOOP_16_modExp_1_while_C_22 = 11'd1618,
    COMP_LOOP_16_modExp_1_while_C_23 = 11'd1619,
    COMP_LOOP_16_modExp_1_while_C_24 = 11'd1620,
    COMP_LOOP_16_modExp_1_while_C_25 = 11'd1621,
    COMP_LOOP_16_modExp_1_while_C_26 = 11'd1622,
    COMP_LOOP_16_modExp_1_while_C_27 = 11'd1623,
    COMP_LOOP_16_modExp_1_while_C_28 = 11'd1624,
    COMP_LOOP_16_modExp_1_while_C_29 = 11'd1625,
    COMP_LOOP_16_modExp_1_while_C_30 = 11'd1626,
    COMP_LOOP_16_modExp_1_while_C_31 = 11'd1627,
    COMP_LOOP_16_modExp_1_while_C_32 = 11'd1628,
    COMP_LOOP_16_modExp_1_while_C_33 = 11'd1629,
    COMP_LOOP_16_modExp_1_while_C_34 = 11'd1630,
    COMP_LOOP_16_modExp_1_while_C_35 = 11'd1631,
    COMP_LOOP_16_modExp_1_while_C_36 = 11'd1632,
    COMP_LOOP_16_modExp_1_while_C_37 = 11'd1633,
    COMP_LOOP_16_modExp_1_while_C_38 = 11'd1634,
    COMP_LOOP_C_962 = 11'd1635,
    COMP_LOOP_C_963 = 11'd1636,
    COMP_LOOP_C_964 = 11'd1637,
    COMP_LOOP_C_965 = 11'd1638,
    COMP_LOOP_C_966 = 11'd1639,
    COMP_LOOP_C_967 = 11'd1640,
    COMP_LOOP_C_968 = 11'd1641,
    COMP_LOOP_C_969 = 11'd1642,
    COMP_LOOP_C_970 = 11'd1643,
    COMP_LOOP_C_971 = 11'd1644,
    COMP_LOOP_C_972 = 11'd1645,
    COMP_LOOP_C_973 = 11'd1646,
    COMP_LOOP_C_974 = 11'd1647,
    COMP_LOOP_C_975 = 11'd1648,
    COMP_LOOP_C_976 = 11'd1649,
    COMP_LOOP_C_977 = 11'd1650,
    COMP_LOOP_C_978 = 11'd1651,
    COMP_LOOP_C_979 = 11'd1652,
    COMP_LOOP_C_980 = 11'd1653,
    COMP_LOOP_C_981 = 11'd1654,
    COMP_LOOP_C_982 = 11'd1655,
    COMP_LOOP_C_983 = 11'd1656,
    COMP_LOOP_C_984 = 11'd1657,
    COMP_LOOP_C_985 = 11'd1658,
    COMP_LOOP_C_986 = 11'd1659,
    COMP_LOOP_C_987 = 11'd1660,
    COMP_LOOP_C_988 = 11'd1661,
    COMP_LOOP_C_989 = 11'd1662,
    COMP_LOOP_C_990 = 11'd1663,
    COMP_LOOP_C_991 = 11'd1664,
    COMP_LOOP_C_992 = 11'd1665,
    COMP_LOOP_C_993 = 11'd1666,
    COMP_LOOP_C_994 = 11'd1667,
    COMP_LOOP_C_995 = 11'd1668,
    COMP_LOOP_C_996 = 11'd1669,
    COMP_LOOP_C_997 = 11'd1670,
    COMP_LOOP_C_998 = 11'd1671,
    COMP_LOOP_C_999 = 11'd1672,
    COMP_LOOP_C_1000 = 11'd1673,
    COMP_LOOP_C_1001 = 11'd1674,
    COMP_LOOP_C_1002 = 11'd1675,
    COMP_LOOP_C_1003 = 11'd1676,
    COMP_LOOP_C_1004 = 11'd1677,
    COMP_LOOP_C_1005 = 11'd1678,
    COMP_LOOP_C_1006 = 11'd1679,
    COMP_LOOP_C_1007 = 11'd1680,
    COMP_LOOP_C_1008 = 11'd1681,
    COMP_LOOP_C_1009 = 11'd1682,
    COMP_LOOP_C_1010 = 11'd1683,
    COMP_LOOP_C_1011 = 11'd1684,
    COMP_LOOP_C_1012 = 11'd1685,
    COMP_LOOP_C_1013 = 11'd1686,
    COMP_LOOP_C_1014 = 11'd1687,
    COMP_LOOP_C_1015 = 11'd1688,
    COMP_LOOP_C_1016 = 11'd1689,
    COMP_LOOP_C_1017 = 11'd1690,
    COMP_LOOP_C_1018 = 11'd1691,
    COMP_LOOP_C_1019 = 11'd1692,
    COMP_LOOP_C_1020 = 11'd1693,
    COMP_LOOP_C_1021 = 11'd1694,
    COMP_LOOP_C_1022 = 11'd1695,
    COMP_LOOP_C_1023 = 11'd1696,
    COMP_LOOP_C_1024 = 11'd1697,
    VEC_LOOP_C_0 = 11'd1698,
    STAGE_LOOP_C_9 = 11'd1699,
    main_C_1 = 11'd1700;

  reg [10:0] state_var;
  reg [10:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : inPlaceNTT_DIT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 11'b00000000001;
        state_var_NS = STAGE_LOOP_C_1;
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = STAGE_LOOP_C_2;
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 11'b00000000011;
        state_var_NS = STAGE_LOOP_C_3;
      end
      STAGE_LOOP_C_3 : begin
        fsm_output = 11'b00000000100;
        state_var_NS = STAGE_LOOP_C_4;
      end
      STAGE_LOOP_C_4 : begin
        fsm_output = 11'b00000000101;
        state_var_NS = STAGE_LOOP_C_5;
      end
      STAGE_LOOP_C_5 : begin
        fsm_output = 11'b00000000110;
        state_var_NS = STAGE_LOOP_C_6;
      end
      STAGE_LOOP_C_6 : begin
        fsm_output = 11'b00000000111;
        state_var_NS = STAGE_LOOP_C_7;
      end
      STAGE_LOOP_C_7 : begin
        fsm_output = 11'b00000001000;
        state_var_NS = STAGE_LOOP_C_8;
      end
      STAGE_LOOP_C_8 : begin
        fsm_output = 11'b00000001001;
        if ( STAGE_LOOP_C_8_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      modExp_while_C_0 : begin
        fsm_output = 11'b00000001010;
        state_var_NS = modExp_while_C_1;
      end
      modExp_while_C_1 : begin
        fsm_output = 11'b00000001011;
        state_var_NS = modExp_while_C_2;
      end
      modExp_while_C_2 : begin
        fsm_output = 11'b00000001100;
        state_var_NS = modExp_while_C_3;
      end
      modExp_while_C_3 : begin
        fsm_output = 11'b00000001101;
        state_var_NS = modExp_while_C_4;
      end
      modExp_while_C_4 : begin
        fsm_output = 11'b00000001110;
        state_var_NS = modExp_while_C_5;
      end
      modExp_while_C_5 : begin
        fsm_output = 11'b00000001111;
        state_var_NS = modExp_while_C_6;
      end
      modExp_while_C_6 : begin
        fsm_output = 11'b00000010000;
        state_var_NS = modExp_while_C_7;
      end
      modExp_while_C_7 : begin
        fsm_output = 11'b00000010001;
        state_var_NS = modExp_while_C_8;
      end
      modExp_while_C_8 : begin
        fsm_output = 11'b00000010010;
        state_var_NS = modExp_while_C_9;
      end
      modExp_while_C_9 : begin
        fsm_output = 11'b00000010011;
        state_var_NS = modExp_while_C_10;
      end
      modExp_while_C_10 : begin
        fsm_output = 11'b00000010100;
        state_var_NS = modExp_while_C_11;
      end
      modExp_while_C_11 : begin
        fsm_output = 11'b00000010101;
        state_var_NS = modExp_while_C_12;
      end
      modExp_while_C_12 : begin
        fsm_output = 11'b00000010110;
        state_var_NS = modExp_while_C_13;
      end
      modExp_while_C_13 : begin
        fsm_output = 11'b00000010111;
        state_var_NS = modExp_while_C_14;
      end
      modExp_while_C_14 : begin
        fsm_output = 11'b00000011000;
        state_var_NS = modExp_while_C_15;
      end
      modExp_while_C_15 : begin
        fsm_output = 11'b00000011001;
        state_var_NS = modExp_while_C_16;
      end
      modExp_while_C_16 : begin
        fsm_output = 11'b00000011010;
        state_var_NS = modExp_while_C_17;
      end
      modExp_while_C_17 : begin
        fsm_output = 11'b00000011011;
        state_var_NS = modExp_while_C_18;
      end
      modExp_while_C_18 : begin
        fsm_output = 11'b00000011100;
        state_var_NS = modExp_while_C_19;
      end
      modExp_while_C_19 : begin
        fsm_output = 11'b00000011101;
        state_var_NS = modExp_while_C_20;
      end
      modExp_while_C_20 : begin
        fsm_output = 11'b00000011110;
        state_var_NS = modExp_while_C_21;
      end
      modExp_while_C_21 : begin
        fsm_output = 11'b00000011111;
        state_var_NS = modExp_while_C_22;
      end
      modExp_while_C_22 : begin
        fsm_output = 11'b00000100000;
        state_var_NS = modExp_while_C_23;
      end
      modExp_while_C_23 : begin
        fsm_output = 11'b00000100001;
        state_var_NS = modExp_while_C_24;
      end
      modExp_while_C_24 : begin
        fsm_output = 11'b00000100010;
        state_var_NS = modExp_while_C_25;
      end
      modExp_while_C_25 : begin
        fsm_output = 11'b00000100011;
        state_var_NS = modExp_while_C_26;
      end
      modExp_while_C_26 : begin
        fsm_output = 11'b00000100100;
        state_var_NS = modExp_while_C_27;
      end
      modExp_while_C_27 : begin
        fsm_output = 11'b00000100101;
        state_var_NS = modExp_while_C_28;
      end
      modExp_while_C_28 : begin
        fsm_output = 11'b00000100110;
        state_var_NS = modExp_while_C_29;
      end
      modExp_while_C_29 : begin
        fsm_output = 11'b00000100111;
        state_var_NS = modExp_while_C_30;
      end
      modExp_while_C_30 : begin
        fsm_output = 11'b00000101000;
        state_var_NS = modExp_while_C_31;
      end
      modExp_while_C_31 : begin
        fsm_output = 11'b00000101001;
        state_var_NS = modExp_while_C_32;
      end
      modExp_while_C_32 : begin
        fsm_output = 11'b00000101010;
        state_var_NS = modExp_while_C_33;
      end
      modExp_while_C_33 : begin
        fsm_output = 11'b00000101011;
        state_var_NS = modExp_while_C_34;
      end
      modExp_while_C_34 : begin
        fsm_output = 11'b00000101100;
        state_var_NS = modExp_while_C_35;
      end
      modExp_while_C_35 : begin
        fsm_output = 11'b00000101101;
        state_var_NS = modExp_while_C_36;
      end
      modExp_while_C_36 : begin
        fsm_output = 11'b00000101110;
        state_var_NS = modExp_while_C_37;
      end
      modExp_while_C_37 : begin
        fsm_output = 11'b00000101111;
        state_var_NS = modExp_while_C_38;
      end
      modExp_while_C_38 : begin
        fsm_output = 11'b00000110000;
        if ( modExp_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_0;
        end
        else begin
          state_var_NS = modExp_while_C_0;
        end
      end
      COMP_LOOP_C_0 : begin
        fsm_output = 11'b00000110001;
        state_var_NS = COMP_LOOP_C_1;
      end
      COMP_LOOP_C_1 : begin
        fsm_output = 11'b00000110010;
        if ( COMP_LOOP_C_1_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_1_modExp_1_while_C_0 : begin
        fsm_output = 11'b00000110011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_1;
      end
      COMP_LOOP_1_modExp_1_while_C_1 : begin
        fsm_output = 11'b00000110100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_2;
      end
      COMP_LOOP_1_modExp_1_while_C_2 : begin
        fsm_output = 11'b00000110101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_3;
      end
      COMP_LOOP_1_modExp_1_while_C_3 : begin
        fsm_output = 11'b00000110110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_4;
      end
      COMP_LOOP_1_modExp_1_while_C_4 : begin
        fsm_output = 11'b00000110111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_5;
      end
      COMP_LOOP_1_modExp_1_while_C_5 : begin
        fsm_output = 11'b00000111000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_6;
      end
      COMP_LOOP_1_modExp_1_while_C_6 : begin
        fsm_output = 11'b00000111001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_7;
      end
      COMP_LOOP_1_modExp_1_while_C_7 : begin
        fsm_output = 11'b00000111010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_8;
      end
      COMP_LOOP_1_modExp_1_while_C_8 : begin
        fsm_output = 11'b00000111011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_9;
      end
      COMP_LOOP_1_modExp_1_while_C_9 : begin
        fsm_output = 11'b00000111100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_10;
      end
      COMP_LOOP_1_modExp_1_while_C_10 : begin
        fsm_output = 11'b00000111101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_11;
      end
      COMP_LOOP_1_modExp_1_while_C_11 : begin
        fsm_output = 11'b00000111110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_12;
      end
      COMP_LOOP_1_modExp_1_while_C_12 : begin
        fsm_output = 11'b00000111111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_13;
      end
      COMP_LOOP_1_modExp_1_while_C_13 : begin
        fsm_output = 11'b00001000000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_14;
      end
      COMP_LOOP_1_modExp_1_while_C_14 : begin
        fsm_output = 11'b00001000001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_15;
      end
      COMP_LOOP_1_modExp_1_while_C_15 : begin
        fsm_output = 11'b00001000010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_16;
      end
      COMP_LOOP_1_modExp_1_while_C_16 : begin
        fsm_output = 11'b00001000011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_17;
      end
      COMP_LOOP_1_modExp_1_while_C_17 : begin
        fsm_output = 11'b00001000100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_18;
      end
      COMP_LOOP_1_modExp_1_while_C_18 : begin
        fsm_output = 11'b00001000101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_19;
      end
      COMP_LOOP_1_modExp_1_while_C_19 : begin
        fsm_output = 11'b00001000110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_20;
      end
      COMP_LOOP_1_modExp_1_while_C_20 : begin
        fsm_output = 11'b00001000111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_21;
      end
      COMP_LOOP_1_modExp_1_while_C_21 : begin
        fsm_output = 11'b00001001000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_22;
      end
      COMP_LOOP_1_modExp_1_while_C_22 : begin
        fsm_output = 11'b00001001001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_23;
      end
      COMP_LOOP_1_modExp_1_while_C_23 : begin
        fsm_output = 11'b00001001010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_24;
      end
      COMP_LOOP_1_modExp_1_while_C_24 : begin
        fsm_output = 11'b00001001011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_25;
      end
      COMP_LOOP_1_modExp_1_while_C_25 : begin
        fsm_output = 11'b00001001100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_26;
      end
      COMP_LOOP_1_modExp_1_while_C_26 : begin
        fsm_output = 11'b00001001101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_27;
      end
      COMP_LOOP_1_modExp_1_while_C_27 : begin
        fsm_output = 11'b00001001110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_28;
      end
      COMP_LOOP_1_modExp_1_while_C_28 : begin
        fsm_output = 11'b00001001111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_29;
      end
      COMP_LOOP_1_modExp_1_while_C_29 : begin
        fsm_output = 11'b00001010000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_30;
      end
      COMP_LOOP_1_modExp_1_while_C_30 : begin
        fsm_output = 11'b00001010001;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_31;
      end
      COMP_LOOP_1_modExp_1_while_C_31 : begin
        fsm_output = 11'b00001010010;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_32;
      end
      COMP_LOOP_1_modExp_1_while_C_32 : begin
        fsm_output = 11'b00001010011;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_33;
      end
      COMP_LOOP_1_modExp_1_while_C_33 : begin
        fsm_output = 11'b00001010100;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_34;
      end
      COMP_LOOP_1_modExp_1_while_C_34 : begin
        fsm_output = 11'b00001010101;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_35;
      end
      COMP_LOOP_1_modExp_1_while_C_35 : begin
        fsm_output = 11'b00001010110;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_36;
      end
      COMP_LOOP_1_modExp_1_while_C_36 : begin
        fsm_output = 11'b00001010111;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_37;
      end
      COMP_LOOP_1_modExp_1_while_C_37 : begin
        fsm_output = 11'b00001011000;
        state_var_NS = COMP_LOOP_1_modExp_1_while_C_38;
      end
      COMP_LOOP_1_modExp_1_while_C_38 : begin
        fsm_output = 11'b00001011001;
        if ( COMP_LOOP_1_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_2;
        end
        else begin
          state_var_NS = COMP_LOOP_1_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_2 : begin
        fsm_output = 11'b00001011010;
        state_var_NS = COMP_LOOP_C_3;
      end
      COMP_LOOP_C_3 : begin
        fsm_output = 11'b00001011011;
        state_var_NS = COMP_LOOP_C_4;
      end
      COMP_LOOP_C_4 : begin
        fsm_output = 11'b00001011100;
        state_var_NS = COMP_LOOP_C_5;
      end
      COMP_LOOP_C_5 : begin
        fsm_output = 11'b00001011101;
        state_var_NS = COMP_LOOP_C_6;
      end
      COMP_LOOP_C_6 : begin
        fsm_output = 11'b00001011110;
        state_var_NS = COMP_LOOP_C_7;
      end
      COMP_LOOP_C_7 : begin
        fsm_output = 11'b00001011111;
        state_var_NS = COMP_LOOP_C_8;
      end
      COMP_LOOP_C_8 : begin
        fsm_output = 11'b00001100000;
        state_var_NS = COMP_LOOP_C_9;
      end
      COMP_LOOP_C_9 : begin
        fsm_output = 11'b00001100001;
        state_var_NS = COMP_LOOP_C_10;
      end
      COMP_LOOP_C_10 : begin
        fsm_output = 11'b00001100010;
        state_var_NS = COMP_LOOP_C_11;
      end
      COMP_LOOP_C_11 : begin
        fsm_output = 11'b00001100011;
        state_var_NS = COMP_LOOP_C_12;
      end
      COMP_LOOP_C_12 : begin
        fsm_output = 11'b00001100100;
        state_var_NS = COMP_LOOP_C_13;
      end
      COMP_LOOP_C_13 : begin
        fsm_output = 11'b00001100101;
        state_var_NS = COMP_LOOP_C_14;
      end
      COMP_LOOP_C_14 : begin
        fsm_output = 11'b00001100110;
        state_var_NS = COMP_LOOP_C_15;
      end
      COMP_LOOP_C_15 : begin
        fsm_output = 11'b00001100111;
        state_var_NS = COMP_LOOP_C_16;
      end
      COMP_LOOP_C_16 : begin
        fsm_output = 11'b00001101000;
        state_var_NS = COMP_LOOP_C_17;
      end
      COMP_LOOP_C_17 : begin
        fsm_output = 11'b00001101001;
        state_var_NS = COMP_LOOP_C_18;
      end
      COMP_LOOP_C_18 : begin
        fsm_output = 11'b00001101010;
        state_var_NS = COMP_LOOP_C_19;
      end
      COMP_LOOP_C_19 : begin
        fsm_output = 11'b00001101011;
        state_var_NS = COMP_LOOP_C_20;
      end
      COMP_LOOP_C_20 : begin
        fsm_output = 11'b00001101100;
        state_var_NS = COMP_LOOP_C_21;
      end
      COMP_LOOP_C_21 : begin
        fsm_output = 11'b00001101101;
        state_var_NS = COMP_LOOP_C_22;
      end
      COMP_LOOP_C_22 : begin
        fsm_output = 11'b00001101110;
        state_var_NS = COMP_LOOP_C_23;
      end
      COMP_LOOP_C_23 : begin
        fsm_output = 11'b00001101111;
        state_var_NS = COMP_LOOP_C_24;
      end
      COMP_LOOP_C_24 : begin
        fsm_output = 11'b00001110000;
        state_var_NS = COMP_LOOP_C_25;
      end
      COMP_LOOP_C_25 : begin
        fsm_output = 11'b00001110001;
        state_var_NS = COMP_LOOP_C_26;
      end
      COMP_LOOP_C_26 : begin
        fsm_output = 11'b00001110010;
        state_var_NS = COMP_LOOP_C_27;
      end
      COMP_LOOP_C_27 : begin
        fsm_output = 11'b00001110011;
        state_var_NS = COMP_LOOP_C_28;
      end
      COMP_LOOP_C_28 : begin
        fsm_output = 11'b00001110100;
        state_var_NS = COMP_LOOP_C_29;
      end
      COMP_LOOP_C_29 : begin
        fsm_output = 11'b00001110101;
        state_var_NS = COMP_LOOP_C_30;
      end
      COMP_LOOP_C_30 : begin
        fsm_output = 11'b00001110110;
        state_var_NS = COMP_LOOP_C_31;
      end
      COMP_LOOP_C_31 : begin
        fsm_output = 11'b00001110111;
        state_var_NS = COMP_LOOP_C_32;
      end
      COMP_LOOP_C_32 : begin
        fsm_output = 11'b00001111000;
        state_var_NS = COMP_LOOP_C_33;
      end
      COMP_LOOP_C_33 : begin
        fsm_output = 11'b00001111001;
        state_var_NS = COMP_LOOP_C_34;
      end
      COMP_LOOP_C_34 : begin
        fsm_output = 11'b00001111010;
        state_var_NS = COMP_LOOP_C_35;
      end
      COMP_LOOP_C_35 : begin
        fsm_output = 11'b00001111011;
        state_var_NS = COMP_LOOP_C_36;
      end
      COMP_LOOP_C_36 : begin
        fsm_output = 11'b00001111100;
        state_var_NS = COMP_LOOP_C_37;
      end
      COMP_LOOP_C_37 : begin
        fsm_output = 11'b00001111101;
        state_var_NS = COMP_LOOP_C_38;
      end
      COMP_LOOP_C_38 : begin
        fsm_output = 11'b00001111110;
        state_var_NS = COMP_LOOP_C_39;
      end
      COMP_LOOP_C_39 : begin
        fsm_output = 11'b00001111111;
        state_var_NS = COMP_LOOP_C_40;
      end
      COMP_LOOP_C_40 : begin
        fsm_output = 11'b00010000000;
        state_var_NS = COMP_LOOP_C_41;
      end
      COMP_LOOP_C_41 : begin
        fsm_output = 11'b00010000001;
        state_var_NS = COMP_LOOP_C_42;
      end
      COMP_LOOP_C_42 : begin
        fsm_output = 11'b00010000010;
        state_var_NS = COMP_LOOP_C_43;
      end
      COMP_LOOP_C_43 : begin
        fsm_output = 11'b00010000011;
        state_var_NS = COMP_LOOP_C_44;
      end
      COMP_LOOP_C_44 : begin
        fsm_output = 11'b00010000100;
        state_var_NS = COMP_LOOP_C_45;
      end
      COMP_LOOP_C_45 : begin
        fsm_output = 11'b00010000101;
        state_var_NS = COMP_LOOP_C_46;
      end
      COMP_LOOP_C_46 : begin
        fsm_output = 11'b00010000110;
        state_var_NS = COMP_LOOP_C_47;
      end
      COMP_LOOP_C_47 : begin
        fsm_output = 11'b00010000111;
        state_var_NS = COMP_LOOP_C_48;
      end
      COMP_LOOP_C_48 : begin
        fsm_output = 11'b00010001000;
        state_var_NS = COMP_LOOP_C_49;
      end
      COMP_LOOP_C_49 : begin
        fsm_output = 11'b00010001001;
        state_var_NS = COMP_LOOP_C_50;
      end
      COMP_LOOP_C_50 : begin
        fsm_output = 11'b00010001010;
        state_var_NS = COMP_LOOP_C_51;
      end
      COMP_LOOP_C_51 : begin
        fsm_output = 11'b00010001011;
        state_var_NS = COMP_LOOP_C_52;
      end
      COMP_LOOP_C_52 : begin
        fsm_output = 11'b00010001100;
        state_var_NS = COMP_LOOP_C_53;
      end
      COMP_LOOP_C_53 : begin
        fsm_output = 11'b00010001101;
        state_var_NS = COMP_LOOP_C_54;
      end
      COMP_LOOP_C_54 : begin
        fsm_output = 11'b00010001110;
        state_var_NS = COMP_LOOP_C_55;
      end
      COMP_LOOP_C_55 : begin
        fsm_output = 11'b00010001111;
        state_var_NS = COMP_LOOP_C_56;
      end
      COMP_LOOP_C_56 : begin
        fsm_output = 11'b00010010000;
        state_var_NS = COMP_LOOP_C_57;
      end
      COMP_LOOP_C_57 : begin
        fsm_output = 11'b00010010001;
        state_var_NS = COMP_LOOP_C_58;
      end
      COMP_LOOP_C_58 : begin
        fsm_output = 11'b00010010010;
        state_var_NS = COMP_LOOP_C_59;
      end
      COMP_LOOP_C_59 : begin
        fsm_output = 11'b00010010011;
        state_var_NS = COMP_LOOP_C_60;
      end
      COMP_LOOP_C_60 : begin
        fsm_output = 11'b00010010100;
        state_var_NS = COMP_LOOP_C_61;
      end
      COMP_LOOP_C_61 : begin
        fsm_output = 11'b00010010101;
        state_var_NS = COMP_LOOP_C_62;
      end
      COMP_LOOP_C_62 : begin
        fsm_output = 11'b00010010110;
        state_var_NS = COMP_LOOP_C_63;
      end
      COMP_LOOP_C_63 : begin
        fsm_output = 11'b00010010111;
        state_var_NS = COMP_LOOP_C_64;
      end
      COMP_LOOP_C_64 : begin
        fsm_output = 11'b00010011000;
        if ( COMP_LOOP_C_64_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_65;
        end
      end
      COMP_LOOP_C_65 : begin
        fsm_output = 11'b00010011001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
      end
      COMP_LOOP_2_modExp_1_while_C_0 : begin
        fsm_output = 11'b00010011010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_1;
      end
      COMP_LOOP_2_modExp_1_while_C_1 : begin
        fsm_output = 11'b00010011011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_2;
      end
      COMP_LOOP_2_modExp_1_while_C_2 : begin
        fsm_output = 11'b00010011100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_3;
      end
      COMP_LOOP_2_modExp_1_while_C_3 : begin
        fsm_output = 11'b00010011101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_4;
      end
      COMP_LOOP_2_modExp_1_while_C_4 : begin
        fsm_output = 11'b00010011110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_5;
      end
      COMP_LOOP_2_modExp_1_while_C_5 : begin
        fsm_output = 11'b00010011111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_6;
      end
      COMP_LOOP_2_modExp_1_while_C_6 : begin
        fsm_output = 11'b00010100000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_7;
      end
      COMP_LOOP_2_modExp_1_while_C_7 : begin
        fsm_output = 11'b00010100001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_8;
      end
      COMP_LOOP_2_modExp_1_while_C_8 : begin
        fsm_output = 11'b00010100010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_9;
      end
      COMP_LOOP_2_modExp_1_while_C_9 : begin
        fsm_output = 11'b00010100011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_10;
      end
      COMP_LOOP_2_modExp_1_while_C_10 : begin
        fsm_output = 11'b00010100100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_11;
      end
      COMP_LOOP_2_modExp_1_while_C_11 : begin
        fsm_output = 11'b00010100101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_12;
      end
      COMP_LOOP_2_modExp_1_while_C_12 : begin
        fsm_output = 11'b00010100110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_13;
      end
      COMP_LOOP_2_modExp_1_while_C_13 : begin
        fsm_output = 11'b00010100111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_14;
      end
      COMP_LOOP_2_modExp_1_while_C_14 : begin
        fsm_output = 11'b00010101000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_15;
      end
      COMP_LOOP_2_modExp_1_while_C_15 : begin
        fsm_output = 11'b00010101001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_16;
      end
      COMP_LOOP_2_modExp_1_while_C_16 : begin
        fsm_output = 11'b00010101010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_17;
      end
      COMP_LOOP_2_modExp_1_while_C_17 : begin
        fsm_output = 11'b00010101011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_18;
      end
      COMP_LOOP_2_modExp_1_while_C_18 : begin
        fsm_output = 11'b00010101100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_19;
      end
      COMP_LOOP_2_modExp_1_while_C_19 : begin
        fsm_output = 11'b00010101101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_20;
      end
      COMP_LOOP_2_modExp_1_while_C_20 : begin
        fsm_output = 11'b00010101110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_21;
      end
      COMP_LOOP_2_modExp_1_while_C_21 : begin
        fsm_output = 11'b00010101111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_22;
      end
      COMP_LOOP_2_modExp_1_while_C_22 : begin
        fsm_output = 11'b00010110000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_23;
      end
      COMP_LOOP_2_modExp_1_while_C_23 : begin
        fsm_output = 11'b00010110001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_24;
      end
      COMP_LOOP_2_modExp_1_while_C_24 : begin
        fsm_output = 11'b00010110010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_25;
      end
      COMP_LOOP_2_modExp_1_while_C_25 : begin
        fsm_output = 11'b00010110011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_26;
      end
      COMP_LOOP_2_modExp_1_while_C_26 : begin
        fsm_output = 11'b00010110100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_27;
      end
      COMP_LOOP_2_modExp_1_while_C_27 : begin
        fsm_output = 11'b00010110101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_28;
      end
      COMP_LOOP_2_modExp_1_while_C_28 : begin
        fsm_output = 11'b00010110110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_29;
      end
      COMP_LOOP_2_modExp_1_while_C_29 : begin
        fsm_output = 11'b00010110111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_30;
      end
      COMP_LOOP_2_modExp_1_while_C_30 : begin
        fsm_output = 11'b00010111000;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_31;
      end
      COMP_LOOP_2_modExp_1_while_C_31 : begin
        fsm_output = 11'b00010111001;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_32;
      end
      COMP_LOOP_2_modExp_1_while_C_32 : begin
        fsm_output = 11'b00010111010;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_33;
      end
      COMP_LOOP_2_modExp_1_while_C_33 : begin
        fsm_output = 11'b00010111011;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_34;
      end
      COMP_LOOP_2_modExp_1_while_C_34 : begin
        fsm_output = 11'b00010111100;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_35;
      end
      COMP_LOOP_2_modExp_1_while_C_35 : begin
        fsm_output = 11'b00010111101;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_36;
      end
      COMP_LOOP_2_modExp_1_while_C_36 : begin
        fsm_output = 11'b00010111110;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_37;
      end
      COMP_LOOP_2_modExp_1_while_C_37 : begin
        fsm_output = 11'b00010111111;
        state_var_NS = COMP_LOOP_2_modExp_1_while_C_38;
      end
      COMP_LOOP_2_modExp_1_while_C_38 : begin
        fsm_output = 11'b00011000000;
        if ( COMP_LOOP_2_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_66;
        end
        else begin
          state_var_NS = COMP_LOOP_2_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_66 : begin
        fsm_output = 11'b00011000001;
        state_var_NS = COMP_LOOP_C_67;
      end
      COMP_LOOP_C_67 : begin
        fsm_output = 11'b00011000010;
        state_var_NS = COMP_LOOP_C_68;
      end
      COMP_LOOP_C_68 : begin
        fsm_output = 11'b00011000011;
        state_var_NS = COMP_LOOP_C_69;
      end
      COMP_LOOP_C_69 : begin
        fsm_output = 11'b00011000100;
        state_var_NS = COMP_LOOP_C_70;
      end
      COMP_LOOP_C_70 : begin
        fsm_output = 11'b00011000101;
        state_var_NS = COMP_LOOP_C_71;
      end
      COMP_LOOP_C_71 : begin
        fsm_output = 11'b00011000110;
        state_var_NS = COMP_LOOP_C_72;
      end
      COMP_LOOP_C_72 : begin
        fsm_output = 11'b00011000111;
        state_var_NS = COMP_LOOP_C_73;
      end
      COMP_LOOP_C_73 : begin
        fsm_output = 11'b00011001000;
        state_var_NS = COMP_LOOP_C_74;
      end
      COMP_LOOP_C_74 : begin
        fsm_output = 11'b00011001001;
        state_var_NS = COMP_LOOP_C_75;
      end
      COMP_LOOP_C_75 : begin
        fsm_output = 11'b00011001010;
        state_var_NS = COMP_LOOP_C_76;
      end
      COMP_LOOP_C_76 : begin
        fsm_output = 11'b00011001011;
        state_var_NS = COMP_LOOP_C_77;
      end
      COMP_LOOP_C_77 : begin
        fsm_output = 11'b00011001100;
        state_var_NS = COMP_LOOP_C_78;
      end
      COMP_LOOP_C_78 : begin
        fsm_output = 11'b00011001101;
        state_var_NS = COMP_LOOP_C_79;
      end
      COMP_LOOP_C_79 : begin
        fsm_output = 11'b00011001110;
        state_var_NS = COMP_LOOP_C_80;
      end
      COMP_LOOP_C_80 : begin
        fsm_output = 11'b00011001111;
        state_var_NS = COMP_LOOP_C_81;
      end
      COMP_LOOP_C_81 : begin
        fsm_output = 11'b00011010000;
        state_var_NS = COMP_LOOP_C_82;
      end
      COMP_LOOP_C_82 : begin
        fsm_output = 11'b00011010001;
        state_var_NS = COMP_LOOP_C_83;
      end
      COMP_LOOP_C_83 : begin
        fsm_output = 11'b00011010010;
        state_var_NS = COMP_LOOP_C_84;
      end
      COMP_LOOP_C_84 : begin
        fsm_output = 11'b00011010011;
        state_var_NS = COMP_LOOP_C_85;
      end
      COMP_LOOP_C_85 : begin
        fsm_output = 11'b00011010100;
        state_var_NS = COMP_LOOP_C_86;
      end
      COMP_LOOP_C_86 : begin
        fsm_output = 11'b00011010101;
        state_var_NS = COMP_LOOP_C_87;
      end
      COMP_LOOP_C_87 : begin
        fsm_output = 11'b00011010110;
        state_var_NS = COMP_LOOP_C_88;
      end
      COMP_LOOP_C_88 : begin
        fsm_output = 11'b00011010111;
        state_var_NS = COMP_LOOP_C_89;
      end
      COMP_LOOP_C_89 : begin
        fsm_output = 11'b00011011000;
        state_var_NS = COMP_LOOP_C_90;
      end
      COMP_LOOP_C_90 : begin
        fsm_output = 11'b00011011001;
        state_var_NS = COMP_LOOP_C_91;
      end
      COMP_LOOP_C_91 : begin
        fsm_output = 11'b00011011010;
        state_var_NS = COMP_LOOP_C_92;
      end
      COMP_LOOP_C_92 : begin
        fsm_output = 11'b00011011011;
        state_var_NS = COMP_LOOP_C_93;
      end
      COMP_LOOP_C_93 : begin
        fsm_output = 11'b00011011100;
        state_var_NS = COMP_LOOP_C_94;
      end
      COMP_LOOP_C_94 : begin
        fsm_output = 11'b00011011101;
        state_var_NS = COMP_LOOP_C_95;
      end
      COMP_LOOP_C_95 : begin
        fsm_output = 11'b00011011110;
        state_var_NS = COMP_LOOP_C_96;
      end
      COMP_LOOP_C_96 : begin
        fsm_output = 11'b00011011111;
        state_var_NS = COMP_LOOP_C_97;
      end
      COMP_LOOP_C_97 : begin
        fsm_output = 11'b00011100000;
        state_var_NS = COMP_LOOP_C_98;
      end
      COMP_LOOP_C_98 : begin
        fsm_output = 11'b00011100001;
        state_var_NS = COMP_LOOP_C_99;
      end
      COMP_LOOP_C_99 : begin
        fsm_output = 11'b00011100010;
        state_var_NS = COMP_LOOP_C_100;
      end
      COMP_LOOP_C_100 : begin
        fsm_output = 11'b00011100011;
        state_var_NS = COMP_LOOP_C_101;
      end
      COMP_LOOP_C_101 : begin
        fsm_output = 11'b00011100100;
        state_var_NS = COMP_LOOP_C_102;
      end
      COMP_LOOP_C_102 : begin
        fsm_output = 11'b00011100101;
        state_var_NS = COMP_LOOP_C_103;
      end
      COMP_LOOP_C_103 : begin
        fsm_output = 11'b00011100110;
        state_var_NS = COMP_LOOP_C_104;
      end
      COMP_LOOP_C_104 : begin
        fsm_output = 11'b00011100111;
        state_var_NS = COMP_LOOP_C_105;
      end
      COMP_LOOP_C_105 : begin
        fsm_output = 11'b00011101000;
        state_var_NS = COMP_LOOP_C_106;
      end
      COMP_LOOP_C_106 : begin
        fsm_output = 11'b00011101001;
        state_var_NS = COMP_LOOP_C_107;
      end
      COMP_LOOP_C_107 : begin
        fsm_output = 11'b00011101010;
        state_var_NS = COMP_LOOP_C_108;
      end
      COMP_LOOP_C_108 : begin
        fsm_output = 11'b00011101011;
        state_var_NS = COMP_LOOP_C_109;
      end
      COMP_LOOP_C_109 : begin
        fsm_output = 11'b00011101100;
        state_var_NS = COMP_LOOP_C_110;
      end
      COMP_LOOP_C_110 : begin
        fsm_output = 11'b00011101101;
        state_var_NS = COMP_LOOP_C_111;
      end
      COMP_LOOP_C_111 : begin
        fsm_output = 11'b00011101110;
        state_var_NS = COMP_LOOP_C_112;
      end
      COMP_LOOP_C_112 : begin
        fsm_output = 11'b00011101111;
        state_var_NS = COMP_LOOP_C_113;
      end
      COMP_LOOP_C_113 : begin
        fsm_output = 11'b00011110000;
        state_var_NS = COMP_LOOP_C_114;
      end
      COMP_LOOP_C_114 : begin
        fsm_output = 11'b00011110001;
        state_var_NS = COMP_LOOP_C_115;
      end
      COMP_LOOP_C_115 : begin
        fsm_output = 11'b00011110010;
        state_var_NS = COMP_LOOP_C_116;
      end
      COMP_LOOP_C_116 : begin
        fsm_output = 11'b00011110011;
        state_var_NS = COMP_LOOP_C_117;
      end
      COMP_LOOP_C_117 : begin
        fsm_output = 11'b00011110100;
        state_var_NS = COMP_LOOP_C_118;
      end
      COMP_LOOP_C_118 : begin
        fsm_output = 11'b00011110101;
        state_var_NS = COMP_LOOP_C_119;
      end
      COMP_LOOP_C_119 : begin
        fsm_output = 11'b00011110110;
        state_var_NS = COMP_LOOP_C_120;
      end
      COMP_LOOP_C_120 : begin
        fsm_output = 11'b00011110111;
        state_var_NS = COMP_LOOP_C_121;
      end
      COMP_LOOP_C_121 : begin
        fsm_output = 11'b00011111000;
        state_var_NS = COMP_LOOP_C_122;
      end
      COMP_LOOP_C_122 : begin
        fsm_output = 11'b00011111001;
        state_var_NS = COMP_LOOP_C_123;
      end
      COMP_LOOP_C_123 : begin
        fsm_output = 11'b00011111010;
        state_var_NS = COMP_LOOP_C_124;
      end
      COMP_LOOP_C_124 : begin
        fsm_output = 11'b00011111011;
        state_var_NS = COMP_LOOP_C_125;
      end
      COMP_LOOP_C_125 : begin
        fsm_output = 11'b00011111100;
        state_var_NS = COMP_LOOP_C_126;
      end
      COMP_LOOP_C_126 : begin
        fsm_output = 11'b00011111101;
        state_var_NS = COMP_LOOP_C_127;
      end
      COMP_LOOP_C_127 : begin
        fsm_output = 11'b00011111110;
        state_var_NS = COMP_LOOP_C_128;
      end
      COMP_LOOP_C_128 : begin
        fsm_output = 11'b00011111111;
        if ( COMP_LOOP_C_128_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_129;
        end
      end
      COMP_LOOP_C_129 : begin
        fsm_output = 11'b00100000000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
      end
      COMP_LOOP_3_modExp_1_while_C_0 : begin
        fsm_output = 11'b00100000001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_1;
      end
      COMP_LOOP_3_modExp_1_while_C_1 : begin
        fsm_output = 11'b00100000010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_2;
      end
      COMP_LOOP_3_modExp_1_while_C_2 : begin
        fsm_output = 11'b00100000011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_3;
      end
      COMP_LOOP_3_modExp_1_while_C_3 : begin
        fsm_output = 11'b00100000100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_4;
      end
      COMP_LOOP_3_modExp_1_while_C_4 : begin
        fsm_output = 11'b00100000101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_5;
      end
      COMP_LOOP_3_modExp_1_while_C_5 : begin
        fsm_output = 11'b00100000110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_6;
      end
      COMP_LOOP_3_modExp_1_while_C_6 : begin
        fsm_output = 11'b00100000111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_7;
      end
      COMP_LOOP_3_modExp_1_while_C_7 : begin
        fsm_output = 11'b00100001000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_8;
      end
      COMP_LOOP_3_modExp_1_while_C_8 : begin
        fsm_output = 11'b00100001001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_9;
      end
      COMP_LOOP_3_modExp_1_while_C_9 : begin
        fsm_output = 11'b00100001010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_10;
      end
      COMP_LOOP_3_modExp_1_while_C_10 : begin
        fsm_output = 11'b00100001011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_11;
      end
      COMP_LOOP_3_modExp_1_while_C_11 : begin
        fsm_output = 11'b00100001100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_12;
      end
      COMP_LOOP_3_modExp_1_while_C_12 : begin
        fsm_output = 11'b00100001101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_13;
      end
      COMP_LOOP_3_modExp_1_while_C_13 : begin
        fsm_output = 11'b00100001110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_14;
      end
      COMP_LOOP_3_modExp_1_while_C_14 : begin
        fsm_output = 11'b00100001111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_15;
      end
      COMP_LOOP_3_modExp_1_while_C_15 : begin
        fsm_output = 11'b00100010000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_16;
      end
      COMP_LOOP_3_modExp_1_while_C_16 : begin
        fsm_output = 11'b00100010001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_17;
      end
      COMP_LOOP_3_modExp_1_while_C_17 : begin
        fsm_output = 11'b00100010010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_18;
      end
      COMP_LOOP_3_modExp_1_while_C_18 : begin
        fsm_output = 11'b00100010011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_19;
      end
      COMP_LOOP_3_modExp_1_while_C_19 : begin
        fsm_output = 11'b00100010100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_20;
      end
      COMP_LOOP_3_modExp_1_while_C_20 : begin
        fsm_output = 11'b00100010101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_21;
      end
      COMP_LOOP_3_modExp_1_while_C_21 : begin
        fsm_output = 11'b00100010110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_22;
      end
      COMP_LOOP_3_modExp_1_while_C_22 : begin
        fsm_output = 11'b00100010111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_23;
      end
      COMP_LOOP_3_modExp_1_while_C_23 : begin
        fsm_output = 11'b00100011000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_24;
      end
      COMP_LOOP_3_modExp_1_while_C_24 : begin
        fsm_output = 11'b00100011001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_25;
      end
      COMP_LOOP_3_modExp_1_while_C_25 : begin
        fsm_output = 11'b00100011010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_26;
      end
      COMP_LOOP_3_modExp_1_while_C_26 : begin
        fsm_output = 11'b00100011011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_27;
      end
      COMP_LOOP_3_modExp_1_while_C_27 : begin
        fsm_output = 11'b00100011100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_28;
      end
      COMP_LOOP_3_modExp_1_while_C_28 : begin
        fsm_output = 11'b00100011101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_29;
      end
      COMP_LOOP_3_modExp_1_while_C_29 : begin
        fsm_output = 11'b00100011110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_30;
      end
      COMP_LOOP_3_modExp_1_while_C_30 : begin
        fsm_output = 11'b00100011111;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_31;
      end
      COMP_LOOP_3_modExp_1_while_C_31 : begin
        fsm_output = 11'b00100100000;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_32;
      end
      COMP_LOOP_3_modExp_1_while_C_32 : begin
        fsm_output = 11'b00100100001;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_33;
      end
      COMP_LOOP_3_modExp_1_while_C_33 : begin
        fsm_output = 11'b00100100010;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_34;
      end
      COMP_LOOP_3_modExp_1_while_C_34 : begin
        fsm_output = 11'b00100100011;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_35;
      end
      COMP_LOOP_3_modExp_1_while_C_35 : begin
        fsm_output = 11'b00100100100;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_36;
      end
      COMP_LOOP_3_modExp_1_while_C_36 : begin
        fsm_output = 11'b00100100101;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_37;
      end
      COMP_LOOP_3_modExp_1_while_C_37 : begin
        fsm_output = 11'b00100100110;
        state_var_NS = COMP_LOOP_3_modExp_1_while_C_38;
      end
      COMP_LOOP_3_modExp_1_while_C_38 : begin
        fsm_output = 11'b00100100111;
        if ( COMP_LOOP_3_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_130;
        end
        else begin
          state_var_NS = COMP_LOOP_3_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_130 : begin
        fsm_output = 11'b00100101000;
        state_var_NS = COMP_LOOP_C_131;
      end
      COMP_LOOP_C_131 : begin
        fsm_output = 11'b00100101001;
        state_var_NS = COMP_LOOP_C_132;
      end
      COMP_LOOP_C_132 : begin
        fsm_output = 11'b00100101010;
        state_var_NS = COMP_LOOP_C_133;
      end
      COMP_LOOP_C_133 : begin
        fsm_output = 11'b00100101011;
        state_var_NS = COMP_LOOP_C_134;
      end
      COMP_LOOP_C_134 : begin
        fsm_output = 11'b00100101100;
        state_var_NS = COMP_LOOP_C_135;
      end
      COMP_LOOP_C_135 : begin
        fsm_output = 11'b00100101101;
        state_var_NS = COMP_LOOP_C_136;
      end
      COMP_LOOP_C_136 : begin
        fsm_output = 11'b00100101110;
        state_var_NS = COMP_LOOP_C_137;
      end
      COMP_LOOP_C_137 : begin
        fsm_output = 11'b00100101111;
        state_var_NS = COMP_LOOP_C_138;
      end
      COMP_LOOP_C_138 : begin
        fsm_output = 11'b00100110000;
        state_var_NS = COMP_LOOP_C_139;
      end
      COMP_LOOP_C_139 : begin
        fsm_output = 11'b00100110001;
        state_var_NS = COMP_LOOP_C_140;
      end
      COMP_LOOP_C_140 : begin
        fsm_output = 11'b00100110010;
        state_var_NS = COMP_LOOP_C_141;
      end
      COMP_LOOP_C_141 : begin
        fsm_output = 11'b00100110011;
        state_var_NS = COMP_LOOP_C_142;
      end
      COMP_LOOP_C_142 : begin
        fsm_output = 11'b00100110100;
        state_var_NS = COMP_LOOP_C_143;
      end
      COMP_LOOP_C_143 : begin
        fsm_output = 11'b00100110101;
        state_var_NS = COMP_LOOP_C_144;
      end
      COMP_LOOP_C_144 : begin
        fsm_output = 11'b00100110110;
        state_var_NS = COMP_LOOP_C_145;
      end
      COMP_LOOP_C_145 : begin
        fsm_output = 11'b00100110111;
        state_var_NS = COMP_LOOP_C_146;
      end
      COMP_LOOP_C_146 : begin
        fsm_output = 11'b00100111000;
        state_var_NS = COMP_LOOP_C_147;
      end
      COMP_LOOP_C_147 : begin
        fsm_output = 11'b00100111001;
        state_var_NS = COMP_LOOP_C_148;
      end
      COMP_LOOP_C_148 : begin
        fsm_output = 11'b00100111010;
        state_var_NS = COMP_LOOP_C_149;
      end
      COMP_LOOP_C_149 : begin
        fsm_output = 11'b00100111011;
        state_var_NS = COMP_LOOP_C_150;
      end
      COMP_LOOP_C_150 : begin
        fsm_output = 11'b00100111100;
        state_var_NS = COMP_LOOP_C_151;
      end
      COMP_LOOP_C_151 : begin
        fsm_output = 11'b00100111101;
        state_var_NS = COMP_LOOP_C_152;
      end
      COMP_LOOP_C_152 : begin
        fsm_output = 11'b00100111110;
        state_var_NS = COMP_LOOP_C_153;
      end
      COMP_LOOP_C_153 : begin
        fsm_output = 11'b00100111111;
        state_var_NS = COMP_LOOP_C_154;
      end
      COMP_LOOP_C_154 : begin
        fsm_output = 11'b00101000000;
        state_var_NS = COMP_LOOP_C_155;
      end
      COMP_LOOP_C_155 : begin
        fsm_output = 11'b00101000001;
        state_var_NS = COMP_LOOP_C_156;
      end
      COMP_LOOP_C_156 : begin
        fsm_output = 11'b00101000010;
        state_var_NS = COMP_LOOP_C_157;
      end
      COMP_LOOP_C_157 : begin
        fsm_output = 11'b00101000011;
        state_var_NS = COMP_LOOP_C_158;
      end
      COMP_LOOP_C_158 : begin
        fsm_output = 11'b00101000100;
        state_var_NS = COMP_LOOP_C_159;
      end
      COMP_LOOP_C_159 : begin
        fsm_output = 11'b00101000101;
        state_var_NS = COMP_LOOP_C_160;
      end
      COMP_LOOP_C_160 : begin
        fsm_output = 11'b00101000110;
        state_var_NS = COMP_LOOP_C_161;
      end
      COMP_LOOP_C_161 : begin
        fsm_output = 11'b00101000111;
        state_var_NS = COMP_LOOP_C_162;
      end
      COMP_LOOP_C_162 : begin
        fsm_output = 11'b00101001000;
        state_var_NS = COMP_LOOP_C_163;
      end
      COMP_LOOP_C_163 : begin
        fsm_output = 11'b00101001001;
        state_var_NS = COMP_LOOP_C_164;
      end
      COMP_LOOP_C_164 : begin
        fsm_output = 11'b00101001010;
        state_var_NS = COMP_LOOP_C_165;
      end
      COMP_LOOP_C_165 : begin
        fsm_output = 11'b00101001011;
        state_var_NS = COMP_LOOP_C_166;
      end
      COMP_LOOP_C_166 : begin
        fsm_output = 11'b00101001100;
        state_var_NS = COMP_LOOP_C_167;
      end
      COMP_LOOP_C_167 : begin
        fsm_output = 11'b00101001101;
        state_var_NS = COMP_LOOP_C_168;
      end
      COMP_LOOP_C_168 : begin
        fsm_output = 11'b00101001110;
        state_var_NS = COMP_LOOP_C_169;
      end
      COMP_LOOP_C_169 : begin
        fsm_output = 11'b00101001111;
        state_var_NS = COMP_LOOP_C_170;
      end
      COMP_LOOP_C_170 : begin
        fsm_output = 11'b00101010000;
        state_var_NS = COMP_LOOP_C_171;
      end
      COMP_LOOP_C_171 : begin
        fsm_output = 11'b00101010001;
        state_var_NS = COMP_LOOP_C_172;
      end
      COMP_LOOP_C_172 : begin
        fsm_output = 11'b00101010010;
        state_var_NS = COMP_LOOP_C_173;
      end
      COMP_LOOP_C_173 : begin
        fsm_output = 11'b00101010011;
        state_var_NS = COMP_LOOP_C_174;
      end
      COMP_LOOP_C_174 : begin
        fsm_output = 11'b00101010100;
        state_var_NS = COMP_LOOP_C_175;
      end
      COMP_LOOP_C_175 : begin
        fsm_output = 11'b00101010101;
        state_var_NS = COMP_LOOP_C_176;
      end
      COMP_LOOP_C_176 : begin
        fsm_output = 11'b00101010110;
        state_var_NS = COMP_LOOP_C_177;
      end
      COMP_LOOP_C_177 : begin
        fsm_output = 11'b00101010111;
        state_var_NS = COMP_LOOP_C_178;
      end
      COMP_LOOP_C_178 : begin
        fsm_output = 11'b00101011000;
        state_var_NS = COMP_LOOP_C_179;
      end
      COMP_LOOP_C_179 : begin
        fsm_output = 11'b00101011001;
        state_var_NS = COMP_LOOP_C_180;
      end
      COMP_LOOP_C_180 : begin
        fsm_output = 11'b00101011010;
        state_var_NS = COMP_LOOP_C_181;
      end
      COMP_LOOP_C_181 : begin
        fsm_output = 11'b00101011011;
        state_var_NS = COMP_LOOP_C_182;
      end
      COMP_LOOP_C_182 : begin
        fsm_output = 11'b00101011100;
        state_var_NS = COMP_LOOP_C_183;
      end
      COMP_LOOP_C_183 : begin
        fsm_output = 11'b00101011101;
        state_var_NS = COMP_LOOP_C_184;
      end
      COMP_LOOP_C_184 : begin
        fsm_output = 11'b00101011110;
        state_var_NS = COMP_LOOP_C_185;
      end
      COMP_LOOP_C_185 : begin
        fsm_output = 11'b00101011111;
        state_var_NS = COMP_LOOP_C_186;
      end
      COMP_LOOP_C_186 : begin
        fsm_output = 11'b00101100000;
        state_var_NS = COMP_LOOP_C_187;
      end
      COMP_LOOP_C_187 : begin
        fsm_output = 11'b00101100001;
        state_var_NS = COMP_LOOP_C_188;
      end
      COMP_LOOP_C_188 : begin
        fsm_output = 11'b00101100010;
        state_var_NS = COMP_LOOP_C_189;
      end
      COMP_LOOP_C_189 : begin
        fsm_output = 11'b00101100011;
        state_var_NS = COMP_LOOP_C_190;
      end
      COMP_LOOP_C_190 : begin
        fsm_output = 11'b00101100100;
        state_var_NS = COMP_LOOP_C_191;
      end
      COMP_LOOP_C_191 : begin
        fsm_output = 11'b00101100101;
        state_var_NS = COMP_LOOP_C_192;
      end
      COMP_LOOP_C_192 : begin
        fsm_output = 11'b00101100110;
        if ( COMP_LOOP_C_192_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_193;
        end
      end
      COMP_LOOP_C_193 : begin
        fsm_output = 11'b00101100111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
      end
      COMP_LOOP_4_modExp_1_while_C_0 : begin
        fsm_output = 11'b00101101000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_1;
      end
      COMP_LOOP_4_modExp_1_while_C_1 : begin
        fsm_output = 11'b00101101001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_2;
      end
      COMP_LOOP_4_modExp_1_while_C_2 : begin
        fsm_output = 11'b00101101010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_3;
      end
      COMP_LOOP_4_modExp_1_while_C_3 : begin
        fsm_output = 11'b00101101011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_4;
      end
      COMP_LOOP_4_modExp_1_while_C_4 : begin
        fsm_output = 11'b00101101100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_5;
      end
      COMP_LOOP_4_modExp_1_while_C_5 : begin
        fsm_output = 11'b00101101101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_6;
      end
      COMP_LOOP_4_modExp_1_while_C_6 : begin
        fsm_output = 11'b00101101110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_7;
      end
      COMP_LOOP_4_modExp_1_while_C_7 : begin
        fsm_output = 11'b00101101111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_8;
      end
      COMP_LOOP_4_modExp_1_while_C_8 : begin
        fsm_output = 11'b00101110000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_9;
      end
      COMP_LOOP_4_modExp_1_while_C_9 : begin
        fsm_output = 11'b00101110001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_10;
      end
      COMP_LOOP_4_modExp_1_while_C_10 : begin
        fsm_output = 11'b00101110010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_11;
      end
      COMP_LOOP_4_modExp_1_while_C_11 : begin
        fsm_output = 11'b00101110011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_12;
      end
      COMP_LOOP_4_modExp_1_while_C_12 : begin
        fsm_output = 11'b00101110100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_13;
      end
      COMP_LOOP_4_modExp_1_while_C_13 : begin
        fsm_output = 11'b00101110101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_14;
      end
      COMP_LOOP_4_modExp_1_while_C_14 : begin
        fsm_output = 11'b00101110110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_15;
      end
      COMP_LOOP_4_modExp_1_while_C_15 : begin
        fsm_output = 11'b00101110111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_16;
      end
      COMP_LOOP_4_modExp_1_while_C_16 : begin
        fsm_output = 11'b00101111000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_17;
      end
      COMP_LOOP_4_modExp_1_while_C_17 : begin
        fsm_output = 11'b00101111001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_18;
      end
      COMP_LOOP_4_modExp_1_while_C_18 : begin
        fsm_output = 11'b00101111010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_19;
      end
      COMP_LOOP_4_modExp_1_while_C_19 : begin
        fsm_output = 11'b00101111011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_20;
      end
      COMP_LOOP_4_modExp_1_while_C_20 : begin
        fsm_output = 11'b00101111100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_21;
      end
      COMP_LOOP_4_modExp_1_while_C_21 : begin
        fsm_output = 11'b00101111101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_22;
      end
      COMP_LOOP_4_modExp_1_while_C_22 : begin
        fsm_output = 11'b00101111110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_23;
      end
      COMP_LOOP_4_modExp_1_while_C_23 : begin
        fsm_output = 11'b00101111111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_24;
      end
      COMP_LOOP_4_modExp_1_while_C_24 : begin
        fsm_output = 11'b00110000000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_25;
      end
      COMP_LOOP_4_modExp_1_while_C_25 : begin
        fsm_output = 11'b00110000001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_26;
      end
      COMP_LOOP_4_modExp_1_while_C_26 : begin
        fsm_output = 11'b00110000010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_27;
      end
      COMP_LOOP_4_modExp_1_while_C_27 : begin
        fsm_output = 11'b00110000011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_28;
      end
      COMP_LOOP_4_modExp_1_while_C_28 : begin
        fsm_output = 11'b00110000100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_29;
      end
      COMP_LOOP_4_modExp_1_while_C_29 : begin
        fsm_output = 11'b00110000101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_30;
      end
      COMP_LOOP_4_modExp_1_while_C_30 : begin
        fsm_output = 11'b00110000110;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_31;
      end
      COMP_LOOP_4_modExp_1_while_C_31 : begin
        fsm_output = 11'b00110000111;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_32;
      end
      COMP_LOOP_4_modExp_1_while_C_32 : begin
        fsm_output = 11'b00110001000;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_33;
      end
      COMP_LOOP_4_modExp_1_while_C_33 : begin
        fsm_output = 11'b00110001001;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_34;
      end
      COMP_LOOP_4_modExp_1_while_C_34 : begin
        fsm_output = 11'b00110001010;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_35;
      end
      COMP_LOOP_4_modExp_1_while_C_35 : begin
        fsm_output = 11'b00110001011;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_36;
      end
      COMP_LOOP_4_modExp_1_while_C_36 : begin
        fsm_output = 11'b00110001100;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_37;
      end
      COMP_LOOP_4_modExp_1_while_C_37 : begin
        fsm_output = 11'b00110001101;
        state_var_NS = COMP_LOOP_4_modExp_1_while_C_38;
      end
      COMP_LOOP_4_modExp_1_while_C_38 : begin
        fsm_output = 11'b00110001110;
        if ( COMP_LOOP_4_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_194;
        end
        else begin
          state_var_NS = COMP_LOOP_4_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_194 : begin
        fsm_output = 11'b00110001111;
        state_var_NS = COMP_LOOP_C_195;
      end
      COMP_LOOP_C_195 : begin
        fsm_output = 11'b00110010000;
        state_var_NS = COMP_LOOP_C_196;
      end
      COMP_LOOP_C_196 : begin
        fsm_output = 11'b00110010001;
        state_var_NS = COMP_LOOP_C_197;
      end
      COMP_LOOP_C_197 : begin
        fsm_output = 11'b00110010010;
        state_var_NS = COMP_LOOP_C_198;
      end
      COMP_LOOP_C_198 : begin
        fsm_output = 11'b00110010011;
        state_var_NS = COMP_LOOP_C_199;
      end
      COMP_LOOP_C_199 : begin
        fsm_output = 11'b00110010100;
        state_var_NS = COMP_LOOP_C_200;
      end
      COMP_LOOP_C_200 : begin
        fsm_output = 11'b00110010101;
        state_var_NS = COMP_LOOP_C_201;
      end
      COMP_LOOP_C_201 : begin
        fsm_output = 11'b00110010110;
        state_var_NS = COMP_LOOP_C_202;
      end
      COMP_LOOP_C_202 : begin
        fsm_output = 11'b00110010111;
        state_var_NS = COMP_LOOP_C_203;
      end
      COMP_LOOP_C_203 : begin
        fsm_output = 11'b00110011000;
        state_var_NS = COMP_LOOP_C_204;
      end
      COMP_LOOP_C_204 : begin
        fsm_output = 11'b00110011001;
        state_var_NS = COMP_LOOP_C_205;
      end
      COMP_LOOP_C_205 : begin
        fsm_output = 11'b00110011010;
        state_var_NS = COMP_LOOP_C_206;
      end
      COMP_LOOP_C_206 : begin
        fsm_output = 11'b00110011011;
        state_var_NS = COMP_LOOP_C_207;
      end
      COMP_LOOP_C_207 : begin
        fsm_output = 11'b00110011100;
        state_var_NS = COMP_LOOP_C_208;
      end
      COMP_LOOP_C_208 : begin
        fsm_output = 11'b00110011101;
        state_var_NS = COMP_LOOP_C_209;
      end
      COMP_LOOP_C_209 : begin
        fsm_output = 11'b00110011110;
        state_var_NS = COMP_LOOP_C_210;
      end
      COMP_LOOP_C_210 : begin
        fsm_output = 11'b00110011111;
        state_var_NS = COMP_LOOP_C_211;
      end
      COMP_LOOP_C_211 : begin
        fsm_output = 11'b00110100000;
        state_var_NS = COMP_LOOP_C_212;
      end
      COMP_LOOP_C_212 : begin
        fsm_output = 11'b00110100001;
        state_var_NS = COMP_LOOP_C_213;
      end
      COMP_LOOP_C_213 : begin
        fsm_output = 11'b00110100010;
        state_var_NS = COMP_LOOP_C_214;
      end
      COMP_LOOP_C_214 : begin
        fsm_output = 11'b00110100011;
        state_var_NS = COMP_LOOP_C_215;
      end
      COMP_LOOP_C_215 : begin
        fsm_output = 11'b00110100100;
        state_var_NS = COMP_LOOP_C_216;
      end
      COMP_LOOP_C_216 : begin
        fsm_output = 11'b00110100101;
        state_var_NS = COMP_LOOP_C_217;
      end
      COMP_LOOP_C_217 : begin
        fsm_output = 11'b00110100110;
        state_var_NS = COMP_LOOP_C_218;
      end
      COMP_LOOP_C_218 : begin
        fsm_output = 11'b00110100111;
        state_var_NS = COMP_LOOP_C_219;
      end
      COMP_LOOP_C_219 : begin
        fsm_output = 11'b00110101000;
        state_var_NS = COMP_LOOP_C_220;
      end
      COMP_LOOP_C_220 : begin
        fsm_output = 11'b00110101001;
        state_var_NS = COMP_LOOP_C_221;
      end
      COMP_LOOP_C_221 : begin
        fsm_output = 11'b00110101010;
        state_var_NS = COMP_LOOP_C_222;
      end
      COMP_LOOP_C_222 : begin
        fsm_output = 11'b00110101011;
        state_var_NS = COMP_LOOP_C_223;
      end
      COMP_LOOP_C_223 : begin
        fsm_output = 11'b00110101100;
        state_var_NS = COMP_LOOP_C_224;
      end
      COMP_LOOP_C_224 : begin
        fsm_output = 11'b00110101101;
        state_var_NS = COMP_LOOP_C_225;
      end
      COMP_LOOP_C_225 : begin
        fsm_output = 11'b00110101110;
        state_var_NS = COMP_LOOP_C_226;
      end
      COMP_LOOP_C_226 : begin
        fsm_output = 11'b00110101111;
        state_var_NS = COMP_LOOP_C_227;
      end
      COMP_LOOP_C_227 : begin
        fsm_output = 11'b00110110000;
        state_var_NS = COMP_LOOP_C_228;
      end
      COMP_LOOP_C_228 : begin
        fsm_output = 11'b00110110001;
        state_var_NS = COMP_LOOP_C_229;
      end
      COMP_LOOP_C_229 : begin
        fsm_output = 11'b00110110010;
        state_var_NS = COMP_LOOP_C_230;
      end
      COMP_LOOP_C_230 : begin
        fsm_output = 11'b00110110011;
        state_var_NS = COMP_LOOP_C_231;
      end
      COMP_LOOP_C_231 : begin
        fsm_output = 11'b00110110100;
        state_var_NS = COMP_LOOP_C_232;
      end
      COMP_LOOP_C_232 : begin
        fsm_output = 11'b00110110101;
        state_var_NS = COMP_LOOP_C_233;
      end
      COMP_LOOP_C_233 : begin
        fsm_output = 11'b00110110110;
        state_var_NS = COMP_LOOP_C_234;
      end
      COMP_LOOP_C_234 : begin
        fsm_output = 11'b00110110111;
        state_var_NS = COMP_LOOP_C_235;
      end
      COMP_LOOP_C_235 : begin
        fsm_output = 11'b00110111000;
        state_var_NS = COMP_LOOP_C_236;
      end
      COMP_LOOP_C_236 : begin
        fsm_output = 11'b00110111001;
        state_var_NS = COMP_LOOP_C_237;
      end
      COMP_LOOP_C_237 : begin
        fsm_output = 11'b00110111010;
        state_var_NS = COMP_LOOP_C_238;
      end
      COMP_LOOP_C_238 : begin
        fsm_output = 11'b00110111011;
        state_var_NS = COMP_LOOP_C_239;
      end
      COMP_LOOP_C_239 : begin
        fsm_output = 11'b00110111100;
        state_var_NS = COMP_LOOP_C_240;
      end
      COMP_LOOP_C_240 : begin
        fsm_output = 11'b00110111101;
        state_var_NS = COMP_LOOP_C_241;
      end
      COMP_LOOP_C_241 : begin
        fsm_output = 11'b00110111110;
        state_var_NS = COMP_LOOP_C_242;
      end
      COMP_LOOP_C_242 : begin
        fsm_output = 11'b00110111111;
        state_var_NS = COMP_LOOP_C_243;
      end
      COMP_LOOP_C_243 : begin
        fsm_output = 11'b00111000000;
        state_var_NS = COMP_LOOP_C_244;
      end
      COMP_LOOP_C_244 : begin
        fsm_output = 11'b00111000001;
        state_var_NS = COMP_LOOP_C_245;
      end
      COMP_LOOP_C_245 : begin
        fsm_output = 11'b00111000010;
        state_var_NS = COMP_LOOP_C_246;
      end
      COMP_LOOP_C_246 : begin
        fsm_output = 11'b00111000011;
        state_var_NS = COMP_LOOP_C_247;
      end
      COMP_LOOP_C_247 : begin
        fsm_output = 11'b00111000100;
        state_var_NS = COMP_LOOP_C_248;
      end
      COMP_LOOP_C_248 : begin
        fsm_output = 11'b00111000101;
        state_var_NS = COMP_LOOP_C_249;
      end
      COMP_LOOP_C_249 : begin
        fsm_output = 11'b00111000110;
        state_var_NS = COMP_LOOP_C_250;
      end
      COMP_LOOP_C_250 : begin
        fsm_output = 11'b00111000111;
        state_var_NS = COMP_LOOP_C_251;
      end
      COMP_LOOP_C_251 : begin
        fsm_output = 11'b00111001000;
        state_var_NS = COMP_LOOP_C_252;
      end
      COMP_LOOP_C_252 : begin
        fsm_output = 11'b00111001001;
        state_var_NS = COMP_LOOP_C_253;
      end
      COMP_LOOP_C_253 : begin
        fsm_output = 11'b00111001010;
        state_var_NS = COMP_LOOP_C_254;
      end
      COMP_LOOP_C_254 : begin
        fsm_output = 11'b00111001011;
        state_var_NS = COMP_LOOP_C_255;
      end
      COMP_LOOP_C_255 : begin
        fsm_output = 11'b00111001100;
        state_var_NS = COMP_LOOP_C_256;
      end
      COMP_LOOP_C_256 : begin
        fsm_output = 11'b00111001101;
        if ( COMP_LOOP_C_256_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_257;
        end
      end
      COMP_LOOP_C_257 : begin
        fsm_output = 11'b00111001110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
      end
      COMP_LOOP_5_modExp_1_while_C_0 : begin
        fsm_output = 11'b00111001111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_1;
      end
      COMP_LOOP_5_modExp_1_while_C_1 : begin
        fsm_output = 11'b00111010000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_2;
      end
      COMP_LOOP_5_modExp_1_while_C_2 : begin
        fsm_output = 11'b00111010001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_3;
      end
      COMP_LOOP_5_modExp_1_while_C_3 : begin
        fsm_output = 11'b00111010010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_4;
      end
      COMP_LOOP_5_modExp_1_while_C_4 : begin
        fsm_output = 11'b00111010011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_5;
      end
      COMP_LOOP_5_modExp_1_while_C_5 : begin
        fsm_output = 11'b00111010100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_6;
      end
      COMP_LOOP_5_modExp_1_while_C_6 : begin
        fsm_output = 11'b00111010101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_7;
      end
      COMP_LOOP_5_modExp_1_while_C_7 : begin
        fsm_output = 11'b00111010110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_8;
      end
      COMP_LOOP_5_modExp_1_while_C_8 : begin
        fsm_output = 11'b00111010111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_9;
      end
      COMP_LOOP_5_modExp_1_while_C_9 : begin
        fsm_output = 11'b00111011000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_10;
      end
      COMP_LOOP_5_modExp_1_while_C_10 : begin
        fsm_output = 11'b00111011001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_11;
      end
      COMP_LOOP_5_modExp_1_while_C_11 : begin
        fsm_output = 11'b00111011010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_12;
      end
      COMP_LOOP_5_modExp_1_while_C_12 : begin
        fsm_output = 11'b00111011011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_13;
      end
      COMP_LOOP_5_modExp_1_while_C_13 : begin
        fsm_output = 11'b00111011100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_14;
      end
      COMP_LOOP_5_modExp_1_while_C_14 : begin
        fsm_output = 11'b00111011101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_15;
      end
      COMP_LOOP_5_modExp_1_while_C_15 : begin
        fsm_output = 11'b00111011110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_16;
      end
      COMP_LOOP_5_modExp_1_while_C_16 : begin
        fsm_output = 11'b00111011111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_17;
      end
      COMP_LOOP_5_modExp_1_while_C_17 : begin
        fsm_output = 11'b00111100000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_18;
      end
      COMP_LOOP_5_modExp_1_while_C_18 : begin
        fsm_output = 11'b00111100001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_19;
      end
      COMP_LOOP_5_modExp_1_while_C_19 : begin
        fsm_output = 11'b00111100010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_20;
      end
      COMP_LOOP_5_modExp_1_while_C_20 : begin
        fsm_output = 11'b00111100011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_21;
      end
      COMP_LOOP_5_modExp_1_while_C_21 : begin
        fsm_output = 11'b00111100100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_22;
      end
      COMP_LOOP_5_modExp_1_while_C_22 : begin
        fsm_output = 11'b00111100101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_23;
      end
      COMP_LOOP_5_modExp_1_while_C_23 : begin
        fsm_output = 11'b00111100110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_24;
      end
      COMP_LOOP_5_modExp_1_while_C_24 : begin
        fsm_output = 11'b00111100111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_25;
      end
      COMP_LOOP_5_modExp_1_while_C_25 : begin
        fsm_output = 11'b00111101000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_26;
      end
      COMP_LOOP_5_modExp_1_while_C_26 : begin
        fsm_output = 11'b00111101001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_27;
      end
      COMP_LOOP_5_modExp_1_while_C_27 : begin
        fsm_output = 11'b00111101010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_28;
      end
      COMP_LOOP_5_modExp_1_while_C_28 : begin
        fsm_output = 11'b00111101011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_29;
      end
      COMP_LOOP_5_modExp_1_while_C_29 : begin
        fsm_output = 11'b00111101100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_30;
      end
      COMP_LOOP_5_modExp_1_while_C_30 : begin
        fsm_output = 11'b00111101101;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_31;
      end
      COMP_LOOP_5_modExp_1_while_C_31 : begin
        fsm_output = 11'b00111101110;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_32;
      end
      COMP_LOOP_5_modExp_1_while_C_32 : begin
        fsm_output = 11'b00111101111;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_33;
      end
      COMP_LOOP_5_modExp_1_while_C_33 : begin
        fsm_output = 11'b00111110000;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_34;
      end
      COMP_LOOP_5_modExp_1_while_C_34 : begin
        fsm_output = 11'b00111110001;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_35;
      end
      COMP_LOOP_5_modExp_1_while_C_35 : begin
        fsm_output = 11'b00111110010;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_36;
      end
      COMP_LOOP_5_modExp_1_while_C_36 : begin
        fsm_output = 11'b00111110011;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_37;
      end
      COMP_LOOP_5_modExp_1_while_C_37 : begin
        fsm_output = 11'b00111110100;
        state_var_NS = COMP_LOOP_5_modExp_1_while_C_38;
      end
      COMP_LOOP_5_modExp_1_while_C_38 : begin
        fsm_output = 11'b00111110101;
        if ( COMP_LOOP_5_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_258;
        end
        else begin
          state_var_NS = COMP_LOOP_5_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_258 : begin
        fsm_output = 11'b00111110110;
        state_var_NS = COMP_LOOP_C_259;
      end
      COMP_LOOP_C_259 : begin
        fsm_output = 11'b00111110111;
        state_var_NS = COMP_LOOP_C_260;
      end
      COMP_LOOP_C_260 : begin
        fsm_output = 11'b00111111000;
        state_var_NS = COMP_LOOP_C_261;
      end
      COMP_LOOP_C_261 : begin
        fsm_output = 11'b00111111001;
        state_var_NS = COMP_LOOP_C_262;
      end
      COMP_LOOP_C_262 : begin
        fsm_output = 11'b00111111010;
        state_var_NS = COMP_LOOP_C_263;
      end
      COMP_LOOP_C_263 : begin
        fsm_output = 11'b00111111011;
        state_var_NS = COMP_LOOP_C_264;
      end
      COMP_LOOP_C_264 : begin
        fsm_output = 11'b00111111100;
        state_var_NS = COMP_LOOP_C_265;
      end
      COMP_LOOP_C_265 : begin
        fsm_output = 11'b00111111101;
        state_var_NS = COMP_LOOP_C_266;
      end
      COMP_LOOP_C_266 : begin
        fsm_output = 11'b00111111110;
        state_var_NS = COMP_LOOP_C_267;
      end
      COMP_LOOP_C_267 : begin
        fsm_output = 11'b00111111111;
        state_var_NS = COMP_LOOP_C_268;
      end
      COMP_LOOP_C_268 : begin
        fsm_output = 11'b01000000000;
        state_var_NS = COMP_LOOP_C_269;
      end
      COMP_LOOP_C_269 : begin
        fsm_output = 11'b01000000001;
        state_var_NS = COMP_LOOP_C_270;
      end
      COMP_LOOP_C_270 : begin
        fsm_output = 11'b01000000010;
        state_var_NS = COMP_LOOP_C_271;
      end
      COMP_LOOP_C_271 : begin
        fsm_output = 11'b01000000011;
        state_var_NS = COMP_LOOP_C_272;
      end
      COMP_LOOP_C_272 : begin
        fsm_output = 11'b01000000100;
        state_var_NS = COMP_LOOP_C_273;
      end
      COMP_LOOP_C_273 : begin
        fsm_output = 11'b01000000101;
        state_var_NS = COMP_LOOP_C_274;
      end
      COMP_LOOP_C_274 : begin
        fsm_output = 11'b01000000110;
        state_var_NS = COMP_LOOP_C_275;
      end
      COMP_LOOP_C_275 : begin
        fsm_output = 11'b01000000111;
        state_var_NS = COMP_LOOP_C_276;
      end
      COMP_LOOP_C_276 : begin
        fsm_output = 11'b01000001000;
        state_var_NS = COMP_LOOP_C_277;
      end
      COMP_LOOP_C_277 : begin
        fsm_output = 11'b01000001001;
        state_var_NS = COMP_LOOP_C_278;
      end
      COMP_LOOP_C_278 : begin
        fsm_output = 11'b01000001010;
        state_var_NS = COMP_LOOP_C_279;
      end
      COMP_LOOP_C_279 : begin
        fsm_output = 11'b01000001011;
        state_var_NS = COMP_LOOP_C_280;
      end
      COMP_LOOP_C_280 : begin
        fsm_output = 11'b01000001100;
        state_var_NS = COMP_LOOP_C_281;
      end
      COMP_LOOP_C_281 : begin
        fsm_output = 11'b01000001101;
        state_var_NS = COMP_LOOP_C_282;
      end
      COMP_LOOP_C_282 : begin
        fsm_output = 11'b01000001110;
        state_var_NS = COMP_LOOP_C_283;
      end
      COMP_LOOP_C_283 : begin
        fsm_output = 11'b01000001111;
        state_var_NS = COMP_LOOP_C_284;
      end
      COMP_LOOP_C_284 : begin
        fsm_output = 11'b01000010000;
        state_var_NS = COMP_LOOP_C_285;
      end
      COMP_LOOP_C_285 : begin
        fsm_output = 11'b01000010001;
        state_var_NS = COMP_LOOP_C_286;
      end
      COMP_LOOP_C_286 : begin
        fsm_output = 11'b01000010010;
        state_var_NS = COMP_LOOP_C_287;
      end
      COMP_LOOP_C_287 : begin
        fsm_output = 11'b01000010011;
        state_var_NS = COMP_LOOP_C_288;
      end
      COMP_LOOP_C_288 : begin
        fsm_output = 11'b01000010100;
        state_var_NS = COMP_LOOP_C_289;
      end
      COMP_LOOP_C_289 : begin
        fsm_output = 11'b01000010101;
        state_var_NS = COMP_LOOP_C_290;
      end
      COMP_LOOP_C_290 : begin
        fsm_output = 11'b01000010110;
        state_var_NS = COMP_LOOP_C_291;
      end
      COMP_LOOP_C_291 : begin
        fsm_output = 11'b01000010111;
        state_var_NS = COMP_LOOP_C_292;
      end
      COMP_LOOP_C_292 : begin
        fsm_output = 11'b01000011000;
        state_var_NS = COMP_LOOP_C_293;
      end
      COMP_LOOP_C_293 : begin
        fsm_output = 11'b01000011001;
        state_var_NS = COMP_LOOP_C_294;
      end
      COMP_LOOP_C_294 : begin
        fsm_output = 11'b01000011010;
        state_var_NS = COMP_LOOP_C_295;
      end
      COMP_LOOP_C_295 : begin
        fsm_output = 11'b01000011011;
        state_var_NS = COMP_LOOP_C_296;
      end
      COMP_LOOP_C_296 : begin
        fsm_output = 11'b01000011100;
        state_var_NS = COMP_LOOP_C_297;
      end
      COMP_LOOP_C_297 : begin
        fsm_output = 11'b01000011101;
        state_var_NS = COMP_LOOP_C_298;
      end
      COMP_LOOP_C_298 : begin
        fsm_output = 11'b01000011110;
        state_var_NS = COMP_LOOP_C_299;
      end
      COMP_LOOP_C_299 : begin
        fsm_output = 11'b01000011111;
        state_var_NS = COMP_LOOP_C_300;
      end
      COMP_LOOP_C_300 : begin
        fsm_output = 11'b01000100000;
        state_var_NS = COMP_LOOP_C_301;
      end
      COMP_LOOP_C_301 : begin
        fsm_output = 11'b01000100001;
        state_var_NS = COMP_LOOP_C_302;
      end
      COMP_LOOP_C_302 : begin
        fsm_output = 11'b01000100010;
        state_var_NS = COMP_LOOP_C_303;
      end
      COMP_LOOP_C_303 : begin
        fsm_output = 11'b01000100011;
        state_var_NS = COMP_LOOP_C_304;
      end
      COMP_LOOP_C_304 : begin
        fsm_output = 11'b01000100100;
        state_var_NS = COMP_LOOP_C_305;
      end
      COMP_LOOP_C_305 : begin
        fsm_output = 11'b01000100101;
        state_var_NS = COMP_LOOP_C_306;
      end
      COMP_LOOP_C_306 : begin
        fsm_output = 11'b01000100110;
        state_var_NS = COMP_LOOP_C_307;
      end
      COMP_LOOP_C_307 : begin
        fsm_output = 11'b01000100111;
        state_var_NS = COMP_LOOP_C_308;
      end
      COMP_LOOP_C_308 : begin
        fsm_output = 11'b01000101000;
        state_var_NS = COMP_LOOP_C_309;
      end
      COMP_LOOP_C_309 : begin
        fsm_output = 11'b01000101001;
        state_var_NS = COMP_LOOP_C_310;
      end
      COMP_LOOP_C_310 : begin
        fsm_output = 11'b01000101010;
        state_var_NS = COMP_LOOP_C_311;
      end
      COMP_LOOP_C_311 : begin
        fsm_output = 11'b01000101011;
        state_var_NS = COMP_LOOP_C_312;
      end
      COMP_LOOP_C_312 : begin
        fsm_output = 11'b01000101100;
        state_var_NS = COMP_LOOP_C_313;
      end
      COMP_LOOP_C_313 : begin
        fsm_output = 11'b01000101101;
        state_var_NS = COMP_LOOP_C_314;
      end
      COMP_LOOP_C_314 : begin
        fsm_output = 11'b01000101110;
        state_var_NS = COMP_LOOP_C_315;
      end
      COMP_LOOP_C_315 : begin
        fsm_output = 11'b01000101111;
        state_var_NS = COMP_LOOP_C_316;
      end
      COMP_LOOP_C_316 : begin
        fsm_output = 11'b01000110000;
        state_var_NS = COMP_LOOP_C_317;
      end
      COMP_LOOP_C_317 : begin
        fsm_output = 11'b01000110001;
        state_var_NS = COMP_LOOP_C_318;
      end
      COMP_LOOP_C_318 : begin
        fsm_output = 11'b01000110010;
        state_var_NS = COMP_LOOP_C_319;
      end
      COMP_LOOP_C_319 : begin
        fsm_output = 11'b01000110011;
        state_var_NS = COMP_LOOP_C_320;
      end
      COMP_LOOP_C_320 : begin
        fsm_output = 11'b01000110100;
        if ( COMP_LOOP_C_320_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_321;
        end
      end
      COMP_LOOP_C_321 : begin
        fsm_output = 11'b01000110101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
      end
      COMP_LOOP_6_modExp_1_while_C_0 : begin
        fsm_output = 11'b01000110110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_1;
      end
      COMP_LOOP_6_modExp_1_while_C_1 : begin
        fsm_output = 11'b01000110111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_2;
      end
      COMP_LOOP_6_modExp_1_while_C_2 : begin
        fsm_output = 11'b01000111000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_3;
      end
      COMP_LOOP_6_modExp_1_while_C_3 : begin
        fsm_output = 11'b01000111001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_4;
      end
      COMP_LOOP_6_modExp_1_while_C_4 : begin
        fsm_output = 11'b01000111010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_5;
      end
      COMP_LOOP_6_modExp_1_while_C_5 : begin
        fsm_output = 11'b01000111011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_6;
      end
      COMP_LOOP_6_modExp_1_while_C_6 : begin
        fsm_output = 11'b01000111100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_7;
      end
      COMP_LOOP_6_modExp_1_while_C_7 : begin
        fsm_output = 11'b01000111101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_8;
      end
      COMP_LOOP_6_modExp_1_while_C_8 : begin
        fsm_output = 11'b01000111110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_9;
      end
      COMP_LOOP_6_modExp_1_while_C_9 : begin
        fsm_output = 11'b01000111111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_10;
      end
      COMP_LOOP_6_modExp_1_while_C_10 : begin
        fsm_output = 11'b01001000000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_11;
      end
      COMP_LOOP_6_modExp_1_while_C_11 : begin
        fsm_output = 11'b01001000001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_12;
      end
      COMP_LOOP_6_modExp_1_while_C_12 : begin
        fsm_output = 11'b01001000010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_13;
      end
      COMP_LOOP_6_modExp_1_while_C_13 : begin
        fsm_output = 11'b01001000011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_14;
      end
      COMP_LOOP_6_modExp_1_while_C_14 : begin
        fsm_output = 11'b01001000100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_15;
      end
      COMP_LOOP_6_modExp_1_while_C_15 : begin
        fsm_output = 11'b01001000101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_16;
      end
      COMP_LOOP_6_modExp_1_while_C_16 : begin
        fsm_output = 11'b01001000110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_17;
      end
      COMP_LOOP_6_modExp_1_while_C_17 : begin
        fsm_output = 11'b01001000111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_18;
      end
      COMP_LOOP_6_modExp_1_while_C_18 : begin
        fsm_output = 11'b01001001000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_19;
      end
      COMP_LOOP_6_modExp_1_while_C_19 : begin
        fsm_output = 11'b01001001001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_20;
      end
      COMP_LOOP_6_modExp_1_while_C_20 : begin
        fsm_output = 11'b01001001010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_21;
      end
      COMP_LOOP_6_modExp_1_while_C_21 : begin
        fsm_output = 11'b01001001011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_22;
      end
      COMP_LOOP_6_modExp_1_while_C_22 : begin
        fsm_output = 11'b01001001100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_23;
      end
      COMP_LOOP_6_modExp_1_while_C_23 : begin
        fsm_output = 11'b01001001101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_24;
      end
      COMP_LOOP_6_modExp_1_while_C_24 : begin
        fsm_output = 11'b01001001110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_25;
      end
      COMP_LOOP_6_modExp_1_while_C_25 : begin
        fsm_output = 11'b01001001111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_26;
      end
      COMP_LOOP_6_modExp_1_while_C_26 : begin
        fsm_output = 11'b01001010000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_27;
      end
      COMP_LOOP_6_modExp_1_while_C_27 : begin
        fsm_output = 11'b01001010001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_28;
      end
      COMP_LOOP_6_modExp_1_while_C_28 : begin
        fsm_output = 11'b01001010010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_29;
      end
      COMP_LOOP_6_modExp_1_while_C_29 : begin
        fsm_output = 11'b01001010011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_30;
      end
      COMP_LOOP_6_modExp_1_while_C_30 : begin
        fsm_output = 11'b01001010100;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_31;
      end
      COMP_LOOP_6_modExp_1_while_C_31 : begin
        fsm_output = 11'b01001010101;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_32;
      end
      COMP_LOOP_6_modExp_1_while_C_32 : begin
        fsm_output = 11'b01001010110;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_33;
      end
      COMP_LOOP_6_modExp_1_while_C_33 : begin
        fsm_output = 11'b01001010111;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_34;
      end
      COMP_LOOP_6_modExp_1_while_C_34 : begin
        fsm_output = 11'b01001011000;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_35;
      end
      COMP_LOOP_6_modExp_1_while_C_35 : begin
        fsm_output = 11'b01001011001;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_36;
      end
      COMP_LOOP_6_modExp_1_while_C_36 : begin
        fsm_output = 11'b01001011010;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_37;
      end
      COMP_LOOP_6_modExp_1_while_C_37 : begin
        fsm_output = 11'b01001011011;
        state_var_NS = COMP_LOOP_6_modExp_1_while_C_38;
      end
      COMP_LOOP_6_modExp_1_while_C_38 : begin
        fsm_output = 11'b01001011100;
        if ( COMP_LOOP_6_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_322;
        end
        else begin
          state_var_NS = COMP_LOOP_6_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_322 : begin
        fsm_output = 11'b01001011101;
        state_var_NS = COMP_LOOP_C_323;
      end
      COMP_LOOP_C_323 : begin
        fsm_output = 11'b01001011110;
        state_var_NS = COMP_LOOP_C_324;
      end
      COMP_LOOP_C_324 : begin
        fsm_output = 11'b01001011111;
        state_var_NS = COMP_LOOP_C_325;
      end
      COMP_LOOP_C_325 : begin
        fsm_output = 11'b01001100000;
        state_var_NS = COMP_LOOP_C_326;
      end
      COMP_LOOP_C_326 : begin
        fsm_output = 11'b01001100001;
        state_var_NS = COMP_LOOP_C_327;
      end
      COMP_LOOP_C_327 : begin
        fsm_output = 11'b01001100010;
        state_var_NS = COMP_LOOP_C_328;
      end
      COMP_LOOP_C_328 : begin
        fsm_output = 11'b01001100011;
        state_var_NS = COMP_LOOP_C_329;
      end
      COMP_LOOP_C_329 : begin
        fsm_output = 11'b01001100100;
        state_var_NS = COMP_LOOP_C_330;
      end
      COMP_LOOP_C_330 : begin
        fsm_output = 11'b01001100101;
        state_var_NS = COMP_LOOP_C_331;
      end
      COMP_LOOP_C_331 : begin
        fsm_output = 11'b01001100110;
        state_var_NS = COMP_LOOP_C_332;
      end
      COMP_LOOP_C_332 : begin
        fsm_output = 11'b01001100111;
        state_var_NS = COMP_LOOP_C_333;
      end
      COMP_LOOP_C_333 : begin
        fsm_output = 11'b01001101000;
        state_var_NS = COMP_LOOP_C_334;
      end
      COMP_LOOP_C_334 : begin
        fsm_output = 11'b01001101001;
        state_var_NS = COMP_LOOP_C_335;
      end
      COMP_LOOP_C_335 : begin
        fsm_output = 11'b01001101010;
        state_var_NS = COMP_LOOP_C_336;
      end
      COMP_LOOP_C_336 : begin
        fsm_output = 11'b01001101011;
        state_var_NS = COMP_LOOP_C_337;
      end
      COMP_LOOP_C_337 : begin
        fsm_output = 11'b01001101100;
        state_var_NS = COMP_LOOP_C_338;
      end
      COMP_LOOP_C_338 : begin
        fsm_output = 11'b01001101101;
        state_var_NS = COMP_LOOP_C_339;
      end
      COMP_LOOP_C_339 : begin
        fsm_output = 11'b01001101110;
        state_var_NS = COMP_LOOP_C_340;
      end
      COMP_LOOP_C_340 : begin
        fsm_output = 11'b01001101111;
        state_var_NS = COMP_LOOP_C_341;
      end
      COMP_LOOP_C_341 : begin
        fsm_output = 11'b01001110000;
        state_var_NS = COMP_LOOP_C_342;
      end
      COMP_LOOP_C_342 : begin
        fsm_output = 11'b01001110001;
        state_var_NS = COMP_LOOP_C_343;
      end
      COMP_LOOP_C_343 : begin
        fsm_output = 11'b01001110010;
        state_var_NS = COMP_LOOP_C_344;
      end
      COMP_LOOP_C_344 : begin
        fsm_output = 11'b01001110011;
        state_var_NS = COMP_LOOP_C_345;
      end
      COMP_LOOP_C_345 : begin
        fsm_output = 11'b01001110100;
        state_var_NS = COMP_LOOP_C_346;
      end
      COMP_LOOP_C_346 : begin
        fsm_output = 11'b01001110101;
        state_var_NS = COMP_LOOP_C_347;
      end
      COMP_LOOP_C_347 : begin
        fsm_output = 11'b01001110110;
        state_var_NS = COMP_LOOP_C_348;
      end
      COMP_LOOP_C_348 : begin
        fsm_output = 11'b01001110111;
        state_var_NS = COMP_LOOP_C_349;
      end
      COMP_LOOP_C_349 : begin
        fsm_output = 11'b01001111000;
        state_var_NS = COMP_LOOP_C_350;
      end
      COMP_LOOP_C_350 : begin
        fsm_output = 11'b01001111001;
        state_var_NS = COMP_LOOP_C_351;
      end
      COMP_LOOP_C_351 : begin
        fsm_output = 11'b01001111010;
        state_var_NS = COMP_LOOP_C_352;
      end
      COMP_LOOP_C_352 : begin
        fsm_output = 11'b01001111011;
        state_var_NS = COMP_LOOP_C_353;
      end
      COMP_LOOP_C_353 : begin
        fsm_output = 11'b01001111100;
        state_var_NS = COMP_LOOP_C_354;
      end
      COMP_LOOP_C_354 : begin
        fsm_output = 11'b01001111101;
        state_var_NS = COMP_LOOP_C_355;
      end
      COMP_LOOP_C_355 : begin
        fsm_output = 11'b01001111110;
        state_var_NS = COMP_LOOP_C_356;
      end
      COMP_LOOP_C_356 : begin
        fsm_output = 11'b01001111111;
        state_var_NS = COMP_LOOP_C_357;
      end
      COMP_LOOP_C_357 : begin
        fsm_output = 11'b01010000000;
        state_var_NS = COMP_LOOP_C_358;
      end
      COMP_LOOP_C_358 : begin
        fsm_output = 11'b01010000001;
        state_var_NS = COMP_LOOP_C_359;
      end
      COMP_LOOP_C_359 : begin
        fsm_output = 11'b01010000010;
        state_var_NS = COMP_LOOP_C_360;
      end
      COMP_LOOP_C_360 : begin
        fsm_output = 11'b01010000011;
        state_var_NS = COMP_LOOP_C_361;
      end
      COMP_LOOP_C_361 : begin
        fsm_output = 11'b01010000100;
        state_var_NS = COMP_LOOP_C_362;
      end
      COMP_LOOP_C_362 : begin
        fsm_output = 11'b01010000101;
        state_var_NS = COMP_LOOP_C_363;
      end
      COMP_LOOP_C_363 : begin
        fsm_output = 11'b01010000110;
        state_var_NS = COMP_LOOP_C_364;
      end
      COMP_LOOP_C_364 : begin
        fsm_output = 11'b01010000111;
        state_var_NS = COMP_LOOP_C_365;
      end
      COMP_LOOP_C_365 : begin
        fsm_output = 11'b01010001000;
        state_var_NS = COMP_LOOP_C_366;
      end
      COMP_LOOP_C_366 : begin
        fsm_output = 11'b01010001001;
        state_var_NS = COMP_LOOP_C_367;
      end
      COMP_LOOP_C_367 : begin
        fsm_output = 11'b01010001010;
        state_var_NS = COMP_LOOP_C_368;
      end
      COMP_LOOP_C_368 : begin
        fsm_output = 11'b01010001011;
        state_var_NS = COMP_LOOP_C_369;
      end
      COMP_LOOP_C_369 : begin
        fsm_output = 11'b01010001100;
        state_var_NS = COMP_LOOP_C_370;
      end
      COMP_LOOP_C_370 : begin
        fsm_output = 11'b01010001101;
        state_var_NS = COMP_LOOP_C_371;
      end
      COMP_LOOP_C_371 : begin
        fsm_output = 11'b01010001110;
        state_var_NS = COMP_LOOP_C_372;
      end
      COMP_LOOP_C_372 : begin
        fsm_output = 11'b01010001111;
        state_var_NS = COMP_LOOP_C_373;
      end
      COMP_LOOP_C_373 : begin
        fsm_output = 11'b01010010000;
        state_var_NS = COMP_LOOP_C_374;
      end
      COMP_LOOP_C_374 : begin
        fsm_output = 11'b01010010001;
        state_var_NS = COMP_LOOP_C_375;
      end
      COMP_LOOP_C_375 : begin
        fsm_output = 11'b01010010010;
        state_var_NS = COMP_LOOP_C_376;
      end
      COMP_LOOP_C_376 : begin
        fsm_output = 11'b01010010011;
        state_var_NS = COMP_LOOP_C_377;
      end
      COMP_LOOP_C_377 : begin
        fsm_output = 11'b01010010100;
        state_var_NS = COMP_LOOP_C_378;
      end
      COMP_LOOP_C_378 : begin
        fsm_output = 11'b01010010101;
        state_var_NS = COMP_LOOP_C_379;
      end
      COMP_LOOP_C_379 : begin
        fsm_output = 11'b01010010110;
        state_var_NS = COMP_LOOP_C_380;
      end
      COMP_LOOP_C_380 : begin
        fsm_output = 11'b01010010111;
        state_var_NS = COMP_LOOP_C_381;
      end
      COMP_LOOP_C_381 : begin
        fsm_output = 11'b01010011000;
        state_var_NS = COMP_LOOP_C_382;
      end
      COMP_LOOP_C_382 : begin
        fsm_output = 11'b01010011001;
        state_var_NS = COMP_LOOP_C_383;
      end
      COMP_LOOP_C_383 : begin
        fsm_output = 11'b01010011010;
        state_var_NS = COMP_LOOP_C_384;
      end
      COMP_LOOP_C_384 : begin
        fsm_output = 11'b01010011011;
        if ( COMP_LOOP_C_384_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_385;
        end
      end
      COMP_LOOP_C_385 : begin
        fsm_output = 11'b01010011100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
      end
      COMP_LOOP_7_modExp_1_while_C_0 : begin
        fsm_output = 11'b01010011101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_1;
      end
      COMP_LOOP_7_modExp_1_while_C_1 : begin
        fsm_output = 11'b01010011110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_2;
      end
      COMP_LOOP_7_modExp_1_while_C_2 : begin
        fsm_output = 11'b01010011111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_3;
      end
      COMP_LOOP_7_modExp_1_while_C_3 : begin
        fsm_output = 11'b01010100000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_4;
      end
      COMP_LOOP_7_modExp_1_while_C_4 : begin
        fsm_output = 11'b01010100001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_5;
      end
      COMP_LOOP_7_modExp_1_while_C_5 : begin
        fsm_output = 11'b01010100010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_6;
      end
      COMP_LOOP_7_modExp_1_while_C_6 : begin
        fsm_output = 11'b01010100011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_7;
      end
      COMP_LOOP_7_modExp_1_while_C_7 : begin
        fsm_output = 11'b01010100100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_8;
      end
      COMP_LOOP_7_modExp_1_while_C_8 : begin
        fsm_output = 11'b01010100101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_9;
      end
      COMP_LOOP_7_modExp_1_while_C_9 : begin
        fsm_output = 11'b01010100110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_10;
      end
      COMP_LOOP_7_modExp_1_while_C_10 : begin
        fsm_output = 11'b01010100111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_11;
      end
      COMP_LOOP_7_modExp_1_while_C_11 : begin
        fsm_output = 11'b01010101000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_12;
      end
      COMP_LOOP_7_modExp_1_while_C_12 : begin
        fsm_output = 11'b01010101001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_13;
      end
      COMP_LOOP_7_modExp_1_while_C_13 : begin
        fsm_output = 11'b01010101010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_14;
      end
      COMP_LOOP_7_modExp_1_while_C_14 : begin
        fsm_output = 11'b01010101011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_15;
      end
      COMP_LOOP_7_modExp_1_while_C_15 : begin
        fsm_output = 11'b01010101100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_16;
      end
      COMP_LOOP_7_modExp_1_while_C_16 : begin
        fsm_output = 11'b01010101101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_17;
      end
      COMP_LOOP_7_modExp_1_while_C_17 : begin
        fsm_output = 11'b01010101110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_18;
      end
      COMP_LOOP_7_modExp_1_while_C_18 : begin
        fsm_output = 11'b01010101111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_19;
      end
      COMP_LOOP_7_modExp_1_while_C_19 : begin
        fsm_output = 11'b01010110000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_20;
      end
      COMP_LOOP_7_modExp_1_while_C_20 : begin
        fsm_output = 11'b01010110001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_21;
      end
      COMP_LOOP_7_modExp_1_while_C_21 : begin
        fsm_output = 11'b01010110010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_22;
      end
      COMP_LOOP_7_modExp_1_while_C_22 : begin
        fsm_output = 11'b01010110011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_23;
      end
      COMP_LOOP_7_modExp_1_while_C_23 : begin
        fsm_output = 11'b01010110100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_24;
      end
      COMP_LOOP_7_modExp_1_while_C_24 : begin
        fsm_output = 11'b01010110101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_25;
      end
      COMP_LOOP_7_modExp_1_while_C_25 : begin
        fsm_output = 11'b01010110110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_26;
      end
      COMP_LOOP_7_modExp_1_while_C_26 : begin
        fsm_output = 11'b01010110111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_27;
      end
      COMP_LOOP_7_modExp_1_while_C_27 : begin
        fsm_output = 11'b01010111000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_28;
      end
      COMP_LOOP_7_modExp_1_while_C_28 : begin
        fsm_output = 11'b01010111001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_29;
      end
      COMP_LOOP_7_modExp_1_while_C_29 : begin
        fsm_output = 11'b01010111010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_30;
      end
      COMP_LOOP_7_modExp_1_while_C_30 : begin
        fsm_output = 11'b01010111011;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_31;
      end
      COMP_LOOP_7_modExp_1_while_C_31 : begin
        fsm_output = 11'b01010111100;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_32;
      end
      COMP_LOOP_7_modExp_1_while_C_32 : begin
        fsm_output = 11'b01010111101;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_33;
      end
      COMP_LOOP_7_modExp_1_while_C_33 : begin
        fsm_output = 11'b01010111110;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_34;
      end
      COMP_LOOP_7_modExp_1_while_C_34 : begin
        fsm_output = 11'b01010111111;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_35;
      end
      COMP_LOOP_7_modExp_1_while_C_35 : begin
        fsm_output = 11'b01011000000;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_36;
      end
      COMP_LOOP_7_modExp_1_while_C_36 : begin
        fsm_output = 11'b01011000001;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_37;
      end
      COMP_LOOP_7_modExp_1_while_C_37 : begin
        fsm_output = 11'b01011000010;
        state_var_NS = COMP_LOOP_7_modExp_1_while_C_38;
      end
      COMP_LOOP_7_modExp_1_while_C_38 : begin
        fsm_output = 11'b01011000011;
        if ( COMP_LOOP_7_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_386;
        end
        else begin
          state_var_NS = COMP_LOOP_7_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_386 : begin
        fsm_output = 11'b01011000100;
        state_var_NS = COMP_LOOP_C_387;
      end
      COMP_LOOP_C_387 : begin
        fsm_output = 11'b01011000101;
        state_var_NS = COMP_LOOP_C_388;
      end
      COMP_LOOP_C_388 : begin
        fsm_output = 11'b01011000110;
        state_var_NS = COMP_LOOP_C_389;
      end
      COMP_LOOP_C_389 : begin
        fsm_output = 11'b01011000111;
        state_var_NS = COMP_LOOP_C_390;
      end
      COMP_LOOP_C_390 : begin
        fsm_output = 11'b01011001000;
        state_var_NS = COMP_LOOP_C_391;
      end
      COMP_LOOP_C_391 : begin
        fsm_output = 11'b01011001001;
        state_var_NS = COMP_LOOP_C_392;
      end
      COMP_LOOP_C_392 : begin
        fsm_output = 11'b01011001010;
        state_var_NS = COMP_LOOP_C_393;
      end
      COMP_LOOP_C_393 : begin
        fsm_output = 11'b01011001011;
        state_var_NS = COMP_LOOP_C_394;
      end
      COMP_LOOP_C_394 : begin
        fsm_output = 11'b01011001100;
        state_var_NS = COMP_LOOP_C_395;
      end
      COMP_LOOP_C_395 : begin
        fsm_output = 11'b01011001101;
        state_var_NS = COMP_LOOP_C_396;
      end
      COMP_LOOP_C_396 : begin
        fsm_output = 11'b01011001110;
        state_var_NS = COMP_LOOP_C_397;
      end
      COMP_LOOP_C_397 : begin
        fsm_output = 11'b01011001111;
        state_var_NS = COMP_LOOP_C_398;
      end
      COMP_LOOP_C_398 : begin
        fsm_output = 11'b01011010000;
        state_var_NS = COMP_LOOP_C_399;
      end
      COMP_LOOP_C_399 : begin
        fsm_output = 11'b01011010001;
        state_var_NS = COMP_LOOP_C_400;
      end
      COMP_LOOP_C_400 : begin
        fsm_output = 11'b01011010010;
        state_var_NS = COMP_LOOP_C_401;
      end
      COMP_LOOP_C_401 : begin
        fsm_output = 11'b01011010011;
        state_var_NS = COMP_LOOP_C_402;
      end
      COMP_LOOP_C_402 : begin
        fsm_output = 11'b01011010100;
        state_var_NS = COMP_LOOP_C_403;
      end
      COMP_LOOP_C_403 : begin
        fsm_output = 11'b01011010101;
        state_var_NS = COMP_LOOP_C_404;
      end
      COMP_LOOP_C_404 : begin
        fsm_output = 11'b01011010110;
        state_var_NS = COMP_LOOP_C_405;
      end
      COMP_LOOP_C_405 : begin
        fsm_output = 11'b01011010111;
        state_var_NS = COMP_LOOP_C_406;
      end
      COMP_LOOP_C_406 : begin
        fsm_output = 11'b01011011000;
        state_var_NS = COMP_LOOP_C_407;
      end
      COMP_LOOP_C_407 : begin
        fsm_output = 11'b01011011001;
        state_var_NS = COMP_LOOP_C_408;
      end
      COMP_LOOP_C_408 : begin
        fsm_output = 11'b01011011010;
        state_var_NS = COMP_LOOP_C_409;
      end
      COMP_LOOP_C_409 : begin
        fsm_output = 11'b01011011011;
        state_var_NS = COMP_LOOP_C_410;
      end
      COMP_LOOP_C_410 : begin
        fsm_output = 11'b01011011100;
        state_var_NS = COMP_LOOP_C_411;
      end
      COMP_LOOP_C_411 : begin
        fsm_output = 11'b01011011101;
        state_var_NS = COMP_LOOP_C_412;
      end
      COMP_LOOP_C_412 : begin
        fsm_output = 11'b01011011110;
        state_var_NS = COMP_LOOP_C_413;
      end
      COMP_LOOP_C_413 : begin
        fsm_output = 11'b01011011111;
        state_var_NS = COMP_LOOP_C_414;
      end
      COMP_LOOP_C_414 : begin
        fsm_output = 11'b01011100000;
        state_var_NS = COMP_LOOP_C_415;
      end
      COMP_LOOP_C_415 : begin
        fsm_output = 11'b01011100001;
        state_var_NS = COMP_LOOP_C_416;
      end
      COMP_LOOP_C_416 : begin
        fsm_output = 11'b01011100010;
        state_var_NS = COMP_LOOP_C_417;
      end
      COMP_LOOP_C_417 : begin
        fsm_output = 11'b01011100011;
        state_var_NS = COMP_LOOP_C_418;
      end
      COMP_LOOP_C_418 : begin
        fsm_output = 11'b01011100100;
        state_var_NS = COMP_LOOP_C_419;
      end
      COMP_LOOP_C_419 : begin
        fsm_output = 11'b01011100101;
        state_var_NS = COMP_LOOP_C_420;
      end
      COMP_LOOP_C_420 : begin
        fsm_output = 11'b01011100110;
        state_var_NS = COMP_LOOP_C_421;
      end
      COMP_LOOP_C_421 : begin
        fsm_output = 11'b01011100111;
        state_var_NS = COMP_LOOP_C_422;
      end
      COMP_LOOP_C_422 : begin
        fsm_output = 11'b01011101000;
        state_var_NS = COMP_LOOP_C_423;
      end
      COMP_LOOP_C_423 : begin
        fsm_output = 11'b01011101001;
        state_var_NS = COMP_LOOP_C_424;
      end
      COMP_LOOP_C_424 : begin
        fsm_output = 11'b01011101010;
        state_var_NS = COMP_LOOP_C_425;
      end
      COMP_LOOP_C_425 : begin
        fsm_output = 11'b01011101011;
        state_var_NS = COMP_LOOP_C_426;
      end
      COMP_LOOP_C_426 : begin
        fsm_output = 11'b01011101100;
        state_var_NS = COMP_LOOP_C_427;
      end
      COMP_LOOP_C_427 : begin
        fsm_output = 11'b01011101101;
        state_var_NS = COMP_LOOP_C_428;
      end
      COMP_LOOP_C_428 : begin
        fsm_output = 11'b01011101110;
        state_var_NS = COMP_LOOP_C_429;
      end
      COMP_LOOP_C_429 : begin
        fsm_output = 11'b01011101111;
        state_var_NS = COMP_LOOP_C_430;
      end
      COMP_LOOP_C_430 : begin
        fsm_output = 11'b01011110000;
        state_var_NS = COMP_LOOP_C_431;
      end
      COMP_LOOP_C_431 : begin
        fsm_output = 11'b01011110001;
        state_var_NS = COMP_LOOP_C_432;
      end
      COMP_LOOP_C_432 : begin
        fsm_output = 11'b01011110010;
        state_var_NS = COMP_LOOP_C_433;
      end
      COMP_LOOP_C_433 : begin
        fsm_output = 11'b01011110011;
        state_var_NS = COMP_LOOP_C_434;
      end
      COMP_LOOP_C_434 : begin
        fsm_output = 11'b01011110100;
        state_var_NS = COMP_LOOP_C_435;
      end
      COMP_LOOP_C_435 : begin
        fsm_output = 11'b01011110101;
        state_var_NS = COMP_LOOP_C_436;
      end
      COMP_LOOP_C_436 : begin
        fsm_output = 11'b01011110110;
        state_var_NS = COMP_LOOP_C_437;
      end
      COMP_LOOP_C_437 : begin
        fsm_output = 11'b01011110111;
        state_var_NS = COMP_LOOP_C_438;
      end
      COMP_LOOP_C_438 : begin
        fsm_output = 11'b01011111000;
        state_var_NS = COMP_LOOP_C_439;
      end
      COMP_LOOP_C_439 : begin
        fsm_output = 11'b01011111001;
        state_var_NS = COMP_LOOP_C_440;
      end
      COMP_LOOP_C_440 : begin
        fsm_output = 11'b01011111010;
        state_var_NS = COMP_LOOP_C_441;
      end
      COMP_LOOP_C_441 : begin
        fsm_output = 11'b01011111011;
        state_var_NS = COMP_LOOP_C_442;
      end
      COMP_LOOP_C_442 : begin
        fsm_output = 11'b01011111100;
        state_var_NS = COMP_LOOP_C_443;
      end
      COMP_LOOP_C_443 : begin
        fsm_output = 11'b01011111101;
        state_var_NS = COMP_LOOP_C_444;
      end
      COMP_LOOP_C_444 : begin
        fsm_output = 11'b01011111110;
        state_var_NS = COMP_LOOP_C_445;
      end
      COMP_LOOP_C_445 : begin
        fsm_output = 11'b01011111111;
        state_var_NS = COMP_LOOP_C_446;
      end
      COMP_LOOP_C_446 : begin
        fsm_output = 11'b01100000000;
        state_var_NS = COMP_LOOP_C_447;
      end
      COMP_LOOP_C_447 : begin
        fsm_output = 11'b01100000001;
        state_var_NS = COMP_LOOP_C_448;
      end
      COMP_LOOP_C_448 : begin
        fsm_output = 11'b01100000010;
        if ( COMP_LOOP_C_448_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_449;
        end
      end
      COMP_LOOP_C_449 : begin
        fsm_output = 11'b01100000011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
      end
      COMP_LOOP_8_modExp_1_while_C_0 : begin
        fsm_output = 11'b01100000100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_1;
      end
      COMP_LOOP_8_modExp_1_while_C_1 : begin
        fsm_output = 11'b01100000101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_2;
      end
      COMP_LOOP_8_modExp_1_while_C_2 : begin
        fsm_output = 11'b01100000110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_3;
      end
      COMP_LOOP_8_modExp_1_while_C_3 : begin
        fsm_output = 11'b01100000111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_4;
      end
      COMP_LOOP_8_modExp_1_while_C_4 : begin
        fsm_output = 11'b01100001000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_5;
      end
      COMP_LOOP_8_modExp_1_while_C_5 : begin
        fsm_output = 11'b01100001001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_6;
      end
      COMP_LOOP_8_modExp_1_while_C_6 : begin
        fsm_output = 11'b01100001010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_7;
      end
      COMP_LOOP_8_modExp_1_while_C_7 : begin
        fsm_output = 11'b01100001011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_8;
      end
      COMP_LOOP_8_modExp_1_while_C_8 : begin
        fsm_output = 11'b01100001100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_9;
      end
      COMP_LOOP_8_modExp_1_while_C_9 : begin
        fsm_output = 11'b01100001101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_10;
      end
      COMP_LOOP_8_modExp_1_while_C_10 : begin
        fsm_output = 11'b01100001110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_11;
      end
      COMP_LOOP_8_modExp_1_while_C_11 : begin
        fsm_output = 11'b01100001111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_12;
      end
      COMP_LOOP_8_modExp_1_while_C_12 : begin
        fsm_output = 11'b01100010000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_13;
      end
      COMP_LOOP_8_modExp_1_while_C_13 : begin
        fsm_output = 11'b01100010001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_14;
      end
      COMP_LOOP_8_modExp_1_while_C_14 : begin
        fsm_output = 11'b01100010010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_15;
      end
      COMP_LOOP_8_modExp_1_while_C_15 : begin
        fsm_output = 11'b01100010011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_16;
      end
      COMP_LOOP_8_modExp_1_while_C_16 : begin
        fsm_output = 11'b01100010100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_17;
      end
      COMP_LOOP_8_modExp_1_while_C_17 : begin
        fsm_output = 11'b01100010101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_18;
      end
      COMP_LOOP_8_modExp_1_while_C_18 : begin
        fsm_output = 11'b01100010110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_19;
      end
      COMP_LOOP_8_modExp_1_while_C_19 : begin
        fsm_output = 11'b01100010111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_20;
      end
      COMP_LOOP_8_modExp_1_while_C_20 : begin
        fsm_output = 11'b01100011000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_21;
      end
      COMP_LOOP_8_modExp_1_while_C_21 : begin
        fsm_output = 11'b01100011001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_22;
      end
      COMP_LOOP_8_modExp_1_while_C_22 : begin
        fsm_output = 11'b01100011010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_23;
      end
      COMP_LOOP_8_modExp_1_while_C_23 : begin
        fsm_output = 11'b01100011011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_24;
      end
      COMP_LOOP_8_modExp_1_while_C_24 : begin
        fsm_output = 11'b01100011100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_25;
      end
      COMP_LOOP_8_modExp_1_while_C_25 : begin
        fsm_output = 11'b01100011101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_26;
      end
      COMP_LOOP_8_modExp_1_while_C_26 : begin
        fsm_output = 11'b01100011110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_27;
      end
      COMP_LOOP_8_modExp_1_while_C_27 : begin
        fsm_output = 11'b01100011111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_28;
      end
      COMP_LOOP_8_modExp_1_while_C_28 : begin
        fsm_output = 11'b01100100000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_29;
      end
      COMP_LOOP_8_modExp_1_while_C_29 : begin
        fsm_output = 11'b01100100001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_30;
      end
      COMP_LOOP_8_modExp_1_while_C_30 : begin
        fsm_output = 11'b01100100010;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_31;
      end
      COMP_LOOP_8_modExp_1_while_C_31 : begin
        fsm_output = 11'b01100100011;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_32;
      end
      COMP_LOOP_8_modExp_1_while_C_32 : begin
        fsm_output = 11'b01100100100;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_33;
      end
      COMP_LOOP_8_modExp_1_while_C_33 : begin
        fsm_output = 11'b01100100101;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_34;
      end
      COMP_LOOP_8_modExp_1_while_C_34 : begin
        fsm_output = 11'b01100100110;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_35;
      end
      COMP_LOOP_8_modExp_1_while_C_35 : begin
        fsm_output = 11'b01100100111;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_36;
      end
      COMP_LOOP_8_modExp_1_while_C_36 : begin
        fsm_output = 11'b01100101000;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_37;
      end
      COMP_LOOP_8_modExp_1_while_C_37 : begin
        fsm_output = 11'b01100101001;
        state_var_NS = COMP_LOOP_8_modExp_1_while_C_38;
      end
      COMP_LOOP_8_modExp_1_while_C_38 : begin
        fsm_output = 11'b01100101010;
        if ( COMP_LOOP_8_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_450;
        end
        else begin
          state_var_NS = COMP_LOOP_8_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_450 : begin
        fsm_output = 11'b01100101011;
        state_var_NS = COMP_LOOP_C_451;
      end
      COMP_LOOP_C_451 : begin
        fsm_output = 11'b01100101100;
        state_var_NS = COMP_LOOP_C_452;
      end
      COMP_LOOP_C_452 : begin
        fsm_output = 11'b01100101101;
        state_var_NS = COMP_LOOP_C_453;
      end
      COMP_LOOP_C_453 : begin
        fsm_output = 11'b01100101110;
        state_var_NS = COMP_LOOP_C_454;
      end
      COMP_LOOP_C_454 : begin
        fsm_output = 11'b01100101111;
        state_var_NS = COMP_LOOP_C_455;
      end
      COMP_LOOP_C_455 : begin
        fsm_output = 11'b01100110000;
        state_var_NS = COMP_LOOP_C_456;
      end
      COMP_LOOP_C_456 : begin
        fsm_output = 11'b01100110001;
        state_var_NS = COMP_LOOP_C_457;
      end
      COMP_LOOP_C_457 : begin
        fsm_output = 11'b01100110010;
        state_var_NS = COMP_LOOP_C_458;
      end
      COMP_LOOP_C_458 : begin
        fsm_output = 11'b01100110011;
        state_var_NS = COMP_LOOP_C_459;
      end
      COMP_LOOP_C_459 : begin
        fsm_output = 11'b01100110100;
        state_var_NS = COMP_LOOP_C_460;
      end
      COMP_LOOP_C_460 : begin
        fsm_output = 11'b01100110101;
        state_var_NS = COMP_LOOP_C_461;
      end
      COMP_LOOP_C_461 : begin
        fsm_output = 11'b01100110110;
        state_var_NS = COMP_LOOP_C_462;
      end
      COMP_LOOP_C_462 : begin
        fsm_output = 11'b01100110111;
        state_var_NS = COMP_LOOP_C_463;
      end
      COMP_LOOP_C_463 : begin
        fsm_output = 11'b01100111000;
        state_var_NS = COMP_LOOP_C_464;
      end
      COMP_LOOP_C_464 : begin
        fsm_output = 11'b01100111001;
        state_var_NS = COMP_LOOP_C_465;
      end
      COMP_LOOP_C_465 : begin
        fsm_output = 11'b01100111010;
        state_var_NS = COMP_LOOP_C_466;
      end
      COMP_LOOP_C_466 : begin
        fsm_output = 11'b01100111011;
        state_var_NS = COMP_LOOP_C_467;
      end
      COMP_LOOP_C_467 : begin
        fsm_output = 11'b01100111100;
        state_var_NS = COMP_LOOP_C_468;
      end
      COMP_LOOP_C_468 : begin
        fsm_output = 11'b01100111101;
        state_var_NS = COMP_LOOP_C_469;
      end
      COMP_LOOP_C_469 : begin
        fsm_output = 11'b01100111110;
        state_var_NS = COMP_LOOP_C_470;
      end
      COMP_LOOP_C_470 : begin
        fsm_output = 11'b01100111111;
        state_var_NS = COMP_LOOP_C_471;
      end
      COMP_LOOP_C_471 : begin
        fsm_output = 11'b01101000000;
        state_var_NS = COMP_LOOP_C_472;
      end
      COMP_LOOP_C_472 : begin
        fsm_output = 11'b01101000001;
        state_var_NS = COMP_LOOP_C_473;
      end
      COMP_LOOP_C_473 : begin
        fsm_output = 11'b01101000010;
        state_var_NS = COMP_LOOP_C_474;
      end
      COMP_LOOP_C_474 : begin
        fsm_output = 11'b01101000011;
        state_var_NS = COMP_LOOP_C_475;
      end
      COMP_LOOP_C_475 : begin
        fsm_output = 11'b01101000100;
        state_var_NS = COMP_LOOP_C_476;
      end
      COMP_LOOP_C_476 : begin
        fsm_output = 11'b01101000101;
        state_var_NS = COMP_LOOP_C_477;
      end
      COMP_LOOP_C_477 : begin
        fsm_output = 11'b01101000110;
        state_var_NS = COMP_LOOP_C_478;
      end
      COMP_LOOP_C_478 : begin
        fsm_output = 11'b01101000111;
        state_var_NS = COMP_LOOP_C_479;
      end
      COMP_LOOP_C_479 : begin
        fsm_output = 11'b01101001000;
        state_var_NS = COMP_LOOP_C_480;
      end
      COMP_LOOP_C_480 : begin
        fsm_output = 11'b01101001001;
        state_var_NS = COMP_LOOP_C_481;
      end
      COMP_LOOP_C_481 : begin
        fsm_output = 11'b01101001010;
        state_var_NS = COMP_LOOP_C_482;
      end
      COMP_LOOP_C_482 : begin
        fsm_output = 11'b01101001011;
        state_var_NS = COMP_LOOP_C_483;
      end
      COMP_LOOP_C_483 : begin
        fsm_output = 11'b01101001100;
        state_var_NS = COMP_LOOP_C_484;
      end
      COMP_LOOP_C_484 : begin
        fsm_output = 11'b01101001101;
        state_var_NS = COMP_LOOP_C_485;
      end
      COMP_LOOP_C_485 : begin
        fsm_output = 11'b01101001110;
        state_var_NS = COMP_LOOP_C_486;
      end
      COMP_LOOP_C_486 : begin
        fsm_output = 11'b01101001111;
        state_var_NS = COMP_LOOP_C_487;
      end
      COMP_LOOP_C_487 : begin
        fsm_output = 11'b01101010000;
        state_var_NS = COMP_LOOP_C_488;
      end
      COMP_LOOP_C_488 : begin
        fsm_output = 11'b01101010001;
        state_var_NS = COMP_LOOP_C_489;
      end
      COMP_LOOP_C_489 : begin
        fsm_output = 11'b01101010010;
        state_var_NS = COMP_LOOP_C_490;
      end
      COMP_LOOP_C_490 : begin
        fsm_output = 11'b01101010011;
        state_var_NS = COMP_LOOP_C_491;
      end
      COMP_LOOP_C_491 : begin
        fsm_output = 11'b01101010100;
        state_var_NS = COMP_LOOP_C_492;
      end
      COMP_LOOP_C_492 : begin
        fsm_output = 11'b01101010101;
        state_var_NS = COMP_LOOP_C_493;
      end
      COMP_LOOP_C_493 : begin
        fsm_output = 11'b01101010110;
        state_var_NS = COMP_LOOP_C_494;
      end
      COMP_LOOP_C_494 : begin
        fsm_output = 11'b01101010111;
        state_var_NS = COMP_LOOP_C_495;
      end
      COMP_LOOP_C_495 : begin
        fsm_output = 11'b01101011000;
        state_var_NS = COMP_LOOP_C_496;
      end
      COMP_LOOP_C_496 : begin
        fsm_output = 11'b01101011001;
        state_var_NS = COMP_LOOP_C_497;
      end
      COMP_LOOP_C_497 : begin
        fsm_output = 11'b01101011010;
        state_var_NS = COMP_LOOP_C_498;
      end
      COMP_LOOP_C_498 : begin
        fsm_output = 11'b01101011011;
        state_var_NS = COMP_LOOP_C_499;
      end
      COMP_LOOP_C_499 : begin
        fsm_output = 11'b01101011100;
        state_var_NS = COMP_LOOP_C_500;
      end
      COMP_LOOP_C_500 : begin
        fsm_output = 11'b01101011101;
        state_var_NS = COMP_LOOP_C_501;
      end
      COMP_LOOP_C_501 : begin
        fsm_output = 11'b01101011110;
        state_var_NS = COMP_LOOP_C_502;
      end
      COMP_LOOP_C_502 : begin
        fsm_output = 11'b01101011111;
        state_var_NS = COMP_LOOP_C_503;
      end
      COMP_LOOP_C_503 : begin
        fsm_output = 11'b01101100000;
        state_var_NS = COMP_LOOP_C_504;
      end
      COMP_LOOP_C_504 : begin
        fsm_output = 11'b01101100001;
        state_var_NS = COMP_LOOP_C_505;
      end
      COMP_LOOP_C_505 : begin
        fsm_output = 11'b01101100010;
        state_var_NS = COMP_LOOP_C_506;
      end
      COMP_LOOP_C_506 : begin
        fsm_output = 11'b01101100011;
        state_var_NS = COMP_LOOP_C_507;
      end
      COMP_LOOP_C_507 : begin
        fsm_output = 11'b01101100100;
        state_var_NS = COMP_LOOP_C_508;
      end
      COMP_LOOP_C_508 : begin
        fsm_output = 11'b01101100101;
        state_var_NS = COMP_LOOP_C_509;
      end
      COMP_LOOP_C_509 : begin
        fsm_output = 11'b01101100110;
        state_var_NS = COMP_LOOP_C_510;
      end
      COMP_LOOP_C_510 : begin
        fsm_output = 11'b01101100111;
        state_var_NS = COMP_LOOP_C_511;
      end
      COMP_LOOP_C_511 : begin
        fsm_output = 11'b01101101000;
        state_var_NS = COMP_LOOP_C_512;
      end
      COMP_LOOP_C_512 : begin
        fsm_output = 11'b01101101001;
        if ( COMP_LOOP_C_512_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_513;
        end
      end
      COMP_LOOP_C_513 : begin
        fsm_output = 11'b01101101010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_0;
      end
      COMP_LOOP_9_modExp_1_while_C_0 : begin
        fsm_output = 11'b01101101011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_1;
      end
      COMP_LOOP_9_modExp_1_while_C_1 : begin
        fsm_output = 11'b01101101100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_2;
      end
      COMP_LOOP_9_modExp_1_while_C_2 : begin
        fsm_output = 11'b01101101101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_3;
      end
      COMP_LOOP_9_modExp_1_while_C_3 : begin
        fsm_output = 11'b01101101110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_4;
      end
      COMP_LOOP_9_modExp_1_while_C_4 : begin
        fsm_output = 11'b01101101111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_5;
      end
      COMP_LOOP_9_modExp_1_while_C_5 : begin
        fsm_output = 11'b01101110000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_6;
      end
      COMP_LOOP_9_modExp_1_while_C_6 : begin
        fsm_output = 11'b01101110001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_7;
      end
      COMP_LOOP_9_modExp_1_while_C_7 : begin
        fsm_output = 11'b01101110010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_8;
      end
      COMP_LOOP_9_modExp_1_while_C_8 : begin
        fsm_output = 11'b01101110011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_9;
      end
      COMP_LOOP_9_modExp_1_while_C_9 : begin
        fsm_output = 11'b01101110100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_10;
      end
      COMP_LOOP_9_modExp_1_while_C_10 : begin
        fsm_output = 11'b01101110101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_11;
      end
      COMP_LOOP_9_modExp_1_while_C_11 : begin
        fsm_output = 11'b01101110110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_12;
      end
      COMP_LOOP_9_modExp_1_while_C_12 : begin
        fsm_output = 11'b01101110111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_13;
      end
      COMP_LOOP_9_modExp_1_while_C_13 : begin
        fsm_output = 11'b01101111000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_14;
      end
      COMP_LOOP_9_modExp_1_while_C_14 : begin
        fsm_output = 11'b01101111001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_15;
      end
      COMP_LOOP_9_modExp_1_while_C_15 : begin
        fsm_output = 11'b01101111010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_16;
      end
      COMP_LOOP_9_modExp_1_while_C_16 : begin
        fsm_output = 11'b01101111011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_17;
      end
      COMP_LOOP_9_modExp_1_while_C_17 : begin
        fsm_output = 11'b01101111100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_18;
      end
      COMP_LOOP_9_modExp_1_while_C_18 : begin
        fsm_output = 11'b01101111101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_19;
      end
      COMP_LOOP_9_modExp_1_while_C_19 : begin
        fsm_output = 11'b01101111110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_20;
      end
      COMP_LOOP_9_modExp_1_while_C_20 : begin
        fsm_output = 11'b01101111111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_21;
      end
      COMP_LOOP_9_modExp_1_while_C_21 : begin
        fsm_output = 11'b01110000000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_22;
      end
      COMP_LOOP_9_modExp_1_while_C_22 : begin
        fsm_output = 11'b01110000001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_23;
      end
      COMP_LOOP_9_modExp_1_while_C_23 : begin
        fsm_output = 11'b01110000010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_24;
      end
      COMP_LOOP_9_modExp_1_while_C_24 : begin
        fsm_output = 11'b01110000011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_25;
      end
      COMP_LOOP_9_modExp_1_while_C_25 : begin
        fsm_output = 11'b01110000100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_26;
      end
      COMP_LOOP_9_modExp_1_while_C_26 : begin
        fsm_output = 11'b01110000101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_27;
      end
      COMP_LOOP_9_modExp_1_while_C_27 : begin
        fsm_output = 11'b01110000110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_28;
      end
      COMP_LOOP_9_modExp_1_while_C_28 : begin
        fsm_output = 11'b01110000111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_29;
      end
      COMP_LOOP_9_modExp_1_while_C_29 : begin
        fsm_output = 11'b01110001000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_30;
      end
      COMP_LOOP_9_modExp_1_while_C_30 : begin
        fsm_output = 11'b01110001001;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_31;
      end
      COMP_LOOP_9_modExp_1_while_C_31 : begin
        fsm_output = 11'b01110001010;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_32;
      end
      COMP_LOOP_9_modExp_1_while_C_32 : begin
        fsm_output = 11'b01110001011;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_33;
      end
      COMP_LOOP_9_modExp_1_while_C_33 : begin
        fsm_output = 11'b01110001100;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_34;
      end
      COMP_LOOP_9_modExp_1_while_C_34 : begin
        fsm_output = 11'b01110001101;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_35;
      end
      COMP_LOOP_9_modExp_1_while_C_35 : begin
        fsm_output = 11'b01110001110;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_36;
      end
      COMP_LOOP_9_modExp_1_while_C_36 : begin
        fsm_output = 11'b01110001111;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_37;
      end
      COMP_LOOP_9_modExp_1_while_C_37 : begin
        fsm_output = 11'b01110010000;
        state_var_NS = COMP_LOOP_9_modExp_1_while_C_38;
      end
      COMP_LOOP_9_modExp_1_while_C_38 : begin
        fsm_output = 11'b01110010001;
        if ( COMP_LOOP_9_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_514;
        end
        else begin
          state_var_NS = COMP_LOOP_9_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_514 : begin
        fsm_output = 11'b01110010010;
        state_var_NS = COMP_LOOP_C_515;
      end
      COMP_LOOP_C_515 : begin
        fsm_output = 11'b01110010011;
        state_var_NS = COMP_LOOP_C_516;
      end
      COMP_LOOP_C_516 : begin
        fsm_output = 11'b01110010100;
        state_var_NS = COMP_LOOP_C_517;
      end
      COMP_LOOP_C_517 : begin
        fsm_output = 11'b01110010101;
        state_var_NS = COMP_LOOP_C_518;
      end
      COMP_LOOP_C_518 : begin
        fsm_output = 11'b01110010110;
        state_var_NS = COMP_LOOP_C_519;
      end
      COMP_LOOP_C_519 : begin
        fsm_output = 11'b01110010111;
        state_var_NS = COMP_LOOP_C_520;
      end
      COMP_LOOP_C_520 : begin
        fsm_output = 11'b01110011000;
        state_var_NS = COMP_LOOP_C_521;
      end
      COMP_LOOP_C_521 : begin
        fsm_output = 11'b01110011001;
        state_var_NS = COMP_LOOP_C_522;
      end
      COMP_LOOP_C_522 : begin
        fsm_output = 11'b01110011010;
        state_var_NS = COMP_LOOP_C_523;
      end
      COMP_LOOP_C_523 : begin
        fsm_output = 11'b01110011011;
        state_var_NS = COMP_LOOP_C_524;
      end
      COMP_LOOP_C_524 : begin
        fsm_output = 11'b01110011100;
        state_var_NS = COMP_LOOP_C_525;
      end
      COMP_LOOP_C_525 : begin
        fsm_output = 11'b01110011101;
        state_var_NS = COMP_LOOP_C_526;
      end
      COMP_LOOP_C_526 : begin
        fsm_output = 11'b01110011110;
        state_var_NS = COMP_LOOP_C_527;
      end
      COMP_LOOP_C_527 : begin
        fsm_output = 11'b01110011111;
        state_var_NS = COMP_LOOP_C_528;
      end
      COMP_LOOP_C_528 : begin
        fsm_output = 11'b01110100000;
        state_var_NS = COMP_LOOP_C_529;
      end
      COMP_LOOP_C_529 : begin
        fsm_output = 11'b01110100001;
        state_var_NS = COMP_LOOP_C_530;
      end
      COMP_LOOP_C_530 : begin
        fsm_output = 11'b01110100010;
        state_var_NS = COMP_LOOP_C_531;
      end
      COMP_LOOP_C_531 : begin
        fsm_output = 11'b01110100011;
        state_var_NS = COMP_LOOP_C_532;
      end
      COMP_LOOP_C_532 : begin
        fsm_output = 11'b01110100100;
        state_var_NS = COMP_LOOP_C_533;
      end
      COMP_LOOP_C_533 : begin
        fsm_output = 11'b01110100101;
        state_var_NS = COMP_LOOP_C_534;
      end
      COMP_LOOP_C_534 : begin
        fsm_output = 11'b01110100110;
        state_var_NS = COMP_LOOP_C_535;
      end
      COMP_LOOP_C_535 : begin
        fsm_output = 11'b01110100111;
        state_var_NS = COMP_LOOP_C_536;
      end
      COMP_LOOP_C_536 : begin
        fsm_output = 11'b01110101000;
        state_var_NS = COMP_LOOP_C_537;
      end
      COMP_LOOP_C_537 : begin
        fsm_output = 11'b01110101001;
        state_var_NS = COMP_LOOP_C_538;
      end
      COMP_LOOP_C_538 : begin
        fsm_output = 11'b01110101010;
        state_var_NS = COMP_LOOP_C_539;
      end
      COMP_LOOP_C_539 : begin
        fsm_output = 11'b01110101011;
        state_var_NS = COMP_LOOP_C_540;
      end
      COMP_LOOP_C_540 : begin
        fsm_output = 11'b01110101100;
        state_var_NS = COMP_LOOP_C_541;
      end
      COMP_LOOP_C_541 : begin
        fsm_output = 11'b01110101101;
        state_var_NS = COMP_LOOP_C_542;
      end
      COMP_LOOP_C_542 : begin
        fsm_output = 11'b01110101110;
        state_var_NS = COMP_LOOP_C_543;
      end
      COMP_LOOP_C_543 : begin
        fsm_output = 11'b01110101111;
        state_var_NS = COMP_LOOP_C_544;
      end
      COMP_LOOP_C_544 : begin
        fsm_output = 11'b01110110000;
        state_var_NS = COMP_LOOP_C_545;
      end
      COMP_LOOP_C_545 : begin
        fsm_output = 11'b01110110001;
        state_var_NS = COMP_LOOP_C_546;
      end
      COMP_LOOP_C_546 : begin
        fsm_output = 11'b01110110010;
        state_var_NS = COMP_LOOP_C_547;
      end
      COMP_LOOP_C_547 : begin
        fsm_output = 11'b01110110011;
        state_var_NS = COMP_LOOP_C_548;
      end
      COMP_LOOP_C_548 : begin
        fsm_output = 11'b01110110100;
        state_var_NS = COMP_LOOP_C_549;
      end
      COMP_LOOP_C_549 : begin
        fsm_output = 11'b01110110101;
        state_var_NS = COMP_LOOP_C_550;
      end
      COMP_LOOP_C_550 : begin
        fsm_output = 11'b01110110110;
        state_var_NS = COMP_LOOP_C_551;
      end
      COMP_LOOP_C_551 : begin
        fsm_output = 11'b01110110111;
        state_var_NS = COMP_LOOP_C_552;
      end
      COMP_LOOP_C_552 : begin
        fsm_output = 11'b01110111000;
        state_var_NS = COMP_LOOP_C_553;
      end
      COMP_LOOP_C_553 : begin
        fsm_output = 11'b01110111001;
        state_var_NS = COMP_LOOP_C_554;
      end
      COMP_LOOP_C_554 : begin
        fsm_output = 11'b01110111010;
        state_var_NS = COMP_LOOP_C_555;
      end
      COMP_LOOP_C_555 : begin
        fsm_output = 11'b01110111011;
        state_var_NS = COMP_LOOP_C_556;
      end
      COMP_LOOP_C_556 : begin
        fsm_output = 11'b01110111100;
        state_var_NS = COMP_LOOP_C_557;
      end
      COMP_LOOP_C_557 : begin
        fsm_output = 11'b01110111101;
        state_var_NS = COMP_LOOP_C_558;
      end
      COMP_LOOP_C_558 : begin
        fsm_output = 11'b01110111110;
        state_var_NS = COMP_LOOP_C_559;
      end
      COMP_LOOP_C_559 : begin
        fsm_output = 11'b01110111111;
        state_var_NS = COMP_LOOP_C_560;
      end
      COMP_LOOP_C_560 : begin
        fsm_output = 11'b01111000000;
        state_var_NS = COMP_LOOP_C_561;
      end
      COMP_LOOP_C_561 : begin
        fsm_output = 11'b01111000001;
        state_var_NS = COMP_LOOP_C_562;
      end
      COMP_LOOP_C_562 : begin
        fsm_output = 11'b01111000010;
        state_var_NS = COMP_LOOP_C_563;
      end
      COMP_LOOP_C_563 : begin
        fsm_output = 11'b01111000011;
        state_var_NS = COMP_LOOP_C_564;
      end
      COMP_LOOP_C_564 : begin
        fsm_output = 11'b01111000100;
        state_var_NS = COMP_LOOP_C_565;
      end
      COMP_LOOP_C_565 : begin
        fsm_output = 11'b01111000101;
        state_var_NS = COMP_LOOP_C_566;
      end
      COMP_LOOP_C_566 : begin
        fsm_output = 11'b01111000110;
        state_var_NS = COMP_LOOP_C_567;
      end
      COMP_LOOP_C_567 : begin
        fsm_output = 11'b01111000111;
        state_var_NS = COMP_LOOP_C_568;
      end
      COMP_LOOP_C_568 : begin
        fsm_output = 11'b01111001000;
        state_var_NS = COMP_LOOP_C_569;
      end
      COMP_LOOP_C_569 : begin
        fsm_output = 11'b01111001001;
        state_var_NS = COMP_LOOP_C_570;
      end
      COMP_LOOP_C_570 : begin
        fsm_output = 11'b01111001010;
        state_var_NS = COMP_LOOP_C_571;
      end
      COMP_LOOP_C_571 : begin
        fsm_output = 11'b01111001011;
        state_var_NS = COMP_LOOP_C_572;
      end
      COMP_LOOP_C_572 : begin
        fsm_output = 11'b01111001100;
        state_var_NS = COMP_LOOP_C_573;
      end
      COMP_LOOP_C_573 : begin
        fsm_output = 11'b01111001101;
        state_var_NS = COMP_LOOP_C_574;
      end
      COMP_LOOP_C_574 : begin
        fsm_output = 11'b01111001110;
        state_var_NS = COMP_LOOP_C_575;
      end
      COMP_LOOP_C_575 : begin
        fsm_output = 11'b01111001111;
        state_var_NS = COMP_LOOP_C_576;
      end
      COMP_LOOP_C_576 : begin
        fsm_output = 11'b01111010000;
        if ( COMP_LOOP_C_576_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_577;
        end
      end
      COMP_LOOP_C_577 : begin
        fsm_output = 11'b01111010001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_0;
      end
      COMP_LOOP_10_modExp_1_while_C_0 : begin
        fsm_output = 11'b01111010010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_1;
      end
      COMP_LOOP_10_modExp_1_while_C_1 : begin
        fsm_output = 11'b01111010011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_2;
      end
      COMP_LOOP_10_modExp_1_while_C_2 : begin
        fsm_output = 11'b01111010100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_3;
      end
      COMP_LOOP_10_modExp_1_while_C_3 : begin
        fsm_output = 11'b01111010101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_4;
      end
      COMP_LOOP_10_modExp_1_while_C_4 : begin
        fsm_output = 11'b01111010110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_5;
      end
      COMP_LOOP_10_modExp_1_while_C_5 : begin
        fsm_output = 11'b01111010111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_6;
      end
      COMP_LOOP_10_modExp_1_while_C_6 : begin
        fsm_output = 11'b01111011000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_7;
      end
      COMP_LOOP_10_modExp_1_while_C_7 : begin
        fsm_output = 11'b01111011001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_8;
      end
      COMP_LOOP_10_modExp_1_while_C_8 : begin
        fsm_output = 11'b01111011010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_9;
      end
      COMP_LOOP_10_modExp_1_while_C_9 : begin
        fsm_output = 11'b01111011011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_10;
      end
      COMP_LOOP_10_modExp_1_while_C_10 : begin
        fsm_output = 11'b01111011100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_11;
      end
      COMP_LOOP_10_modExp_1_while_C_11 : begin
        fsm_output = 11'b01111011101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_12;
      end
      COMP_LOOP_10_modExp_1_while_C_12 : begin
        fsm_output = 11'b01111011110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_13;
      end
      COMP_LOOP_10_modExp_1_while_C_13 : begin
        fsm_output = 11'b01111011111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_14;
      end
      COMP_LOOP_10_modExp_1_while_C_14 : begin
        fsm_output = 11'b01111100000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_15;
      end
      COMP_LOOP_10_modExp_1_while_C_15 : begin
        fsm_output = 11'b01111100001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_16;
      end
      COMP_LOOP_10_modExp_1_while_C_16 : begin
        fsm_output = 11'b01111100010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_17;
      end
      COMP_LOOP_10_modExp_1_while_C_17 : begin
        fsm_output = 11'b01111100011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_18;
      end
      COMP_LOOP_10_modExp_1_while_C_18 : begin
        fsm_output = 11'b01111100100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_19;
      end
      COMP_LOOP_10_modExp_1_while_C_19 : begin
        fsm_output = 11'b01111100101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_20;
      end
      COMP_LOOP_10_modExp_1_while_C_20 : begin
        fsm_output = 11'b01111100110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_21;
      end
      COMP_LOOP_10_modExp_1_while_C_21 : begin
        fsm_output = 11'b01111100111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_22;
      end
      COMP_LOOP_10_modExp_1_while_C_22 : begin
        fsm_output = 11'b01111101000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_23;
      end
      COMP_LOOP_10_modExp_1_while_C_23 : begin
        fsm_output = 11'b01111101001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_24;
      end
      COMP_LOOP_10_modExp_1_while_C_24 : begin
        fsm_output = 11'b01111101010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_25;
      end
      COMP_LOOP_10_modExp_1_while_C_25 : begin
        fsm_output = 11'b01111101011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_26;
      end
      COMP_LOOP_10_modExp_1_while_C_26 : begin
        fsm_output = 11'b01111101100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_27;
      end
      COMP_LOOP_10_modExp_1_while_C_27 : begin
        fsm_output = 11'b01111101101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_28;
      end
      COMP_LOOP_10_modExp_1_while_C_28 : begin
        fsm_output = 11'b01111101110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_29;
      end
      COMP_LOOP_10_modExp_1_while_C_29 : begin
        fsm_output = 11'b01111101111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_30;
      end
      COMP_LOOP_10_modExp_1_while_C_30 : begin
        fsm_output = 11'b01111110000;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_31;
      end
      COMP_LOOP_10_modExp_1_while_C_31 : begin
        fsm_output = 11'b01111110001;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_32;
      end
      COMP_LOOP_10_modExp_1_while_C_32 : begin
        fsm_output = 11'b01111110010;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_33;
      end
      COMP_LOOP_10_modExp_1_while_C_33 : begin
        fsm_output = 11'b01111110011;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_34;
      end
      COMP_LOOP_10_modExp_1_while_C_34 : begin
        fsm_output = 11'b01111110100;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_35;
      end
      COMP_LOOP_10_modExp_1_while_C_35 : begin
        fsm_output = 11'b01111110101;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_36;
      end
      COMP_LOOP_10_modExp_1_while_C_36 : begin
        fsm_output = 11'b01111110110;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_37;
      end
      COMP_LOOP_10_modExp_1_while_C_37 : begin
        fsm_output = 11'b01111110111;
        state_var_NS = COMP_LOOP_10_modExp_1_while_C_38;
      end
      COMP_LOOP_10_modExp_1_while_C_38 : begin
        fsm_output = 11'b01111111000;
        if ( COMP_LOOP_10_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_578;
        end
        else begin
          state_var_NS = COMP_LOOP_10_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_578 : begin
        fsm_output = 11'b01111111001;
        state_var_NS = COMP_LOOP_C_579;
      end
      COMP_LOOP_C_579 : begin
        fsm_output = 11'b01111111010;
        state_var_NS = COMP_LOOP_C_580;
      end
      COMP_LOOP_C_580 : begin
        fsm_output = 11'b01111111011;
        state_var_NS = COMP_LOOP_C_581;
      end
      COMP_LOOP_C_581 : begin
        fsm_output = 11'b01111111100;
        state_var_NS = COMP_LOOP_C_582;
      end
      COMP_LOOP_C_582 : begin
        fsm_output = 11'b01111111101;
        state_var_NS = COMP_LOOP_C_583;
      end
      COMP_LOOP_C_583 : begin
        fsm_output = 11'b01111111110;
        state_var_NS = COMP_LOOP_C_584;
      end
      COMP_LOOP_C_584 : begin
        fsm_output = 11'b01111111111;
        state_var_NS = COMP_LOOP_C_585;
      end
      COMP_LOOP_C_585 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = COMP_LOOP_C_586;
      end
      COMP_LOOP_C_586 : begin
        fsm_output = 11'b10000000001;
        state_var_NS = COMP_LOOP_C_587;
      end
      COMP_LOOP_C_587 : begin
        fsm_output = 11'b10000000010;
        state_var_NS = COMP_LOOP_C_588;
      end
      COMP_LOOP_C_588 : begin
        fsm_output = 11'b10000000011;
        state_var_NS = COMP_LOOP_C_589;
      end
      COMP_LOOP_C_589 : begin
        fsm_output = 11'b10000000100;
        state_var_NS = COMP_LOOP_C_590;
      end
      COMP_LOOP_C_590 : begin
        fsm_output = 11'b10000000101;
        state_var_NS = COMP_LOOP_C_591;
      end
      COMP_LOOP_C_591 : begin
        fsm_output = 11'b10000000110;
        state_var_NS = COMP_LOOP_C_592;
      end
      COMP_LOOP_C_592 : begin
        fsm_output = 11'b10000000111;
        state_var_NS = COMP_LOOP_C_593;
      end
      COMP_LOOP_C_593 : begin
        fsm_output = 11'b10000001000;
        state_var_NS = COMP_LOOP_C_594;
      end
      COMP_LOOP_C_594 : begin
        fsm_output = 11'b10000001001;
        state_var_NS = COMP_LOOP_C_595;
      end
      COMP_LOOP_C_595 : begin
        fsm_output = 11'b10000001010;
        state_var_NS = COMP_LOOP_C_596;
      end
      COMP_LOOP_C_596 : begin
        fsm_output = 11'b10000001011;
        state_var_NS = COMP_LOOP_C_597;
      end
      COMP_LOOP_C_597 : begin
        fsm_output = 11'b10000001100;
        state_var_NS = COMP_LOOP_C_598;
      end
      COMP_LOOP_C_598 : begin
        fsm_output = 11'b10000001101;
        state_var_NS = COMP_LOOP_C_599;
      end
      COMP_LOOP_C_599 : begin
        fsm_output = 11'b10000001110;
        state_var_NS = COMP_LOOP_C_600;
      end
      COMP_LOOP_C_600 : begin
        fsm_output = 11'b10000001111;
        state_var_NS = COMP_LOOP_C_601;
      end
      COMP_LOOP_C_601 : begin
        fsm_output = 11'b10000010000;
        state_var_NS = COMP_LOOP_C_602;
      end
      COMP_LOOP_C_602 : begin
        fsm_output = 11'b10000010001;
        state_var_NS = COMP_LOOP_C_603;
      end
      COMP_LOOP_C_603 : begin
        fsm_output = 11'b10000010010;
        state_var_NS = COMP_LOOP_C_604;
      end
      COMP_LOOP_C_604 : begin
        fsm_output = 11'b10000010011;
        state_var_NS = COMP_LOOP_C_605;
      end
      COMP_LOOP_C_605 : begin
        fsm_output = 11'b10000010100;
        state_var_NS = COMP_LOOP_C_606;
      end
      COMP_LOOP_C_606 : begin
        fsm_output = 11'b10000010101;
        state_var_NS = COMP_LOOP_C_607;
      end
      COMP_LOOP_C_607 : begin
        fsm_output = 11'b10000010110;
        state_var_NS = COMP_LOOP_C_608;
      end
      COMP_LOOP_C_608 : begin
        fsm_output = 11'b10000010111;
        state_var_NS = COMP_LOOP_C_609;
      end
      COMP_LOOP_C_609 : begin
        fsm_output = 11'b10000011000;
        state_var_NS = COMP_LOOP_C_610;
      end
      COMP_LOOP_C_610 : begin
        fsm_output = 11'b10000011001;
        state_var_NS = COMP_LOOP_C_611;
      end
      COMP_LOOP_C_611 : begin
        fsm_output = 11'b10000011010;
        state_var_NS = COMP_LOOP_C_612;
      end
      COMP_LOOP_C_612 : begin
        fsm_output = 11'b10000011011;
        state_var_NS = COMP_LOOP_C_613;
      end
      COMP_LOOP_C_613 : begin
        fsm_output = 11'b10000011100;
        state_var_NS = COMP_LOOP_C_614;
      end
      COMP_LOOP_C_614 : begin
        fsm_output = 11'b10000011101;
        state_var_NS = COMP_LOOP_C_615;
      end
      COMP_LOOP_C_615 : begin
        fsm_output = 11'b10000011110;
        state_var_NS = COMP_LOOP_C_616;
      end
      COMP_LOOP_C_616 : begin
        fsm_output = 11'b10000011111;
        state_var_NS = COMP_LOOP_C_617;
      end
      COMP_LOOP_C_617 : begin
        fsm_output = 11'b10000100000;
        state_var_NS = COMP_LOOP_C_618;
      end
      COMP_LOOP_C_618 : begin
        fsm_output = 11'b10000100001;
        state_var_NS = COMP_LOOP_C_619;
      end
      COMP_LOOP_C_619 : begin
        fsm_output = 11'b10000100010;
        state_var_NS = COMP_LOOP_C_620;
      end
      COMP_LOOP_C_620 : begin
        fsm_output = 11'b10000100011;
        state_var_NS = COMP_LOOP_C_621;
      end
      COMP_LOOP_C_621 : begin
        fsm_output = 11'b10000100100;
        state_var_NS = COMP_LOOP_C_622;
      end
      COMP_LOOP_C_622 : begin
        fsm_output = 11'b10000100101;
        state_var_NS = COMP_LOOP_C_623;
      end
      COMP_LOOP_C_623 : begin
        fsm_output = 11'b10000100110;
        state_var_NS = COMP_LOOP_C_624;
      end
      COMP_LOOP_C_624 : begin
        fsm_output = 11'b10000100111;
        state_var_NS = COMP_LOOP_C_625;
      end
      COMP_LOOP_C_625 : begin
        fsm_output = 11'b10000101000;
        state_var_NS = COMP_LOOP_C_626;
      end
      COMP_LOOP_C_626 : begin
        fsm_output = 11'b10000101001;
        state_var_NS = COMP_LOOP_C_627;
      end
      COMP_LOOP_C_627 : begin
        fsm_output = 11'b10000101010;
        state_var_NS = COMP_LOOP_C_628;
      end
      COMP_LOOP_C_628 : begin
        fsm_output = 11'b10000101011;
        state_var_NS = COMP_LOOP_C_629;
      end
      COMP_LOOP_C_629 : begin
        fsm_output = 11'b10000101100;
        state_var_NS = COMP_LOOP_C_630;
      end
      COMP_LOOP_C_630 : begin
        fsm_output = 11'b10000101101;
        state_var_NS = COMP_LOOP_C_631;
      end
      COMP_LOOP_C_631 : begin
        fsm_output = 11'b10000101110;
        state_var_NS = COMP_LOOP_C_632;
      end
      COMP_LOOP_C_632 : begin
        fsm_output = 11'b10000101111;
        state_var_NS = COMP_LOOP_C_633;
      end
      COMP_LOOP_C_633 : begin
        fsm_output = 11'b10000110000;
        state_var_NS = COMP_LOOP_C_634;
      end
      COMP_LOOP_C_634 : begin
        fsm_output = 11'b10000110001;
        state_var_NS = COMP_LOOP_C_635;
      end
      COMP_LOOP_C_635 : begin
        fsm_output = 11'b10000110010;
        state_var_NS = COMP_LOOP_C_636;
      end
      COMP_LOOP_C_636 : begin
        fsm_output = 11'b10000110011;
        state_var_NS = COMP_LOOP_C_637;
      end
      COMP_LOOP_C_637 : begin
        fsm_output = 11'b10000110100;
        state_var_NS = COMP_LOOP_C_638;
      end
      COMP_LOOP_C_638 : begin
        fsm_output = 11'b10000110101;
        state_var_NS = COMP_LOOP_C_639;
      end
      COMP_LOOP_C_639 : begin
        fsm_output = 11'b10000110110;
        state_var_NS = COMP_LOOP_C_640;
      end
      COMP_LOOP_C_640 : begin
        fsm_output = 11'b10000110111;
        if ( COMP_LOOP_C_640_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_641;
        end
      end
      COMP_LOOP_C_641 : begin
        fsm_output = 11'b10000111000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_0;
      end
      COMP_LOOP_11_modExp_1_while_C_0 : begin
        fsm_output = 11'b10000111001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_1;
      end
      COMP_LOOP_11_modExp_1_while_C_1 : begin
        fsm_output = 11'b10000111010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_2;
      end
      COMP_LOOP_11_modExp_1_while_C_2 : begin
        fsm_output = 11'b10000111011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_3;
      end
      COMP_LOOP_11_modExp_1_while_C_3 : begin
        fsm_output = 11'b10000111100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_4;
      end
      COMP_LOOP_11_modExp_1_while_C_4 : begin
        fsm_output = 11'b10000111101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_5;
      end
      COMP_LOOP_11_modExp_1_while_C_5 : begin
        fsm_output = 11'b10000111110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_6;
      end
      COMP_LOOP_11_modExp_1_while_C_6 : begin
        fsm_output = 11'b10000111111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_7;
      end
      COMP_LOOP_11_modExp_1_while_C_7 : begin
        fsm_output = 11'b10001000000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_8;
      end
      COMP_LOOP_11_modExp_1_while_C_8 : begin
        fsm_output = 11'b10001000001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_9;
      end
      COMP_LOOP_11_modExp_1_while_C_9 : begin
        fsm_output = 11'b10001000010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_10;
      end
      COMP_LOOP_11_modExp_1_while_C_10 : begin
        fsm_output = 11'b10001000011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_11;
      end
      COMP_LOOP_11_modExp_1_while_C_11 : begin
        fsm_output = 11'b10001000100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_12;
      end
      COMP_LOOP_11_modExp_1_while_C_12 : begin
        fsm_output = 11'b10001000101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_13;
      end
      COMP_LOOP_11_modExp_1_while_C_13 : begin
        fsm_output = 11'b10001000110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_14;
      end
      COMP_LOOP_11_modExp_1_while_C_14 : begin
        fsm_output = 11'b10001000111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_15;
      end
      COMP_LOOP_11_modExp_1_while_C_15 : begin
        fsm_output = 11'b10001001000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_16;
      end
      COMP_LOOP_11_modExp_1_while_C_16 : begin
        fsm_output = 11'b10001001001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_17;
      end
      COMP_LOOP_11_modExp_1_while_C_17 : begin
        fsm_output = 11'b10001001010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_18;
      end
      COMP_LOOP_11_modExp_1_while_C_18 : begin
        fsm_output = 11'b10001001011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_19;
      end
      COMP_LOOP_11_modExp_1_while_C_19 : begin
        fsm_output = 11'b10001001100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_20;
      end
      COMP_LOOP_11_modExp_1_while_C_20 : begin
        fsm_output = 11'b10001001101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_21;
      end
      COMP_LOOP_11_modExp_1_while_C_21 : begin
        fsm_output = 11'b10001001110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_22;
      end
      COMP_LOOP_11_modExp_1_while_C_22 : begin
        fsm_output = 11'b10001001111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_23;
      end
      COMP_LOOP_11_modExp_1_while_C_23 : begin
        fsm_output = 11'b10001010000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_24;
      end
      COMP_LOOP_11_modExp_1_while_C_24 : begin
        fsm_output = 11'b10001010001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_25;
      end
      COMP_LOOP_11_modExp_1_while_C_25 : begin
        fsm_output = 11'b10001010010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_26;
      end
      COMP_LOOP_11_modExp_1_while_C_26 : begin
        fsm_output = 11'b10001010011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_27;
      end
      COMP_LOOP_11_modExp_1_while_C_27 : begin
        fsm_output = 11'b10001010100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_28;
      end
      COMP_LOOP_11_modExp_1_while_C_28 : begin
        fsm_output = 11'b10001010101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_29;
      end
      COMP_LOOP_11_modExp_1_while_C_29 : begin
        fsm_output = 11'b10001010110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_30;
      end
      COMP_LOOP_11_modExp_1_while_C_30 : begin
        fsm_output = 11'b10001010111;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_31;
      end
      COMP_LOOP_11_modExp_1_while_C_31 : begin
        fsm_output = 11'b10001011000;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_32;
      end
      COMP_LOOP_11_modExp_1_while_C_32 : begin
        fsm_output = 11'b10001011001;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_33;
      end
      COMP_LOOP_11_modExp_1_while_C_33 : begin
        fsm_output = 11'b10001011010;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_34;
      end
      COMP_LOOP_11_modExp_1_while_C_34 : begin
        fsm_output = 11'b10001011011;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_35;
      end
      COMP_LOOP_11_modExp_1_while_C_35 : begin
        fsm_output = 11'b10001011100;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_36;
      end
      COMP_LOOP_11_modExp_1_while_C_36 : begin
        fsm_output = 11'b10001011101;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_37;
      end
      COMP_LOOP_11_modExp_1_while_C_37 : begin
        fsm_output = 11'b10001011110;
        state_var_NS = COMP_LOOP_11_modExp_1_while_C_38;
      end
      COMP_LOOP_11_modExp_1_while_C_38 : begin
        fsm_output = 11'b10001011111;
        if ( COMP_LOOP_11_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_642;
        end
        else begin
          state_var_NS = COMP_LOOP_11_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_642 : begin
        fsm_output = 11'b10001100000;
        state_var_NS = COMP_LOOP_C_643;
      end
      COMP_LOOP_C_643 : begin
        fsm_output = 11'b10001100001;
        state_var_NS = COMP_LOOP_C_644;
      end
      COMP_LOOP_C_644 : begin
        fsm_output = 11'b10001100010;
        state_var_NS = COMP_LOOP_C_645;
      end
      COMP_LOOP_C_645 : begin
        fsm_output = 11'b10001100011;
        state_var_NS = COMP_LOOP_C_646;
      end
      COMP_LOOP_C_646 : begin
        fsm_output = 11'b10001100100;
        state_var_NS = COMP_LOOP_C_647;
      end
      COMP_LOOP_C_647 : begin
        fsm_output = 11'b10001100101;
        state_var_NS = COMP_LOOP_C_648;
      end
      COMP_LOOP_C_648 : begin
        fsm_output = 11'b10001100110;
        state_var_NS = COMP_LOOP_C_649;
      end
      COMP_LOOP_C_649 : begin
        fsm_output = 11'b10001100111;
        state_var_NS = COMP_LOOP_C_650;
      end
      COMP_LOOP_C_650 : begin
        fsm_output = 11'b10001101000;
        state_var_NS = COMP_LOOP_C_651;
      end
      COMP_LOOP_C_651 : begin
        fsm_output = 11'b10001101001;
        state_var_NS = COMP_LOOP_C_652;
      end
      COMP_LOOP_C_652 : begin
        fsm_output = 11'b10001101010;
        state_var_NS = COMP_LOOP_C_653;
      end
      COMP_LOOP_C_653 : begin
        fsm_output = 11'b10001101011;
        state_var_NS = COMP_LOOP_C_654;
      end
      COMP_LOOP_C_654 : begin
        fsm_output = 11'b10001101100;
        state_var_NS = COMP_LOOP_C_655;
      end
      COMP_LOOP_C_655 : begin
        fsm_output = 11'b10001101101;
        state_var_NS = COMP_LOOP_C_656;
      end
      COMP_LOOP_C_656 : begin
        fsm_output = 11'b10001101110;
        state_var_NS = COMP_LOOP_C_657;
      end
      COMP_LOOP_C_657 : begin
        fsm_output = 11'b10001101111;
        state_var_NS = COMP_LOOP_C_658;
      end
      COMP_LOOP_C_658 : begin
        fsm_output = 11'b10001110000;
        state_var_NS = COMP_LOOP_C_659;
      end
      COMP_LOOP_C_659 : begin
        fsm_output = 11'b10001110001;
        state_var_NS = COMP_LOOP_C_660;
      end
      COMP_LOOP_C_660 : begin
        fsm_output = 11'b10001110010;
        state_var_NS = COMP_LOOP_C_661;
      end
      COMP_LOOP_C_661 : begin
        fsm_output = 11'b10001110011;
        state_var_NS = COMP_LOOP_C_662;
      end
      COMP_LOOP_C_662 : begin
        fsm_output = 11'b10001110100;
        state_var_NS = COMP_LOOP_C_663;
      end
      COMP_LOOP_C_663 : begin
        fsm_output = 11'b10001110101;
        state_var_NS = COMP_LOOP_C_664;
      end
      COMP_LOOP_C_664 : begin
        fsm_output = 11'b10001110110;
        state_var_NS = COMP_LOOP_C_665;
      end
      COMP_LOOP_C_665 : begin
        fsm_output = 11'b10001110111;
        state_var_NS = COMP_LOOP_C_666;
      end
      COMP_LOOP_C_666 : begin
        fsm_output = 11'b10001111000;
        state_var_NS = COMP_LOOP_C_667;
      end
      COMP_LOOP_C_667 : begin
        fsm_output = 11'b10001111001;
        state_var_NS = COMP_LOOP_C_668;
      end
      COMP_LOOP_C_668 : begin
        fsm_output = 11'b10001111010;
        state_var_NS = COMP_LOOP_C_669;
      end
      COMP_LOOP_C_669 : begin
        fsm_output = 11'b10001111011;
        state_var_NS = COMP_LOOP_C_670;
      end
      COMP_LOOP_C_670 : begin
        fsm_output = 11'b10001111100;
        state_var_NS = COMP_LOOP_C_671;
      end
      COMP_LOOP_C_671 : begin
        fsm_output = 11'b10001111101;
        state_var_NS = COMP_LOOP_C_672;
      end
      COMP_LOOP_C_672 : begin
        fsm_output = 11'b10001111110;
        state_var_NS = COMP_LOOP_C_673;
      end
      COMP_LOOP_C_673 : begin
        fsm_output = 11'b10001111111;
        state_var_NS = COMP_LOOP_C_674;
      end
      COMP_LOOP_C_674 : begin
        fsm_output = 11'b10010000000;
        state_var_NS = COMP_LOOP_C_675;
      end
      COMP_LOOP_C_675 : begin
        fsm_output = 11'b10010000001;
        state_var_NS = COMP_LOOP_C_676;
      end
      COMP_LOOP_C_676 : begin
        fsm_output = 11'b10010000010;
        state_var_NS = COMP_LOOP_C_677;
      end
      COMP_LOOP_C_677 : begin
        fsm_output = 11'b10010000011;
        state_var_NS = COMP_LOOP_C_678;
      end
      COMP_LOOP_C_678 : begin
        fsm_output = 11'b10010000100;
        state_var_NS = COMP_LOOP_C_679;
      end
      COMP_LOOP_C_679 : begin
        fsm_output = 11'b10010000101;
        state_var_NS = COMP_LOOP_C_680;
      end
      COMP_LOOP_C_680 : begin
        fsm_output = 11'b10010000110;
        state_var_NS = COMP_LOOP_C_681;
      end
      COMP_LOOP_C_681 : begin
        fsm_output = 11'b10010000111;
        state_var_NS = COMP_LOOP_C_682;
      end
      COMP_LOOP_C_682 : begin
        fsm_output = 11'b10010001000;
        state_var_NS = COMP_LOOP_C_683;
      end
      COMP_LOOP_C_683 : begin
        fsm_output = 11'b10010001001;
        state_var_NS = COMP_LOOP_C_684;
      end
      COMP_LOOP_C_684 : begin
        fsm_output = 11'b10010001010;
        state_var_NS = COMP_LOOP_C_685;
      end
      COMP_LOOP_C_685 : begin
        fsm_output = 11'b10010001011;
        state_var_NS = COMP_LOOP_C_686;
      end
      COMP_LOOP_C_686 : begin
        fsm_output = 11'b10010001100;
        state_var_NS = COMP_LOOP_C_687;
      end
      COMP_LOOP_C_687 : begin
        fsm_output = 11'b10010001101;
        state_var_NS = COMP_LOOP_C_688;
      end
      COMP_LOOP_C_688 : begin
        fsm_output = 11'b10010001110;
        state_var_NS = COMP_LOOP_C_689;
      end
      COMP_LOOP_C_689 : begin
        fsm_output = 11'b10010001111;
        state_var_NS = COMP_LOOP_C_690;
      end
      COMP_LOOP_C_690 : begin
        fsm_output = 11'b10010010000;
        state_var_NS = COMP_LOOP_C_691;
      end
      COMP_LOOP_C_691 : begin
        fsm_output = 11'b10010010001;
        state_var_NS = COMP_LOOP_C_692;
      end
      COMP_LOOP_C_692 : begin
        fsm_output = 11'b10010010010;
        state_var_NS = COMP_LOOP_C_693;
      end
      COMP_LOOP_C_693 : begin
        fsm_output = 11'b10010010011;
        state_var_NS = COMP_LOOP_C_694;
      end
      COMP_LOOP_C_694 : begin
        fsm_output = 11'b10010010100;
        state_var_NS = COMP_LOOP_C_695;
      end
      COMP_LOOP_C_695 : begin
        fsm_output = 11'b10010010101;
        state_var_NS = COMP_LOOP_C_696;
      end
      COMP_LOOP_C_696 : begin
        fsm_output = 11'b10010010110;
        state_var_NS = COMP_LOOP_C_697;
      end
      COMP_LOOP_C_697 : begin
        fsm_output = 11'b10010010111;
        state_var_NS = COMP_LOOP_C_698;
      end
      COMP_LOOP_C_698 : begin
        fsm_output = 11'b10010011000;
        state_var_NS = COMP_LOOP_C_699;
      end
      COMP_LOOP_C_699 : begin
        fsm_output = 11'b10010011001;
        state_var_NS = COMP_LOOP_C_700;
      end
      COMP_LOOP_C_700 : begin
        fsm_output = 11'b10010011010;
        state_var_NS = COMP_LOOP_C_701;
      end
      COMP_LOOP_C_701 : begin
        fsm_output = 11'b10010011011;
        state_var_NS = COMP_LOOP_C_702;
      end
      COMP_LOOP_C_702 : begin
        fsm_output = 11'b10010011100;
        state_var_NS = COMP_LOOP_C_703;
      end
      COMP_LOOP_C_703 : begin
        fsm_output = 11'b10010011101;
        state_var_NS = COMP_LOOP_C_704;
      end
      COMP_LOOP_C_704 : begin
        fsm_output = 11'b10010011110;
        if ( COMP_LOOP_C_704_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_705;
        end
      end
      COMP_LOOP_C_705 : begin
        fsm_output = 11'b10010011111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_0;
      end
      COMP_LOOP_12_modExp_1_while_C_0 : begin
        fsm_output = 11'b10010100000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_1;
      end
      COMP_LOOP_12_modExp_1_while_C_1 : begin
        fsm_output = 11'b10010100001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_2;
      end
      COMP_LOOP_12_modExp_1_while_C_2 : begin
        fsm_output = 11'b10010100010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_3;
      end
      COMP_LOOP_12_modExp_1_while_C_3 : begin
        fsm_output = 11'b10010100011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_4;
      end
      COMP_LOOP_12_modExp_1_while_C_4 : begin
        fsm_output = 11'b10010100100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_5;
      end
      COMP_LOOP_12_modExp_1_while_C_5 : begin
        fsm_output = 11'b10010100101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_6;
      end
      COMP_LOOP_12_modExp_1_while_C_6 : begin
        fsm_output = 11'b10010100110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_7;
      end
      COMP_LOOP_12_modExp_1_while_C_7 : begin
        fsm_output = 11'b10010100111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_8;
      end
      COMP_LOOP_12_modExp_1_while_C_8 : begin
        fsm_output = 11'b10010101000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_9;
      end
      COMP_LOOP_12_modExp_1_while_C_9 : begin
        fsm_output = 11'b10010101001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_10;
      end
      COMP_LOOP_12_modExp_1_while_C_10 : begin
        fsm_output = 11'b10010101010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_11;
      end
      COMP_LOOP_12_modExp_1_while_C_11 : begin
        fsm_output = 11'b10010101011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_12;
      end
      COMP_LOOP_12_modExp_1_while_C_12 : begin
        fsm_output = 11'b10010101100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_13;
      end
      COMP_LOOP_12_modExp_1_while_C_13 : begin
        fsm_output = 11'b10010101101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_14;
      end
      COMP_LOOP_12_modExp_1_while_C_14 : begin
        fsm_output = 11'b10010101110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_15;
      end
      COMP_LOOP_12_modExp_1_while_C_15 : begin
        fsm_output = 11'b10010101111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_16;
      end
      COMP_LOOP_12_modExp_1_while_C_16 : begin
        fsm_output = 11'b10010110000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_17;
      end
      COMP_LOOP_12_modExp_1_while_C_17 : begin
        fsm_output = 11'b10010110001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_18;
      end
      COMP_LOOP_12_modExp_1_while_C_18 : begin
        fsm_output = 11'b10010110010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_19;
      end
      COMP_LOOP_12_modExp_1_while_C_19 : begin
        fsm_output = 11'b10010110011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_20;
      end
      COMP_LOOP_12_modExp_1_while_C_20 : begin
        fsm_output = 11'b10010110100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_21;
      end
      COMP_LOOP_12_modExp_1_while_C_21 : begin
        fsm_output = 11'b10010110101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_22;
      end
      COMP_LOOP_12_modExp_1_while_C_22 : begin
        fsm_output = 11'b10010110110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_23;
      end
      COMP_LOOP_12_modExp_1_while_C_23 : begin
        fsm_output = 11'b10010110111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_24;
      end
      COMP_LOOP_12_modExp_1_while_C_24 : begin
        fsm_output = 11'b10010111000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_25;
      end
      COMP_LOOP_12_modExp_1_while_C_25 : begin
        fsm_output = 11'b10010111001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_26;
      end
      COMP_LOOP_12_modExp_1_while_C_26 : begin
        fsm_output = 11'b10010111010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_27;
      end
      COMP_LOOP_12_modExp_1_while_C_27 : begin
        fsm_output = 11'b10010111011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_28;
      end
      COMP_LOOP_12_modExp_1_while_C_28 : begin
        fsm_output = 11'b10010111100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_29;
      end
      COMP_LOOP_12_modExp_1_while_C_29 : begin
        fsm_output = 11'b10010111101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_30;
      end
      COMP_LOOP_12_modExp_1_while_C_30 : begin
        fsm_output = 11'b10010111110;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_31;
      end
      COMP_LOOP_12_modExp_1_while_C_31 : begin
        fsm_output = 11'b10010111111;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_32;
      end
      COMP_LOOP_12_modExp_1_while_C_32 : begin
        fsm_output = 11'b10011000000;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_33;
      end
      COMP_LOOP_12_modExp_1_while_C_33 : begin
        fsm_output = 11'b10011000001;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_34;
      end
      COMP_LOOP_12_modExp_1_while_C_34 : begin
        fsm_output = 11'b10011000010;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_35;
      end
      COMP_LOOP_12_modExp_1_while_C_35 : begin
        fsm_output = 11'b10011000011;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_36;
      end
      COMP_LOOP_12_modExp_1_while_C_36 : begin
        fsm_output = 11'b10011000100;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_37;
      end
      COMP_LOOP_12_modExp_1_while_C_37 : begin
        fsm_output = 11'b10011000101;
        state_var_NS = COMP_LOOP_12_modExp_1_while_C_38;
      end
      COMP_LOOP_12_modExp_1_while_C_38 : begin
        fsm_output = 11'b10011000110;
        if ( COMP_LOOP_12_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_706;
        end
        else begin
          state_var_NS = COMP_LOOP_12_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_706 : begin
        fsm_output = 11'b10011000111;
        state_var_NS = COMP_LOOP_C_707;
      end
      COMP_LOOP_C_707 : begin
        fsm_output = 11'b10011001000;
        state_var_NS = COMP_LOOP_C_708;
      end
      COMP_LOOP_C_708 : begin
        fsm_output = 11'b10011001001;
        state_var_NS = COMP_LOOP_C_709;
      end
      COMP_LOOP_C_709 : begin
        fsm_output = 11'b10011001010;
        state_var_NS = COMP_LOOP_C_710;
      end
      COMP_LOOP_C_710 : begin
        fsm_output = 11'b10011001011;
        state_var_NS = COMP_LOOP_C_711;
      end
      COMP_LOOP_C_711 : begin
        fsm_output = 11'b10011001100;
        state_var_NS = COMP_LOOP_C_712;
      end
      COMP_LOOP_C_712 : begin
        fsm_output = 11'b10011001101;
        state_var_NS = COMP_LOOP_C_713;
      end
      COMP_LOOP_C_713 : begin
        fsm_output = 11'b10011001110;
        state_var_NS = COMP_LOOP_C_714;
      end
      COMP_LOOP_C_714 : begin
        fsm_output = 11'b10011001111;
        state_var_NS = COMP_LOOP_C_715;
      end
      COMP_LOOP_C_715 : begin
        fsm_output = 11'b10011010000;
        state_var_NS = COMP_LOOP_C_716;
      end
      COMP_LOOP_C_716 : begin
        fsm_output = 11'b10011010001;
        state_var_NS = COMP_LOOP_C_717;
      end
      COMP_LOOP_C_717 : begin
        fsm_output = 11'b10011010010;
        state_var_NS = COMP_LOOP_C_718;
      end
      COMP_LOOP_C_718 : begin
        fsm_output = 11'b10011010011;
        state_var_NS = COMP_LOOP_C_719;
      end
      COMP_LOOP_C_719 : begin
        fsm_output = 11'b10011010100;
        state_var_NS = COMP_LOOP_C_720;
      end
      COMP_LOOP_C_720 : begin
        fsm_output = 11'b10011010101;
        state_var_NS = COMP_LOOP_C_721;
      end
      COMP_LOOP_C_721 : begin
        fsm_output = 11'b10011010110;
        state_var_NS = COMP_LOOP_C_722;
      end
      COMP_LOOP_C_722 : begin
        fsm_output = 11'b10011010111;
        state_var_NS = COMP_LOOP_C_723;
      end
      COMP_LOOP_C_723 : begin
        fsm_output = 11'b10011011000;
        state_var_NS = COMP_LOOP_C_724;
      end
      COMP_LOOP_C_724 : begin
        fsm_output = 11'b10011011001;
        state_var_NS = COMP_LOOP_C_725;
      end
      COMP_LOOP_C_725 : begin
        fsm_output = 11'b10011011010;
        state_var_NS = COMP_LOOP_C_726;
      end
      COMP_LOOP_C_726 : begin
        fsm_output = 11'b10011011011;
        state_var_NS = COMP_LOOP_C_727;
      end
      COMP_LOOP_C_727 : begin
        fsm_output = 11'b10011011100;
        state_var_NS = COMP_LOOP_C_728;
      end
      COMP_LOOP_C_728 : begin
        fsm_output = 11'b10011011101;
        state_var_NS = COMP_LOOP_C_729;
      end
      COMP_LOOP_C_729 : begin
        fsm_output = 11'b10011011110;
        state_var_NS = COMP_LOOP_C_730;
      end
      COMP_LOOP_C_730 : begin
        fsm_output = 11'b10011011111;
        state_var_NS = COMP_LOOP_C_731;
      end
      COMP_LOOP_C_731 : begin
        fsm_output = 11'b10011100000;
        state_var_NS = COMP_LOOP_C_732;
      end
      COMP_LOOP_C_732 : begin
        fsm_output = 11'b10011100001;
        state_var_NS = COMP_LOOP_C_733;
      end
      COMP_LOOP_C_733 : begin
        fsm_output = 11'b10011100010;
        state_var_NS = COMP_LOOP_C_734;
      end
      COMP_LOOP_C_734 : begin
        fsm_output = 11'b10011100011;
        state_var_NS = COMP_LOOP_C_735;
      end
      COMP_LOOP_C_735 : begin
        fsm_output = 11'b10011100100;
        state_var_NS = COMP_LOOP_C_736;
      end
      COMP_LOOP_C_736 : begin
        fsm_output = 11'b10011100101;
        state_var_NS = COMP_LOOP_C_737;
      end
      COMP_LOOP_C_737 : begin
        fsm_output = 11'b10011100110;
        state_var_NS = COMP_LOOP_C_738;
      end
      COMP_LOOP_C_738 : begin
        fsm_output = 11'b10011100111;
        state_var_NS = COMP_LOOP_C_739;
      end
      COMP_LOOP_C_739 : begin
        fsm_output = 11'b10011101000;
        state_var_NS = COMP_LOOP_C_740;
      end
      COMP_LOOP_C_740 : begin
        fsm_output = 11'b10011101001;
        state_var_NS = COMP_LOOP_C_741;
      end
      COMP_LOOP_C_741 : begin
        fsm_output = 11'b10011101010;
        state_var_NS = COMP_LOOP_C_742;
      end
      COMP_LOOP_C_742 : begin
        fsm_output = 11'b10011101011;
        state_var_NS = COMP_LOOP_C_743;
      end
      COMP_LOOP_C_743 : begin
        fsm_output = 11'b10011101100;
        state_var_NS = COMP_LOOP_C_744;
      end
      COMP_LOOP_C_744 : begin
        fsm_output = 11'b10011101101;
        state_var_NS = COMP_LOOP_C_745;
      end
      COMP_LOOP_C_745 : begin
        fsm_output = 11'b10011101110;
        state_var_NS = COMP_LOOP_C_746;
      end
      COMP_LOOP_C_746 : begin
        fsm_output = 11'b10011101111;
        state_var_NS = COMP_LOOP_C_747;
      end
      COMP_LOOP_C_747 : begin
        fsm_output = 11'b10011110000;
        state_var_NS = COMP_LOOP_C_748;
      end
      COMP_LOOP_C_748 : begin
        fsm_output = 11'b10011110001;
        state_var_NS = COMP_LOOP_C_749;
      end
      COMP_LOOP_C_749 : begin
        fsm_output = 11'b10011110010;
        state_var_NS = COMP_LOOP_C_750;
      end
      COMP_LOOP_C_750 : begin
        fsm_output = 11'b10011110011;
        state_var_NS = COMP_LOOP_C_751;
      end
      COMP_LOOP_C_751 : begin
        fsm_output = 11'b10011110100;
        state_var_NS = COMP_LOOP_C_752;
      end
      COMP_LOOP_C_752 : begin
        fsm_output = 11'b10011110101;
        state_var_NS = COMP_LOOP_C_753;
      end
      COMP_LOOP_C_753 : begin
        fsm_output = 11'b10011110110;
        state_var_NS = COMP_LOOP_C_754;
      end
      COMP_LOOP_C_754 : begin
        fsm_output = 11'b10011110111;
        state_var_NS = COMP_LOOP_C_755;
      end
      COMP_LOOP_C_755 : begin
        fsm_output = 11'b10011111000;
        state_var_NS = COMP_LOOP_C_756;
      end
      COMP_LOOP_C_756 : begin
        fsm_output = 11'b10011111001;
        state_var_NS = COMP_LOOP_C_757;
      end
      COMP_LOOP_C_757 : begin
        fsm_output = 11'b10011111010;
        state_var_NS = COMP_LOOP_C_758;
      end
      COMP_LOOP_C_758 : begin
        fsm_output = 11'b10011111011;
        state_var_NS = COMP_LOOP_C_759;
      end
      COMP_LOOP_C_759 : begin
        fsm_output = 11'b10011111100;
        state_var_NS = COMP_LOOP_C_760;
      end
      COMP_LOOP_C_760 : begin
        fsm_output = 11'b10011111101;
        state_var_NS = COMP_LOOP_C_761;
      end
      COMP_LOOP_C_761 : begin
        fsm_output = 11'b10011111110;
        state_var_NS = COMP_LOOP_C_762;
      end
      COMP_LOOP_C_762 : begin
        fsm_output = 11'b10011111111;
        state_var_NS = COMP_LOOP_C_763;
      end
      COMP_LOOP_C_763 : begin
        fsm_output = 11'b10100000000;
        state_var_NS = COMP_LOOP_C_764;
      end
      COMP_LOOP_C_764 : begin
        fsm_output = 11'b10100000001;
        state_var_NS = COMP_LOOP_C_765;
      end
      COMP_LOOP_C_765 : begin
        fsm_output = 11'b10100000010;
        state_var_NS = COMP_LOOP_C_766;
      end
      COMP_LOOP_C_766 : begin
        fsm_output = 11'b10100000011;
        state_var_NS = COMP_LOOP_C_767;
      end
      COMP_LOOP_C_767 : begin
        fsm_output = 11'b10100000100;
        state_var_NS = COMP_LOOP_C_768;
      end
      COMP_LOOP_C_768 : begin
        fsm_output = 11'b10100000101;
        if ( COMP_LOOP_C_768_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_769;
        end
      end
      COMP_LOOP_C_769 : begin
        fsm_output = 11'b10100000110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_0;
      end
      COMP_LOOP_13_modExp_1_while_C_0 : begin
        fsm_output = 11'b10100000111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_1;
      end
      COMP_LOOP_13_modExp_1_while_C_1 : begin
        fsm_output = 11'b10100001000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_2;
      end
      COMP_LOOP_13_modExp_1_while_C_2 : begin
        fsm_output = 11'b10100001001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_3;
      end
      COMP_LOOP_13_modExp_1_while_C_3 : begin
        fsm_output = 11'b10100001010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_4;
      end
      COMP_LOOP_13_modExp_1_while_C_4 : begin
        fsm_output = 11'b10100001011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_5;
      end
      COMP_LOOP_13_modExp_1_while_C_5 : begin
        fsm_output = 11'b10100001100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_6;
      end
      COMP_LOOP_13_modExp_1_while_C_6 : begin
        fsm_output = 11'b10100001101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_7;
      end
      COMP_LOOP_13_modExp_1_while_C_7 : begin
        fsm_output = 11'b10100001110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_8;
      end
      COMP_LOOP_13_modExp_1_while_C_8 : begin
        fsm_output = 11'b10100001111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_9;
      end
      COMP_LOOP_13_modExp_1_while_C_9 : begin
        fsm_output = 11'b10100010000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_10;
      end
      COMP_LOOP_13_modExp_1_while_C_10 : begin
        fsm_output = 11'b10100010001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_11;
      end
      COMP_LOOP_13_modExp_1_while_C_11 : begin
        fsm_output = 11'b10100010010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_12;
      end
      COMP_LOOP_13_modExp_1_while_C_12 : begin
        fsm_output = 11'b10100010011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_13;
      end
      COMP_LOOP_13_modExp_1_while_C_13 : begin
        fsm_output = 11'b10100010100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_14;
      end
      COMP_LOOP_13_modExp_1_while_C_14 : begin
        fsm_output = 11'b10100010101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_15;
      end
      COMP_LOOP_13_modExp_1_while_C_15 : begin
        fsm_output = 11'b10100010110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_16;
      end
      COMP_LOOP_13_modExp_1_while_C_16 : begin
        fsm_output = 11'b10100010111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_17;
      end
      COMP_LOOP_13_modExp_1_while_C_17 : begin
        fsm_output = 11'b10100011000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_18;
      end
      COMP_LOOP_13_modExp_1_while_C_18 : begin
        fsm_output = 11'b10100011001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_19;
      end
      COMP_LOOP_13_modExp_1_while_C_19 : begin
        fsm_output = 11'b10100011010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_20;
      end
      COMP_LOOP_13_modExp_1_while_C_20 : begin
        fsm_output = 11'b10100011011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_21;
      end
      COMP_LOOP_13_modExp_1_while_C_21 : begin
        fsm_output = 11'b10100011100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_22;
      end
      COMP_LOOP_13_modExp_1_while_C_22 : begin
        fsm_output = 11'b10100011101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_23;
      end
      COMP_LOOP_13_modExp_1_while_C_23 : begin
        fsm_output = 11'b10100011110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_24;
      end
      COMP_LOOP_13_modExp_1_while_C_24 : begin
        fsm_output = 11'b10100011111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_25;
      end
      COMP_LOOP_13_modExp_1_while_C_25 : begin
        fsm_output = 11'b10100100000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_26;
      end
      COMP_LOOP_13_modExp_1_while_C_26 : begin
        fsm_output = 11'b10100100001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_27;
      end
      COMP_LOOP_13_modExp_1_while_C_27 : begin
        fsm_output = 11'b10100100010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_28;
      end
      COMP_LOOP_13_modExp_1_while_C_28 : begin
        fsm_output = 11'b10100100011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_29;
      end
      COMP_LOOP_13_modExp_1_while_C_29 : begin
        fsm_output = 11'b10100100100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_30;
      end
      COMP_LOOP_13_modExp_1_while_C_30 : begin
        fsm_output = 11'b10100100101;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_31;
      end
      COMP_LOOP_13_modExp_1_while_C_31 : begin
        fsm_output = 11'b10100100110;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_32;
      end
      COMP_LOOP_13_modExp_1_while_C_32 : begin
        fsm_output = 11'b10100100111;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_33;
      end
      COMP_LOOP_13_modExp_1_while_C_33 : begin
        fsm_output = 11'b10100101000;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_34;
      end
      COMP_LOOP_13_modExp_1_while_C_34 : begin
        fsm_output = 11'b10100101001;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_35;
      end
      COMP_LOOP_13_modExp_1_while_C_35 : begin
        fsm_output = 11'b10100101010;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_36;
      end
      COMP_LOOP_13_modExp_1_while_C_36 : begin
        fsm_output = 11'b10100101011;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_37;
      end
      COMP_LOOP_13_modExp_1_while_C_37 : begin
        fsm_output = 11'b10100101100;
        state_var_NS = COMP_LOOP_13_modExp_1_while_C_38;
      end
      COMP_LOOP_13_modExp_1_while_C_38 : begin
        fsm_output = 11'b10100101101;
        if ( COMP_LOOP_13_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_770;
        end
        else begin
          state_var_NS = COMP_LOOP_13_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_770 : begin
        fsm_output = 11'b10100101110;
        state_var_NS = COMP_LOOP_C_771;
      end
      COMP_LOOP_C_771 : begin
        fsm_output = 11'b10100101111;
        state_var_NS = COMP_LOOP_C_772;
      end
      COMP_LOOP_C_772 : begin
        fsm_output = 11'b10100110000;
        state_var_NS = COMP_LOOP_C_773;
      end
      COMP_LOOP_C_773 : begin
        fsm_output = 11'b10100110001;
        state_var_NS = COMP_LOOP_C_774;
      end
      COMP_LOOP_C_774 : begin
        fsm_output = 11'b10100110010;
        state_var_NS = COMP_LOOP_C_775;
      end
      COMP_LOOP_C_775 : begin
        fsm_output = 11'b10100110011;
        state_var_NS = COMP_LOOP_C_776;
      end
      COMP_LOOP_C_776 : begin
        fsm_output = 11'b10100110100;
        state_var_NS = COMP_LOOP_C_777;
      end
      COMP_LOOP_C_777 : begin
        fsm_output = 11'b10100110101;
        state_var_NS = COMP_LOOP_C_778;
      end
      COMP_LOOP_C_778 : begin
        fsm_output = 11'b10100110110;
        state_var_NS = COMP_LOOP_C_779;
      end
      COMP_LOOP_C_779 : begin
        fsm_output = 11'b10100110111;
        state_var_NS = COMP_LOOP_C_780;
      end
      COMP_LOOP_C_780 : begin
        fsm_output = 11'b10100111000;
        state_var_NS = COMP_LOOP_C_781;
      end
      COMP_LOOP_C_781 : begin
        fsm_output = 11'b10100111001;
        state_var_NS = COMP_LOOP_C_782;
      end
      COMP_LOOP_C_782 : begin
        fsm_output = 11'b10100111010;
        state_var_NS = COMP_LOOP_C_783;
      end
      COMP_LOOP_C_783 : begin
        fsm_output = 11'b10100111011;
        state_var_NS = COMP_LOOP_C_784;
      end
      COMP_LOOP_C_784 : begin
        fsm_output = 11'b10100111100;
        state_var_NS = COMP_LOOP_C_785;
      end
      COMP_LOOP_C_785 : begin
        fsm_output = 11'b10100111101;
        state_var_NS = COMP_LOOP_C_786;
      end
      COMP_LOOP_C_786 : begin
        fsm_output = 11'b10100111110;
        state_var_NS = COMP_LOOP_C_787;
      end
      COMP_LOOP_C_787 : begin
        fsm_output = 11'b10100111111;
        state_var_NS = COMP_LOOP_C_788;
      end
      COMP_LOOP_C_788 : begin
        fsm_output = 11'b10101000000;
        state_var_NS = COMP_LOOP_C_789;
      end
      COMP_LOOP_C_789 : begin
        fsm_output = 11'b10101000001;
        state_var_NS = COMP_LOOP_C_790;
      end
      COMP_LOOP_C_790 : begin
        fsm_output = 11'b10101000010;
        state_var_NS = COMP_LOOP_C_791;
      end
      COMP_LOOP_C_791 : begin
        fsm_output = 11'b10101000011;
        state_var_NS = COMP_LOOP_C_792;
      end
      COMP_LOOP_C_792 : begin
        fsm_output = 11'b10101000100;
        state_var_NS = COMP_LOOP_C_793;
      end
      COMP_LOOP_C_793 : begin
        fsm_output = 11'b10101000101;
        state_var_NS = COMP_LOOP_C_794;
      end
      COMP_LOOP_C_794 : begin
        fsm_output = 11'b10101000110;
        state_var_NS = COMP_LOOP_C_795;
      end
      COMP_LOOP_C_795 : begin
        fsm_output = 11'b10101000111;
        state_var_NS = COMP_LOOP_C_796;
      end
      COMP_LOOP_C_796 : begin
        fsm_output = 11'b10101001000;
        state_var_NS = COMP_LOOP_C_797;
      end
      COMP_LOOP_C_797 : begin
        fsm_output = 11'b10101001001;
        state_var_NS = COMP_LOOP_C_798;
      end
      COMP_LOOP_C_798 : begin
        fsm_output = 11'b10101001010;
        state_var_NS = COMP_LOOP_C_799;
      end
      COMP_LOOP_C_799 : begin
        fsm_output = 11'b10101001011;
        state_var_NS = COMP_LOOP_C_800;
      end
      COMP_LOOP_C_800 : begin
        fsm_output = 11'b10101001100;
        state_var_NS = COMP_LOOP_C_801;
      end
      COMP_LOOP_C_801 : begin
        fsm_output = 11'b10101001101;
        state_var_NS = COMP_LOOP_C_802;
      end
      COMP_LOOP_C_802 : begin
        fsm_output = 11'b10101001110;
        state_var_NS = COMP_LOOP_C_803;
      end
      COMP_LOOP_C_803 : begin
        fsm_output = 11'b10101001111;
        state_var_NS = COMP_LOOP_C_804;
      end
      COMP_LOOP_C_804 : begin
        fsm_output = 11'b10101010000;
        state_var_NS = COMP_LOOP_C_805;
      end
      COMP_LOOP_C_805 : begin
        fsm_output = 11'b10101010001;
        state_var_NS = COMP_LOOP_C_806;
      end
      COMP_LOOP_C_806 : begin
        fsm_output = 11'b10101010010;
        state_var_NS = COMP_LOOP_C_807;
      end
      COMP_LOOP_C_807 : begin
        fsm_output = 11'b10101010011;
        state_var_NS = COMP_LOOP_C_808;
      end
      COMP_LOOP_C_808 : begin
        fsm_output = 11'b10101010100;
        state_var_NS = COMP_LOOP_C_809;
      end
      COMP_LOOP_C_809 : begin
        fsm_output = 11'b10101010101;
        state_var_NS = COMP_LOOP_C_810;
      end
      COMP_LOOP_C_810 : begin
        fsm_output = 11'b10101010110;
        state_var_NS = COMP_LOOP_C_811;
      end
      COMP_LOOP_C_811 : begin
        fsm_output = 11'b10101010111;
        state_var_NS = COMP_LOOP_C_812;
      end
      COMP_LOOP_C_812 : begin
        fsm_output = 11'b10101011000;
        state_var_NS = COMP_LOOP_C_813;
      end
      COMP_LOOP_C_813 : begin
        fsm_output = 11'b10101011001;
        state_var_NS = COMP_LOOP_C_814;
      end
      COMP_LOOP_C_814 : begin
        fsm_output = 11'b10101011010;
        state_var_NS = COMP_LOOP_C_815;
      end
      COMP_LOOP_C_815 : begin
        fsm_output = 11'b10101011011;
        state_var_NS = COMP_LOOP_C_816;
      end
      COMP_LOOP_C_816 : begin
        fsm_output = 11'b10101011100;
        state_var_NS = COMP_LOOP_C_817;
      end
      COMP_LOOP_C_817 : begin
        fsm_output = 11'b10101011101;
        state_var_NS = COMP_LOOP_C_818;
      end
      COMP_LOOP_C_818 : begin
        fsm_output = 11'b10101011110;
        state_var_NS = COMP_LOOP_C_819;
      end
      COMP_LOOP_C_819 : begin
        fsm_output = 11'b10101011111;
        state_var_NS = COMP_LOOP_C_820;
      end
      COMP_LOOP_C_820 : begin
        fsm_output = 11'b10101100000;
        state_var_NS = COMP_LOOP_C_821;
      end
      COMP_LOOP_C_821 : begin
        fsm_output = 11'b10101100001;
        state_var_NS = COMP_LOOP_C_822;
      end
      COMP_LOOP_C_822 : begin
        fsm_output = 11'b10101100010;
        state_var_NS = COMP_LOOP_C_823;
      end
      COMP_LOOP_C_823 : begin
        fsm_output = 11'b10101100011;
        state_var_NS = COMP_LOOP_C_824;
      end
      COMP_LOOP_C_824 : begin
        fsm_output = 11'b10101100100;
        state_var_NS = COMP_LOOP_C_825;
      end
      COMP_LOOP_C_825 : begin
        fsm_output = 11'b10101100101;
        state_var_NS = COMP_LOOP_C_826;
      end
      COMP_LOOP_C_826 : begin
        fsm_output = 11'b10101100110;
        state_var_NS = COMP_LOOP_C_827;
      end
      COMP_LOOP_C_827 : begin
        fsm_output = 11'b10101100111;
        state_var_NS = COMP_LOOP_C_828;
      end
      COMP_LOOP_C_828 : begin
        fsm_output = 11'b10101101000;
        state_var_NS = COMP_LOOP_C_829;
      end
      COMP_LOOP_C_829 : begin
        fsm_output = 11'b10101101001;
        state_var_NS = COMP_LOOP_C_830;
      end
      COMP_LOOP_C_830 : begin
        fsm_output = 11'b10101101010;
        state_var_NS = COMP_LOOP_C_831;
      end
      COMP_LOOP_C_831 : begin
        fsm_output = 11'b10101101011;
        state_var_NS = COMP_LOOP_C_832;
      end
      COMP_LOOP_C_832 : begin
        fsm_output = 11'b10101101100;
        if ( COMP_LOOP_C_832_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_833;
        end
      end
      COMP_LOOP_C_833 : begin
        fsm_output = 11'b10101101101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_0;
      end
      COMP_LOOP_14_modExp_1_while_C_0 : begin
        fsm_output = 11'b10101101110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_1;
      end
      COMP_LOOP_14_modExp_1_while_C_1 : begin
        fsm_output = 11'b10101101111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_2;
      end
      COMP_LOOP_14_modExp_1_while_C_2 : begin
        fsm_output = 11'b10101110000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_3;
      end
      COMP_LOOP_14_modExp_1_while_C_3 : begin
        fsm_output = 11'b10101110001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_4;
      end
      COMP_LOOP_14_modExp_1_while_C_4 : begin
        fsm_output = 11'b10101110010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_5;
      end
      COMP_LOOP_14_modExp_1_while_C_5 : begin
        fsm_output = 11'b10101110011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_6;
      end
      COMP_LOOP_14_modExp_1_while_C_6 : begin
        fsm_output = 11'b10101110100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_7;
      end
      COMP_LOOP_14_modExp_1_while_C_7 : begin
        fsm_output = 11'b10101110101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_8;
      end
      COMP_LOOP_14_modExp_1_while_C_8 : begin
        fsm_output = 11'b10101110110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_9;
      end
      COMP_LOOP_14_modExp_1_while_C_9 : begin
        fsm_output = 11'b10101110111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_10;
      end
      COMP_LOOP_14_modExp_1_while_C_10 : begin
        fsm_output = 11'b10101111000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_11;
      end
      COMP_LOOP_14_modExp_1_while_C_11 : begin
        fsm_output = 11'b10101111001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_12;
      end
      COMP_LOOP_14_modExp_1_while_C_12 : begin
        fsm_output = 11'b10101111010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_13;
      end
      COMP_LOOP_14_modExp_1_while_C_13 : begin
        fsm_output = 11'b10101111011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_14;
      end
      COMP_LOOP_14_modExp_1_while_C_14 : begin
        fsm_output = 11'b10101111100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_15;
      end
      COMP_LOOP_14_modExp_1_while_C_15 : begin
        fsm_output = 11'b10101111101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_16;
      end
      COMP_LOOP_14_modExp_1_while_C_16 : begin
        fsm_output = 11'b10101111110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_17;
      end
      COMP_LOOP_14_modExp_1_while_C_17 : begin
        fsm_output = 11'b10101111111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_18;
      end
      COMP_LOOP_14_modExp_1_while_C_18 : begin
        fsm_output = 11'b10110000000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_19;
      end
      COMP_LOOP_14_modExp_1_while_C_19 : begin
        fsm_output = 11'b10110000001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_20;
      end
      COMP_LOOP_14_modExp_1_while_C_20 : begin
        fsm_output = 11'b10110000010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_21;
      end
      COMP_LOOP_14_modExp_1_while_C_21 : begin
        fsm_output = 11'b10110000011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_22;
      end
      COMP_LOOP_14_modExp_1_while_C_22 : begin
        fsm_output = 11'b10110000100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_23;
      end
      COMP_LOOP_14_modExp_1_while_C_23 : begin
        fsm_output = 11'b10110000101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_24;
      end
      COMP_LOOP_14_modExp_1_while_C_24 : begin
        fsm_output = 11'b10110000110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_25;
      end
      COMP_LOOP_14_modExp_1_while_C_25 : begin
        fsm_output = 11'b10110000111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_26;
      end
      COMP_LOOP_14_modExp_1_while_C_26 : begin
        fsm_output = 11'b10110001000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_27;
      end
      COMP_LOOP_14_modExp_1_while_C_27 : begin
        fsm_output = 11'b10110001001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_28;
      end
      COMP_LOOP_14_modExp_1_while_C_28 : begin
        fsm_output = 11'b10110001010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_29;
      end
      COMP_LOOP_14_modExp_1_while_C_29 : begin
        fsm_output = 11'b10110001011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_30;
      end
      COMP_LOOP_14_modExp_1_while_C_30 : begin
        fsm_output = 11'b10110001100;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_31;
      end
      COMP_LOOP_14_modExp_1_while_C_31 : begin
        fsm_output = 11'b10110001101;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_32;
      end
      COMP_LOOP_14_modExp_1_while_C_32 : begin
        fsm_output = 11'b10110001110;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_33;
      end
      COMP_LOOP_14_modExp_1_while_C_33 : begin
        fsm_output = 11'b10110001111;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_34;
      end
      COMP_LOOP_14_modExp_1_while_C_34 : begin
        fsm_output = 11'b10110010000;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_35;
      end
      COMP_LOOP_14_modExp_1_while_C_35 : begin
        fsm_output = 11'b10110010001;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_36;
      end
      COMP_LOOP_14_modExp_1_while_C_36 : begin
        fsm_output = 11'b10110010010;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_37;
      end
      COMP_LOOP_14_modExp_1_while_C_37 : begin
        fsm_output = 11'b10110010011;
        state_var_NS = COMP_LOOP_14_modExp_1_while_C_38;
      end
      COMP_LOOP_14_modExp_1_while_C_38 : begin
        fsm_output = 11'b10110010100;
        if ( COMP_LOOP_14_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_834;
        end
        else begin
          state_var_NS = COMP_LOOP_14_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_834 : begin
        fsm_output = 11'b10110010101;
        state_var_NS = COMP_LOOP_C_835;
      end
      COMP_LOOP_C_835 : begin
        fsm_output = 11'b10110010110;
        state_var_NS = COMP_LOOP_C_836;
      end
      COMP_LOOP_C_836 : begin
        fsm_output = 11'b10110010111;
        state_var_NS = COMP_LOOP_C_837;
      end
      COMP_LOOP_C_837 : begin
        fsm_output = 11'b10110011000;
        state_var_NS = COMP_LOOP_C_838;
      end
      COMP_LOOP_C_838 : begin
        fsm_output = 11'b10110011001;
        state_var_NS = COMP_LOOP_C_839;
      end
      COMP_LOOP_C_839 : begin
        fsm_output = 11'b10110011010;
        state_var_NS = COMP_LOOP_C_840;
      end
      COMP_LOOP_C_840 : begin
        fsm_output = 11'b10110011011;
        state_var_NS = COMP_LOOP_C_841;
      end
      COMP_LOOP_C_841 : begin
        fsm_output = 11'b10110011100;
        state_var_NS = COMP_LOOP_C_842;
      end
      COMP_LOOP_C_842 : begin
        fsm_output = 11'b10110011101;
        state_var_NS = COMP_LOOP_C_843;
      end
      COMP_LOOP_C_843 : begin
        fsm_output = 11'b10110011110;
        state_var_NS = COMP_LOOP_C_844;
      end
      COMP_LOOP_C_844 : begin
        fsm_output = 11'b10110011111;
        state_var_NS = COMP_LOOP_C_845;
      end
      COMP_LOOP_C_845 : begin
        fsm_output = 11'b10110100000;
        state_var_NS = COMP_LOOP_C_846;
      end
      COMP_LOOP_C_846 : begin
        fsm_output = 11'b10110100001;
        state_var_NS = COMP_LOOP_C_847;
      end
      COMP_LOOP_C_847 : begin
        fsm_output = 11'b10110100010;
        state_var_NS = COMP_LOOP_C_848;
      end
      COMP_LOOP_C_848 : begin
        fsm_output = 11'b10110100011;
        state_var_NS = COMP_LOOP_C_849;
      end
      COMP_LOOP_C_849 : begin
        fsm_output = 11'b10110100100;
        state_var_NS = COMP_LOOP_C_850;
      end
      COMP_LOOP_C_850 : begin
        fsm_output = 11'b10110100101;
        state_var_NS = COMP_LOOP_C_851;
      end
      COMP_LOOP_C_851 : begin
        fsm_output = 11'b10110100110;
        state_var_NS = COMP_LOOP_C_852;
      end
      COMP_LOOP_C_852 : begin
        fsm_output = 11'b10110100111;
        state_var_NS = COMP_LOOP_C_853;
      end
      COMP_LOOP_C_853 : begin
        fsm_output = 11'b10110101000;
        state_var_NS = COMP_LOOP_C_854;
      end
      COMP_LOOP_C_854 : begin
        fsm_output = 11'b10110101001;
        state_var_NS = COMP_LOOP_C_855;
      end
      COMP_LOOP_C_855 : begin
        fsm_output = 11'b10110101010;
        state_var_NS = COMP_LOOP_C_856;
      end
      COMP_LOOP_C_856 : begin
        fsm_output = 11'b10110101011;
        state_var_NS = COMP_LOOP_C_857;
      end
      COMP_LOOP_C_857 : begin
        fsm_output = 11'b10110101100;
        state_var_NS = COMP_LOOP_C_858;
      end
      COMP_LOOP_C_858 : begin
        fsm_output = 11'b10110101101;
        state_var_NS = COMP_LOOP_C_859;
      end
      COMP_LOOP_C_859 : begin
        fsm_output = 11'b10110101110;
        state_var_NS = COMP_LOOP_C_860;
      end
      COMP_LOOP_C_860 : begin
        fsm_output = 11'b10110101111;
        state_var_NS = COMP_LOOP_C_861;
      end
      COMP_LOOP_C_861 : begin
        fsm_output = 11'b10110110000;
        state_var_NS = COMP_LOOP_C_862;
      end
      COMP_LOOP_C_862 : begin
        fsm_output = 11'b10110110001;
        state_var_NS = COMP_LOOP_C_863;
      end
      COMP_LOOP_C_863 : begin
        fsm_output = 11'b10110110010;
        state_var_NS = COMP_LOOP_C_864;
      end
      COMP_LOOP_C_864 : begin
        fsm_output = 11'b10110110011;
        state_var_NS = COMP_LOOP_C_865;
      end
      COMP_LOOP_C_865 : begin
        fsm_output = 11'b10110110100;
        state_var_NS = COMP_LOOP_C_866;
      end
      COMP_LOOP_C_866 : begin
        fsm_output = 11'b10110110101;
        state_var_NS = COMP_LOOP_C_867;
      end
      COMP_LOOP_C_867 : begin
        fsm_output = 11'b10110110110;
        state_var_NS = COMP_LOOP_C_868;
      end
      COMP_LOOP_C_868 : begin
        fsm_output = 11'b10110110111;
        state_var_NS = COMP_LOOP_C_869;
      end
      COMP_LOOP_C_869 : begin
        fsm_output = 11'b10110111000;
        state_var_NS = COMP_LOOP_C_870;
      end
      COMP_LOOP_C_870 : begin
        fsm_output = 11'b10110111001;
        state_var_NS = COMP_LOOP_C_871;
      end
      COMP_LOOP_C_871 : begin
        fsm_output = 11'b10110111010;
        state_var_NS = COMP_LOOP_C_872;
      end
      COMP_LOOP_C_872 : begin
        fsm_output = 11'b10110111011;
        state_var_NS = COMP_LOOP_C_873;
      end
      COMP_LOOP_C_873 : begin
        fsm_output = 11'b10110111100;
        state_var_NS = COMP_LOOP_C_874;
      end
      COMP_LOOP_C_874 : begin
        fsm_output = 11'b10110111101;
        state_var_NS = COMP_LOOP_C_875;
      end
      COMP_LOOP_C_875 : begin
        fsm_output = 11'b10110111110;
        state_var_NS = COMP_LOOP_C_876;
      end
      COMP_LOOP_C_876 : begin
        fsm_output = 11'b10110111111;
        state_var_NS = COMP_LOOP_C_877;
      end
      COMP_LOOP_C_877 : begin
        fsm_output = 11'b10111000000;
        state_var_NS = COMP_LOOP_C_878;
      end
      COMP_LOOP_C_878 : begin
        fsm_output = 11'b10111000001;
        state_var_NS = COMP_LOOP_C_879;
      end
      COMP_LOOP_C_879 : begin
        fsm_output = 11'b10111000010;
        state_var_NS = COMP_LOOP_C_880;
      end
      COMP_LOOP_C_880 : begin
        fsm_output = 11'b10111000011;
        state_var_NS = COMP_LOOP_C_881;
      end
      COMP_LOOP_C_881 : begin
        fsm_output = 11'b10111000100;
        state_var_NS = COMP_LOOP_C_882;
      end
      COMP_LOOP_C_882 : begin
        fsm_output = 11'b10111000101;
        state_var_NS = COMP_LOOP_C_883;
      end
      COMP_LOOP_C_883 : begin
        fsm_output = 11'b10111000110;
        state_var_NS = COMP_LOOP_C_884;
      end
      COMP_LOOP_C_884 : begin
        fsm_output = 11'b10111000111;
        state_var_NS = COMP_LOOP_C_885;
      end
      COMP_LOOP_C_885 : begin
        fsm_output = 11'b10111001000;
        state_var_NS = COMP_LOOP_C_886;
      end
      COMP_LOOP_C_886 : begin
        fsm_output = 11'b10111001001;
        state_var_NS = COMP_LOOP_C_887;
      end
      COMP_LOOP_C_887 : begin
        fsm_output = 11'b10111001010;
        state_var_NS = COMP_LOOP_C_888;
      end
      COMP_LOOP_C_888 : begin
        fsm_output = 11'b10111001011;
        state_var_NS = COMP_LOOP_C_889;
      end
      COMP_LOOP_C_889 : begin
        fsm_output = 11'b10111001100;
        state_var_NS = COMP_LOOP_C_890;
      end
      COMP_LOOP_C_890 : begin
        fsm_output = 11'b10111001101;
        state_var_NS = COMP_LOOP_C_891;
      end
      COMP_LOOP_C_891 : begin
        fsm_output = 11'b10111001110;
        state_var_NS = COMP_LOOP_C_892;
      end
      COMP_LOOP_C_892 : begin
        fsm_output = 11'b10111001111;
        state_var_NS = COMP_LOOP_C_893;
      end
      COMP_LOOP_C_893 : begin
        fsm_output = 11'b10111010000;
        state_var_NS = COMP_LOOP_C_894;
      end
      COMP_LOOP_C_894 : begin
        fsm_output = 11'b10111010001;
        state_var_NS = COMP_LOOP_C_895;
      end
      COMP_LOOP_C_895 : begin
        fsm_output = 11'b10111010010;
        state_var_NS = COMP_LOOP_C_896;
      end
      COMP_LOOP_C_896 : begin
        fsm_output = 11'b10111010011;
        if ( COMP_LOOP_C_896_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_897;
        end
      end
      COMP_LOOP_C_897 : begin
        fsm_output = 11'b10111010100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_0;
      end
      COMP_LOOP_15_modExp_1_while_C_0 : begin
        fsm_output = 11'b10111010101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_1;
      end
      COMP_LOOP_15_modExp_1_while_C_1 : begin
        fsm_output = 11'b10111010110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_2;
      end
      COMP_LOOP_15_modExp_1_while_C_2 : begin
        fsm_output = 11'b10111010111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_3;
      end
      COMP_LOOP_15_modExp_1_while_C_3 : begin
        fsm_output = 11'b10111011000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_4;
      end
      COMP_LOOP_15_modExp_1_while_C_4 : begin
        fsm_output = 11'b10111011001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_5;
      end
      COMP_LOOP_15_modExp_1_while_C_5 : begin
        fsm_output = 11'b10111011010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_6;
      end
      COMP_LOOP_15_modExp_1_while_C_6 : begin
        fsm_output = 11'b10111011011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_7;
      end
      COMP_LOOP_15_modExp_1_while_C_7 : begin
        fsm_output = 11'b10111011100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_8;
      end
      COMP_LOOP_15_modExp_1_while_C_8 : begin
        fsm_output = 11'b10111011101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_9;
      end
      COMP_LOOP_15_modExp_1_while_C_9 : begin
        fsm_output = 11'b10111011110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_10;
      end
      COMP_LOOP_15_modExp_1_while_C_10 : begin
        fsm_output = 11'b10111011111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_11;
      end
      COMP_LOOP_15_modExp_1_while_C_11 : begin
        fsm_output = 11'b10111100000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_12;
      end
      COMP_LOOP_15_modExp_1_while_C_12 : begin
        fsm_output = 11'b10111100001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_13;
      end
      COMP_LOOP_15_modExp_1_while_C_13 : begin
        fsm_output = 11'b10111100010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_14;
      end
      COMP_LOOP_15_modExp_1_while_C_14 : begin
        fsm_output = 11'b10111100011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_15;
      end
      COMP_LOOP_15_modExp_1_while_C_15 : begin
        fsm_output = 11'b10111100100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_16;
      end
      COMP_LOOP_15_modExp_1_while_C_16 : begin
        fsm_output = 11'b10111100101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_17;
      end
      COMP_LOOP_15_modExp_1_while_C_17 : begin
        fsm_output = 11'b10111100110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_18;
      end
      COMP_LOOP_15_modExp_1_while_C_18 : begin
        fsm_output = 11'b10111100111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_19;
      end
      COMP_LOOP_15_modExp_1_while_C_19 : begin
        fsm_output = 11'b10111101000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_20;
      end
      COMP_LOOP_15_modExp_1_while_C_20 : begin
        fsm_output = 11'b10111101001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_21;
      end
      COMP_LOOP_15_modExp_1_while_C_21 : begin
        fsm_output = 11'b10111101010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_22;
      end
      COMP_LOOP_15_modExp_1_while_C_22 : begin
        fsm_output = 11'b10111101011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_23;
      end
      COMP_LOOP_15_modExp_1_while_C_23 : begin
        fsm_output = 11'b10111101100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_24;
      end
      COMP_LOOP_15_modExp_1_while_C_24 : begin
        fsm_output = 11'b10111101101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_25;
      end
      COMP_LOOP_15_modExp_1_while_C_25 : begin
        fsm_output = 11'b10111101110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_26;
      end
      COMP_LOOP_15_modExp_1_while_C_26 : begin
        fsm_output = 11'b10111101111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_27;
      end
      COMP_LOOP_15_modExp_1_while_C_27 : begin
        fsm_output = 11'b10111110000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_28;
      end
      COMP_LOOP_15_modExp_1_while_C_28 : begin
        fsm_output = 11'b10111110001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_29;
      end
      COMP_LOOP_15_modExp_1_while_C_29 : begin
        fsm_output = 11'b10111110010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_30;
      end
      COMP_LOOP_15_modExp_1_while_C_30 : begin
        fsm_output = 11'b10111110011;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_31;
      end
      COMP_LOOP_15_modExp_1_while_C_31 : begin
        fsm_output = 11'b10111110100;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_32;
      end
      COMP_LOOP_15_modExp_1_while_C_32 : begin
        fsm_output = 11'b10111110101;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_33;
      end
      COMP_LOOP_15_modExp_1_while_C_33 : begin
        fsm_output = 11'b10111110110;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_34;
      end
      COMP_LOOP_15_modExp_1_while_C_34 : begin
        fsm_output = 11'b10111110111;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_35;
      end
      COMP_LOOP_15_modExp_1_while_C_35 : begin
        fsm_output = 11'b10111111000;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_36;
      end
      COMP_LOOP_15_modExp_1_while_C_36 : begin
        fsm_output = 11'b10111111001;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_37;
      end
      COMP_LOOP_15_modExp_1_while_C_37 : begin
        fsm_output = 11'b10111111010;
        state_var_NS = COMP_LOOP_15_modExp_1_while_C_38;
      end
      COMP_LOOP_15_modExp_1_while_C_38 : begin
        fsm_output = 11'b10111111011;
        if ( COMP_LOOP_15_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_898;
        end
        else begin
          state_var_NS = COMP_LOOP_15_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_898 : begin
        fsm_output = 11'b10111111100;
        state_var_NS = COMP_LOOP_C_899;
      end
      COMP_LOOP_C_899 : begin
        fsm_output = 11'b10111111101;
        state_var_NS = COMP_LOOP_C_900;
      end
      COMP_LOOP_C_900 : begin
        fsm_output = 11'b10111111110;
        state_var_NS = COMP_LOOP_C_901;
      end
      COMP_LOOP_C_901 : begin
        fsm_output = 11'b10111111111;
        state_var_NS = COMP_LOOP_C_902;
      end
      COMP_LOOP_C_902 : begin
        fsm_output = 11'b11000000000;
        state_var_NS = COMP_LOOP_C_903;
      end
      COMP_LOOP_C_903 : begin
        fsm_output = 11'b11000000001;
        state_var_NS = COMP_LOOP_C_904;
      end
      COMP_LOOP_C_904 : begin
        fsm_output = 11'b11000000010;
        state_var_NS = COMP_LOOP_C_905;
      end
      COMP_LOOP_C_905 : begin
        fsm_output = 11'b11000000011;
        state_var_NS = COMP_LOOP_C_906;
      end
      COMP_LOOP_C_906 : begin
        fsm_output = 11'b11000000100;
        state_var_NS = COMP_LOOP_C_907;
      end
      COMP_LOOP_C_907 : begin
        fsm_output = 11'b11000000101;
        state_var_NS = COMP_LOOP_C_908;
      end
      COMP_LOOP_C_908 : begin
        fsm_output = 11'b11000000110;
        state_var_NS = COMP_LOOP_C_909;
      end
      COMP_LOOP_C_909 : begin
        fsm_output = 11'b11000000111;
        state_var_NS = COMP_LOOP_C_910;
      end
      COMP_LOOP_C_910 : begin
        fsm_output = 11'b11000001000;
        state_var_NS = COMP_LOOP_C_911;
      end
      COMP_LOOP_C_911 : begin
        fsm_output = 11'b11000001001;
        state_var_NS = COMP_LOOP_C_912;
      end
      COMP_LOOP_C_912 : begin
        fsm_output = 11'b11000001010;
        state_var_NS = COMP_LOOP_C_913;
      end
      COMP_LOOP_C_913 : begin
        fsm_output = 11'b11000001011;
        state_var_NS = COMP_LOOP_C_914;
      end
      COMP_LOOP_C_914 : begin
        fsm_output = 11'b11000001100;
        state_var_NS = COMP_LOOP_C_915;
      end
      COMP_LOOP_C_915 : begin
        fsm_output = 11'b11000001101;
        state_var_NS = COMP_LOOP_C_916;
      end
      COMP_LOOP_C_916 : begin
        fsm_output = 11'b11000001110;
        state_var_NS = COMP_LOOP_C_917;
      end
      COMP_LOOP_C_917 : begin
        fsm_output = 11'b11000001111;
        state_var_NS = COMP_LOOP_C_918;
      end
      COMP_LOOP_C_918 : begin
        fsm_output = 11'b11000010000;
        state_var_NS = COMP_LOOP_C_919;
      end
      COMP_LOOP_C_919 : begin
        fsm_output = 11'b11000010001;
        state_var_NS = COMP_LOOP_C_920;
      end
      COMP_LOOP_C_920 : begin
        fsm_output = 11'b11000010010;
        state_var_NS = COMP_LOOP_C_921;
      end
      COMP_LOOP_C_921 : begin
        fsm_output = 11'b11000010011;
        state_var_NS = COMP_LOOP_C_922;
      end
      COMP_LOOP_C_922 : begin
        fsm_output = 11'b11000010100;
        state_var_NS = COMP_LOOP_C_923;
      end
      COMP_LOOP_C_923 : begin
        fsm_output = 11'b11000010101;
        state_var_NS = COMP_LOOP_C_924;
      end
      COMP_LOOP_C_924 : begin
        fsm_output = 11'b11000010110;
        state_var_NS = COMP_LOOP_C_925;
      end
      COMP_LOOP_C_925 : begin
        fsm_output = 11'b11000010111;
        state_var_NS = COMP_LOOP_C_926;
      end
      COMP_LOOP_C_926 : begin
        fsm_output = 11'b11000011000;
        state_var_NS = COMP_LOOP_C_927;
      end
      COMP_LOOP_C_927 : begin
        fsm_output = 11'b11000011001;
        state_var_NS = COMP_LOOP_C_928;
      end
      COMP_LOOP_C_928 : begin
        fsm_output = 11'b11000011010;
        state_var_NS = COMP_LOOP_C_929;
      end
      COMP_LOOP_C_929 : begin
        fsm_output = 11'b11000011011;
        state_var_NS = COMP_LOOP_C_930;
      end
      COMP_LOOP_C_930 : begin
        fsm_output = 11'b11000011100;
        state_var_NS = COMP_LOOP_C_931;
      end
      COMP_LOOP_C_931 : begin
        fsm_output = 11'b11000011101;
        state_var_NS = COMP_LOOP_C_932;
      end
      COMP_LOOP_C_932 : begin
        fsm_output = 11'b11000011110;
        state_var_NS = COMP_LOOP_C_933;
      end
      COMP_LOOP_C_933 : begin
        fsm_output = 11'b11000011111;
        state_var_NS = COMP_LOOP_C_934;
      end
      COMP_LOOP_C_934 : begin
        fsm_output = 11'b11000100000;
        state_var_NS = COMP_LOOP_C_935;
      end
      COMP_LOOP_C_935 : begin
        fsm_output = 11'b11000100001;
        state_var_NS = COMP_LOOP_C_936;
      end
      COMP_LOOP_C_936 : begin
        fsm_output = 11'b11000100010;
        state_var_NS = COMP_LOOP_C_937;
      end
      COMP_LOOP_C_937 : begin
        fsm_output = 11'b11000100011;
        state_var_NS = COMP_LOOP_C_938;
      end
      COMP_LOOP_C_938 : begin
        fsm_output = 11'b11000100100;
        state_var_NS = COMP_LOOP_C_939;
      end
      COMP_LOOP_C_939 : begin
        fsm_output = 11'b11000100101;
        state_var_NS = COMP_LOOP_C_940;
      end
      COMP_LOOP_C_940 : begin
        fsm_output = 11'b11000100110;
        state_var_NS = COMP_LOOP_C_941;
      end
      COMP_LOOP_C_941 : begin
        fsm_output = 11'b11000100111;
        state_var_NS = COMP_LOOP_C_942;
      end
      COMP_LOOP_C_942 : begin
        fsm_output = 11'b11000101000;
        state_var_NS = COMP_LOOP_C_943;
      end
      COMP_LOOP_C_943 : begin
        fsm_output = 11'b11000101001;
        state_var_NS = COMP_LOOP_C_944;
      end
      COMP_LOOP_C_944 : begin
        fsm_output = 11'b11000101010;
        state_var_NS = COMP_LOOP_C_945;
      end
      COMP_LOOP_C_945 : begin
        fsm_output = 11'b11000101011;
        state_var_NS = COMP_LOOP_C_946;
      end
      COMP_LOOP_C_946 : begin
        fsm_output = 11'b11000101100;
        state_var_NS = COMP_LOOP_C_947;
      end
      COMP_LOOP_C_947 : begin
        fsm_output = 11'b11000101101;
        state_var_NS = COMP_LOOP_C_948;
      end
      COMP_LOOP_C_948 : begin
        fsm_output = 11'b11000101110;
        state_var_NS = COMP_LOOP_C_949;
      end
      COMP_LOOP_C_949 : begin
        fsm_output = 11'b11000101111;
        state_var_NS = COMP_LOOP_C_950;
      end
      COMP_LOOP_C_950 : begin
        fsm_output = 11'b11000110000;
        state_var_NS = COMP_LOOP_C_951;
      end
      COMP_LOOP_C_951 : begin
        fsm_output = 11'b11000110001;
        state_var_NS = COMP_LOOP_C_952;
      end
      COMP_LOOP_C_952 : begin
        fsm_output = 11'b11000110010;
        state_var_NS = COMP_LOOP_C_953;
      end
      COMP_LOOP_C_953 : begin
        fsm_output = 11'b11000110011;
        state_var_NS = COMP_LOOP_C_954;
      end
      COMP_LOOP_C_954 : begin
        fsm_output = 11'b11000110100;
        state_var_NS = COMP_LOOP_C_955;
      end
      COMP_LOOP_C_955 : begin
        fsm_output = 11'b11000110101;
        state_var_NS = COMP_LOOP_C_956;
      end
      COMP_LOOP_C_956 : begin
        fsm_output = 11'b11000110110;
        state_var_NS = COMP_LOOP_C_957;
      end
      COMP_LOOP_C_957 : begin
        fsm_output = 11'b11000110111;
        state_var_NS = COMP_LOOP_C_958;
      end
      COMP_LOOP_C_958 : begin
        fsm_output = 11'b11000111000;
        state_var_NS = COMP_LOOP_C_959;
      end
      COMP_LOOP_C_959 : begin
        fsm_output = 11'b11000111001;
        state_var_NS = COMP_LOOP_C_960;
      end
      COMP_LOOP_C_960 : begin
        fsm_output = 11'b11000111010;
        if ( COMP_LOOP_C_960_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_961;
        end
      end
      COMP_LOOP_C_961 : begin
        fsm_output = 11'b11000111011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_0;
      end
      COMP_LOOP_16_modExp_1_while_C_0 : begin
        fsm_output = 11'b11000111100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_1;
      end
      COMP_LOOP_16_modExp_1_while_C_1 : begin
        fsm_output = 11'b11000111101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_2;
      end
      COMP_LOOP_16_modExp_1_while_C_2 : begin
        fsm_output = 11'b11000111110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_3;
      end
      COMP_LOOP_16_modExp_1_while_C_3 : begin
        fsm_output = 11'b11000111111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_4;
      end
      COMP_LOOP_16_modExp_1_while_C_4 : begin
        fsm_output = 11'b11001000000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_5;
      end
      COMP_LOOP_16_modExp_1_while_C_5 : begin
        fsm_output = 11'b11001000001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_6;
      end
      COMP_LOOP_16_modExp_1_while_C_6 : begin
        fsm_output = 11'b11001000010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_7;
      end
      COMP_LOOP_16_modExp_1_while_C_7 : begin
        fsm_output = 11'b11001000011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_8;
      end
      COMP_LOOP_16_modExp_1_while_C_8 : begin
        fsm_output = 11'b11001000100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_9;
      end
      COMP_LOOP_16_modExp_1_while_C_9 : begin
        fsm_output = 11'b11001000101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_10;
      end
      COMP_LOOP_16_modExp_1_while_C_10 : begin
        fsm_output = 11'b11001000110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_11;
      end
      COMP_LOOP_16_modExp_1_while_C_11 : begin
        fsm_output = 11'b11001000111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_12;
      end
      COMP_LOOP_16_modExp_1_while_C_12 : begin
        fsm_output = 11'b11001001000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_13;
      end
      COMP_LOOP_16_modExp_1_while_C_13 : begin
        fsm_output = 11'b11001001001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_14;
      end
      COMP_LOOP_16_modExp_1_while_C_14 : begin
        fsm_output = 11'b11001001010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_15;
      end
      COMP_LOOP_16_modExp_1_while_C_15 : begin
        fsm_output = 11'b11001001011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_16;
      end
      COMP_LOOP_16_modExp_1_while_C_16 : begin
        fsm_output = 11'b11001001100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_17;
      end
      COMP_LOOP_16_modExp_1_while_C_17 : begin
        fsm_output = 11'b11001001101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_18;
      end
      COMP_LOOP_16_modExp_1_while_C_18 : begin
        fsm_output = 11'b11001001110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_19;
      end
      COMP_LOOP_16_modExp_1_while_C_19 : begin
        fsm_output = 11'b11001001111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_20;
      end
      COMP_LOOP_16_modExp_1_while_C_20 : begin
        fsm_output = 11'b11001010000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_21;
      end
      COMP_LOOP_16_modExp_1_while_C_21 : begin
        fsm_output = 11'b11001010001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_22;
      end
      COMP_LOOP_16_modExp_1_while_C_22 : begin
        fsm_output = 11'b11001010010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_23;
      end
      COMP_LOOP_16_modExp_1_while_C_23 : begin
        fsm_output = 11'b11001010011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_24;
      end
      COMP_LOOP_16_modExp_1_while_C_24 : begin
        fsm_output = 11'b11001010100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_25;
      end
      COMP_LOOP_16_modExp_1_while_C_25 : begin
        fsm_output = 11'b11001010101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_26;
      end
      COMP_LOOP_16_modExp_1_while_C_26 : begin
        fsm_output = 11'b11001010110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_27;
      end
      COMP_LOOP_16_modExp_1_while_C_27 : begin
        fsm_output = 11'b11001010111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_28;
      end
      COMP_LOOP_16_modExp_1_while_C_28 : begin
        fsm_output = 11'b11001011000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_29;
      end
      COMP_LOOP_16_modExp_1_while_C_29 : begin
        fsm_output = 11'b11001011001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_30;
      end
      COMP_LOOP_16_modExp_1_while_C_30 : begin
        fsm_output = 11'b11001011010;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_31;
      end
      COMP_LOOP_16_modExp_1_while_C_31 : begin
        fsm_output = 11'b11001011011;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_32;
      end
      COMP_LOOP_16_modExp_1_while_C_32 : begin
        fsm_output = 11'b11001011100;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_33;
      end
      COMP_LOOP_16_modExp_1_while_C_33 : begin
        fsm_output = 11'b11001011101;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_34;
      end
      COMP_LOOP_16_modExp_1_while_C_34 : begin
        fsm_output = 11'b11001011110;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_35;
      end
      COMP_LOOP_16_modExp_1_while_C_35 : begin
        fsm_output = 11'b11001011111;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_36;
      end
      COMP_LOOP_16_modExp_1_while_C_36 : begin
        fsm_output = 11'b11001100000;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_37;
      end
      COMP_LOOP_16_modExp_1_while_C_37 : begin
        fsm_output = 11'b11001100001;
        state_var_NS = COMP_LOOP_16_modExp_1_while_C_38;
      end
      COMP_LOOP_16_modExp_1_while_C_38 : begin
        fsm_output = 11'b11001100010;
        if ( COMP_LOOP_16_modExp_1_while_C_38_tr0 ) begin
          state_var_NS = COMP_LOOP_C_962;
        end
        else begin
          state_var_NS = COMP_LOOP_16_modExp_1_while_C_0;
        end
      end
      COMP_LOOP_C_962 : begin
        fsm_output = 11'b11001100011;
        state_var_NS = COMP_LOOP_C_963;
      end
      COMP_LOOP_C_963 : begin
        fsm_output = 11'b11001100100;
        state_var_NS = COMP_LOOP_C_964;
      end
      COMP_LOOP_C_964 : begin
        fsm_output = 11'b11001100101;
        state_var_NS = COMP_LOOP_C_965;
      end
      COMP_LOOP_C_965 : begin
        fsm_output = 11'b11001100110;
        state_var_NS = COMP_LOOP_C_966;
      end
      COMP_LOOP_C_966 : begin
        fsm_output = 11'b11001100111;
        state_var_NS = COMP_LOOP_C_967;
      end
      COMP_LOOP_C_967 : begin
        fsm_output = 11'b11001101000;
        state_var_NS = COMP_LOOP_C_968;
      end
      COMP_LOOP_C_968 : begin
        fsm_output = 11'b11001101001;
        state_var_NS = COMP_LOOP_C_969;
      end
      COMP_LOOP_C_969 : begin
        fsm_output = 11'b11001101010;
        state_var_NS = COMP_LOOP_C_970;
      end
      COMP_LOOP_C_970 : begin
        fsm_output = 11'b11001101011;
        state_var_NS = COMP_LOOP_C_971;
      end
      COMP_LOOP_C_971 : begin
        fsm_output = 11'b11001101100;
        state_var_NS = COMP_LOOP_C_972;
      end
      COMP_LOOP_C_972 : begin
        fsm_output = 11'b11001101101;
        state_var_NS = COMP_LOOP_C_973;
      end
      COMP_LOOP_C_973 : begin
        fsm_output = 11'b11001101110;
        state_var_NS = COMP_LOOP_C_974;
      end
      COMP_LOOP_C_974 : begin
        fsm_output = 11'b11001101111;
        state_var_NS = COMP_LOOP_C_975;
      end
      COMP_LOOP_C_975 : begin
        fsm_output = 11'b11001110000;
        state_var_NS = COMP_LOOP_C_976;
      end
      COMP_LOOP_C_976 : begin
        fsm_output = 11'b11001110001;
        state_var_NS = COMP_LOOP_C_977;
      end
      COMP_LOOP_C_977 : begin
        fsm_output = 11'b11001110010;
        state_var_NS = COMP_LOOP_C_978;
      end
      COMP_LOOP_C_978 : begin
        fsm_output = 11'b11001110011;
        state_var_NS = COMP_LOOP_C_979;
      end
      COMP_LOOP_C_979 : begin
        fsm_output = 11'b11001110100;
        state_var_NS = COMP_LOOP_C_980;
      end
      COMP_LOOP_C_980 : begin
        fsm_output = 11'b11001110101;
        state_var_NS = COMP_LOOP_C_981;
      end
      COMP_LOOP_C_981 : begin
        fsm_output = 11'b11001110110;
        state_var_NS = COMP_LOOP_C_982;
      end
      COMP_LOOP_C_982 : begin
        fsm_output = 11'b11001110111;
        state_var_NS = COMP_LOOP_C_983;
      end
      COMP_LOOP_C_983 : begin
        fsm_output = 11'b11001111000;
        state_var_NS = COMP_LOOP_C_984;
      end
      COMP_LOOP_C_984 : begin
        fsm_output = 11'b11001111001;
        state_var_NS = COMP_LOOP_C_985;
      end
      COMP_LOOP_C_985 : begin
        fsm_output = 11'b11001111010;
        state_var_NS = COMP_LOOP_C_986;
      end
      COMP_LOOP_C_986 : begin
        fsm_output = 11'b11001111011;
        state_var_NS = COMP_LOOP_C_987;
      end
      COMP_LOOP_C_987 : begin
        fsm_output = 11'b11001111100;
        state_var_NS = COMP_LOOP_C_988;
      end
      COMP_LOOP_C_988 : begin
        fsm_output = 11'b11001111101;
        state_var_NS = COMP_LOOP_C_989;
      end
      COMP_LOOP_C_989 : begin
        fsm_output = 11'b11001111110;
        state_var_NS = COMP_LOOP_C_990;
      end
      COMP_LOOP_C_990 : begin
        fsm_output = 11'b11001111111;
        state_var_NS = COMP_LOOP_C_991;
      end
      COMP_LOOP_C_991 : begin
        fsm_output = 11'b11010000000;
        state_var_NS = COMP_LOOP_C_992;
      end
      COMP_LOOP_C_992 : begin
        fsm_output = 11'b11010000001;
        state_var_NS = COMP_LOOP_C_993;
      end
      COMP_LOOP_C_993 : begin
        fsm_output = 11'b11010000010;
        state_var_NS = COMP_LOOP_C_994;
      end
      COMP_LOOP_C_994 : begin
        fsm_output = 11'b11010000011;
        state_var_NS = COMP_LOOP_C_995;
      end
      COMP_LOOP_C_995 : begin
        fsm_output = 11'b11010000100;
        state_var_NS = COMP_LOOP_C_996;
      end
      COMP_LOOP_C_996 : begin
        fsm_output = 11'b11010000101;
        state_var_NS = COMP_LOOP_C_997;
      end
      COMP_LOOP_C_997 : begin
        fsm_output = 11'b11010000110;
        state_var_NS = COMP_LOOP_C_998;
      end
      COMP_LOOP_C_998 : begin
        fsm_output = 11'b11010000111;
        state_var_NS = COMP_LOOP_C_999;
      end
      COMP_LOOP_C_999 : begin
        fsm_output = 11'b11010001000;
        state_var_NS = COMP_LOOP_C_1000;
      end
      COMP_LOOP_C_1000 : begin
        fsm_output = 11'b11010001001;
        state_var_NS = COMP_LOOP_C_1001;
      end
      COMP_LOOP_C_1001 : begin
        fsm_output = 11'b11010001010;
        state_var_NS = COMP_LOOP_C_1002;
      end
      COMP_LOOP_C_1002 : begin
        fsm_output = 11'b11010001011;
        state_var_NS = COMP_LOOP_C_1003;
      end
      COMP_LOOP_C_1003 : begin
        fsm_output = 11'b11010001100;
        state_var_NS = COMP_LOOP_C_1004;
      end
      COMP_LOOP_C_1004 : begin
        fsm_output = 11'b11010001101;
        state_var_NS = COMP_LOOP_C_1005;
      end
      COMP_LOOP_C_1005 : begin
        fsm_output = 11'b11010001110;
        state_var_NS = COMP_LOOP_C_1006;
      end
      COMP_LOOP_C_1006 : begin
        fsm_output = 11'b11010001111;
        state_var_NS = COMP_LOOP_C_1007;
      end
      COMP_LOOP_C_1007 : begin
        fsm_output = 11'b11010010000;
        state_var_NS = COMP_LOOP_C_1008;
      end
      COMP_LOOP_C_1008 : begin
        fsm_output = 11'b11010010001;
        state_var_NS = COMP_LOOP_C_1009;
      end
      COMP_LOOP_C_1009 : begin
        fsm_output = 11'b11010010010;
        state_var_NS = COMP_LOOP_C_1010;
      end
      COMP_LOOP_C_1010 : begin
        fsm_output = 11'b11010010011;
        state_var_NS = COMP_LOOP_C_1011;
      end
      COMP_LOOP_C_1011 : begin
        fsm_output = 11'b11010010100;
        state_var_NS = COMP_LOOP_C_1012;
      end
      COMP_LOOP_C_1012 : begin
        fsm_output = 11'b11010010101;
        state_var_NS = COMP_LOOP_C_1013;
      end
      COMP_LOOP_C_1013 : begin
        fsm_output = 11'b11010010110;
        state_var_NS = COMP_LOOP_C_1014;
      end
      COMP_LOOP_C_1014 : begin
        fsm_output = 11'b11010010111;
        state_var_NS = COMP_LOOP_C_1015;
      end
      COMP_LOOP_C_1015 : begin
        fsm_output = 11'b11010011000;
        state_var_NS = COMP_LOOP_C_1016;
      end
      COMP_LOOP_C_1016 : begin
        fsm_output = 11'b11010011001;
        state_var_NS = COMP_LOOP_C_1017;
      end
      COMP_LOOP_C_1017 : begin
        fsm_output = 11'b11010011010;
        state_var_NS = COMP_LOOP_C_1018;
      end
      COMP_LOOP_C_1018 : begin
        fsm_output = 11'b11010011011;
        state_var_NS = COMP_LOOP_C_1019;
      end
      COMP_LOOP_C_1019 : begin
        fsm_output = 11'b11010011100;
        state_var_NS = COMP_LOOP_C_1020;
      end
      COMP_LOOP_C_1020 : begin
        fsm_output = 11'b11010011101;
        state_var_NS = COMP_LOOP_C_1021;
      end
      COMP_LOOP_C_1021 : begin
        fsm_output = 11'b11010011110;
        state_var_NS = COMP_LOOP_C_1022;
      end
      COMP_LOOP_C_1022 : begin
        fsm_output = 11'b11010011111;
        state_var_NS = COMP_LOOP_C_1023;
      end
      COMP_LOOP_C_1023 : begin
        fsm_output = 11'b11010100000;
        state_var_NS = COMP_LOOP_C_1024;
      end
      COMP_LOOP_C_1024 : begin
        fsm_output = 11'b11010100001;
        if ( COMP_LOOP_C_1024_tr0 ) begin
          state_var_NS = VEC_LOOP_C_0;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      VEC_LOOP_C_0 : begin
        fsm_output = 11'b11010100010;
        if ( VEC_LOOP_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_9;
        end
        else begin
          state_var_NS = COMP_LOOP_C_0;
        end
      end
      STAGE_LOOP_C_9 : begin
        fsm_output = 11'b11010100011;
        if ( STAGE_LOOP_C_9_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 11'b11010100100;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 11'b00000000000;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT_core
// ------------------------------------------------------------------


module inPlaceNTT_DIT_core (
  clk, rst, vec_rsc_triosy_0_0_lz, vec_rsc_triosy_0_1_lz, vec_rsc_triosy_0_2_lz,
      vec_rsc_triosy_0_3_lz, vec_rsc_triosy_0_4_lz, vec_rsc_triosy_0_5_lz, vec_rsc_triosy_0_6_lz,
      vec_rsc_triosy_0_7_lz, vec_rsc_triosy_0_8_lz, vec_rsc_triosy_0_9_lz, vec_rsc_triosy_0_10_lz,
      vec_rsc_triosy_0_11_lz, vec_rsc_triosy_0_12_lz, vec_rsc_triosy_0_13_lz, vec_rsc_triosy_0_14_lz,
      vec_rsc_triosy_0_15_lz, p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz,
      vec_rsc_0_0_i_qa_d, vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_1_i_qa_d,
      vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_3_i_qa_d, vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_4_i_qa_d,
      vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_6_i_qa_d, vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_7_i_qa_d,
      vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_9_i_qa_d, vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_10_i_qa_d,
      vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_11_i_qa_d, vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_12_i_qa_d, vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_13_i_qa_d,
      vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      vec_rsc_0_15_i_qa_d, vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d, vec_rsc_0_0_i_adra_d_pff,
      vec_rsc_0_0_i_da_d_pff, vec_rsc_0_0_i_wea_d_pff, vec_rsc_0_1_i_wea_d_pff, vec_rsc_0_2_i_wea_d_pff,
      vec_rsc_0_3_i_wea_d_pff, vec_rsc_0_4_i_wea_d_pff, vec_rsc_0_5_i_wea_d_pff,
      vec_rsc_0_6_i_wea_d_pff, vec_rsc_0_7_i_wea_d_pff, vec_rsc_0_8_i_wea_d_pff,
      vec_rsc_0_9_i_wea_d_pff, vec_rsc_0_10_i_wea_d_pff, vec_rsc_0_11_i_wea_d_pff,
      vec_rsc_0_12_i_wea_d_pff, vec_rsc_0_13_i_wea_d_pff, vec_rsc_0_14_i_wea_d_pff,
      vec_rsc_0_15_i_wea_d_pff
);
  input clk;
  input rst;
  output vec_rsc_triosy_0_0_lz;
  output vec_rsc_triosy_0_1_lz;
  output vec_rsc_triosy_0_2_lz;
  output vec_rsc_triosy_0_3_lz;
  output vec_rsc_triosy_0_4_lz;
  output vec_rsc_triosy_0_5_lz;
  output vec_rsc_triosy_0_6_lz;
  output vec_rsc_triosy_0_7_lz;
  output vec_rsc_triosy_0_8_lz;
  output vec_rsc_triosy_0_9_lz;
  output vec_rsc_triosy_0_10_lz;
  output vec_rsc_triosy_0_11_lz;
  output vec_rsc_triosy_0_12_lz;
  output vec_rsc_triosy_0_13_lz;
  output vec_rsc_triosy_0_14_lz;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  input [63:0] vec_rsc_0_0_i_qa_d;
  output vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_1_i_qa_d;
  output vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_2_i_qa_d;
  output vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_3_i_qa_d;
  output vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_4_i_qa_d;
  output vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_5_i_qa_d;
  output vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_6_i_qa_d;
  output vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_7_i_qa_d;
  output vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_8_i_qa_d;
  output vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_9_i_qa_d;
  output vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_10_i_qa_d;
  output vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_11_i_qa_d;
  output vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_12_i_qa_d;
  output vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_13_i_qa_d;
  output vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_14_i_qa_d;
  output vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  input [63:0] vec_rsc_0_15_i_qa_d;
  output vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] vec_rsc_0_0_i_adra_d_pff;
  output [63:0] vec_rsc_0_0_i_da_d_pff;
  output vec_rsc_0_0_i_wea_d_pff;
  output vec_rsc_0_1_i_wea_d_pff;
  output vec_rsc_0_2_i_wea_d_pff;
  output vec_rsc_0_3_i_wea_d_pff;
  output vec_rsc_0_4_i_wea_d_pff;
  output vec_rsc_0_5_i_wea_d_pff;
  output vec_rsc_0_6_i_wea_d_pff;
  output vec_rsc_0_7_i_wea_d_pff;
  output vec_rsc_0_8_i_wea_d_pff;
  output vec_rsc_0_9_i_wea_d_pff;
  output vec_rsc_0_10_i_wea_d_pff;
  output vec_rsc_0_11_i_wea_d_pff;
  output vec_rsc_0_12_i_wea_d_pff;
  output vec_rsc_0_13_i_wea_d_pff;
  output vec_rsc_0_14_i_wea_d_pff;
  output vec_rsc_0_15_i_wea_d_pff;


  // Interconnect Declarations
  wire [63:0] p_rsci_idat;
  wire [63:0] r_rsci_idat;
  reg [63:0] modulo_result_rem_cmp_a;
  reg [63:0] modulo_result_rem_cmp_b;
  wire [63:0] modulo_result_rem_cmp_z;
  reg [64:0] operator_66_true_div_cmp_a;
  wire [64:0] operator_66_true_div_cmp_z;
  reg [9:0] operator_66_true_div_cmp_b_9_0;
  wire [10:0] fsm_output;
  wire nor_tmp_4;
  wire mux_tmp_14;
  wire not_tmp_39;
  wire or_tmp_68;
  wire not_tmp_49;
  wire mux_tmp_119;
  wire or_tmp_88;
  wire mux_tmp_130;
  wire mux_tmp_131;
  wire or_tmp_93;
  wire nand_tmp_4;
  wire or_tmp_94;
  wire mux_tmp_139;
  wire mux_tmp_141;
  wire or_tmp_96;
  wire mux_tmp_165;
  wire or_tmp_104;
  wire mux_tmp_214;
  wire mux_tmp_215;
  wire nand_tmp_7;
  wire mux_tmp_227;
  wire nor_tmp_23;
  wire mux_tmp_228;
  wire mux_tmp_231;
  wire mux_tmp_236;
  wire or_tmp_114;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire and_dcpl_4;
  wire and_dcpl_5;
  wire and_dcpl_6;
  wire not_tmp_90;
  wire or_tmp_167;
  wire nor_tmp_48;
  wire or_tmp_222;
  wire not_tmp_133;
  wire nor_tmp_82;
  wire or_tmp_258;
  wire and_dcpl_19;
  wire and_dcpl_26;
  wire and_dcpl_27;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_44;
  wire and_dcpl_48;
  wire and_dcpl_55;
  wire and_dcpl_59;
  wire not_tmp_208;
  wire and_dcpl_87;
  wire and_dcpl_88;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_98;
  wire and_dcpl_103;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire and_dcpl_111;
  wire and_dcpl_112;
  wire and_dcpl_113;
  wire and_dcpl_114;
  wire and_dcpl_115;
  wire and_dcpl_117;
  wire and_dcpl_118;
  wire or_tmp_453;
  wire mux_tmp_1082;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire and_dcpl_130;
  wire and_dcpl_135;
  wire and_dcpl_136;
  wire and_dcpl_139;
  wire and_dcpl_140;
  wire and_dcpl_144;
  wire and_dcpl_146;
  wire and_dcpl_147;
  wire and_dcpl_149;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_155;
  wire and_dcpl_162;
  wire and_dcpl_164;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_185;
  wire and_dcpl_189;
  wire and_dcpl_191;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_202;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_211;
  wire and_dcpl_219;
  wire and_dcpl_224;
  wire and_dcpl_226;
  wire and_dcpl_231;
  wire not_tmp_248;
  wire mux_tmp_1116;
  wire or_tmp_532;
  wire not_tmp_253;
  wire mux_tmp_1180;
  wire or_tmp_643;
  wire mux_tmp_1244;
  wire or_tmp_756;
  wire mux_tmp_1308;
  wire or_tmp_866;
  wire mux_tmp_1372;
  wire or_tmp_974;
  wire mux_tmp_1436;
  wire or_tmp_1085;
  wire mux_tmp_1500;
  wire or_tmp_1198;
  wire mux_tmp_1564;
  wire or_tmp_1308;
  wire not_tmp_318;
  wire mux_tmp_1628;
  wire or_tmp_1416;
  wire mux_tmp_1692;
  wire or_tmp_1527;
  wire mux_tmp_1756;
  wire or_tmp_1640;
  wire mux_tmp_1820;
  wire or_tmp_1750;
  wire not_tmp_357;
  wire mux_tmp_1884;
  wire or_tmp_1858;
  wire mux_tmp_1948;
  wire or_tmp_1969;
  wire not_tmp_377;
  wire mux_tmp_2012;
  wire or_tmp_2082;
  wire not_tmp_387;
  wire mux_tmp_2076;
  wire not_tmp_390;
  wire or_tmp_2192;
  wire nor_tmp_265;
  wire and_dcpl_235;
  wire and_dcpl_236;
  wire and_dcpl_237;
  wire or_tmp_2274;
  wire or_tmp_2276;
  wire or_tmp_2277;
  wire or_tmp_2280;
  wire or_tmp_2281;
  wire mux_tmp_2159;
  wire or_tmp_2294;
  wire mux_tmp_2172;
  wire or_tmp_2297;
  wire mux_tmp_2176;
  wire mux_tmp_2178;
  wire or_tmp_2302;
  wire mux_tmp_2235;
  wire mux_tmp_2241;
  wire or_tmp_2340;
  wire or_tmp_2341;
  wire mux_tmp_2262;
  wire mux_tmp_2287;
  wire mux_tmp_2289;
  wire mux_tmp_2293;
  wire or_tmp_2360;
  wire mux_tmp_2311;
  wire or_tmp_2376;
  wire or_tmp_2389;
  wire mux_tmp_2347;
  wire or_tmp_2390;
  wire mux_tmp_2348;
  wire mux_tmp_2350;
  wire not_tmp_431;
  wire mux_tmp_2353;
  wire or_tmp_2393;
  wire or_tmp_2394;
  wire mux_tmp_2355;
  wire mux_tmp_2356;
  wire or_tmp_2396;
  wire or_tmp_2397;
  wire or_tmp_2399;
  wire mux_tmp_2359;
  wire mux_tmp_2361;
  wire mux_tmp_2363;
  wire mux_tmp_2364;
  wire or_tmp_2404;
  wire mux_tmp_2365;
  wire nand_tmp_54;
  wire or_tmp_2405;
  wire mux_tmp_2369;
  wire mux_tmp_2370;
  wire mux_tmp_2371;
  wire mux_tmp_2376;
  wire mux_tmp_2377;
  wire mux_tmp_2378;
  wire mux_tmp_2382;
  wire or_tmp_2407;
  wire mux_tmp_2386;
  wire mux_tmp_2389;
  wire mux_tmp_2424;
  wire not_tmp_441;
  wire or_tmp_2436;
  wire not_tmp_446;
  wire and_dcpl_241;
  wire and_dcpl_245;
  wire and_dcpl_247;
  wire nor_tmp_324;
  wire or_tmp_2474;
  wire mux_tmp_2640;
  wire mux_tmp_2659;
  wire and_dcpl_256;
  wire mux_tmp_2669;
  wire mux_tmp_2672;
  wire mux_tmp_2675;
  wire not_tmp_500;
  wire mux_tmp_2682;
  wire mux_tmp_2690;
  wire mux_tmp_2691;
  wire mux_tmp_2693;
  wire or_tmp_2603;
  wire or_tmp_2604;
  wire mux_tmp_2700;
  wire mux_tmp_2702;
  wire mux_tmp_2703;
  wire mux_tmp_2706;
  wire mux_tmp_2709;
  wire mux_tmp_2715;
  wire mux_tmp_2736;
  wire and_dcpl_257;
  wire and_dcpl_260;
  wire and_dcpl_262;
  wire and_dcpl_270;
  wire and_dcpl_278;
  wire and_dcpl_280;
  wire mux_tmp_2745;
  wire mux_tmp_2760;
  wire or_tmp_2651;
  wire or_tmp_2682;
  wire or_tmp_2683;
  wire or_tmp_2690;
  wire or_tmp_2693;
  wire or_tmp_2696;
  wire or_tmp_2697;
  wire mux_tmp_2796;
  wire or_tmp_2701;
  wire or_tmp_2703;
  wire or_tmp_2704;
  wire or_tmp_2706;
  wire or_tmp_2709;
  wire or_tmp_2714;
  wire mux_tmp_2841;
  wire or_tmp_2729;
  wire or_tmp_2731;
  wire mux_tmp_2843;
  wire mux_tmp_2844;
  wire or_tmp_2734;
  wire mux_tmp_2848;
  wire mux_tmp_2850;
  wire or_tmp_2736;
  wire mux_tmp_2851;
  wire mux_tmp_2856;
  wire nand_tmp_67;
  wire mux_tmp_2862;
  wire mux_tmp_2863;
  wire or_tmp_2739;
  wire mux_tmp_2867;
  wire or_tmp_2740;
  wire mux_tmp_2876;
  wire mux_tmp_2878;
  wire mux_tmp_2879;
  wire or_tmp_2742;
  wire mux_tmp_2880;
  wire mux_tmp_2886;
  wire mux_tmp_2888;
  wire mux_tmp_2890;
  wire or_tmp_2743;
  wire nand_tmp_68;
  wire mux_tmp_2895;
  wire or_tmp_2745;
  wire or_tmp_2746;
  wire nand_tmp_69;
  wire mux_tmp_2906;
  wire mux_tmp_2910;
  wire nand_tmp_70;
  wire mux_tmp_2912;
  wire nand_tmp_71;
  wire mux_tmp_2916;
  wire mux_tmp_2920;
  wire or_tmp_2749;
  wire or_tmp_2774;
  wire mux_tmp_2996;
  wire not_tmp_557;
  wire nor_tmp_405;
  wire mux_tmp_3007;
  wire mux_tmp_3008;
  wire or_tmp_2791;
  wire mux_tmp_3014;
  wire or_tmp_2795;
  wire or_tmp_2802;
  wire or_tmp_2803;
  wire mux_tmp_3024;
  wire mux_tmp_3032;
  wire mux_tmp_3049;
  wire or_tmp_2814;
  wire nor_tmp_410;
  wire and_dcpl_304;
  wire not_tmp_619;
  wire mux_tmp_3329;
  wire nor_tmp_457;
  wire mux_tmp_3341;
  wire mux_tmp_3343;
  wire mux_tmp_3361;
  wire or_tmp_2988;
  wire mux_tmp_3378;
  wire not_tmp_647;
  wire mux_tmp_3410;
  wire mux_tmp_3414;
  wire mux_tmp_3415;
  wire mux_tmp_3417;
  wire or_tmp_3023;
  wire mux_tmp_3418;
  wire mux_tmp_3420;
  wire mux_tmp_3421;
  wire mux_tmp_3423;
  wire mux_tmp_3424;
  wire mux_tmp_3425;
  wire not_tmp_663;
  wire mux_tmp_3429;
  wire mux_tmp_3432;
  wire mux_tmp_3434;
  wire mux_tmp_3435;
  wire not_tmp_665;
  wire mux_tmp_3453;
  wire mux_tmp_3456;
  wire mux_tmp_3457;
  wire mux_tmp_3458;
  wire mux_tmp_3459;
  wire not_tmp_672;
  wire mux_tmp_3463;
  wire mux_tmp_3464;
  wire mux_tmp_3472;
  wire mux_tmp_3473;
  wire mux_tmp_3474;
  wire mux_tmp_3477;
  wire mux_tmp_3481;
  wire mux_tmp_3491;
  wire not_tmp_688;
  wire or_tmp_3053;
  wire mux_tmp_3529;
  wire not_tmp_701;
  wire or_tmp_3095;
  wire mux_tmp_3547;
  wire mux_tmp_3551;
  wire mux_tmp_3574;
  wire mux_tmp_3576;
  wire mux_tmp_3577;
  wire mux_tmp_3618;
  wire or_tmp_3135;
  wire mux_tmp_3632;
  wire or_tmp_3176;
  wire or_tmp_3190;
  wire mux_tmp_3673;
  wire mux_tmp_3674;
  wire mux_tmp_3679;
  wire mux_tmp_3681;
  wire and_tmp_28;
  wire mux_tmp_3691;
  wire or_tmp_3224;
  wire mux_tmp_3698;
  wire mux_tmp_3701;
  wire mux_tmp_3705;
  wire mux_tmp_3720;
  wire mux_tmp_3724;
  wire mux_tmp_3736;
  wire mux_tmp_3737;
  wire mux_tmp_3739;
  wire mux_tmp_3753;
  reg COMP_LOOP_COMP_LOOP_and_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_10_itm;
  reg COMP_LOOP_nor_11_itm;
  wire [11:0] COMP_LOOP_acc_1_cse_6_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_6_sva_1;
  reg [11:0] VEC_LOOP_j_sva_11_0;
  reg [4:0] COMP_LOOP_k_9_4_sva_4_0;
  reg COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  reg COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  reg [11:0] COMP_LOOP_acc_10_cse_12_1_1_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_14_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_14_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_2_sva;
  reg [10:0] COMP_LOOP_acc_14_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_14_psp_sva;
  reg [10:0] COMP_LOOP_acc_17_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_17_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_6_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_10_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_10_sva;
  reg [10:0] COMP_LOOP_acc_11_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_11_psp_sva;
  reg [10:0] COMP_LOOP_acc_20_psp_sva;
  wire [11:0] nl_COMP_LOOP_acc_20_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_4_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_sva;
  reg [9:0] COMP_LOOP_acc_19_psp_sva;
  reg [8:0] COMP_LOOP_acc_16_psp_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_8_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_8_sva;
  reg [11:0] COMP_LOOP_acc_1_cse_12_sva;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_12_sva;
  reg [9:0] COMP_LOOP_acc_13_psp_sva;
  reg [63:0] tmp_10_lpi_4_dfm;
  wire [11:0] COMP_LOOP_acc_1_cse_2_sva_1;
  wire [12:0] nl_COMP_LOOP_acc_1_cse_2_sva_1;
  wire mux_2771_m1c;
  wire and_279_m1c;
  wire and_281_m1c;
  wire and_284_m1c;
  wire and_286_m1c;
  wire and_288_m1c;
  wire and_291_m1c;
  wire and_292_m1c;
  wire and_295_m1c;
  wire and_297_m1c;
  wire and_299_m1c;
  wire and_302_m1c;
  wire and_304_m1c;
  wire and_307_m1c;
  wire and_309_m1c;
  wire and_311_m1c;
  wire and_273_m1c;
  wire nor_1445_cse;
  wire mux_1157_cse;
  wire nand_332_cse;
  wire mux_1413_cse;
  wire nand_324_cse;
  wire mux_1669_cse;
  wire mux_1925_cse;
  reg reg_vec_rsc_triosy_0_15_obj_ld_cse;
  wire and_527_cse;
  wire or_2377_cse;
  wire or_2368_cse;
  wire and_529_cse;
  wire and_526_cse;
  wire or_3388_cse;
  wire nor_758_cse;
  wire nand_196_cse;
  wire or_2419_cse;
  wire nor_297_cse;
  wire nor_303_cse;
  wire mux_125_cse;
  wire nand_356_cse;
  wire or_491_cse;
  wire nand_357_cse;
  wire nand_358_cse;
  wire or_2921_cse;
  wire or_2918_cse;
  wire and_536_cse;
  wire nor_753_cse;
  wire nand_159_cse;
  wire or_2387_cse;
  wire or_2912_cse;
  wire mux_554_cse;
  wire or_181_cse;
  wire and_458_cse;
  wire and_407_cse;
  wire or_3039_cse;
  wire and_459_cse;
  wire or_2644_cse;
  wire or_470_cse;
  wire and_672_cse;
  wire and_395_cse;
  wire and_676_cse;
  wire or_361_cse;
  wire or_2414_cse;
  wire or_3063_cse;
  wire and_756_cse;
  wire nand_142_cse;
  wire and_366_cse;
  wire and_350_cse;
  wire or_3427_cse;
  wire or_2991_cse;
  wire nand_138_cse;
  wire or_2407_cse;
  wire or_2998_cse;
  wire or_469_cse;
  wire and_757_cse;
  wire nor_609_cse;
  wire or_352_cse;
  wire and_404_cse;
  wire and_707_cse;
  wire or_259_cse;
  wire nor_1580_cse;
  wire or_586_cse;
  wire or_591_cse;
  wire nand_334_cse;
  wire or_702_cse;
  wire nor_209_cse;
  wire nand_337_cse;
  wire or_1028_cse;
  wire nor_223_cse;
  wire or_1470_cse;
  wire nor_239_cse;
  wire or_1912_cse;
  wire and_564_cse;
  wire mux_2926_cse;
  wire mux_2486_cse;
  wire or_2540_cse;
  wire nor_694_cse;
  wire or_70_cse;
  wire or_56_cse;
  wire nor_657_cse;
  wire nand_367_cse;
  wire or_2947_cse;
  wire or_2905_cse;
  wire or_3079_cse;
  wire and_524_cse;
  wire or_3074_cse;
  wire nand_183_cse;
  wire nor_667_cse;
  wire or_163_cse;
  wire or_3417_cse;
  wire and_465_cse;
  wire mux_1149_cse;
  wire mux_1277_cse;
  wire mux_1405_cse;
  wire mux_1533_cse;
  wire mux_1661_cse;
  wire mux_1789_cse;
  wire mux_1917_cse;
  wire mux_2045_cse;
  wire nor_697_cse;
  wire nor_653_cse;
  wire mux_3254_cse;
  wire mux_3555_cse;
  wire or_3008_cse;
  wire mux_155_cse;
  wire mux_171_cse;
  wire mux_1036_cse;
  wire mux_981_cse;
  wire nand_386_cse;
  wire mux_2465_cse;
  wire or_2528_cse;
  wire or_2534_cse;
  wire nand_173_cse;
  wire or_2541_cse;
  wire mux_2516_cse;
  wire mux_2494_cse;
  wire mux_2515_cse;
  wire mux_544_cse;
  wire mux_2171_cse;
  wire mux_2203_cse;
  wire mux_3281_cse;
  wire mux_648_cse;
  wire mux_2998_cse;
  wire or_2835_cse;
  wire mux_259_cse;
  wire mux_3245_cse;
  wire mux_498_cse;
  wire mux_161_cse;
  wire mux_340_cse;
  wire mux_375_cse;
  wire mux_2643_cse;
  wire [7:0] COMP_LOOP_acc_psp_sva_1;
  wire [8:0] nl_COMP_LOOP_acc_psp_sva_1;
  reg [7:0] COMP_LOOP_acc_psp_sva;
  reg [63:0] COMP_LOOP_10_mul_mut;
  wire mux_2698_itm;
  wire mux_2757_itm;
  wire mux_2840_itm;
  wire mux_3485_itm;
  wire mux_3494_itm;
  wire and_dcpl_332;
  wire [12:0] z_out;
  wire [13:0] nl_z_out;
  wire and_dcpl_333;
  wire and_dcpl_338;
  wire and_dcpl_340;
  wire and_dcpl_342;
  wire and_dcpl_344;
  wire and_dcpl_345;
  wire and_dcpl_349;
  wire and_dcpl_350;
  wire and_dcpl_356;
  wire and_dcpl_359;
  wire [64:0] z_out_1;
  wire [65:0] nl_z_out_1;
  wire and_dcpl_367;
  wire and_dcpl_371;
  wire and_dcpl_383;
  wire and_dcpl_390;
  wire and_dcpl_393;
  wire and_dcpl_403;
  wire and_dcpl_411;
  wire and_dcpl_412;
  wire and_dcpl_422;
  wire and_dcpl_428;
  wire and_dcpl_432;
  wire and_dcpl_446;
  wire and_dcpl_453;
  wire and_dcpl_460;
  wire and_dcpl_468;
  wire and_dcpl_472;
  wire and_dcpl_473;
  wire and_dcpl_475;
  wire and_dcpl_481;
  wire and_dcpl_486;
  wire and_dcpl_488;
  wire and_dcpl_493;
  wire and_dcpl_494;
  wire and_dcpl_495;
  wire and_dcpl_500;
  wire and_dcpl_503;
  wire and_dcpl_505;
  wire and_dcpl_507;
  wire and_dcpl_510;
  wire and_dcpl_513;
  wire [9:0] z_out_3;
  wire and_dcpl_531;
  wire and_dcpl_539;
  wire and_dcpl_540;
  wire and_dcpl_544;
  wire and_dcpl_551;
  wire and_dcpl_553;
  wire and_dcpl_557;
  wire and_dcpl_561;
  wire [9:0] z_out_4;
  wire [10:0] nl_z_out_4;
  wire and_dcpl_567;
  wire and_dcpl_568;
  wire and_dcpl_569;
  wire and_dcpl_594;
  wire [9:0] z_out_5;
  wire [10:0] nl_z_out_5;
  wire and_dcpl_627;
  wire and_dcpl_628;
  wire and_dcpl_631;
  wire and_dcpl_636;
  wire and_dcpl_642;
  wire or_tmp_3282;
  wire not_tmp_834;
  wire not_tmp_835;
  wire not_tmp_838;
  wire and_dcpl_647;
  wire and_dcpl_650;
  wire [64:0] z_out_6;
  wire and_dcpl_660;
  wire and_dcpl_669;
  wire and_dcpl_678;
  wire and_dcpl_686;
  wire [6:0] z_out_7;
  wire or_tmp_3307;
  wire or_tmp_3312;
  wire or_tmp_3326;
  wire [63:0] z_out_8;
  wire signed [128:0] nl_z_out_8;
  reg [63:0] p_sva;
  reg [63:0] r_sva;
  reg [3:0] STAGE_LOOP_i_3_0_sva;
  reg [9:0] STAGE_LOOP_lshift_psp_sva;
  reg [63:0] modExp_result_sva;
  reg modExp_exp_1_7_1_sva;
  reg modExp_exp_1_6_1_sva;
  reg modExp_exp_1_5_1_sva;
  reg modExp_exp_1_4_1_sva;
  reg COMP_LOOP_COMP_LOOP_nor_itm;
  reg COMP_LOOP_COMP_LOOP_and_2_itm;
  reg COMP_LOOP_COMP_LOOP_and_4_itm;
  reg COMP_LOOP_COMP_LOOP_and_5_itm;
  reg COMP_LOOP_COMP_LOOP_and_6_itm;
  reg COMP_LOOP_COMP_LOOP_and_8_itm;
  reg COMP_LOOP_COMP_LOOP_and_9_itm;
  reg COMP_LOOP_COMP_LOOP_and_11_itm;
  reg COMP_LOOP_COMP_LOOP_and_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_13_itm;
  reg COMP_LOOP_COMP_LOOP_and_14_itm;
  reg COMP_LOOP_COMP_LOOP_nor_1_itm;
  reg COMP_LOOP_nor_12_itm;
  reg COMP_LOOP_COMP_LOOP_and_62_itm;
  reg COMP_LOOP_COMP_LOOP_and_64_itm;
  reg COMP_LOOP_COMP_LOOP_and_68_itm;
  reg COMP_LOOP_COMP_LOOP_and_139_itm;
  reg COMP_LOOP_COMP_LOOP_and_140_itm;
  reg COMP_LOOP_COMP_LOOP_and_141_itm;
  reg COMP_LOOP_COMP_LOOP_and_143_itm;
  reg COMP_LOOP_COMP_LOOP_and_144_itm;
  reg COMP_LOOP_COMP_LOOP_and_145_itm;
  reg COMP_LOOP_COMP_LOOP_and_146_itm;
  reg COMP_LOOP_COMP_LOOP_and_147_itm;
  reg COMP_LOOP_COMP_LOOP_and_148_itm;
  reg COMP_LOOP_COMP_LOOP_and_149_itm;
  reg COMP_LOOP_nor_134_itm;
  reg COMP_LOOP_nor_137_itm;
  reg COMP_LOOP_COMP_LOOP_and_305_itm;
  reg [63:0] COMP_LOOP_10_acc_8_itm;
  wire STAGE_LOOP_i_3_0_sva_mx0c1;
  wire [3:0] STAGE_LOOP_i_3_0_sva_2;
  wire [4:0] nl_STAGE_LOOP_i_3_0_sva_2;
  wire [63:0] COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [64:0] nl_COMP_LOOP_1_acc_5_mut_mx0w5;
  wire [63:0] COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
  wire signed [127:0] nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1;
  wire [9:0] STAGE_LOOP_lshift_psp_sva_mx0w0;
  wire VEC_LOOP_j_sva_11_0_mx0c1;
  wire modExp_result_sva_mx0c0;
  wire [62:0] operator_64_false_slc_modExp_exp_63_1_3;
  wire [63:0] modulo_qr_sva_1_mx0w6;
  wire [64:0] nl_modulo_qr_sva_1_mx0w6;
  wire modExp_while_and_3;
  wire modExp_while_and_5;
  wire and_317_m1c;
  wire modExp_result_and_rgt;
  wire modExp_result_and_1_rgt;
  wire and_978_ssc;
  wire COMP_LOOP_or_32_cse;
  wire or_80_cse;
  wire and_816_cse;
  wire and_815_cse;
  wire and_825_cse;
  wire nor_1670_cse;
  wire and_824_ssc;
  wire COMP_LOOP_or_54_ssc;
  wire COMP_LOOP_or_55_ssc;
  wire and_872_ssc;
  wire and_820_cse;
  wire and_830_cse;
  wire and_842_cse;
  wire and_849_cse;
  wire and_870_cse;
  wire and_873_cse;
  wire and_827_cse;
  wire and_835_cse;
  wire mux_tmp_3828;
  wire mux_tmp_3830;
  wire nor_tmp_549;
  wire or_tmp_3337;
  wire or_tmp_3339;
  wire mux_tmp_3839;
  wire mux_tmp_3841;
  wire or_tmp_3344;
  wire nor_tmp_552;
  wire or_tmp_3347;
  wire mux_tmp_3848;
  wire nor_tmp_554;
  wire or_tmp_3352;
  wire mux_tmp_3856;
  wire mux_tmp_3864;
  wire or_tmp_3357;
  wire or_tmp_3381;
  wire or_tmp_3382;
  wire or_tmp_3384;
  wire mux_tmp_3892;
  wire not_tmp_882;
  wire not_tmp_883;
  wire or_tmp_3402;
  wire mux_tmp_3903;
  wire or_tmp_3403;
  wire mux_tmp_3906;
  wire mux_tmp_3907;
  wire or_tmp_3409;
  wire [64:0] operator_64_false_mux1h_2_rgt;
  reg operator_64_false_acc_mut_64;
  reg [63:0] operator_64_false_acc_mut_63_0;
  wire or_2914_cse;
  wire or_2400_cse;
  wire and_521_cse;
  wire nor_1704_cse;
  wire or_2855_cse;
  wire or_2965_cse;
  wire mux_3935_cse;
  wire or_3532_cse;
  wire or_2421_cse;
  wire COMP_LOOP_or_61_itm;
  wire COMP_LOOP_or_24_itm;
  wire COMP_LOOP_nor_633_itm;
  wire COMP_LOOP_nor_685_itm;
  wire COMP_LOOP_or_65_itm;
  wire COMP_LOOP_nor_687_itm;
  wire STAGE_LOOP_acc_itm_2_1;
  wire [11:0] z_out_2_12_1;
  wire nor_1657_cse;

  wire[0:0] or_651_nl;
  wire[0:0] or_650_nl;
  wire[0:0] or_638_nl;
  wire[0:0] or_637_nl;
  wire[0:0] or_859_nl;
  wire[0:0] or_858_nl;
  wire[0:0] or_1093_nl;
  wire[0:0] or_1092_nl;
  wire[0:0] or_1080_nl;
  wire[0:0] or_1079_nl;
  wire[0:0] or_1301_nl;
  wire[0:0] or_1300_nl;
  wire[0:0] or_1535_nl;
  wire[0:0] or_1534_nl;
  wire[0:0] or_1522_nl;
  wire[0:0] or_1521_nl;
  wire[0:0] or_1743_nl;
  wire[0:0] or_1742_nl;
  wire[0:0] nand_259_nl;
  wire[0:0] or_1976_nl;
  wire[0:0] or_1964_nl;
  wire[0:0] or_1963_nl;
  wire[0:0] nand_231_nl;
  wire[0:0] or_2184_nl;
  wire[0:0] nor_1584_nl;
  wire[0:0] and_739_nl;
  wire[0:0] modulo_result_or_nl;
  wire[0:0] mux_2231_nl;
  wire[0:0] mux_2230_nl;
  wire[0:0] mux_2229_nl;
  wire[0:0] mux_2228_nl;
  wire[0:0] mux_2227_nl;
  wire[0:0] mux_2226_nl;
  wire[0:0] mux_2225_nl;
  wire[0:0] mux_2224_nl;
  wire[0:0] nand_195_nl;
  wire[0:0] mux_2223_nl;
  wire[0:0] mux_2222_nl;
  wire[0:0] mux_2221_nl;
  wire[0:0] or_2375_nl;
  wire[0:0] mux_2220_nl;
  wire[0:0] mux_2219_nl;
  wire[0:0] mux_2218_nl;
  wire[0:0] mux_2217_nl;
  wire[0:0] mux_2216_nl;
  wire[0:0] or_2373_nl;
  wire[0:0] or_2371_nl;
  wire[0:0] mux_2215_nl;
  wire[0:0] mux_2214_nl;
  wire[0:0] mux_2213_nl;
  wire[0:0] mux_2212_nl;
  wire[0:0] mux_2211_nl;
  wire[0:0] mux_2210_nl;
  wire[0:0] mux_2209_nl;
  wire[0:0] or_2367_nl;
  wire[0:0] mux_2208_nl;
  wire[0:0] mux_2207_nl;
  wire[0:0] mux_2206_nl;
  wire[0:0] mux_2205_nl;
  wire[0:0] mux_2204_nl;
  wire[0:0] mux_2202_nl;
  wire[0:0] mux_2201_nl;
  wire[0:0] mux_2200_nl;
  wire[0:0] or_2364_nl;
  wire[0:0] mux_2199_nl;
  wire[0:0] mux_2198_nl;
  wire[0:0] mux_2197_nl;
  wire[0:0] or_2362_nl;
  wire[0:0] or_2360_nl;
  wire[0:0] mux_2196_nl;
  wire[0:0] mux_2195_nl;
  wire[0:0] mux_2194_nl;
  wire[0:0] mux_2193_nl;
  wire[0:0] mux_2192_nl;
  wire[0:0] mux_2191_nl;
  wire[0:0] mux_2190_nl;
  wire[0:0] mux_2189_nl;
  wire[0:0] mux_2188_nl;
  wire[0:0] mux_2187_nl;
  wire[0:0] mux_2186_nl;
  wire[0:0] mux_2185_nl;
  wire[0:0] mux_2184_nl;
  wire[0:0] mux_2183_nl;
  wire[0:0] mux_2182_nl;
  wire[0:0] mux_2181_nl;
  wire[0:0] mux_2180_nl;
  wire[0:0] mux_2179_nl;
  wire[0:0] or_2357_nl;
  wire[0:0] mux_2177_nl;
  wire[0:0] or_2355_nl;
  wire[0:0] mux_2174_nl;
  wire[0:0] mux_2173_nl;
  wire[0:0] mux_2170_nl;
  wire[0:0] mux_2169_nl;
  wire[0:0] or_2351_nl;
  wire[0:0] mux_2168_nl;
  wire[0:0] mux_2167_nl;
  wire[0:0] or_2347_nl;
  wire[0:0] mux_2166_nl;
  wire[0:0] mux_2165_nl;
  wire[0:0] mux_2164_nl;
  wire[0:0] mux_2163_nl;
  wire[0:0] mux_2162_nl;
  wire[0:0] mux_2161_nl;
  wire[0:0] mux_2160_nl;
  wire[0:0] or_2343_nl;
  wire[0:0] mux_2158_nl;
  wire[0:0] mux_2157_nl;
  wire[0:0] mux_2156_nl;
  wire[0:0] mux_2155_nl;
  wire[0:0] mux_2154_nl;
  wire[0:0] mux_2153_nl;
  wire[0:0] mux_2152_nl;
  wire[0:0] mux_2151_nl;
  wire[0:0] mux_2150_nl;
  wire[0:0] mux_2149_nl;
  wire[0:0] mux_2148_nl;
  wire[0:0] mux_2147_nl;
  wire[0:0] mux_2146_nl;
  wire[0:0] or_2339_nl;
  wire[0:0] mux_2144_nl;
  wire[0:0] mux_2143_nl;
  wire[0:0] mux_2142_nl;
  wire[0:0] mux_2141_nl;
  wire[0:0] mux_2140_nl;
  wire[0:0] mux_2139_nl;
  wire[0:0] or_2335_nl;
  wire[0:0] mux_2138_nl;
  wire[0:0] mux_2137_nl;
  wire[0:0] mux_2136_nl;
  wire[0:0] nand_197_nl;
  wire[0:0] mux_2135_nl;
  wire[0:0] mux_2134_nl;
  wire[0:0] mux_2133_nl;
  wire[0:0] mux_2331_nl;
  wire[0:0] mux_2330_nl;
  wire[0:0] mux_2329_nl;
  wire[0:0] mux_2328_nl;
  wire[0:0] mux_2327_nl;
  wire[0:0] mux_2326_nl;
  wire[0:0] mux_2325_nl;
  wire[0:0] mux_2324_nl;
  wire[0:0] mux_2323_nl;
  wire[0:0] mux_2322_nl;
  wire[0:0] and_519_nl;
  wire[0:0] mux_2321_nl;
  wire[0:0] mux_2320_nl;
  wire[0:0] mux_2319_nl;
  wire[0:0] mux_2318_nl;
  wire[0:0] mux_2317_nl;
  wire[0:0] mux_2316_nl;
  wire[0:0] mux_2315_nl;
  wire[0:0] mux_2314_nl;
  wire[0:0] mux_2313_nl;
  wire[0:0] mux_2312_nl;
  wire[0:0] mux_2310_nl;
  wire[0:0] mux_2309_nl;
  wire[0:0] or_2418_nl;
  wire[0:0] mux_2308_nl;
  wire[0:0] mux_2307_nl;
  wire[0:0] mux_2306_nl;
  wire[0:0] mux_2305_nl;
  wire[0:0] mux_2304_nl;
  wire[0:0] mux_2303_nl;
  wire[0:0] mux_2302_nl;
  wire[0:0] mux_2301_nl;
  wire[0:0] mux_2300_nl;
  wire[0:0] mux_2299_nl;
  wire[0:0] mux_2298_nl;
  wire[0:0] mux_2297_nl;
  wire[0:0] mux_2296_nl;
  wire[0:0] mux_2295_nl;
  wire[0:0] mux_2294_nl;
  wire[0:0] or_2408_nl;
  wire[0:0] mux_2292_nl;
  wire[0:0] mux_2291_nl;
  wire[0:0] mux_2290_nl;
  wire[0:0] mux_2288_nl;
  wire[0:0] mux_2286_nl;
  wire[0:0] mux_2285_nl;
  wire[0:0] or_2406_nl;
  wire[0:0] or_2404_nl;
  wire[0:0] mux_2284_nl;
  wire[0:0] mux_2283_nl;
  wire[0:0] mux_2282_nl;
  wire[0:0] mux_2281_nl;
  wire[0:0] mux_2280_nl;
  wire[0:0] or_2403_nl;
  wire[0:0] mux_2279_nl;
  wire[0:0] mux_2278_nl;
  wire[0:0] or_2402_nl;
  wire[0:0] mux_2277_nl;
  wire[0:0] mux_2276_nl;
  wire[0:0] mux_2275_nl;
  wire[0:0] mux_2274_nl;
  wire[0:0] mux_2273_nl;
  wire[0:0] mux_2272_nl;
  wire[0:0] nor_295_nl;
  wire[0:0] mux_2271_nl;
  wire[0:0] mux_2270_nl;
  wire[0:0] mux_2269_nl;
  wire[0:0] mux_2268_nl;
  wire[0:0] mux_2267_nl;
  wire[0:0] or_2398_nl;
  wire[0:0] mux_2266_nl;
  wire[0:0] mux_2265_nl;
  wire[0:0] mux_2264_nl;
  wire[0:0] mux_2263_nl;
  wire[0:0] mux_2261_nl;
  wire[0:0] mux_2260_nl;
  wire[0:0] mux_2259_nl;
  wire[0:0] or_2395_nl;
  wire[0:0] mux_2257_nl;
  wire[0:0] mux_2256_nl;
  wire[0:0] mux_2255_nl;
  wire[0:0] mux_2254_nl;
  wire[0:0] mux_2253_nl;
  wire[0:0] mux_2251_nl;
  wire[0:0] mux_2250_nl;
  wire[0:0] mux_2249_nl;
  wire[0:0] or_2392_nl;
  wire[0:0] mux_2248_nl;
  wire[0:0] mux_2247_nl;
  wire[0:0] mux_2246_nl;
  wire[0:0] mux_2245_nl;
  wire[0:0] or_2390_nl;
  wire[0:0] mux_2244_nl;
  wire[0:0] or_2385_nl;
  wire[0:0] mux_2243_nl;
  wire[0:0] mux_2237_nl;
  wire[0:0] nand_51_nl;
  wire[0:0] mux_2236_nl;
  wire[0:0] mux_2346_nl;
  wire[0:0] mux_2345_nl;
  wire[0:0] mux_2344_nl;
  wire[0:0] nand_189_nl;
  wire[0:0] mux_2343_nl;
  wire[0:0] and_517_nl;
  wire[0:0] nor_752_nl;
  wire[0:0] mux_2341_nl;
  wire[0:0] or_3386_nl;
  wire[0:0] nand_190_nl;
  wire[0:0] or_2438_nl;
  wire[0:0] mux_2340_nl;
  wire[0:0] or_2437_nl;
  wire[0:0] mux_2339_nl;
  wire[0:0] mux_2338_nl;
  wire[0:0] mux_2337_nl;
  wire[0:0] mux_2336_nl;
  wire[0:0] mux_2335_nl;
  wire[0:0] or_2435_nl;
  wire[0:0] or_2433_nl;
  wire[0:0] or_2431_nl;
  wire[0:0] or_2430_nl;
  wire[0:0] mux_2334_nl;
  wire[0:0] nand_191_nl;
  wire[0:0] mux_2333_nl;
  wire[0:0] or_2427_nl;
  wire[0:0] or_2426_nl;
  wire[0:0] mux_2418_nl;
  wire[0:0] mux_2417_nl;
  wire[0:0] mux_2416_nl;
  wire[0:0] mux_2415_nl;
  wire[0:0] mux_2414_nl;
  wire[0:0] mux_2413_nl;
  wire[0:0] mux_2412_nl;
  wire[0:0] mux_2411_nl;
  wire[0:0] mux_2410_nl;
  wire[0:0] mux_2409_nl;
  wire[0:0] mux_2408_nl;
  wire[0:0] mux_2407_nl;
  wire[0:0] mux_2406_nl;
  wire[0:0] mux_2405_nl;
  wire[0:0] mux_2404_nl;
  wire[0:0] mux_2403_nl;
  wire[0:0] mux_2402_nl;
  wire[0:0] mux_2401_nl;
  wire[0:0] mux_2400_nl;
  wire[0:0] mux_2399_nl;
  wire[0:0] mux_2398_nl;
  wire[0:0] mux_2397_nl;
  wire[0:0] mux_2396_nl;
  wire[0:0] mux_2395_nl;
  wire[0:0] mux_2394_nl;
  wire[0:0] mux_2393_nl;
  wire[0:0] mux_2392_nl;
  wire[0:0] mux_2391_nl;
  wire[0:0] mux_2390_nl;
  wire[0:0] mux_2384_nl;
  wire[0:0] mux_2383_nl;
  wire[0:0] mux_2381_nl;
  wire[0:0] mux_2380_nl;
  wire[0:0] mux_2379_nl;
  wire[0:0] mux_2374_nl;
  wire[0:0] mux_2373_nl;
  wire[0:0] mux_2372_nl;
  wire[0:0] mux_2368_nl;
  wire[0:0] mux_2367_nl;
  wire[0:0] mux_2366_nl;
  wire[0:0] mux_2362_nl;
  wire[0:0] mux_2360_nl;
  wire[0:0] mux_2358_nl;
  wire[0:0] mux_2357_nl;
  wire[0:0] mux_2354_nl;
  wire[0:0] mux_2351_nl;
  wire[0:0] mux_2349_nl;
  wire[0:0] mux_2452_nl;
  wire[0:0] mux_2451_nl;
  wire[0:0] mux_2450_nl;
  wire[0:0] mux_2449_nl;
  wire[0:0] or_3396_nl;
  wire[0:0] nand_175_nl;
  wire[63:0] modExp_while_if_mux1h_nl;
  wire[0:0] and_323_nl;
  wire[0:0] mux_3257_nl;
  wire[0:0] mux_3256_nl;
  wire[0:0] nor_640_nl;
  wire[0:0] mux_3255_nl;
  wire[0:0] or_2920_nl;
  wire[0:0] mux_3253_nl;
  wire[0:0] and_421_nl;
  wire[0:0] mux_3252_nl;
  wire[0:0] nor_641_nl;
  wire[0:0] mux_3251_nl;
  wire[0:0] nand_85_nl;
  wire[0:0] mux_3250_nl;
  wire[0:0] nor_642_nl;
  wire[0:0] nor_643_nl;
  wire[0:0] mux_3249_nl;
  wire[0:0] mux_3248_nl;
  wire[0:0] and_422_nl;
  wire[0:0] mux_3247_nl;
  wire[0:0] and_423_nl;
  wire[0:0] mux_3246_nl;
  wire[0:0] or_2910_nl;
  wire[0:0] nor_644_nl;
  wire[0:0] nor_645_nl;
  wire[0:0] modExp_while_if_and_nl;
  wire[0:0] modExp_while_if_and_1_nl;
  wire[0:0] and_261_nl;
  wire[0:0] mux_2545_nl;
  wire[0:0] mux_2544_nl;
  wire[0:0] mux_2543_nl;
  wire[0:0] mux_2542_nl;
  wire[0:0] mux_2541_nl;
  wire[0:0] mux_2540_nl;
  wire[0:0] or_2578_nl;
  wire[0:0] mux_2630_nl;
  wire[0:0] mux_2629_nl;
  wire[0:0] mux_2628_nl;
  wire[0:0] mux_2610_nl;
  wire[0:0] mux_2609_nl;
  wire[0:0] or_2624_nl;
  wire[0:0] mux_2608_nl;
  wire[0:0] mux_2607_nl;
  wire[0:0] or_2622_nl;
  wire[0:0] mux_2532_nl;
  wire[0:0] mux_2617_nl;
  wire[0:0] mux_2616_nl;
  wire[0:0] mux_2615_nl;
  wire[0:0] mux_2614_nl;
  wire[0:0] nor_696_nl;
  wire[0:0] or_2627_nl;
  wire[0:0] mux_2600_nl;
  wire[0:0] mux_2599_nl;
  wire[0:0] mux_2598_nl;
  wire[0:0] mux_2524_nl;
  wire[0:0] mux_2523_nl;
  wire[0:0] mux_2522_nl;
  wire[0:0] mux_2521_nl;
  wire[0:0] mux_2520_nl;
  wire[0:0] mux_2624_nl;
  wire[0:0] mux_2623_nl;
  wire[0:0] mux_2622_nl;
  wire[0:0] mux_2620_nl;
  wire[0:0] mux_2619_nl;
  wire[0:0] mux_2604_nl;
  wire[0:0] mux_2603_nl;
  wire[0:0] mux_2602_nl;
  wire[0:0] mux_2586_nl;
  wire[0:0] or_2620_nl;
  wire[0:0] mux_2508_nl;
  wire[0:0] mux_2613_nl;
  wire[0:0] or_2625_nl;
  wire[0:0] mux_2597_nl;
  wire[0:0] mux_2596_nl;
  wire[0:0] mux_2595_nl;
  wire[0:0] mux_2594_nl;
  wire[0:0] or_2616_nl;
  wire[0:0] mux_2593_nl;
  wire[0:0] nor_704_nl;
  wire[0:0] or_2612_nl;
  wire[0:0] mux_2501_nl;
  wire[0:0] mux_2500_nl;
  wire[0:0] mux_2499_nl;
  wire[0:0] mux_2498_nl;
  wire[0:0] mux_2497_nl;
  wire[0:0] mux_2496_nl;
  wire[0:0] mux_2495_nl;
  wire[0:0] mux_2561_nl;
  wire[0:0] mux_2560_nl;
  wire[0:0] nor_707_nl;
  wire[0:0] or_2591_nl;
  wire[0:0] mux_2559_nl;
  wire[0:0] or_2589_nl;
  wire[0:0] mux_2490_nl;
  wire[0:0] mux_2576_nl;
  wire[0:0] mux_2575_nl;
  wire[0:0] mux_2574_nl;
  wire[0:0] mux_2572_nl;
  wire[0:0] mux_2571_nl;
  wire[0:0] mux_2570_nl;
  wire[0:0] or_2602_nl;
  wire[0:0] mux_2553_nl;
  wire[0:0] mux_2552_nl;
  wire[0:0] nor_709_nl;
  wire[0:0] mux_2551_nl;
  wire[0:0] mux_2550_nl;
  wire[0:0] mux_2478_nl;
  wire[0:0] mux_2477_nl;
  wire[0:0] mux_2585_nl;
  wire[0:0] mux_2584_nl;
  wire[0:0] mux_2583_nl;
  wire[0:0] mux_2582_nl;
  wire[0:0] mux_2581_nl;
  wire[0:0] mux_2580_nl;
  wire[0:0] mux_2579_nl;
  wire[0:0] mux_2578_nl;
  wire[0:0] or_2608_nl;
  wire[0:0] or_2606_nl;
  wire[0:0] mux_2558_nl;
  wire[0:0] mux_2557_nl;
  wire[0:0] mux_2556_nl;
  wire[0:0] mux_2464_nl;
  wire[0:0] mux_2569_nl;
  wire[0:0] mux_2568_nl;
  wire[0:0] mux_2567_nl;
  wire[0:0] mux_2566_nl;
  wire[0:0] or_2598_nl;
  wire[0:0] mux_2565_nl;
  wire[0:0] mux_2564_nl;
  wire[0:0] mux_2549_nl;
  wire[0:0] mux_2548_nl;
  wire[0:0] or_2582_nl;
  wire[0:0] mux_2547_nl;
  wire[0:0] mux_2546_nl;
  wire[0:0] or_2580_nl;
  wire[0:0] mux_3889_nl;
  wire[0:0] mux_3888_nl;
  wire[0:0] mux_3887_nl;
  wire[0:0] mux_3886_nl;
  wire[0:0] nor_1705_nl;
  wire[0:0] mux_3885_nl;
  wire[0:0] or_3549_nl;
  wire[0:0] mux_3884_nl;
  wire[0:0] mux_3883_nl;
  wire[0:0] nor_1706_nl;
  wire[0:0] and_1165_nl;
  wire[0:0] and_1166_nl;
  wire[0:0] mux_3882_nl;
  wire[0:0] mux_3881_nl;
  wire[0:0] or_3619_nl;
  wire[0:0] or_3620_nl;
  wire[0:0] mux_3880_nl;
  wire[0:0] or_3543_nl;
  wire[0:0] mux_3879_nl;
  wire[0:0] mux_3878_nl;
  wire[0:0] mux_3877_nl;
  wire[0:0] or_3541_nl;
  wire[0:0] mux_3876_nl;
  wire[0:0] nor_1708_nl;
  wire[0:0] mux_3875_nl;
  wire[0:0] mux_3874_nl;
  wire[0:0] mux_3873_nl;
  wire[0:0] mux_3872_nl;
  wire[0:0] mux_3871_nl;
  wire[0:0] or_3537_nl;
  wire[0:0] mux_3870_nl;
  wire[0:0] mux_3869_nl;
  wire[0:0] mux_3868_nl;
  wire[0:0] or_3534_nl;
  wire[0:0] mux_3867_nl;
  wire[0:0] nand_417_nl;
  wire[0:0] mux_3865_nl;
  wire[0:0] mux_3864_nl;
  wire[0:0] and_1168_nl;
  wire[0:0] mux_3863_nl;
  wire[0:0] mux_3862_nl;
  wire[0:0] mux_3861_nl;
  wire[0:0] mux_3860_nl;
  wire[0:0] mux_3859_nl;
  wire[0:0] mux_3857_nl;
  wire[0:0] or_3529_nl;
  wire[0:0] mux_3856_nl;
  wire[0:0] mux_3855_nl;
  wire[0:0] mux_3854_nl;
  wire[0:0] mux_3853_nl;
  wire[0:0] mux_3852_nl;
  wire[0:0] mux_3851_nl;
  wire[0:0] mux_3848_nl;
  wire[0:0] mux_3847_nl;
  wire[0:0] mux_3846_nl;
  wire[0:0] mux_3845_nl;
  wire[0:0] mux_3844_nl;
  wire[0:0] or_3522_nl;
  wire[0:0] mux_3840_nl;
  wire[0:0] mux_3839_nl;
  wire[0:0] mux_3838_nl;
  wire[0:0] nand_416_nl;
  wire[0:0] mux_3837_nl;
  wire[0:0] mux_3836_nl;
  wire[0:0] mux_3835_nl;
  wire[0:0] mux_3834_nl;
  wire[0:0] mux_3833_nl;
  wire[0:0] or_3513_nl;
  wire[0:0] mux_3831_nl;
  wire[0:0] or_3609_nl;
  wire[0:0] mux_3943_nl;
  wire[0:0] mux_3942_nl;
  wire[0:0] mux_3941_nl;
  wire[0:0] mux_3940_nl;
  wire[0:0] mux_3939_nl;
  wire[0:0] mux_3938_nl;
  wire[0:0] or_3612_nl;
  wire[0:0] or_3611_nl;
  wire[0:0] mux_3937_nl;
  wire[0:0] mux_3936_nl;
  wire[0:0] or_3608_nl;
  wire[0:0] mux_3934_nl;
  wire[0:0] mux_3933_nl;
  wire[0:0] or_3606_nl;
  wire[0:0] mux_3932_nl;
  wire[0:0] or_3604_nl;
  wire[0:0] nand_423_nl;
  wire[0:0] mux_3931_nl;
  wire[0:0] mux_3930_nl;
  wire[0:0] mux_3929_nl;
  wire[0:0] or_3601_nl;
  wire[0:0] mux_3928_nl;
  wire[0:0] or_3600_nl;
  wire[0:0] mux_3927_nl;
  wire[0:0] mux_3926_nl;
  wire[0:0] mux_3925_nl;
  wire[0:0] mux_3924_nl;
  wire[0:0] mux_3923_nl;
  wire[0:0] or_3599_nl;
  wire[0:0] or_3598_nl;
  wire[0:0] mux_3922_nl;
  wire[0:0] nand_420_nl;
  wire[0:0] or_3597_nl;
  wire[0:0] mux_3921_nl;
  wire[0:0] mux_3920_nl;
  wire[0:0] or_3595_nl;
  wire[0:0] mux_3919_nl;
  wire[0:0] mux_3918_nl;
  wire[0:0] or_3594_nl;
  wire[0:0] or_3593_nl;
  wire[0:0] or_3591_nl;
  wire[0:0] or_3590_nl;
  wire[0:0] mux_3917_nl;
  wire[0:0] or_3589_nl;
  wire[0:0] mux_3916_nl;
  wire[0:0] mux_3915_nl;
  wire[0:0] mux_3914_nl;
  wire[0:0] mux_3913_nl;
  wire[0:0] mux_3912_nl;
  wire[0:0] mux_3911_nl;
  wire[0:0] mux_3910_nl;
  wire[0:0] mux_3906_nl;
  wire[0:0] or_3578_nl;
  wire[0:0] or_3576_nl;
  wire[0:0] mux_3903_nl;
  wire[0:0] or_3575_nl;
  wire[0:0] mux_3902_nl;
  wire[0:0] mux_3901_nl;
  wire[0:0] or_3573_nl;
  wire[0:0] or_3572_nl;
  wire[0:0] mux_3900_nl;
  wire[0:0] mux_3899_nl;
  wire[0:0] or_3571_nl;
  wire[0:0] mux_3898_nl;
  wire[0:0] or_3569_nl;
  wire[0:0] mux_3897_nl;
  wire[0:0] or_3568_nl;
  wire[0:0] mux_3896_nl;
  wire[0:0] or_3565_nl;
  wire[0:0] mux_3895_nl;
  wire[0:0] mux_3892_nl;
  wire[0:0] or_3556_nl;
  wire[0:0] mux_3891_nl;
  wire[0:0] or_3554_nl;
  wire[0:0] mux_3890_nl;
  wire[0:0] or_3553_nl;
  wire[0:0] or_3551_nl;
  wire[0:0] or_3508_nl;
  wire[0:0] mux_2639_nl;
  wire[0:0] or_2642_nl;
  wire[0:0] mux_2638_nl;
  wire[0:0] or_2641_nl;
  wire[0:0] or_2640_nl;
  wire[0:0] or_2638_nl;
  wire[0:0] mux_3946_nl;
  wire[0:0] nor_1700_nl;
  wire[0:0] nor_1701_nl;
  wire[0:0] mux_3945_nl;
  wire[0:0] mux_3944_nl;
  wire[0:0] or_3616_nl;
  wire[0:0] or_3615_nl;
  wire[0:0] or_3613_nl;
  wire[0:0] mux_2668_nl;
  wire[0:0] mux_2667_nl;
  wire[0:0] mux_2666_nl;
  wire[0:0] mux_2665_nl;
  wire[0:0] mux_2664_nl;
  wire[0:0] mux_2663_nl;
  wire[0:0] nor_690_nl;
  wire[0:0] mux_2662_nl;
  wire[0:0] mux_2661_nl;
  wire[0:0] mux_2660_nl;
  wire[0:0] nand_170_nl;
  wire[0:0] COMP_LOOP_or_8_nl;
  wire[0:0] COMP_LOOP_or_9_nl;
  wire[0:0] COMP_LOOP_or_10_nl;
  wire[0:0] COMP_LOOP_or_11_nl;
  wire[0:0] COMP_LOOP_or_12_nl;
  wire[0:0] COMP_LOOP_or_13_nl;
  wire[0:0] COMP_LOOP_or_14_nl;
  wire[0:0] COMP_LOOP_or_15_nl;
  wire[0:0] COMP_LOOP_or_16_nl;
  wire[0:0] COMP_LOOP_or_17_nl;
  wire[0:0] COMP_LOOP_or_18_nl;
  wire[0:0] COMP_LOOP_or_19_nl;
  wire[0:0] COMP_LOOP_or_20_nl;
  wire[0:0] COMP_LOOP_or_21_nl;
  wire[0:0] COMP_LOOP_or_22_nl;
  wire[0:0] COMP_LOOP_or_23_nl;
  wire[0:0] mux_2741_nl;
  wire[0:0] mux_2740_nl;
  wire[0:0] mux_2739_nl;
  wire[0:0] mux_2738_nl;
  wire[0:0] mux_2737_nl;
  wire[0:0] and_276_nl;
  wire[0:0] mux_2735_nl;
  wire[0:0] mux_2734_nl;
  wire[0:0] nor_687_nl;
  wire[0:0] mux_2733_nl;
  wire[0:0] mux_2732_nl;
  wire[0:0] mux_2731_nl;
  wire[0:0] mux_2730_nl;
  wire[0:0] mux_2729_nl;
  wire[0:0] mux_2728_nl;
  wire[0:0] or_2666_nl;
  wire[0:0] mux_2727_nl;
  wire[0:0] and_454_nl;
  wire[0:0] mux_2726_nl;
  wire[0:0] mux_2725_nl;
  wire[0:0] mux_2724_nl;
  wire[0:0] mux_2723_nl;
  wire[0:0] mux_2722_nl;
  wire[0:0] mux_2721_nl;
  wire[0:0] mux_2720_nl;
  wire[0:0] mux_2719_nl;
  wire[0:0] mux_2718_nl;
  wire[0:0] mux_2717_nl;
  wire[0:0] mux_2716_nl;
  wire[0:0] mux_2714_nl;
  wire[0:0] mux_2713_nl;
  wire[0:0] mux_2712_nl;
  wire[0:0] mux_2711_nl;
  wire[0:0] mux_2710_nl;
  wire[0:0] mux_2707_nl;
  wire[0:0] mux_2705_nl;
  wire[0:0] mux_2704_nl;
  wire[0:0] mux_2701_nl;
  wire[0:0] mux_2699_nl;
  wire[0:0] mux_2697_nl;
  wire[0:0] mux_2696_nl;
  wire[0:0] mux_2695_nl;
  wire[0:0] mux_2694_nl;
  wire[0:0] mux_2692_nl;
  wire[0:0] mux_2689_nl;
  wire[0:0] mux_2688_nl;
  wire[0:0] mux_2687_nl;
  wire[0:0] mux_2686_nl;
  wire[0:0] mux_2685_nl;
  wire[0:0] mux_2684_nl;
  wire[0:0] mux_2683_nl;
  wire[0:0] mux_2680_nl;
  wire[0:0] mux_2679_nl;
  wire[0:0] mux_2678_nl;
  wire[0:0] or_2658_nl;
  wire[0:0] mux_2674_nl;
  wire[0:0] mux_2673_nl;
  wire[0:0] mux_2671_nl;
  wire[0:0] mux_2770_nl;
  wire[0:0] nor_678_nl;
  wire[0:0] mux_2769_nl;
  wire[0:0] nand_166_nl;
  wire[0:0] nor_679_nl;
  wire[0:0] mux_2768_nl;
  wire[0:0] or_2717_nl;
  wire[0:0] mux_2767_nl;
  wire[0:0] or_2716_nl;
  wire[0:0] or_2714_nl;
  wire[0:0] nand_58_nl;
  wire[0:0] mux_2766_nl;
  wire[0:0] mux_2765_nl;
  wire[0:0] mux_2764_nl;
  wire[0:0] nor_680_nl;
  wire[0:0] mux_2763_nl;
  wire[0:0] mux_2762_nl;
  wire[0:0] or_2708_nl;
  wire[0:0] nor_681_nl;
  wire[0:0] mux_2761_nl;
  wire[0:0] or_2702_nl;
  wire[0:0] and_451_nl;
  wire[0:0] mux_2759_nl;
  wire[0:0] nor_682_nl;
  wire[0:0] mux_2758_nl;
  wire[0:0] nor_683_nl;
  wire[0:0] nor_684_nl;
  wire[0:0] mux_2743_nl;
  wire[0:0] nor_685_nl;
  wire[0:0] nor_686_nl;
  wire[0:0] and_312_nl;
  wire[0:0] COMP_LOOP_or_29_nl;
  wire[0:0] COMP_LOOP_or_30_nl;
  wire[0:0] COMP_LOOP_and_277_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_932_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_934_nl;
  wire[0:0] COMP_LOOP_and_1_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_936_nl;
  wire[0:0] COMP_LOOP_and_2_nl;
  wire[0:0] COMP_LOOP_and_3_nl;
  wire[0:0] COMP_LOOP_and_4_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_930_nl;
  wire[0:0] COMP_LOOP_and_5_nl;
  wire[0:0] COMP_LOOP_and_6_nl;
  wire[0:0] COMP_LOOP_and_7_nl;
  wire[0:0] COMP_LOOP_and_8_nl;
  wire[0:0] COMP_LOOP_and_9_nl;
  wire[0:0] COMP_LOOP_and_10_nl;
  wire[0:0] COMP_LOOP_and_11_nl;
  wire[0:0] mux_129_nl;
  wire[0:0] mux_128_nl;
  wire[0:0] nand_3_nl;
  wire[0:0] mux_127_nl;
  wire[0:0] mux_126_nl;
  wire[0:0] nand_2_nl;
  wire[0:0] or_92_nl;
  wire[0:0] mux_124_nl;
  wire[0:0] mux_123_nl;
  wire[0:0] or_91_nl;
  wire[0:0] or_89_nl;
  wire[0:0] or_88_nl;
  wire[0:0] mux_122_nl;
  wire[0:0] mux_121_nl;
  wire[0:0] mux_120_nl;
  wire[0:0] or_87_nl;
  wire[0:0] or_85_nl;
  wire[0:0] or_81_nl;
  wire[0:0] mux_118_nl;
  wire[0:0] mux_117_nl;
  wire[0:0] or_79_nl;
  wire[0:0] mux_116_nl;
  wire[0:0] nand_373_nl;
  wire[0:0] mux_2981_nl;
  wire[0:0] mux_2980_nl;
  wire[0:0] mux_2979_nl;
  wire[0:0] mux_2978_nl;
  wire[0:0] mux_2977_nl;
  wire[0:0] mux_2976_nl;
  wire[0:0] mux_2975_nl;
  wire[0:0] mux_2974_nl;
  wire[0:0] mux_2973_nl;
  wire[0:0] mux_2972_nl;
  wire[0:0] mux_2971_nl;
  wire[0:0] mux_2970_nl;
  wire[0:0] mux_2969_nl;
  wire[0:0] mux_2968_nl;
  wire[0:0] mux_2967_nl;
  wire[0:0] mux_2966_nl;
  wire[0:0] mux_2965_nl;
  wire[0:0] mux_2964_nl;
  wire[0:0] mux_2963_nl;
  wire[0:0] mux_2962_nl;
  wire[0:0] mux_2961_nl;
  wire[0:0] mux_2960_nl;
  wire[0:0] or_2810_nl;
  wire[0:0] mux_2959_nl;
  wire[0:0] nand_72_nl;
  wire[0:0] mux_2958_nl;
  wire[0:0] mux_2957_nl;
  wire[0:0] mux_2956_nl;
  wire[0:0] mux_2955_nl;
  wire[0:0] mux_2954_nl;
  wire[0:0] mux_2953_nl;
  wire[0:0] mux_2952_nl;
  wire[0:0] mux_2951_nl;
  wire[0:0] mux_2950_nl;
  wire[0:0] mux_2949_nl;
  wire[0:0] mux_2948_nl;
  wire[0:0] or_2809_nl;
  wire[0:0] mux_2947_nl;
  wire[0:0] mux_2946_nl;
  wire[0:0] mux_2945_nl;
  wire[0:0] mux_2944_nl;
  wire[0:0] mux_2943_nl;
  wire[0:0] mux_2942_nl;
  wire[0:0] mux_2941_nl;
  wire[0:0] mux_2940_nl;
  wire[0:0] mux_2939_nl;
  wire[0:0] mux_2938_nl;
  wire[0:0] mux_2937_nl;
  wire[0:0] mux_2936_nl;
  wire[0:0] mux_2935_nl;
  wire[0:0] mux_2934_nl;
  wire[0:0] mux_2933_nl;
  wire[0:0] mux_2932_nl;
  wire[0:0] mux_2931_nl;
  wire[0:0] mux_2930_nl;
  wire[0:0] mux_2929_nl;
  wire[0:0] mux_2928_nl;
  wire[0:0] or_2807_nl;
  wire[0:0] mux_2927_nl;
  wire[0:0] mux_2925_nl;
  wire[0:0] mux_2924_nl;
  wire[0:0] mux_2923_nl;
  wire[0:0] mux_2922_nl;
  wire[0:0] mux_2921_nl;
  wire[0:0] mux_2919_nl;
  wire[0:0] mux_2918_nl;
  wire[0:0] mux_2917_nl;
  wire[0:0] mux_2915_nl;
  wire[0:0] mux_2914_nl;
  wire[0:0] mux_2913_nl;
  wire[0:0] mux_2911_nl;
  wire[0:0] mux_2908_nl;
  wire[0:0] mux_2907_nl;
  wire[0:0] mux_2905_nl;
  wire[0:0] mux_2904_nl;
  wire[0:0] mux_2903_nl;
  wire[0:0] mux_2902_nl;
  wire[0:0] mux_2900_nl;
  wire[0:0] mux_2899_nl;
  wire[0:0] mux_2898_nl;
  wire[0:0] mux_2897_nl;
  wire[0:0] mux_2896_nl;
  wire[0:0] mux_2894_nl;
  wire[0:0] mux_2893_nl;
  wire[0:0] mux_2892_nl;
  wire[0:0] mux_2891_nl;
  wire[0:0] mux_2889_nl;
  wire[0:0] mux_2887_nl;
  wire[0:0] mux_2885_nl;
  wire[0:0] mux_2884_nl;
  wire[0:0] mux_2883_nl;
  wire[0:0] mux_2882_nl;
  wire[0:0] mux_2881_nl;
  wire[0:0] mux_2877_nl;
  wire[0:0] mux_2874_nl;
  wire[0:0] mux_2873_nl;
  wire[0:0] mux_2872_nl;
  wire[0:0] mux_2871_nl;
  wire[0:0] mux_2870_nl;
  wire[0:0] mux_2869_nl;
  wire[0:0] mux_2868_nl;
  wire[0:0] mux_2865_nl;
  wire[0:0] mux_2864_nl;
  wire[0:0] mux_2861_nl;
  wire[0:0] mux_2860_nl;
  wire[0:0] mux_2859_nl;
  wire[0:0] or_2797_nl;
  wire[0:0] mux_2857_nl;
  wire[0:0] nand_66_nl;
  wire[0:0] mux_2855_nl;
  wire[0:0] mux_2854_nl;
  wire[0:0] mux_2853_nl;
  wire[0:0] mux_2852_nl;
  wire[0:0] mux_2847_nl;
  wire[0:0] mux_2845_nl;
  wire[0:0] mux_2842_nl;
  wire[0:0] COMP_LOOP_mux1h_428_nl;
  wire[0:0] COMP_LOOP_nor_11_nl;
  wire[0:0] COMP_LOOP_and_274_nl;
  wire[0:0] mux_3070_nl;
  wire[0:0] mux_3069_nl;
  wire[0:0] mux_3068_nl;
  wire[0:0] mux_3067_nl;
  wire[0:0] mux_3066_nl;
  wire[0:0] mux_3065_nl;
  wire[0:0] or_2881_nl;
  wire[0:0] mux_3064_nl;
  wire[0:0] mux_3063_nl;
  wire[0:0] mux_3062_nl;
  wire[0:0] mux_3061_nl;
  wire[0:0] mux_3060_nl;
  wire[0:0] mux_3059_nl;
  wire[0:0] or_449_nl;
  wire[0:0] or_2876_nl;
  wire[0:0] mux_3058_nl;
  wire[0:0] mux_3057_nl;
  wire[0:0] mux_3056_nl;
  wire[0:0] nor_407_nl;
  wire[0:0] mux_3055_nl;
  wire[0:0] mux_3054_nl;
  wire[0:0] mux_3053_nl;
  wire[0:0] mux_3052_nl;
  wire[0:0] mux_3051_nl;
  wire[0:0] or_439_nl;
  wire[0:0] mux_3050_nl;
  wire[0:0] mux_3048_nl;
  wire[0:0] mux_3047_nl;
  wire[0:0] or_2870_nl;
  wire[0:0] mux_3046_nl;
  wire[0:0] mux_3045_nl;
  wire[0:0] mux_3044_nl;
  wire[0:0] mux_3043_nl;
  wire[0:0] mux_3042_nl;
  wire[0:0] mux_3041_nl;
  wire[0:0] mux_3040_nl;
  wire[0:0] mux_3039_nl;
  wire[0:0] mux_3038_nl;
  wire[0:0] mux_3036_nl;
  wire[0:0] mux_3035_nl;
  wire[0:0] mux_3034_nl;
  wire[0:0] mux_3033_nl;
  wire[0:0] mux_3030_nl;
  wire[0:0] or_2866_nl;
  wire[0:0] or_2865_nl;
  wire[0:0] mux_3029_nl;
  wire[0:0] mux_3028_nl;
  wire[0:0] mux_3027_nl;
  wire[0:0] mux_3026_nl;
  wire[0:0] mux_3025_nl;
  wire[0:0] mux_3023_nl;
  wire[0:0] or_2859_nl;
  wire[0:0] mux_3021_nl;
  wire[0:0] mux_3020_nl;
  wire[0:0] mux_3019_nl;
  wire[0:0] mux_3018_nl;
  wire[0:0] mux_3017_nl;
  wire[0:0] mux_3016_nl;
  wire[0:0] mux_3015_nl;
  wire[0:0] mux_3013_nl;
  wire[0:0] or_2851_nl;
  wire[0:0] mux_3012_nl;
  wire[0:0] mux_3011_nl;
  wire[0:0] mux_3010_nl;
  wire[0:0] mux_3009_nl;
  wire[0:0] mux_3005_nl;
  wire[0:0] or_2846_nl;
  wire[0:0] mux_2989_nl;
  wire[0:0] or_3440_nl;
  wire[0:0] mux_2988_nl;
  wire[0:0] or_2821_nl;
  wire[0:0] mux_2987_nl;
  wire[0:0] nand_74_nl;
  wire[0:0] mux_2986_nl;
  wire[0:0] nor_671_nl;
  wire[0:0] nor_672_nl;
  wire[0:0] or_2818_nl;
  wire[0:0] mux_2985_nl;
  wire[0:0] or_3441_nl;
  wire[0:0] or_3442_nl;
  wire[0:0] mux_2984_nl;
  wire[0:0] nand_73_nl;
  wire[0:0] mux_2983_nl;
  wire[0:0] and_447_nl;
  wire[0:0] nor_675_nl;
  wire[0:0] or_2811_nl;
  wire[0:0] mux_3077_nl;
  wire[0:0] mux_3076_nl;
  wire[0:0] nor_646_nl;
  wire[0:0] mux_3075_nl;
  wire[0:0] nor_647_nl;
  wire[0:0] and_439_nl;
  wire[0:0] mux_3074_nl;
  wire[0:0] nor_648_nl;
  wire[0:0] nor_649_nl;
  wire[0:0] mux_3073_nl;
  wire[0:0] and_440_nl;
  wire[0:0] mux_3072_nl;
  wire[0:0] nor_650_nl;
  wire[0:0] mux_3071_nl;
  wire[0:0] nor_651_nl;
  wire[0:0] nor_652_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_17_nl;
  wire[0:0] or_2962_nl;
  wire[0:0] or_2961_nl;
  wire[63:0] COMP_LOOP_1_acc_8_nl;
  wire[64:0] nl_COMP_LOOP_1_acc_8_nl;
  wire[0:0] mux_3288_nl;
  wire[0:0] mux_3287_nl;
  wire[0:0] mux_3286_nl;
  wire[0:0] mux_3285_nl;
  wire[0:0] nor_631_nl;
  wire[0:0] nor_632_nl;
  wire[0:0] mux_3284_nl;
  wire[0:0] and_417_nl;
  wire[0:0] nor_633_nl;
  wire[0:0] mux_3280_nl;
  wire[0:0] or_2959_nl;
  wire[0:0] mux_3279_nl;
  wire[0:0] or_2958_nl;
  wire[0:0] or_2957_nl;
  wire[0:0] mux_3278_nl;
  wire[0:0] or_2954_nl;
  wire[0:0] mux_3277_nl;
  wire[0:0] mux_3276_nl;
  wire[0:0] and_418_nl;
  wire[0:0] nor_634_nl;
  wire[0:0] nor_635_nl;
  wire[0:0] mux_3275_nl;
  wire[0:0] nand_92_nl;
  wire[0:0] or_2945_nl;
  wire[0:0] mux_3273_nl;
  wire[0:0] or_2943_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_and_10_nl;
  wire[9:0] COMP_LOOP_1_acc_nl;
  wire[10:0] nl_COMP_LOOP_1_acc_nl;
  wire[0:0] mux_3334_nl;
  wire[0:0] mux_3333_nl;
  wire[0:0] mux_3332_nl;
  wire[0:0] mux_3331_nl;
  wire[0:0] mux_3330_nl;
  wire[0:0] mux_2642_nl;
  wire[0:0] or_2647_nl;
  wire[0:0] mux_3327_nl;
  wire[0:0] mux_3326_nl;
  wire[0:0] or_3032_nl;
  wire[0:0] and_410_nl;
  wire[0:0] mux_3325_nl;
  wire[0:0] and_411_nl;
  wire[0:0] mux_3340_nl;
  wire[0:0] mux_3339_nl;
  wire[0:0] mux_3338_nl;
  wire[0:0] mux_3337_nl;
  wire[0:0] or_3037_nl;
  wire[0:0] mux_3336_nl;
  wire[0:0] and_408_nl;
  wire[0:0] or_3036_nl;
  wire[0:0] mux_3350_nl;
  wire[0:0] mux_3349_nl;
  wire[0:0] mux_3348_nl;
  wire[0:0] mux_3347_nl;
  wire[0:0] mux_3346_nl;
  wire[0:0] mux_3345_nl;
  wire[0:0] mux_3344_nl;
  wire[0:0] mux_3355_nl;
  wire[0:0] mux_3354_nl;
  wire[0:0] mux_3353_nl;
  wire[0:0] mux_3351_nl;
  wire[0:0] nor_623_nl;
  wire[0:0] mux_3359_nl;
  wire[0:0] mux_3358_nl;
  wire[0:0] mux_3357_nl;
  wire[0:0] mux_3356_nl;
  wire[0:0] and_401_nl;
  wire[0:0] and_402_nl;
  wire[0:0] mux_3364_nl;
  wire[0:0] mux_3363_nl;
  wire[0:0] mux_3362_nl;
  wire[0:0] or_3045_nl;
  wire[0:0] mux_3360_nl;
  wire[0:0] mux_3367_nl;
  wire[0:0] mux_3366_nl;
  wire[0:0] nor_621_nl;
  wire[0:0] mux_3365_nl;
  wire[0:0] or_3048_nl;
  wire[0:0] and_334_nl;
  wire[0:0] mux_3372_nl;
  wire[0:0] mux_3371_nl;
  wire[0:0] mux_3370_nl;
  wire[0:0] nor_619_nl;
  wire[0:0] nor_620_nl;
  wire[0:0] mux_3369_nl;
  wire[0:0] and_337_nl;
  wire[0:0] mux_3368_nl;
  wire[0:0] and_30_nl;
  wire[0:0] mux_3375_nl;
  wire[0:0] mux_3374_nl;
  wire[0:0] nor_1596_nl;
  wire[0:0] mux_3373_nl;
  wire[0:0] nor_1597_nl;
  wire[0:0] and_749_nl;
  wire[0:0] and_750_nl;
  wire[0:0] mux_3381_nl;
  wire[0:0] mux_3380_nl;
  wire[0:0] mux_3379_nl;
  wire[0:0] or_3060_nl;
  wire[0:0] mux_3377_nl;
  wire[0:0] mux_3376_nl;
  wire[0:0] or_3058_nl;
  wire[0:0] mux_3386_nl;
  wire[0:0] mux_3385_nl;
  wire[0:0] mux_3384_nl;
  wire[0:0] or_3065_nl;
  wire[0:0] mux_3383_nl;
  wire[0:0] and_394_nl;
  wire[0:0] mux_3391_nl;
  wire[0:0] mux_3390_nl;
  wire[0:0] mux_3389_nl;
  wire[0:0] mux_3388_nl;
  wire[0:0] nor_615_nl;
  wire[0:0] and_391_nl;
  wire[0:0] mux_3396_nl;
  wire[0:0] mux_3395_nl;
  wire[0:0] mux_3394_nl;
  wire[0:0] nor_613_nl;
  wire[0:0] nor_614_nl;
  wire[0:0] mux_3393_nl;
  wire[0:0] and_388_nl;
  wire[0:0] mux_3400_nl;
  wire[0:0] mux_3399_nl;
  wire[0:0] nor_611_nl;
  wire[0:0] mux_3398_nl;
  wire[0:0] nor_612_nl;
  wire[0:0] and_384_nl;
  wire[0:0] and_386_nl;
  wire[0:0] nor_1680_nl;
  wire[0:0] mux_3403_nl;
  wire[0:0] or_3078_nl;
  wire[0:0] and_1162_nl;
  wire[0:0] mux_3402_nl;
  wire[0:0] or_3076_nl;
  wire[0:0] mux_3408_nl;
  wire[0:0] mux_3407_nl;
  wire[0:0] mux_3406_nl;
  wire[0:0] nor_610_nl;
  wire[0:0] mux_3405_nl;
  wire[0:0] and_341_nl;
  wire[0:0] COMP_LOOP_mux1h_464_nl;
  wire[0:0] mux_3521_nl;
  wire[0:0] mux_3520_nl;
  wire[0:0] mux_3519_nl;
  wire[0:0] mux_3518_nl;
  wire[0:0] or_3501_nl;
  wire[0:0] mux_3517_nl;
  wire[0:0] or_3502_nl;
  wire[0:0] or_3503_nl;
  wire[0:0] or_3504_nl;
  wire[0:0] mux_3516_nl;
  wire[0:0] mux_3515_nl;
  wire[0:0] or_3133_nl;
  wire[0:0] mux_3514_nl;
  wire[0:0] or_3131_nl;
  wire[0:0] or_3130_nl;
  wire[0:0] mux_3513_nl;
  wire[0:0] mux_3512_nl;
  wire[0:0] or_3505_nl;
  wire[0:0] nand_412_nl;
  wire[0:0] mux_3511_nl;
  wire[0:0] nor_600_nl;
  wire[0:0] nor_601_nl;
  wire[0:0] mux_3510_nl;
  wire[0:0] or_3506_nl;
  wire[0:0] mux_3509_nl;
  wire[0:0] or_3124_nl;
  wire[0:0] or_3123_nl;
  wire[0:0] nand_413_nl;
  wire[0:0] mux_3508_nl;
  wire[0:0] or_3120_nl;
  wire[0:0] COMP_LOOP_mux1h_474_nl;
  wire[0:0] COMP_LOOP_nor_12_nl;
  wire[0:0] mux_3616_nl;
  wire[0:0] mux_3615_nl;
  wire[0:0] mux_3614_nl;
  wire[0:0] mux_3613_nl;
  wire[0:0] mux_3612_nl;
  wire[0:0] mux_3611_nl;
  wire[0:0] mux_3610_nl;
  wire[0:0] mux_3609_nl;
  wire[0:0] mux_3608_nl;
  wire[0:0] mux_3607_nl;
  wire[0:0] mux_3606_nl;
  wire[0:0] mux_3605_nl;
  wire[0:0] mux_3604_nl;
  wire[0:0] mux_3603_nl;
  wire[0:0] mux_3602_nl;
  wire[0:0] mux_3601_nl;
  wire[0:0] mux_3600_nl;
  wire[0:0] mux_3599_nl;
  wire[0:0] or_3192_nl;
  wire[0:0] mux_3598_nl;
  wire[0:0] mux_3597_nl;
  wire[0:0] mux_3596_nl;
  wire[0:0] mux_3595_nl;
  wire[0:0] mux_493_nl;
  wire[0:0] mux_3592_nl;
  wire[0:0] mux_3591_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] mux_3588_nl;
  wire[0:0] mux_3586_nl;
  wire[0:0] mux_3585_nl;
  wire[0:0] mux_3584_nl;
  wire[0:0] mux_3583_nl;
  wire[0:0] and_364_nl;
  wire[0:0] mux_3582_nl;
  wire[0:0] mux_3581_nl;
  wire[0:0] mux_3580_nl;
  wire[0:0] mux_3579_nl;
  wire[0:0] mux_3578_nl;
  wire[0:0] mux_3572_nl;
  wire[0:0] mux_3571_nl;
  wire[0:0] mux_3570_nl;
  wire[0:0] mux_3569_nl;
  wire[0:0] mux_481_nl;
  wire[0:0] mux_3566_nl;
  wire[0:0] mux_3565_nl;
  wire[0:0] mux_3563_nl;
  wire[0:0] mux_3562_nl;
  wire[0:0] mux_3560_nl;
  wire[0:0] mux_3559_nl;
  wire[0:0] mux_3558_nl;
  wire[0:0] mux_3557_nl;
  wire[0:0] and_365_nl;
  wire[0:0] mux_3556_nl;
  wire[0:0] mux_3554_nl;
  wire[0:0] mux_3553_nl;
  wire[0:0] mux_3552_nl;
  wire[0:0] mux_3548_nl;
  wire[0:0] mux_3546_nl;
  wire[0:0] or_3177_nl;
  wire[0:0] mux_3545_nl;
  wire[0:0] mux_3630_nl;
  wire[0:0] mux_3629_nl;
  wire[0:0] mux_3628_nl;
  wire[0:0] nor_565_nl;
  wire[0:0] mux_3627_nl;
  wire[0:0] nor_566_nl;
  wire[0:0] mux_3626_nl;
  wire[0:0] or_3213_nl;
  wire[0:0] or_3211_nl;
  wire[0:0] mux_3625_nl;
  wire[0:0] nor_567_nl;
  wire[0:0] mux_3624_nl;
  wire[0:0] nor_568_nl;
  wire[0:0] nor_569_nl;
  wire[0:0] mux_3623_nl;
  wire[0:0] mux_3622_nl;
  wire[0:0] nor_570_nl;
  wire[0:0] mux_3621_nl;
  wire[0:0] or_3203_nl;
  wire[0:0] nor_571_nl;
  wire[0:0] mux_3620_nl;
  wire[0:0] mux_3619_nl;
  wire[0:0] nor_572_nl;
  wire[0:0] and_362_nl;
  wire[0:0] mux_3617_nl;
  wire[0:0] nor_573_nl;
  wire[0:0] nor_574_nl;
  wire[0:0] nor_575_nl;
  wire[0:0] mux_3542_nl;
  wire[0:0] nand_411_nl;
  wire[0:0] mux_3541_nl;
  wire[0:0] nor_578_nl;
  wire[0:0] mux_3540_nl;
  wire[0:0] or_3171_nl;
  wire[0:0] mux_3539_nl;
  wire[0:0] nor_579_nl;
  wire[0:0] nor_580_nl;
  wire[0:0] or_3499_nl;
  wire[0:0] mux_3538_nl;
  wire[0:0] or_3166_nl;
  wire[0:0] mux_3537_nl;
  wire[0:0] nand_139_nl;
  wire[0:0] nand_104_nl;
  wire[0:0] mux_3536_nl;
  wire[0:0] nor_582_nl;
  wire[0:0] nor_583_nl;
  wire[0:0] mux_3636_nl;
  wire[0:0] nor_562_nl;
  wire[0:0] mux_3635_nl;
  wire[0:0] or_3228_nl;
  wire[0:0] mux_3634_nl;
  wire[0:0] or_3226_nl;
  wire[0:0] or_3224_nl;
  wire[0:0] and_361_nl;
  wire[0:0] mux_3633_nl;
  wire[0:0] nor_563_nl;
  wire[0:0] nor_564_nl;
  wire[0:0] mux_3631_nl;
  wire[0:0] or_3217_nl;
  wire[0:0] or_3215_nl;
  wire[0:0] COMP_LOOP_mux1h_477_nl;
  wire[0:0] COMP_LOOP_nor_14_nl;
  wire[0:0] mux_3642_nl;
  wire[0:0] mux_3641_nl;
  wire[0:0] mux_3640_nl;
  wire[0:0] mux_3639_nl;
  wire[0:0] mux_3638_nl;
  wire[0:0] mux_3637_nl;
  wire[0:0] mux_3649_nl;
  wire[0:0] or_3497_nl;
  wire[0:0] mux_3648_nl;
  wire[0:0] or_3241_nl;
  wire[0:0] mux_3647_nl;
  wire[0:0] or_3240_nl;
  wire[0:0] or_3239_nl;
  wire[0:0] mux_3646_nl;
  wire[0:0] or_3236_nl;
  wire[0:0] mux_3645_nl;
  wire[0:0] or_3235_nl;
  wire[0:0] or_3234_nl;
  wire[0:0] mux_3644_nl;
  wire[0:0] or_3498_nl;
  wire[0:0] nand_410_nl;
  wire[0:0] mux_3643_nl;
  wire[0:0] nor_560_nl;
  wire[0:0] nor_561_nl;
  wire[0:0] mux_3656_nl;
  wire[0:0] mux_3655_nl;
  wire[0:0] nor_555_nl;
  wire[0:0] nor_556_nl;
  wire[0:0] mux_3654_nl;
  wire[0:0] mux_3653_nl;
  wire[0:0] or_3253_nl;
  wire[0:0] or_3251_nl;
  wire[0:0] nor_557_nl;
  wire[0:0] mux_3652_nl;
  wire[0:0] or_3249_nl;
  wire[0:0] mux_3651_nl;
  wire[0:0] nand_383_nl;
  wire[0:0] or_3246_nl;
  wire[0:0] mux_3650_nl;
  wire[0:0] or_3244_nl;
  wire[0:0] COMP_LOOP_mux1h_479_nl;
  wire[0:0] COMP_LOOP_nor_17_nl;
  wire[0:0] mux_3663_nl;
  wire[0:0] nand_389_nl;
  wire[0:0] mux_3662_nl;
  wire[0:0] nor_552_nl;
  wire[0:0] mux_3661_nl;
  wire[0:0] mux_3660_nl;
  wire[0:0] or_3266_nl;
  wire[0:0] nand_130_nl;
  wire[0:0] nor_553_nl;
  wire[0:0] or_3443_nl;
  wire[0:0] mux_3659_nl;
  wire[0:0] or_3353_nl;
  wire[0:0] mux_3658_nl;
  wire[0:0] or_3261_nl;
  wire[0:0] or_3260_nl;
  wire[0:0] mux_3657_nl;
  wire[0:0] mux_3670_nl;
  wire[0:0] mux_3669_nl;
  wire[0:0] nor_547_nl;
  wire[0:0] and_357_nl;
  wire[0:0] mux_3668_nl;
  wire[0:0] nor_548_nl;
  wire[0:0] mux_3667_nl;
  wire[0:0] or_3282_nl;
  wire[0:0] nand_382_nl;
  wire[0:0] and_358_nl;
  wire[0:0] mux_3666_nl;
  wire[0:0] nor_549_nl;
  wire[0:0] nor_550_nl;
  wire[0:0] nor_551_nl;
  wire[0:0] mux_3665_nl;
  wire[0:0] or_3274_nl;
  wire[0:0] mux_3664_nl;
  wire[0:0] or_3273_nl;
  wire[0:0] or_3271_nl;
  wire[0:0] or_3269_nl;
  wire[0:0] COMP_LOOP_mux1h_480_nl;
  wire[0:0] mux_3766_nl;
  wire[0:0] mux_3765_nl;
  wire[0:0] mux_3764_nl;
  wire[0:0] mux_3763_nl;
  wire[0:0] mux_3762_nl;
  wire[0:0] mux_3761_nl;
  wire[0:0] mux_3760_nl;
  wire[0:0] mux_3759_nl;
  wire[0:0] mux_3758_nl;
  wire[0:0] mux_3757_nl;
  wire[0:0] mux_3756_nl;
  wire[0:0] mux_3755_nl;
  wire[0:0] mux_3754_nl;
  wire[0:0] mux_3752_nl;
  wire[0:0] mux_3751_nl;
  wire[0:0] mux_3750_nl;
  wire[0:0] or_3302_nl;
  wire[0:0] mux_3749_nl;
  wire[0:0] mux_3748_nl;
  wire[0:0] mux_3747_nl;
  wire[0:0] mux_3746_nl;
  wire[0:0] mux_3745_nl;
  wire[0:0] mux_3744_nl;
  wire[0:0] mux_3743_nl;
  wire[0:0] nor_546_nl;
  wire[0:0] mux_3742_nl;
  wire[0:0] mux_3741_nl;
  wire[0:0] mux_3740_nl;
  wire[0:0] mux_3735_nl;
  wire[0:0] mux_3734_nl;
  wire[0:0] mux_3733_nl;
  wire[0:0] or_3298_nl;
  wire[0:0] mux_3732_nl;
  wire[0:0] mux_3731_nl;
  wire[0:0] and_349_nl;
  wire[0:0] mux_3730_nl;
  wire[0:0] mux_3729_nl;
  wire[0:0] mux_3728_nl;
  wire[0:0] mux_3727_nl;
  wire[0:0] mux_3726_nl;
  wire[0:0] mux_3725_nl;
  wire[0:0] mux_3723_nl;
  wire[0:0] mux_3722_nl;
  wire[0:0] mux_3721_nl;
  wire[0:0] mux_3719_nl;
  wire[0:0] mux_3717_nl;
  wire[0:0] mux_3716_nl;
  wire[0:0] mux_3715_nl;
  wire[0:0] mux_3714_nl;
  wire[0:0] mux_3713_nl;
  wire[0:0] mux_3711_nl;
  wire[0:0] mux_3710_nl;
  wire[0:0] mux_3709_nl;
  wire[0:0] mux_3708_nl;
  wire[0:0] mux_3707_nl;
  wire[0:0] mux_3706_nl;
  wire[0:0] or_3295_nl;
  wire[0:0] mux_3703_nl;
  wire[0:0] mux_3702_nl;
  wire[0:0] mux_3699_nl;
  wire[0:0] mux_3695_nl;
  wire[0:0] mux_3694_nl;
  wire[0:0] mux_3693_nl;
  wire[0:0] mux_3692_nl;
  wire[0:0] mux_3690_nl;
  wire[0:0] mux_3689_nl;
  wire[0:0] mux_3688_nl;
  wire[0:0] mux_3687_nl;
  wire[0:0] nand_380_nl;
  wire[0:0] mux_3686_nl;
  wire[0:0] mux_3685_nl;
  wire[0:0] mux_3684_nl;
  wire[0:0] mux_3683_nl;
  wire[0:0] mux_3682_nl;
  wire[0:0] mux_3680_nl;
  wire[0:0] mux_3678_nl;
  wire[0:0] nor_527_nl;
  wire[0:0] mux_3677_nl;
  wire[0:0] mux_3676_nl;
  wire[0:0] mux_3675_nl;
  wire[0:0] COMP_LOOP_or_28_nl;
  wire[0:0] or_18_nl;
  wire[0:0] or_84_nl;
  wire[0:0] or_83_nl;
  wire[0:0] or_108_nl;
  wire[0:0] mux_1078_nl;
  wire[0:0] mux_1077_nl;
  wire[0:0] or_3394_nl;
  wire[0:0] or_510_nl;
  wire[0:0] mux_1081_nl;
  wire[0:0] or_508_nl;
  wire[0:0] or_580_nl;
  wire[0:0] or_579_nl;
  wire[0:0] or_691_nl;
  wire[0:0] or_690_nl;
  wire[0:0] or_802_nl;
  wire[0:0] or_801_nl;
  wire[0:0] or_912_nl;
  wire[0:0] or_911_nl;
  wire[0:0] or_1022_nl;
  wire[0:0] or_1021_nl;
  wire[0:0] or_1133_nl;
  wire[0:0] or_1132_nl;
  wire[0:0] or_1244_nl;
  wire[0:0] or_1243_nl;
  wire[0:0] or_1354_nl;
  wire[0:0] or_1353_nl;
  wire[0:0] or_1464_nl;
  wire[0:0] or_1463_nl;
  wire[0:0] or_1575_nl;
  wire[0:0] or_1574_nl;
  wire[0:0] or_1686_nl;
  wire[0:0] or_1685_nl;
  wire[0:0] or_1796_nl;
  wire[0:0] or_1795_nl;
  wire[0:0] or_1906_nl;
  wire[0:0] or_1905_nl;
  wire[0:0] or_2017_nl;
  wire[0:0] or_2016_nl;
  wire[0:0] or_2128_nl;
  wire[0:0] or_2127_nl;
  wire[0:0] nand_225_nl;
  wire[0:0] or_2237_nl;
  wire[0:0] mux_2175_nl;
  wire[0:0] mux_2234_nl;
  wire[0:0] mux_2239_nl;
  wire[0:0] nand_188_nl;
  wire[0:0] or_2447_nl;
  wire[0:0] mux_2352_nl;
  wire[0:0] or_2448_nl;
  wire[0:0] or_2451_nl;
  wire[0:0] or_2457_nl;
  wire[0:0] or_2459_nl;
  wire[0:0] mux_2375_nl;
  wire[0:0] or_2462_nl;
  wire[0:0] mux_2385_nl;
  wire[0:0] mux_2388_nl;
  wire[0:0] mux_2387_nl;
  wire[0:0] or_2475_nl;
  wire[0:0] or_2474_nl;
  wire[0:0] mux_2431_nl;
  wire[0:0] nor_741_nl;
  wire[0:0] mux_2430_nl;
  wire[0:0] or_2488_nl;
  wire[0:0] or_2487_nl;
  wire[0:0] mux_2429_nl;
  wire[0:0] mux_2428_nl;
  wire[0:0] nor_742_nl;
  wire[0:0] mux_2427_nl;
  wire[0:0] or_2484_nl;
  wire[0:0] nand_182_nl;
  wire[0:0] nor_743_nl;
  wire[0:0] mux_2426_nl;
  wire[0:0] nor_744_nl;
  wire[0:0] mux_2425_nl;
  wire[0:0] or_2479_nl;
  wire[0:0] or_2478_nl;
  wire[0:0] nor_745_nl;
  wire[0:0] mux_2423_nl;
  wire[0:0] mux_2422_nl;
  wire[0:0] mux_2421_nl;
  wire[0:0] nor_746_nl;
  wire[0:0] nor_747_nl;
  wire[0:0] mux_2420_nl;
  wire[0:0] nor_748_nl;
  wire[0:0] nor_749_nl;
  wire[0:0] mux_2419_nl;
  wire[0:0] nand_388_nl;
  wire[0:0] or_2465_nl;
  wire[0:0] nor_750_nl;
  wire[0:0] mux_2445_nl;
  wire[0:0] mux_2444_nl;
  wire[0:0] mux_2443_nl;
  wire[0:0] nor_729_nl;
  wire[0:0] mux_2442_nl;
  wire[0:0] or_2512_nl;
  wire[0:0] nor_730_nl;
  wire[0:0] nor_1628_nl;
  wire[0:0] mux_2441_nl;
  wire[0:0] nor_732_nl;
  wire[0:0] mux_2440_nl;
  wire[0:0] nor_733_nl;
  wire[0:0] mux_2439_nl;
  wire[0:0] nor_734_nl;
  wire[0:0] nor_735_nl;
  wire[0:0] mux_2438_nl;
  wire[0:0] mux_2437_nl;
  wire[0:0] nor_736_nl;
  wire[0:0] mux_2436_nl;
  wire[0:0] mux_2435_nl;
  wire[0:0] nor_737_nl;
  wire[0:0] nor_738_nl;
  wire[0:0] nor_739_nl;
  wire[0:0] nor_740_nl;
  wire[0:0] mux_2434_nl;
  wire[0:0] or_2495_nl;
  wire[0:0] mux_2433_nl;
  wire[0:0] or_2494_nl;
  wire[0:0] or_2490_nl;
  wire[0:0] mux_2448_nl;
  wire[0:0] mux_2447_nl;
  wire[0:0] nor_1612_nl;
  wire[0:0] mux_2453_nl;
  wire[0:0] nor_726_nl;
  wire[0:0] nor_727_nl;
  wire[0:0] mux_2681_nl;
  wire[0:0] mux_2708_nl;
  wire[0:0] nor_1575_nl;
  wire[0:0] or_2678_nl;
  wire[0:0] or_2677_nl;
  wire[0:0] mux_2756_nl;
  wire[0:0] or_2696_nl;
  wire[0:0] mux_2755_nl;
  wire[0:0] or_2695_nl;
  wire[0:0] mux_2754_nl;
  wire[0:0] or_2694_nl;
  wire[0:0] or_2693_nl;
  wire[0:0] mux_2753_nl;
  wire[0:0] mux_2752_nl;
  wire[0:0] or_2690_nl;
  wire[0:0] mux_2751_nl;
  wire[0:0] mux_2750_nl;
  wire[0:0] or_2689_nl;
  wire[0:0] or_2687_nl;
  wire[0:0] mux_2749_nl;
  wire[0:0] or_2686_nl;
  wire[0:0] or_2684_nl;
  wire[0:0] or_2682_nl;
  wire[0:0] mux_2748_nl;
  wire[0:0] mux_2747_nl;
  wire[0:0] or_2681_nl;
  wire[0:0] mux_2746_nl;
  wire[0:0] or_2676_nl;
  wire[0:0] mux_2744_nl;
  wire[0:0] or_2675_nl;
  wire[0:0] or_2674_nl;
  wire[0:0] or_2705_nl;
  wire[0:0] or_2704_nl;
  wire[0:0] mux_2839_nl;
  wire[0:0] mux_2838_nl;
  wire[0:0] mux_2837_nl;
  wire[0:0] or_2785_nl;
  wire[0:0] mux_2836_nl;
  wire[0:0] or_2784_nl;
  wire[0:0] mux_2835_nl;
  wire[0:0] mux_2834_nl;
  wire[0:0] mux_2833_nl;
  wire[0:0] mux_2832_nl;
  wire[0:0] mux_2831_nl;
  wire[0:0] mux_2830_nl;
  wire[0:0] nand_65_nl;
  wire[0:0] mux_2829_nl;
  wire[0:0] nand_394_nl;
  wire[0:0] mux_2828_nl;
  wire[0:0] mux_2827_nl;
  wire[0:0] or_2780_nl;
  wire[0:0] mux_2826_nl;
  wire[0:0] mux_2825_nl;
  wire[0:0] mux_2824_nl;
  wire[0:0] or_2778_nl;
  wire[0:0] mux_2823_nl;
  wire[0:0] mux_2822_nl;
  wire[0:0] mux_2821_nl;
  wire[0:0] mux_2820_nl;
  wire[0:0] or_2776_nl;
  wire[0:0] mux_2819_nl;
  wire[0:0] mux_2818_nl;
  wire[0:0] mux_2817_nl;
  wire[0:0] or_2775_nl;
  wire[0:0] mux_2816_nl;
  wire[0:0] or_2774_nl;
  wire[0:0] nand_64_nl;
  wire[0:0] mux_2815_nl;
  wire[0:0] mux_2814_nl;
  wire[0:0] mux_2813_nl;
  wire[0:0] or_2771_nl;
  wire[0:0] mux_2812_nl;
  wire[0:0] mux_2811_nl;
  wire[0:0] or_2770_nl;
  wire[0:0] mux_2810_nl;
  wire[0:0] mux_2809_nl;
  wire[0:0] mux_2808_nl;
  wire[0:0] mux_2807_nl;
  wire[0:0] nand_63_nl;
  wire[0:0] mux_2806_nl;
  wire[0:0] mux_2805_nl;
  wire[0:0] mux_2804_nl;
  wire[0:0] mux_2803_nl;
  wire[0:0] mux_2802_nl;
  wire[0:0] mux_2801_nl;
  wire[0:0] mux_2800_nl;
  wire[0:0] mux_2799_nl;
  wire[0:0] or_2759_nl;
  wire[0:0] mux_2798_nl;
  wire[0:0] mux_2797_nl;
  wire[0:0] mux_2795_nl;
  wire[0:0] nand_62_nl;
  wire[0:0] mux_2794_nl;
  wire[0:0] or_2754_nl;
  wire[0:0] mux_2793_nl;
  wire[0:0] mux_2792_nl;
  wire[0:0] mux_2791_nl;
  wire[0:0] or_2751_nl;
  wire[0:0] mux_2790_nl;
  wire[0:0] mux_2789_nl;
  wire[0:0] or_2747_nl;
  wire[0:0] mux_2788_nl;
  wire[0:0] or_2743_nl;
  wire[0:0] mux_2787_nl;
  wire[0:0] mux_2786_nl;
  wire[0:0] or_2740_nl;
  wire[0:0] mux_2858_nl;
  wire[0:0] mux_2875_nl;
  wire[0:0] or_2800_nl;
  wire[0:0] mux_2901_nl;
  wire[0:0] mux_2909_nl;
  wire[0:0] or_2840_nl;
  wire[0:0] mux_3002_nl;
  wire[0:0] mux_3001_nl;
  wire[0:0] nor_661_nl;
  wire[0:0] mux_3000_nl;
  wire[0:0] nor_662_nl;
  wire[0:0] mux_2999_nl;
  wire[0:0] or_2842_nl;
  wire[0:0] nor_663_nl;
  wire[0:0] nor_664_nl;
  wire[0:0] mux_2997_nl;
  wire[0:0] or_2836_nl;
  wire[0:0] or_2831_nl;
  wire[0:0] mux_2995_nl;
  wire[0:0] mux_2994_nl;
  wire[0:0] and_445_nl;
  wire[0:0] mux_2993_nl;
  wire[0:0] nor_665_nl;
  wire[0:0] mux_2992_nl;
  wire[0:0] nor_666_nl;
  wire[0:0] mux_2991_nl;
  wire[0:0] mux_2990_nl;
  wire[0:0] and_446_nl;
  wire[0:0] nor_668_nl;
  wire[0:0] nor_669_nl;
  wire[0:0] mux_3799_nl;
  wire[0:0] mux_3006_nl;
  wire[0:0] or_2848_nl;
  wire[0:0] or_2863_nl;
  wire[0:0] mux_3031_nl;
  wire[0:0] or_3367_nl;
  wire[0:0] mux_3321_nl;
  wire[0:0] or_3025_nl;
  wire[0:0] nand_149_nl;
  wire[0:0] mux_3320_nl;
  wire[0:0] mux_3319_nl;
  wire[0:0] or_3023_nl;
  wire[0:0] or_3022_nl;
  wire[0:0] mux_3342_nl;
  wire[0:0] or_3061_nl;
  wire[0:0] or_3087_nl;
  wire[0:0] or_12_nl;
  wire[0:0] mux_3416_nl;
  wire[0:0] mux_3427_nl;
  wire[0:0] mux_3426_nl;
  wire[0:0] mux_3422_nl;
  wire[0:0] mux_3431_nl;
  wire[0:0] mux_3430_nl;
  wire[0:0] mux_3433_nl;
  wire[0:0] mux_3436_nl;
  wire[0:0] mux_3452_nl;
  wire[0:0] mux_3451_nl;
  wire[0:0] mux_3450_nl;
  wire[0:0] mux_3449_nl;
  wire[0:0] mux_3448_nl;
  wire[0:0] mux_3447_nl;
  wire[0:0] mux_3446_nl;
  wire[0:0] mux_3445_nl;
  wire[0:0] mux_3444_nl;
  wire[0:0] mux_3443_nl;
  wire[0:0] mux_3442_nl;
  wire[0:0] mux_3441_nl;
  wire[0:0] mux_3440_nl;
  wire[0:0] mux_3439_nl;
  wire[0:0] mux_3438_nl;
  wire[0:0] mux_3413_nl;
  wire[0:0] mux_3412_nl;
  wire[0:0] or_3090_nl;
  wire[0:0] mux_3411_nl;
  wire[0:0] or_3088_nl;
  wire[0:0] mux_3455_nl;
  wire[0:0] mux_3454_nl;
  wire[0:0] mux_3460_nl;
  wire[0:0] mux_3462_nl;
  wire[0:0] mux_3471_nl;
  wire[0:0] mux_3470_nl;
  wire[0:0] mux_3469_nl;
  wire[0:0] mux_3468_nl;
  wire[0:0] mux_3467_nl;
  wire[0:0] mux_3466_nl;
  wire[0:0] mux_3465_nl;
  wire[0:0] or_3095_nl;
  wire[0:0] mux_3476_nl;
  wire[0:0] mux_3475_nl;
  wire[0:0] mux_3480_nl;
  wire[0:0] mux_3479_nl;
  wire[0:0] mux_3478_nl;
  wire[0:0] mux_3484_nl;
  wire[0:0] mux_3490_nl;
  wire[0:0] mux_3489_nl;
  wire[0:0] mux_3488_nl;
  wire[0:0] mux_3493_nl;
  wire[0:0] mux_3492_nl;
  wire[0:0] mux_3487_nl;
  wire[0:0] mux_3486_nl;
  wire[0:0] mux_3483_nl;
  wire[0:0] mux_3482_nl;
  wire[0:0] mux_3506_nl;
  wire[0:0] nor_603_nl;
  wire[0:0] mux_3505_nl;
  wire[0:0] or_3117_nl;
  wire[0:0] mux_3504_nl;
  wire[0:0] or_3116_nl;
  wire[0:0] or_3115_nl;
  wire[0:0] mux_3503_nl;
  wire[0:0] and_376_nl;
  wire[0:0] mux_3502_nl;
  wire[0:0] mux_3501_nl;
  wire[0:0] nor_604_nl;
  wire[0:0] nor_605_nl;
  wire[0:0] mux_3500_nl;
  wire[0:0] nor_606_nl;
  wire[0:0] nor_607_nl;
  wire[0:0] nor_608_nl;
  wire[0:0] mux_3499_nl;
  wire[0:0] mux_3498_nl;
  wire[0:0] or_3104_nl;
  wire[0:0] mux_3497_nl;
  wire[0:0] or_3099_nl;
  wire[0:0] mux_3495_nl;
  wire[0:0] or_3098_nl;
  wire[0:0] or_3097_nl;
  wire[0:0] or_3154_nl;
  wire[0:0] mux_3534_nl;
  wire[0:0] mux_3533_nl;
  wire[0:0] nor_584_nl;
  wire[0:0] nor_585_nl;
  wire[0:0] mux_3532_nl;
  wire[0:0] nand_103_nl;
  wire[0:0] or_3157_nl;
  wire[0:0] mux_3531_nl;
  wire[0:0] and_371_nl;
  wire[0:0] mux_3530_nl;
  wire[0:0] nor_586_nl;
  wire[0:0] nor_587_nl;
  wire[0:0] nor_588_nl;
  wire[0:0] mux_3528_nl;
  wire[0:0] mux_3527_nl;
  wire[0:0] and_372_nl;
  wire[0:0] mux_3526_nl;
  wire[0:0] nor_589_nl;
  wire[0:0] and_373_nl;
  wire[0:0] mux_3525_nl;
  wire[0:0] nor_590_nl;
  wire[0:0] mux_3524_nl;
  wire[0:0] nor_591_nl;
  wire[0:0] nor_593_nl;
  wire[0:0] mux_3522_nl;
  wire[0:0] or_3142_nl;
  wire[0:0] or_3141_nl;
  wire[0:0] or_3178_nl;
  wire[0:0] mux_460_nl;
  wire[0:0] or_3199_nl;
  wire[0:0] or_3222_nl;
  wire[0:0] or_3221_nl;
  wire[0:0] or_127_nl;
  wire[0:0] or_134_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] mux_3738_nl;
  wire[0:0] mux_2657_nl;
  wire[0:0] mux_2656_nl;
  wire[0:0] mux_2655_nl;
  wire[0:0] mux_2654_nl;
  wire[0:0] nor_693_nl;
  wire[0:0] mux_2653_nl;
  wire[0:0] and_467_nl;
  wire[2:0] STAGE_LOOP_acc_nl;
  wire[3:0] nl_STAGE_LOOP_acc_nl;
  wire[0:0] and_139_nl;
  wire[0:0] mux_1093_nl;
  wire[0:0] mux_1092_nl;
  wire[0:0] mux_1091_nl;
  wire[0:0] or_522_nl;
  wire[0:0] or_520_nl;
  wire[0:0] mux_1090_nl;
  wire[0:0] mux_1089_nl;
  wire[0:0] or_518_nl;
  wire[0:0] mux_1088_nl;
  wire[0:0] or_516_nl;
  wire[0:0] mux_1087_nl;
  wire[0:0] or_515_nl;
  wire[0:0] or_513_nl;
  wire[0:0] mux_1086_nl;
  wire[0:0] mux_1085_nl;
  wire[0:0] mux_1084_nl;
  wire[0:0] or_512_nl;
  wire[0:0] or_511_nl;
  wire[0:0] mux_1083_nl;
  wire[0:0] or_506_nl;
  wire[0:0] or_504_nl;
  wire[0:0] and_144_nl;
  wire[0:0] mux_1094_nl;
  wire[0:0] nor_1513_nl;
  wire[0:0] nor_1514_nl;
  wire[0:0] and_153_nl;
  wire[0:0] mux_1095_nl;
  wire[0:0] nor_1511_nl;
  wire[0:0] nor_1512_nl;
  wire[0:0] and_162_nl;
  wire[0:0] mux_1096_nl;
  wire[0:0] nor_1509_nl;
  wire[0:0] nor_1510_nl;
  wire[0:0] and_170_nl;
  wire[0:0] mux_1097_nl;
  wire[0:0] and_758_nl;
  wire[0:0] nor_1508_nl;
  wire[0:0] and_180_nl;
  wire[0:0] mux_1098_nl;
  wire[0:0] nor_1505_nl;
  wire[0:0] nor_1506_nl;
  wire[0:0] and_187_nl;
  wire[0:0] mux_1099_nl;
  wire[0:0] nor_1503_nl;
  wire[0:0] nor_1504_nl;
  wire[0:0] and_195_nl;
  wire[0:0] mux_1100_nl;
  wire[0:0] nor_1501_nl;
  wire[0:0] nor_1502_nl;
  wire[0:0] and_201_nl;
  wire[0:0] mux_1101_nl;
  wire[0:0] nor_1499_nl;
  wire[0:0] nor_1500_nl;
  wire[0:0] nor_1625_nl;
  wire[0:0] mux_1102_nl;
  wire[0:0] or_3445_nl;
  wire[0:0] or_3446_nl;
  wire[0:0] and_213_nl;
  wire[0:0] mux_1103_nl;
  wire[0:0] nor_1495_nl;
  wire[0:0] nor_1496_nl;
  wire[0:0] and_219_nl;
  wire[0:0] mux_1104_nl;
  wire[0:0] nor_1493_nl;
  wire[0:0] nor_1494_nl;
  wire[0:0] and_225_nl;
  wire[0:0] mux_1105_nl;
  wire[0:0] and_760_nl;
  wire[0:0] nor_1492_nl;
  wire[0:0] and_235_nl;
  wire[0:0] mux_1106_nl;
  wire[0:0] nor_1489_nl;
  wire[0:0] and_748_nl;
  wire[0:0] and_241_nl;
  wire[0:0] mux_1107_nl;
  wire[0:0] and_627_nl;
  wire[0:0] nor_1488_nl;
  wire[0:0] and_249_nl;
  wire[0:0] mux_1108_nl;
  wire[0:0] nor_1486_nl;
  wire[0:0] nor_1487_nl;
  wire[0:0] mux_1138_nl;
  wire[0:0] mux_1137_nl;
  wire[0:0] mux_1136_nl;
  wire[0:0] nor_1471_nl;
  wire[0:0] mux_1135_nl;
  wire[0:0] mux_1134_nl;
  wire[0:0] or_618_nl;
  wire[0:0] or_617_nl;
  wire[0:0] or_615_nl;
  wire[0:0] nor_1472_nl;
  wire[0:0] mux_1133_nl;
  wire[0:0] nor_1473_nl;
  wire[0:0] mux_1132_nl;
  wire[0:0] nor_1474_nl;
  wire[0:0] mux_1131_nl;
  wire[0:0] nor_1475_nl;
  wire[0:0] nor_1476_nl;
  wire[0:0] mux_1130_nl;
  wire[0:0] and_626_nl;
  wire[0:0] mux_1129_nl;
  wire[0:0] or_606_nl;
  wire[0:0] mux_1128_nl;
  wire[0:0] or_605_nl;
  wire[0:0] mux_1127_nl;
  wire[0:0] nor_1477_nl;
  wire[0:0] mux_1126_nl;
  wire[0:0] or_602_nl;
  wire[0:0] mux_1125_nl;
  wire[0:0] or_600_nl;
  wire[0:0] nor_1478_nl;
  wire[0:0] mux_1124_nl;
  wire[0:0] mux_1123_nl;
  wire[0:0] mux_1122_nl;
  wire[0:0] nor_1479_nl;
  wire[0:0] mux_1121_nl;
  wire[0:0] or_596_nl;
  wire[0:0] or_594_nl;
  wire[0:0] nor_1480_nl;
  wire[0:0] mux_1120_nl;
  wire[0:0] mux_1119_nl;
  wire[0:0] or_590_nl;
  wire[0:0] nor_1481_nl;
  wire[0:0] mux_1118_nl;
  wire[0:0] mux_1117_nl;
  wire[0:0] or_583_nl;
  wire[0:0] or_581_nl;
  wire[0:0] mux_1115_nl;
  wire[0:0] nor_1482_nl;
  wire[0:0] mux_1114_nl;
  wire[0:0] mux_1113_nl;
  wire[0:0] or_576_nl;
  wire[0:0] or_574_nl;
  wire[0:0] mux_1112_nl;
  wire[0:0] or_573_nl;
  wire[0:0] or_572_nl;
  wire[0:0] mux_1111_nl;
  wire[0:0] nor_1483_nl;
  wire[0:0] mux_1110_nl;
  wire[0:0] nor_1484_nl;
  wire[0:0] nor_1485_nl;
  wire[0:0] mux_1109_nl;
  wire[0:0] or_567_nl;
  wire[0:0] or_565_nl;
  wire[0:0] mux_1171_nl;
  wire[0:0] and_623_nl;
  wire[0:0] mux_1170_nl;
  wire[0:0] nor_1440_nl;
  wire[0:0] mux_1169_nl;
  wire[0:0] or_674_nl;
  wire[0:0] or_673_nl;
  wire[0:0] mux_1168_nl;
  wire[0:0] nor_1441_nl;
  wire[0:0] mux_1167_nl;
  wire[0:0] nor_1442_nl;
  wire[0:0] nor_1443_nl;
  wire[0:0] mux_1166_nl;
  wire[0:0] mux_1165_nl;
  wire[0:0] mux_1164_nl;
  wire[0:0] nor_1444_nl;
  wire[0:0] mux_1163_nl;
  wire[0:0] mux_1162_nl;
  wire[0:0] nor_1446_nl;
  wire[0:0] nor_1447_nl;
  wire[0:0] or_660_nl;
  wire[0:0] mux_1161_nl;
  wire[0:0] nor_1448_nl;
  wire[0:0] mux_1160_nl;
  wire[0:0] nor_1449_nl;
  wire[0:0] nor_1450_nl;
  wire[0:0] mux_1159_nl;
  wire[0:0] mux_1158_nl;
  wire[0:0] nor_1451_nl;
  wire[0:0] nor_1452_nl;
  wire[0:0] nor_1453_nl;
  wire[0:0] mux_1156_nl;
  wire[0:0] mux_1155_nl;
  wire[0:0] mux_1154_nl;
  wire[0:0] mux_1153_nl;
  wire[0:0] and_624_nl;
  wire[0:0] mux_1152_nl;
  wire[0:0] nor_1454_nl;
  wire[0:0] nor_1455_nl;
  wire[0:0] and_625_nl;
  wire[0:0] mux_1151_nl;
  wire[0:0] nor_1456_nl;
  wire[0:0] nor_1457_nl;
  wire[0:0] mux_1150_nl;
  wire[0:0] nor_1458_nl;
  wire[0:0] nor_1459_nl;
  wire[0:0] mux_1148_nl;
  wire[0:0] nor_1460_nl;
  wire[0:0] mux_1147_nl;
  wire[0:0] nor_1461_nl;
  wire[0:0] nor_1462_nl;
  wire[0:0] mux_1146_nl;
  wire[0:0] mux_1145_nl;
  wire[0:0] nor_1463_nl;
  wire[0:0] nor_1464_nl;
  wire[0:0] mux_1144_nl;
  wire[0:0] mux_1143_nl;
  wire[0:0] mux_1142_nl;
  wire[0:0] nor_1465_nl;
  wire[0:0] mux_1141_nl;
  wire[0:0] nor_1466_nl;
  wire[0:0] nor_1467_nl;
  wire[0:0] nor_1468_nl;
  wire[0:0] mux_1140_nl;
  wire[0:0] nor_1469_nl;
  wire[0:0] nor_1470_nl;
  wire[0:0] mux_1202_nl;
  wire[0:0] mux_1201_nl;
  wire[0:0] mux_1200_nl;
  wire[0:0] nor_1425_nl;
  wire[0:0] mux_1199_nl;
  wire[0:0] mux_1198_nl;
  wire[0:0] or_729_nl;
  wire[0:0] or_728_nl;
  wire[0:0] or_726_nl;
  wire[0:0] nor_1426_nl;
  wire[0:0] mux_1197_nl;
  wire[0:0] nor_1427_nl;
  wire[0:0] mux_1196_nl;
  wire[0:0] nor_1428_nl;
  wire[0:0] mux_1195_nl;
  wire[0:0] nor_1429_nl;
  wire[0:0] nor_1430_nl;
  wire[0:0] mux_1194_nl;
  wire[0:0] and_622_nl;
  wire[0:0] mux_1193_nl;
  wire[0:0] or_717_nl;
  wire[0:0] mux_1192_nl;
  wire[0:0] or_716_nl;
  wire[0:0] mux_1191_nl;
  wire[0:0] nor_1431_nl;
  wire[0:0] mux_1190_nl;
  wire[0:0] or_713_nl;
  wire[0:0] mux_1189_nl;
  wire[0:0] or_711_nl;
  wire[0:0] nor_1432_nl;
  wire[0:0] mux_1188_nl;
  wire[0:0] mux_1187_nl;
  wire[0:0] mux_1186_nl;
  wire[0:0] nor_1433_nl;
  wire[0:0] mux_1185_nl;
  wire[0:0] or_707_nl;
  wire[0:0] or_705_nl;
  wire[0:0] nor_1434_nl;
  wire[0:0] mux_1184_nl;
  wire[0:0] mux_1183_nl;
  wire[0:0] or_701_nl;
  wire[0:0] nor_1435_nl;
  wire[0:0] mux_1182_nl;
  wire[0:0] mux_1181_nl;
  wire[0:0] or_694_nl;
  wire[0:0] or_692_nl;
  wire[0:0] mux_1179_nl;
  wire[0:0] nor_1436_nl;
  wire[0:0] mux_1178_nl;
  wire[0:0] mux_1177_nl;
  wire[0:0] or_687_nl;
  wire[0:0] or_685_nl;
  wire[0:0] mux_1176_nl;
  wire[0:0] or_684_nl;
  wire[0:0] or_683_nl;
  wire[0:0] mux_1175_nl;
  wire[0:0] nor_1437_nl;
  wire[0:0] mux_1174_nl;
  wire[0:0] nor_1438_nl;
  wire[0:0] nor_1439_nl;
  wire[0:0] mux_1173_nl;
  wire[0:0] or_678_nl;
  wire[0:0] or_676_nl;
  wire[0:0] mux_1235_nl;
  wire[0:0] and_619_nl;
  wire[0:0] mux_1234_nl;
  wire[0:0] nor_1394_nl;
  wire[0:0] mux_1233_nl;
  wire[0:0] or_785_nl;
  wire[0:0] or_784_nl;
  wire[0:0] mux_1232_nl;
  wire[0:0] nor_1395_nl;
  wire[0:0] mux_1231_nl;
  wire[0:0] nor_1396_nl;
  wire[0:0] nor_1397_nl;
  wire[0:0] mux_1230_nl;
  wire[0:0] mux_1229_nl;
  wire[0:0] mux_1228_nl;
  wire[0:0] nor_1398_nl;
  wire[0:0] mux_1227_nl;
  wire[0:0] mux_1226_nl;
  wire[0:0] nor_1400_nl;
  wire[0:0] nor_1401_nl;
  wire[0:0] or_771_nl;
  wire[0:0] mux_1225_nl;
  wire[0:0] nor_1402_nl;
  wire[0:0] mux_1224_nl;
  wire[0:0] nor_1403_nl;
  wire[0:0] nor_1404_nl;
  wire[0:0] mux_1223_nl;
  wire[0:0] mux_1222_nl;
  wire[0:0] nor_1405_nl;
  wire[0:0] nor_1406_nl;
  wire[0:0] nor_1407_nl;
  wire[0:0] mux_1220_nl;
  wire[0:0] mux_1219_nl;
  wire[0:0] mux_1218_nl;
  wire[0:0] mux_1217_nl;
  wire[0:0] and_620_nl;
  wire[0:0] mux_1216_nl;
  wire[0:0] nor_1408_nl;
  wire[0:0] nor_1409_nl;
  wire[0:0] and_621_nl;
  wire[0:0] mux_1215_nl;
  wire[0:0] nor_1410_nl;
  wire[0:0] nor_1411_nl;
  wire[0:0] mux_1214_nl;
  wire[0:0] nor_1412_nl;
  wire[0:0] nor_1413_nl;
  wire[0:0] mux_1212_nl;
  wire[0:0] nor_1414_nl;
  wire[0:0] mux_1211_nl;
  wire[0:0] nor_1415_nl;
  wire[0:0] nor_1416_nl;
  wire[0:0] mux_1210_nl;
  wire[0:0] mux_1209_nl;
  wire[0:0] nor_1417_nl;
  wire[0:0] nor_1418_nl;
  wire[0:0] mux_1208_nl;
  wire[0:0] mux_1207_nl;
  wire[0:0] mux_1206_nl;
  wire[0:0] nor_1419_nl;
  wire[0:0] mux_1205_nl;
  wire[0:0] nor_1420_nl;
  wire[0:0] nor_1421_nl;
  wire[0:0] nor_1422_nl;
  wire[0:0] mux_1204_nl;
  wire[0:0] nor_1423_nl;
  wire[0:0] nor_1424_nl;
  wire[0:0] mux_1266_nl;
  wire[0:0] mux_1265_nl;
  wire[0:0] mux_1264_nl;
  wire[0:0] nor_1379_nl;
  wire[0:0] mux_1263_nl;
  wire[0:0] mux_1262_nl;
  wire[0:0] or_839_nl;
  wire[0:0] or_838_nl;
  wire[0:0] or_836_nl;
  wire[0:0] nor_1380_nl;
  wire[0:0] mux_1261_nl;
  wire[0:0] nor_1381_nl;
  wire[0:0] mux_1260_nl;
  wire[0:0] nor_1382_nl;
  wire[0:0] mux_1259_nl;
  wire[0:0] nor_1383_nl;
  wire[0:0] nor_1384_nl;
  wire[0:0] mux_1258_nl;
  wire[0:0] and_618_nl;
  wire[0:0] mux_1257_nl;
  wire[0:0] or_827_nl;
  wire[0:0] mux_1256_nl;
  wire[0:0] or_826_nl;
  wire[0:0] mux_1255_nl;
  wire[0:0] nor_1385_nl;
  wire[0:0] mux_1254_nl;
  wire[0:0] or_823_nl;
  wire[0:0] mux_1253_nl;
  wire[0:0] or_821_nl;
  wire[0:0] nor_1386_nl;
  wire[0:0] mux_1252_nl;
  wire[0:0] mux_1251_nl;
  wire[0:0] mux_1250_nl;
  wire[0:0] nor_1387_nl;
  wire[0:0] mux_1249_nl;
  wire[0:0] or_817_nl;
  wire[0:0] or_815_nl;
  wire[0:0] nor_1388_nl;
  wire[0:0] mux_1248_nl;
  wire[0:0] mux_1247_nl;
  wire[0:0] or_809_nl;
  wire[0:0] nor_1389_nl;
  wire[0:0] mux_1246_nl;
  wire[0:0] mux_1245_nl;
  wire[0:0] or_805_nl;
  wire[0:0] or_803_nl;
  wire[0:0] mux_1243_nl;
  wire[0:0] nor_1390_nl;
  wire[0:0] mux_1242_nl;
  wire[0:0] mux_1241_nl;
  wire[0:0] or_798_nl;
  wire[0:0] or_796_nl;
  wire[0:0] mux_1240_nl;
  wire[0:0] or_795_nl;
  wire[0:0] or_794_nl;
  wire[0:0] mux_1239_nl;
  wire[0:0] nor_1391_nl;
  wire[0:0] mux_1238_nl;
  wire[0:0] nor_1392_nl;
  wire[0:0] nor_1393_nl;
  wire[0:0] mux_1237_nl;
  wire[0:0] or_789_nl;
  wire[0:0] or_787_nl;
  wire[0:0] mux_1299_nl;
  wire[0:0] and_615_nl;
  wire[0:0] mux_1298_nl;
  wire[0:0] nor_1348_nl;
  wire[0:0] mux_1297_nl;
  wire[0:0] or_895_nl;
  wire[0:0] or_894_nl;
  wire[0:0] mux_1296_nl;
  wire[0:0] nor_1349_nl;
  wire[0:0] mux_1295_nl;
  wire[0:0] nor_1350_nl;
  wire[0:0] nor_1351_nl;
  wire[0:0] mux_1294_nl;
  wire[0:0] mux_1293_nl;
  wire[0:0] mux_1292_nl;
  wire[0:0] nor_1352_nl;
  wire[0:0] mux_1291_nl;
  wire[0:0] mux_1290_nl;
  wire[0:0] nor_1354_nl;
  wire[0:0] nor_1355_nl;
  wire[0:0] or_881_nl;
  wire[0:0] mux_1289_nl;
  wire[0:0] nor_1356_nl;
  wire[0:0] mux_1288_nl;
  wire[0:0] nor_1357_nl;
  wire[0:0] nor_1358_nl;
  wire[0:0] mux_1287_nl;
  wire[0:0] mux_1286_nl;
  wire[0:0] nor_1359_nl;
  wire[0:0] nor_1360_nl;
  wire[0:0] nor_1361_nl;
  wire[0:0] mux_1284_nl;
  wire[0:0] mux_1283_nl;
  wire[0:0] mux_1282_nl;
  wire[0:0] mux_1281_nl;
  wire[0:0] and_616_nl;
  wire[0:0] mux_1280_nl;
  wire[0:0] nor_1362_nl;
  wire[0:0] nor_1363_nl;
  wire[0:0] and_617_nl;
  wire[0:0] mux_1279_nl;
  wire[0:0] nor_1364_nl;
  wire[0:0] nor_1365_nl;
  wire[0:0] mux_1278_nl;
  wire[0:0] nor_1366_nl;
  wire[0:0] nor_1367_nl;
  wire[0:0] mux_1276_nl;
  wire[0:0] nor_1368_nl;
  wire[0:0] mux_1275_nl;
  wire[0:0] nor_1369_nl;
  wire[0:0] nor_1370_nl;
  wire[0:0] mux_1274_nl;
  wire[0:0] mux_1273_nl;
  wire[0:0] nor_1371_nl;
  wire[0:0] nor_1372_nl;
  wire[0:0] mux_1272_nl;
  wire[0:0] mux_1271_nl;
  wire[0:0] mux_1270_nl;
  wire[0:0] nor_1373_nl;
  wire[0:0] mux_1269_nl;
  wire[0:0] nor_1374_nl;
  wire[0:0] nor_1375_nl;
  wire[0:0] nor_1376_nl;
  wire[0:0] mux_1268_nl;
  wire[0:0] nor_1377_nl;
  wire[0:0] nor_1378_nl;
  wire[0:0] mux_1330_nl;
  wire[0:0] mux_1329_nl;
  wire[0:0] mux_1328_nl;
  wire[0:0] nor_1333_nl;
  wire[0:0] mux_1327_nl;
  wire[0:0] mux_1326_nl;
  wire[0:0] or_949_nl;
  wire[0:0] nand_404_nl;
  wire[0:0] or_946_nl;
  wire[0:0] nor_1334_nl;
  wire[0:0] mux_1325_nl;
  wire[0:0] nor_1335_nl;
  wire[0:0] mux_1324_nl;
  wire[0:0] nor_1336_nl;
  wire[0:0] mux_1323_nl;
  wire[0:0] nor_1337_nl;
  wire[0:0] nor_1338_nl;
  wire[0:0] mux_1322_nl;
  wire[0:0] and_614_nl;
  wire[0:0] mux_1321_nl;
  wire[0:0] nand_327_nl;
  wire[0:0] mux_1320_nl;
  wire[0:0] or_936_nl;
  wire[0:0] mux_1319_nl;
  wire[0:0] nor_1339_nl;
  wire[0:0] mux_1318_nl;
  wire[0:0] or_933_nl;
  wire[0:0] mux_1317_nl;
  wire[0:0] or_931_nl;
  wire[0:0] nor_1340_nl;
  wire[0:0] mux_1316_nl;
  wire[0:0] mux_1315_nl;
  wire[0:0] mux_1314_nl;
  wire[0:0] nor_1341_nl;
  wire[0:0] mux_1313_nl;
  wire[0:0] or_927_nl;
  wire[0:0] or_925_nl;
  wire[0:0] nor_1342_nl;
  wire[0:0] mux_1312_nl;
  wire[0:0] mux_1311_nl;
  wire[0:0] or_919_nl;
  wire[0:0] nor_1343_nl;
  wire[0:0] mux_1310_nl;
  wire[0:0] mux_1309_nl;
  wire[0:0] or_915_nl;
  wire[0:0] or_913_nl;
  wire[0:0] mux_1307_nl;
  wire[0:0] nor_1344_nl;
  wire[0:0] mux_1306_nl;
  wire[0:0] mux_1305_nl;
  wire[0:0] or_908_nl;
  wire[0:0] or_906_nl;
  wire[0:0] mux_1304_nl;
  wire[0:0] or_905_nl;
  wire[0:0] or_904_nl;
  wire[0:0] mux_1303_nl;
  wire[0:0] nor_1345_nl;
  wire[0:0] mux_1302_nl;
  wire[0:0] nor_1346_nl;
  wire[0:0] nor_1347_nl;
  wire[0:0] mux_1301_nl;
  wire[0:0] or_899_nl;
  wire[0:0] or_897_nl;
  wire[0:0] mux_1363_nl;
  wire[0:0] and_611_nl;
  wire[0:0] mux_1362_nl;
  wire[0:0] nor_1302_nl;
  wire[0:0] mux_1361_nl;
  wire[0:0] or_1005_nl;
  wire[0:0] or_1004_nl;
  wire[0:0] mux_1360_nl;
  wire[0:0] nor_1303_nl;
  wire[0:0] mux_1359_nl;
  wire[0:0] nor_1304_nl;
  wire[0:0] nor_1305_nl;
  wire[0:0] mux_1358_nl;
  wire[0:0] mux_1357_nl;
  wire[0:0] mux_1356_nl;
  wire[0:0] nor_1306_nl;
  wire[0:0] mux_1355_nl;
  wire[0:0] mux_1354_nl;
  wire[0:0] nor_1308_nl;
  wire[0:0] nor_1309_nl;
  wire[0:0] or_991_nl;
  wire[0:0] mux_1353_nl;
  wire[0:0] nor_1310_nl;
  wire[0:0] mux_1352_nl;
  wire[0:0] nor_1311_nl;
  wire[0:0] nor_1312_nl;
  wire[0:0] mux_1351_nl;
  wire[0:0] mux_1350_nl;
  wire[0:0] nor_1313_nl;
  wire[0:0] nor_1314_nl;
  wire[0:0] nor_1315_nl;
  wire[0:0] mux_1348_nl;
  wire[0:0] mux_1347_nl;
  wire[0:0] mux_1346_nl;
  wire[0:0] mux_1345_nl;
  wire[0:0] and_612_nl;
  wire[0:0] mux_1344_nl;
  wire[0:0] nor_1316_nl;
  wire[0:0] nor_1317_nl;
  wire[0:0] and_613_nl;
  wire[0:0] mux_1343_nl;
  wire[0:0] nor_1318_nl;
  wire[0:0] nor_1319_nl;
  wire[0:0] mux_1342_nl;
  wire[0:0] nor_1320_nl;
  wire[0:0] nor_1321_nl;
  wire[0:0] mux_1340_nl;
  wire[0:0] nor_1322_nl;
  wire[0:0] mux_1339_nl;
  wire[0:0] nor_1323_nl;
  wire[0:0] nor_1324_nl;
  wire[0:0] mux_1338_nl;
  wire[0:0] mux_1337_nl;
  wire[0:0] nor_1325_nl;
  wire[0:0] nor_1326_nl;
  wire[0:0] mux_1336_nl;
  wire[0:0] mux_1335_nl;
  wire[0:0] mux_1334_nl;
  wire[0:0] nor_1327_nl;
  wire[0:0] mux_1333_nl;
  wire[0:0] nor_1328_nl;
  wire[0:0] nor_1329_nl;
  wire[0:0] nor_1330_nl;
  wire[0:0] mux_1332_nl;
  wire[0:0] nor_1331_nl;
  wire[0:0] nor_1332_nl;
  wire[0:0] mux_1394_nl;
  wire[0:0] mux_1393_nl;
  wire[0:0] mux_1392_nl;
  wire[0:0] nor_1287_nl;
  wire[0:0] mux_1391_nl;
  wire[0:0] mux_1390_nl;
  wire[0:0] or_1060_nl;
  wire[0:0] or_1059_nl;
  wire[0:0] or_1057_nl;
  wire[0:0] nor_1288_nl;
  wire[0:0] mux_1389_nl;
  wire[0:0] nor_1289_nl;
  wire[0:0] mux_1388_nl;
  wire[0:0] nor_1290_nl;
  wire[0:0] mux_1387_nl;
  wire[0:0] nor_1291_nl;
  wire[0:0] nor_1292_nl;
  wire[0:0] mux_1386_nl;
  wire[0:0] and_610_nl;
  wire[0:0] mux_1385_nl;
  wire[0:0] or_1048_nl;
  wire[0:0] mux_1384_nl;
  wire[0:0] or_1047_nl;
  wire[0:0] mux_1383_nl;
  wire[0:0] nor_1293_nl;
  wire[0:0] mux_1382_nl;
  wire[0:0] or_1044_nl;
  wire[0:0] mux_1381_nl;
  wire[0:0] or_1042_nl;
  wire[0:0] nor_1294_nl;
  wire[0:0] mux_1380_nl;
  wire[0:0] mux_1379_nl;
  wire[0:0] mux_1378_nl;
  wire[0:0] nor_1295_nl;
  wire[0:0] mux_1377_nl;
  wire[0:0] or_1038_nl;
  wire[0:0] or_1036_nl;
  wire[0:0] nor_1296_nl;
  wire[0:0] mux_1376_nl;
  wire[0:0] mux_1375_nl;
  wire[0:0] or_1032_nl;
  wire[0:0] nor_1297_nl;
  wire[0:0] mux_1374_nl;
  wire[0:0] mux_1373_nl;
  wire[0:0] or_1025_nl;
  wire[0:0] or_1023_nl;
  wire[0:0] mux_1371_nl;
  wire[0:0] nor_1298_nl;
  wire[0:0] mux_1370_nl;
  wire[0:0] mux_1369_nl;
  wire[0:0] or_1018_nl;
  wire[0:0] or_1016_nl;
  wire[0:0] mux_1368_nl;
  wire[0:0] or_1015_nl;
  wire[0:0] or_1014_nl;
  wire[0:0] mux_1367_nl;
  wire[0:0] nor_1299_nl;
  wire[0:0] mux_1366_nl;
  wire[0:0] nor_1300_nl;
  wire[0:0] nor_1301_nl;
  wire[0:0] mux_1365_nl;
  wire[0:0] or_1009_nl;
  wire[0:0] or_1007_nl;
  wire[0:0] mux_1427_nl;
  wire[0:0] and_607_nl;
  wire[0:0] mux_1426_nl;
  wire[0:0] nor_1256_nl;
  wire[0:0] mux_1425_nl;
  wire[0:0] or_1116_nl;
  wire[0:0] or_1115_nl;
  wire[0:0] mux_1424_nl;
  wire[0:0] nor_1257_nl;
  wire[0:0] mux_1423_nl;
  wire[0:0] nor_1258_nl;
  wire[0:0] nor_1259_nl;
  wire[0:0] mux_1422_nl;
  wire[0:0] mux_1421_nl;
  wire[0:0] mux_1420_nl;
  wire[0:0] nor_1260_nl;
  wire[0:0] mux_1419_nl;
  wire[0:0] mux_1418_nl;
  wire[0:0] nor_1262_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] or_1102_nl;
  wire[0:0] mux_1417_nl;
  wire[0:0] nor_1264_nl;
  wire[0:0] mux_1416_nl;
  wire[0:0] nor_1265_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] mux_1415_nl;
  wire[0:0] mux_1414_nl;
  wire[0:0] nor_1267_nl;
  wire[0:0] nor_1268_nl;
  wire[0:0] nor_1269_nl;
  wire[0:0] mux_1412_nl;
  wire[0:0] mux_1411_nl;
  wire[0:0] mux_1410_nl;
  wire[0:0] mux_1409_nl;
  wire[0:0] and_608_nl;
  wire[0:0] mux_1408_nl;
  wire[0:0] nor_1270_nl;
  wire[0:0] nor_1271_nl;
  wire[0:0] and_609_nl;
  wire[0:0] mux_1407_nl;
  wire[0:0] nor_1272_nl;
  wire[0:0] nor_1273_nl;
  wire[0:0] mux_1406_nl;
  wire[0:0] nor_1274_nl;
  wire[0:0] nor_1275_nl;
  wire[0:0] mux_1404_nl;
  wire[0:0] nor_1276_nl;
  wire[0:0] mux_1403_nl;
  wire[0:0] nor_1277_nl;
  wire[0:0] nor_1278_nl;
  wire[0:0] mux_1402_nl;
  wire[0:0] mux_1401_nl;
  wire[0:0] nor_1279_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] mux_1400_nl;
  wire[0:0] mux_1399_nl;
  wire[0:0] mux_1398_nl;
  wire[0:0] nor_1281_nl;
  wire[0:0] mux_1397_nl;
  wire[0:0] nor_1282_nl;
  wire[0:0] nor_1283_nl;
  wire[0:0] nor_1284_nl;
  wire[0:0] mux_1396_nl;
  wire[0:0] nor_1285_nl;
  wire[0:0] nor_1286_nl;
  wire[0:0] mux_1458_nl;
  wire[0:0] mux_1457_nl;
  wire[0:0] mux_1456_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] mux_1455_nl;
  wire[0:0] mux_1454_nl;
  wire[0:0] or_1171_nl;
  wire[0:0] nand_403_nl;
  wire[0:0] or_1168_nl;
  wire[0:0] nor_1242_nl;
  wire[0:0] mux_1453_nl;
  wire[0:0] nor_1243_nl;
  wire[0:0] mux_1452_nl;
  wire[0:0] nor_1244_nl;
  wire[0:0] mux_1451_nl;
  wire[0:0] nor_1245_nl;
  wire[0:0] nor_1246_nl;
  wire[0:0] mux_1450_nl;
  wire[0:0] and_606_nl;
  wire[0:0] mux_1449_nl;
  wire[0:0] nand_318_nl;
  wire[0:0] mux_1448_nl;
  wire[0:0] or_1158_nl;
  wire[0:0] mux_1447_nl;
  wire[0:0] nor_1247_nl;
  wire[0:0] mux_1446_nl;
  wire[0:0] or_1155_nl;
  wire[0:0] mux_1445_nl;
  wire[0:0] or_1153_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] mux_1444_nl;
  wire[0:0] mux_1443_nl;
  wire[0:0] mux_1442_nl;
  wire[0:0] nor_1249_nl;
  wire[0:0] mux_1441_nl;
  wire[0:0] or_1149_nl;
  wire[0:0] or_1147_nl;
  wire[0:0] nor_1250_nl;
  wire[0:0] mux_1440_nl;
  wire[0:0] mux_1439_nl;
  wire[0:0] or_1143_nl;
  wire[0:0] nor_1251_nl;
  wire[0:0] mux_1438_nl;
  wire[0:0] mux_1437_nl;
  wire[0:0] or_1136_nl;
  wire[0:0] or_1134_nl;
  wire[0:0] mux_1435_nl;
  wire[0:0] nor_1252_nl;
  wire[0:0] mux_1434_nl;
  wire[0:0] mux_1433_nl;
  wire[0:0] or_1129_nl;
  wire[0:0] or_1127_nl;
  wire[0:0] mux_1432_nl;
  wire[0:0] or_1126_nl;
  wire[0:0] or_1125_nl;
  wire[0:0] mux_1431_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] mux_1430_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] nor_1255_nl;
  wire[0:0] mux_1429_nl;
  wire[0:0] or_1120_nl;
  wire[0:0] or_1118_nl;
  wire[0:0] mux_1491_nl;
  wire[0:0] and_603_nl;
  wire[0:0] mux_1490_nl;
  wire[0:0] nor_1210_nl;
  wire[0:0] mux_1489_nl;
  wire[0:0] or_1227_nl;
  wire[0:0] or_1226_nl;
  wire[0:0] mux_1488_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] mux_1487_nl;
  wire[0:0] nor_1212_nl;
  wire[0:0] nor_1213_nl;
  wire[0:0] mux_1486_nl;
  wire[0:0] mux_1485_nl;
  wire[0:0] mux_1484_nl;
  wire[0:0] nor_1214_nl;
  wire[0:0] mux_1483_nl;
  wire[0:0] mux_1482_nl;
  wire[0:0] nor_1216_nl;
  wire[0:0] nor_1217_nl;
  wire[0:0] or_1213_nl;
  wire[0:0] mux_1481_nl;
  wire[0:0] nor_1218_nl;
  wire[0:0] mux_1480_nl;
  wire[0:0] nor_1219_nl;
  wire[0:0] nor_1220_nl;
  wire[0:0] mux_1479_nl;
  wire[0:0] mux_1478_nl;
  wire[0:0] nor_1221_nl;
  wire[0:0] nor_1222_nl;
  wire[0:0] nor_1223_nl;
  wire[0:0] mux_1476_nl;
  wire[0:0] mux_1475_nl;
  wire[0:0] mux_1474_nl;
  wire[0:0] mux_1473_nl;
  wire[0:0] and_604_nl;
  wire[0:0] mux_1472_nl;
  wire[0:0] nor_1224_nl;
  wire[0:0] nor_1225_nl;
  wire[0:0] and_605_nl;
  wire[0:0] mux_1471_nl;
  wire[0:0] nor_1226_nl;
  wire[0:0] nor_1227_nl;
  wire[0:0] mux_1470_nl;
  wire[0:0] nor_1228_nl;
  wire[0:0] nor_1229_nl;
  wire[0:0] mux_1468_nl;
  wire[0:0] nor_1230_nl;
  wire[0:0] mux_1467_nl;
  wire[0:0] nor_1231_nl;
  wire[0:0] nor_1232_nl;
  wire[0:0] mux_1466_nl;
  wire[0:0] mux_1465_nl;
  wire[0:0] nor_1233_nl;
  wire[0:0] nor_1234_nl;
  wire[0:0] mux_1464_nl;
  wire[0:0] mux_1463_nl;
  wire[0:0] mux_1462_nl;
  wire[0:0] nor_1235_nl;
  wire[0:0] mux_1461_nl;
  wire[0:0] nor_1236_nl;
  wire[0:0] nor_1237_nl;
  wire[0:0] nor_1238_nl;
  wire[0:0] mux_1460_nl;
  wire[0:0] nor_1239_nl;
  wire[0:0] nor_1240_nl;
  wire[0:0] mux_1522_nl;
  wire[0:0] mux_1521_nl;
  wire[0:0] mux_1520_nl;
  wire[0:0] nor_1195_nl;
  wire[0:0] mux_1519_nl;
  wire[0:0] mux_1518_nl;
  wire[0:0] or_1281_nl;
  wire[0:0] nand_402_nl;
  wire[0:0] or_1278_nl;
  wire[0:0] nor_1196_nl;
  wire[0:0] mux_1517_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] mux_1516_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] mux_1515_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] nor_1200_nl;
  wire[0:0] mux_1514_nl;
  wire[0:0] and_602_nl;
  wire[0:0] mux_1513_nl;
  wire[0:0] nand_313_nl;
  wire[0:0] mux_1512_nl;
  wire[0:0] or_1268_nl;
  wire[0:0] mux_1511_nl;
  wire[0:0] nor_1201_nl;
  wire[0:0] mux_1510_nl;
  wire[0:0] or_1265_nl;
  wire[0:0] mux_1509_nl;
  wire[0:0] or_1263_nl;
  wire[0:0] nor_1202_nl;
  wire[0:0] mux_1508_nl;
  wire[0:0] mux_1507_nl;
  wire[0:0] mux_1506_nl;
  wire[0:0] nor_1203_nl;
  wire[0:0] mux_1505_nl;
  wire[0:0] or_1259_nl;
  wire[0:0] or_1257_nl;
  wire[0:0] nor_1204_nl;
  wire[0:0] mux_1504_nl;
  wire[0:0] mux_1503_nl;
  wire[0:0] or_1251_nl;
  wire[0:0] nor_1205_nl;
  wire[0:0] mux_1502_nl;
  wire[0:0] mux_1501_nl;
  wire[0:0] or_1247_nl;
  wire[0:0] or_1245_nl;
  wire[0:0] mux_1499_nl;
  wire[0:0] nor_1206_nl;
  wire[0:0] mux_1498_nl;
  wire[0:0] mux_1497_nl;
  wire[0:0] or_1240_nl;
  wire[0:0] or_1238_nl;
  wire[0:0] mux_1496_nl;
  wire[0:0] or_1237_nl;
  wire[0:0] or_1236_nl;
  wire[0:0] mux_1495_nl;
  wire[0:0] nor_1207_nl;
  wire[0:0] mux_1494_nl;
  wire[0:0] nor_1208_nl;
  wire[0:0] nor_1209_nl;
  wire[0:0] mux_1493_nl;
  wire[0:0] or_1231_nl;
  wire[0:0] or_1229_nl;
  wire[0:0] mux_1555_nl;
  wire[0:0] and_599_nl;
  wire[0:0] mux_1554_nl;
  wire[0:0] nor_1164_nl;
  wire[0:0] mux_1553_nl;
  wire[0:0] or_1337_nl;
  wire[0:0] or_1336_nl;
  wire[0:0] mux_1552_nl;
  wire[0:0] nor_1165_nl;
  wire[0:0] mux_1551_nl;
  wire[0:0] nor_1166_nl;
  wire[0:0] nor_1167_nl;
  wire[0:0] mux_1550_nl;
  wire[0:0] mux_1549_nl;
  wire[0:0] mux_1548_nl;
  wire[0:0] nor_1168_nl;
  wire[0:0] mux_1547_nl;
  wire[0:0] mux_1546_nl;
  wire[0:0] nor_1170_nl;
  wire[0:0] nor_1171_nl;
  wire[0:0] or_1323_nl;
  wire[0:0] mux_1545_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] mux_1544_nl;
  wire[0:0] nor_1173_nl;
  wire[0:0] nor_1174_nl;
  wire[0:0] mux_1543_nl;
  wire[0:0] mux_1542_nl;
  wire[0:0] nor_1175_nl;
  wire[0:0] nor_1176_nl;
  wire[0:0] nor_1177_nl;
  wire[0:0] mux_1540_nl;
  wire[0:0] mux_1539_nl;
  wire[0:0] mux_1538_nl;
  wire[0:0] mux_1537_nl;
  wire[0:0] and_600_nl;
  wire[0:0] mux_1536_nl;
  wire[0:0] nor_1178_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] and_601_nl;
  wire[0:0] mux_1535_nl;
  wire[0:0] nor_1180_nl;
  wire[0:0] nor_1181_nl;
  wire[0:0] mux_1534_nl;
  wire[0:0] nor_1182_nl;
  wire[0:0] nor_1183_nl;
  wire[0:0] mux_1532_nl;
  wire[0:0] nor_1184_nl;
  wire[0:0] mux_1531_nl;
  wire[0:0] nor_1185_nl;
  wire[0:0] nor_1186_nl;
  wire[0:0] mux_1530_nl;
  wire[0:0] mux_1529_nl;
  wire[0:0] nor_1187_nl;
  wire[0:0] nor_1188_nl;
  wire[0:0] mux_1528_nl;
  wire[0:0] mux_1527_nl;
  wire[0:0] mux_1526_nl;
  wire[0:0] nor_1189_nl;
  wire[0:0] mux_1525_nl;
  wire[0:0] nor_1190_nl;
  wire[0:0] nor_1191_nl;
  wire[0:0] nor_1192_nl;
  wire[0:0] mux_1524_nl;
  wire[0:0] nor_1193_nl;
  wire[0:0] nor_1194_nl;
  wire[0:0] mux_1586_nl;
  wire[0:0] mux_1585_nl;
  wire[0:0] mux_1584_nl;
  wire[0:0] nor_1149_nl;
  wire[0:0] mux_1583_nl;
  wire[0:0] mux_1582_nl;
  wire[0:0] nand_302_nl;
  wire[0:0] nand_401_nl;
  wire[0:0] or_1388_nl;
  wire[0:0] nor_1150_nl;
  wire[0:0] mux_1581_nl;
  wire[0:0] and_762_nl;
  wire[0:0] mux_1580_nl;
  wire[0:0] nor_1152_nl;
  wire[0:0] mux_1579_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] nor_1154_nl;
  wire[0:0] mux_1578_nl;
  wire[0:0] and_598_nl;
  wire[0:0] mux_1577_nl;
  wire[0:0] nand_305_nl;
  wire[0:0] mux_1576_nl;
  wire[0:0] or_1378_nl;
  wire[0:0] mux_1575_nl;
  wire[0:0] nor_1155_nl;
  wire[0:0] mux_1574_nl;
  wire[0:0] or_1375_nl;
  wire[0:0] mux_1573_nl;
  wire[0:0] nand_400_nl;
  wire[0:0] nor_1156_nl;
  wire[0:0] mux_1572_nl;
  wire[0:0] mux_1571_nl;
  wire[0:0] mux_1570_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] mux_1569_nl;
  wire[0:0] or_1369_nl;
  wire[0:0] or_1367_nl;
  wire[0:0] nor_1158_nl;
  wire[0:0] mux_1568_nl;
  wire[0:0] mux_1567_nl;
  wire[0:0] or_1361_nl;
  wire[0:0] nor_1159_nl;
  wire[0:0] mux_1566_nl;
  wire[0:0] mux_1565_nl;
  wire[0:0] or_1357_nl;
  wire[0:0] or_1355_nl;
  wire[0:0] mux_1563_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] mux_1562_nl;
  wire[0:0] mux_1561_nl;
  wire[0:0] or_1350_nl;
  wire[0:0] or_1348_nl;
  wire[0:0] mux_1560_nl;
  wire[0:0] nand_310_nl;
  wire[0:0] or_1346_nl;
  wire[0:0] mux_1559_nl;
  wire[0:0] nor_1161_nl;
  wire[0:0] mux_1558_nl;
  wire[0:0] and_763_nl;
  wire[0:0] nor_1163_nl;
  wire[0:0] mux_1557_nl;
  wire[0:0] or_1341_nl;
  wire[0:0] or_1339_nl;
  wire[0:0] mux_1619_nl;
  wire[0:0] and_593_nl;
  wire[0:0] mux_1618_nl;
  wire[0:0] nor_1120_nl;
  wire[0:0] mux_1617_nl;
  wire[0:0] or_1447_nl;
  wire[0:0] or_1446_nl;
  wire[0:0] mux_1616_nl;
  wire[0:0] nor_1121_nl;
  wire[0:0] mux_1615_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] nor_1123_nl;
  wire[0:0] mux_1614_nl;
  wire[0:0] mux_1613_nl;
  wire[0:0] mux_1612_nl;
  wire[0:0] nor_1124_nl;
  wire[0:0] mux_1611_nl;
  wire[0:0] mux_1610_nl;
  wire[0:0] nor_1126_nl;
  wire[0:0] nor_1127_nl;
  wire[0:0] nand_295_nl;
  wire[0:0] mux_1609_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] mux_1608_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] nor_1130_nl;
  wire[0:0] mux_1607_nl;
  wire[0:0] mux_1606_nl;
  wire[0:0] nor_1131_nl;
  wire[0:0] nor_1132_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] mux_1604_nl;
  wire[0:0] mux_1603_nl;
  wire[0:0] mux_1602_nl;
  wire[0:0] mux_1601_nl;
  wire[0:0] and_594_nl;
  wire[0:0] mux_1600_nl;
  wire[0:0] nor_1134_nl;
  wire[0:0] nor_1135_nl;
  wire[0:0] and_595_nl;
  wire[0:0] mux_1599_nl;
  wire[0:0] nor_1136_nl;
  wire[0:0] nor_1137_nl;
  wire[0:0] mux_1598_nl;
  wire[0:0] nor_1138_nl;
  wire[0:0] nor_1139_nl;
  wire[0:0] mux_1596_nl;
  wire[0:0] nor_1140_nl;
  wire[0:0] mux_1595_nl;
  wire[0:0] nor_1141_nl;
  wire[0:0] and_596_nl;
  wire[0:0] mux_1594_nl;
  wire[0:0] mux_1593_nl;
  wire[0:0] nor_1142_nl;
  wire[0:0] nor_1143_nl;
  wire[0:0] mux_1592_nl;
  wire[0:0] mux_1591_nl;
  wire[0:0] mux_1590_nl;
  wire[0:0] nor_1144_nl;
  wire[0:0] mux_1589_nl;
  wire[0:0] nor_1145_nl;
  wire[0:0] nor_1146_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] mux_1588_nl;
  wire[0:0] and_597_nl;
  wire[0:0] nor_1148_nl;
  wire[0:0] mux_1650_nl;
  wire[0:0] mux_1649_nl;
  wire[0:0] mux_1648_nl;
  wire[0:0] nor_1105_nl;
  wire[0:0] mux_1647_nl;
  wire[0:0] mux_1646_nl;
  wire[0:0] or_1502_nl;
  wire[0:0] or_1501_nl;
  wire[0:0] or_1499_nl;
  wire[0:0] nor_1106_nl;
  wire[0:0] mux_1645_nl;
  wire[0:0] nor_1107_nl;
  wire[0:0] mux_1644_nl;
  wire[0:0] nor_1108_nl;
  wire[0:0] mux_1643_nl;
  wire[0:0] nor_1109_nl;
  wire[0:0] nor_1110_nl;
  wire[0:0] mux_1642_nl;
  wire[0:0] and_592_nl;
  wire[0:0] mux_1641_nl;
  wire[0:0] or_1490_nl;
  wire[0:0] mux_1640_nl;
  wire[0:0] or_1489_nl;
  wire[0:0] mux_1639_nl;
  wire[0:0] nor_1111_nl;
  wire[0:0] mux_1638_nl;
  wire[0:0] or_1486_nl;
  wire[0:0] mux_1637_nl;
  wire[0:0] or_1484_nl;
  wire[0:0] nor_1112_nl;
  wire[0:0] mux_1636_nl;
  wire[0:0] mux_1635_nl;
  wire[0:0] mux_1634_nl;
  wire[0:0] nor_1113_nl;
  wire[0:0] mux_1633_nl;
  wire[0:0] or_1480_nl;
  wire[0:0] or_1478_nl;
  wire[0:0] nor_1114_nl;
  wire[0:0] mux_1632_nl;
  wire[0:0] mux_1631_nl;
  wire[0:0] or_1474_nl;
  wire[0:0] nor_1115_nl;
  wire[0:0] mux_1630_nl;
  wire[0:0] mux_1629_nl;
  wire[0:0] or_1467_nl;
  wire[0:0] or_1465_nl;
  wire[0:0] mux_1627_nl;
  wire[0:0] nor_1116_nl;
  wire[0:0] mux_1626_nl;
  wire[0:0] mux_1625_nl;
  wire[0:0] or_1460_nl;
  wire[0:0] or_1458_nl;
  wire[0:0] mux_1624_nl;
  wire[0:0] or_1457_nl;
  wire[0:0] or_1456_nl;
  wire[0:0] mux_1623_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] mux_1622_nl;
  wire[0:0] nor_1118_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] mux_1621_nl;
  wire[0:0] or_1451_nl;
  wire[0:0] or_1449_nl;
  wire[0:0] mux_1683_nl;
  wire[0:0] and_589_nl;
  wire[0:0] mux_1682_nl;
  wire[0:0] nor_1074_nl;
  wire[0:0] mux_1681_nl;
  wire[0:0] or_1558_nl;
  wire[0:0] or_1557_nl;
  wire[0:0] mux_1680_nl;
  wire[0:0] nor_1075_nl;
  wire[0:0] mux_1679_nl;
  wire[0:0] nor_1076_nl;
  wire[0:0] nor_1077_nl;
  wire[0:0] mux_1678_nl;
  wire[0:0] mux_1677_nl;
  wire[0:0] mux_1676_nl;
  wire[0:0] nor_1078_nl;
  wire[0:0] mux_1675_nl;
  wire[0:0] mux_1674_nl;
  wire[0:0] nor_1080_nl;
  wire[0:0] nor_1081_nl;
  wire[0:0] or_1544_nl;
  wire[0:0] mux_1673_nl;
  wire[0:0] nor_1082_nl;
  wire[0:0] mux_1672_nl;
  wire[0:0] nor_1083_nl;
  wire[0:0] nor_1084_nl;
  wire[0:0] mux_1671_nl;
  wire[0:0] mux_1670_nl;
  wire[0:0] nor_1085_nl;
  wire[0:0] nor_1086_nl;
  wire[0:0] nor_1087_nl;
  wire[0:0] mux_1668_nl;
  wire[0:0] mux_1667_nl;
  wire[0:0] mux_1666_nl;
  wire[0:0] mux_1665_nl;
  wire[0:0] and_590_nl;
  wire[0:0] mux_1664_nl;
  wire[0:0] nor_1088_nl;
  wire[0:0] nor_1089_nl;
  wire[0:0] and_591_nl;
  wire[0:0] mux_1663_nl;
  wire[0:0] nor_1090_nl;
  wire[0:0] nor_1091_nl;
  wire[0:0] mux_1662_nl;
  wire[0:0] nor_1092_nl;
  wire[0:0] nor_1093_nl;
  wire[0:0] mux_1660_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] mux_1659_nl;
  wire[0:0] nor_1095_nl;
  wire[0:0] nor_1096_nl;
  wire[0:0] mux_1658_nl;
  wire[0:0] mux_1657_nl;
  wire[0:0] nor_1097_nl;
  wire[0:0] nor_1098_nl;
  wire[0:0] mux_1656_nl;
  wire[0:0] mux_1655_nl;
  wire[0:0] mux_1654_nl;
  wire[0:0] nor_1099_nl;
  wire[0:0] mux_1653_nl;
  wire[0:0] nor_1100_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] nor_1102_nl;
  wire[0:0] mux_1652_nl;
  wire[0:0] nor_1103_nl;
  wire[0:0] nor_1104_nl;
  wire[0:0] mux_1714_nl;
  wire[0:0] mux_1713_nl;
  wire[0:0] mux_1712_nl;
  wire[0:0] nor_1059_nl;
  wire[0:0] mux_1711_nl;
  wire[0:0] mux_1710_nl;
  wire[0:0] or_1613_nl;
  wire[0:0] or_1612_nl;
  wire[0:0] or_1610_nl;
  wire[0:0] nor_1060_nl;
  wire[0:0] mux_1709_nl;
  wire[0:0] nor_1061_nl;
  wire[0:0] mux_1708_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] mux_1707_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] mux_1706_nl;
  wire[0:0] and_588_nl;
  wire[0:0] mux_1705_nl;
  wire[0:0] nand_287_nl;
  wire[0:0] mux_1704_nl;
  wire[0:0] or_1600_nl;
  wire[0:0] mux_1703_nl;
  wire[0:0] nor_1065_nl;
  wire[0:0] mux_1702_nl;
  wire[0:0] or_1597_nl;
  wire[0:0] mux_1701_nl;
  wire[0:0] or_1595_nl;
  wire[0:0] nor_1066_nl;
  wire[0:0] mux_1700_nl;
  wire[0:0] mux_1699_nl;
  wire[0:0] mux_1698_nl;
  wire[0:0] nor_1067_nl;
  wire[0:0] mux_1697_nl;
  wire[0:0] or_1591_nl;
  wire[0:0] or_1589_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] mux_1696_nl;
  wire[0:0] mux_1695_nl;
  wire[0:0] or_1585_nl;
  wire[0:0] nor_1069_nl;
  wire[0:0] mux_1694_nl;
  wire[0:0] mux_1693_nl;
  wire[0:0] or_1578_nl;
  wire[0:0] or_1576_nl;
  wire[0:0] mux_1691_nl;
  wire[0:0] nor_1070_nl;
  wire[0:0] mux_1690_nl;
  wire[0:0] mux_1689_nl;
  wire[0:0] or_1571_nl;
  wire[0:0] or_1569_nl;
  wire[0:0] mux_1688_nl;
  wire[0:0] or_1568_nl;
  wire[0:0] or_1567_nl;
  wire[0:0] mux_1687_nl;
  wire[0:0] nor_1071_nl;
  wire[0:0] mux_1686_nl;
  wire[0:0] nor_1072_nl;
  wire[0:0] nor_1073_nl;
  wire[0:0] mux_1685_nl;
  wire[0:0] or_1562_nl;
  wire[0:0] or_1560_nl;
  wire[0:0] mux_1747_nl;
  wire[0:0] and_585_nl;
  wire[0:0] mux_1746_nl;
  wire[0:0] nor_1028_nl;
  wire[0:0] mux_1745_nl;
  wire[0:0] or_1669_nl;
  wire[0:0] or_1668_nl;
  wire[0:0] mux_1744_nl;
  wire[0:0] nor_1029_nl;
  wire[0:0] mux_1743_nl;
  wire[0:0] nor_1030_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] mux_1742_nl;
  wire[0:0] mux_1741_nl;
  wire[0:0] mux_1740_nl;
  wire[0:0] nor_1032_nl;
  wire[0:0] mux_1739_nl;
  wire[0:0] mux_1738_nl;
  wire[0:0] nor_1034_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] or_1655_nl;
  wire[0:0] mux_1737_nl;
  wire[0:0] nor_1036_nl;
  wire[0:0] mux_1736_nl;
  wire[0:0] nor_1037_nl;
  wire[0:0] nor_1038_nl;
  wire[0:0] mux_1735_nl;
  wire[0:0] mux_1734_nl;
  wire[0:0] nor_1039_nl;
  wire[0:0] nor_1040_nl;
  wire[0:0] nor_1041_nl;
  wire[0:0] mux_1732_nl;
  wire[0:0] mux_1731_nl;
  wire[0:0] mux_1730_nl;
  wire[0:0] mux_1729_nl;
  wire[0:0] and_586_nl;
  wire[0:0] mux_1728_nl;
  wire[0:0] nor_1042_nl;
  wire[0:0] nor_1043_nl;
  wire[0:0] and_587_nl;
  wire[0:0] mux_1727_nl;
  wire[0:0] nor_1044_nl;
  wire[0:0] nor_1045_nl;
  wire[0:0] mux_1726_nl;
  wire[0:0] nor_1046_nl;
  wire[0:0] nor_1047_nl;
  wire[0:0] mux_1724_nl;
  wire[0:0] nor_1048_nl;
  wire[0:0] mux_1723_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] nor_1050_nl;
  wire[0:0] mux_1722_nl;
  wire[0:0] mux_1721_nl;
  wire[0:0] nor_1051_nl;
  wire[0:0] nor_1052_nl;
  wire[0:0] mux_1720_nl;
  wire[0:0] mux_1719_nl;
  wire[0:0] mux_1718_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] mux_1717_nl;
  wire[0:0] nor_1054_nl;
  wire[0:0] nor_1055_nl;
  wire[0:0] nor_1056_nl;
  wire[0:0] mux_1716_nl;
  wire[0:0] nor_1057_nl;
  wire[0:0] nor_1058_nl;
  wire[0:0] mux_1778_nl;
  wire[0:0] mux_1777_nl;
  wire[0:0] mux_1776_nl;
  wire[0:0] nor_1013_nl;
  wire[0:0] mux_1775_nl;
  wire[0:0] mux_1774_nl;
  wire[0:0] or_1723_nl;
  wire[0:0] or_1722_nl;
  wire[0:0] or_1720_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] mux_1773_nl;
  wire[0:0] nor_1015_nl;
  wire[0:0] mux_1772_nl;
  wire[0:0] nor_1016_nl;
  wire[0:0] mux_1771_nl;
  wire[0:0] nor_1017_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] mux_1770_nl;
  wire[0:0] and_584_nl;
  wire[0:0] mux_1769_nl;
  wire[0:0] nand_282_nl;
  wire[0:0] mux_1768_nl;
  wire[0:0] or_1710_nl;
  wire[0:0] mux_1767_nl;
  wire[0:0] nor_1019_nl;
  wire[0:0] mux_1766_nl;
  wire[0:0] or_1707_nl;
  wire[0:0] mux_1765_nl;
  wire[0:0] or_1705_nl;
  wire[0:0] nor_1020_nl;
  wire[0:0] mux_1764_nl;
  wire[0:0] mux_1763_nl;
  wire[0:0] mux_1762_nl;
  wire[0:0] nor_1021_nl;
  wire[0:0] mux_1761_nl;
  wire[0:0] or_1701_nl;
  wire[0:0] or_1699_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] mux_1760_nl;
  wire[0:0] mux_1759_nl;
  wire[0:0] or_1693_nl;
  wire[0:0] nor_1023_nl;
  wire[0:0] mux_1758_nl;
  wire[0:0] mux_1757_nl;
  wire[0:0] or_1689_nl;
  wire[0:0] or_1687_nl;
  wire[0:0] mux_1755_nl;
  wire[0:0] nor_1024_nl;
  wire[0:0] mux_1754_nl;
  wire[0:0] mux_1753_nl;
  wire[0:0] or_1682_nl;
  wire[0:0] or_1680_nl;
  wire[0:0] mux_1752_nl;
  wire[0:0] or_1679_nl;
  wire[0:0] or_1678_nl;
  wire[0:0] mux_1751_nl;
  wire[0:0] nor_1025_nl;
  wire[0:0] mux_1750_nl;
  wire[0:0] and_761_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] mux_1749_nl;
  wire[0:0] or_1673_nl;
  wire[0:0] or_1671_nl;
  wire[0:0] mux_1811_nl;
  wire[0:0] and_581_nl;
  wire[0:0] mux_1810_nl;
  wire[0:0] nor_982_nl;
  wire[0:0] mux_1809_nl;
  wire[0:0] or_1779_nl;
  wire[0:0] or_1778_nl;
  wire[0:0] mux_1808_nl;
  wire[0:0] nor_983_nl;
  wire[0:0] mux_1807_nl;
  wire[0:0] nor_984_nl;
  wire[0:0] nor_985_nl;
  wire[0:0] mux_1806_nl;
  wire[0:0] mux_1805_nl;
  wire[0:0] mux_1804_nl;
  wire[0:0] nor_986_nl;
  wire[0:0] mux_1803_nl;
  wire[0:0] mux_1802_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] nor_989_nl;
  wire[0:0] or_1765_nl;
  wire[0:0] mux_1801_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] mux_1800_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] mux_1799_nl;
  wire[0:0] mux_1798_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] nor_994_nl;
  wire[0:0] nor_995_nl;
  wire[0:0] mux_1796_nl;
  wire[0:0] mux_1795_nl;
  wire[0:0] mux_1794_nl;
  wire[0:0] mux_1793_nl;
  wire[0:0] and_582_nl;
  wire[0:0] mux_1792_nl;
  wire[0:0] nor_996_nl;
  wire[0:0] nor_997_nl;
  wire[0:0] and_583_nl;
  wire[0:0] mux_1791_nl;
  wire[0:0] nor_998_nl;
  wire[0:0] nor_999_nl;
  wire[0:0] mux_1790_nl;
  wire[0:0] nor_1000_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] mux_1788_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] mux_1787_nl;
  wire[0:0] nor_1003_nl;
  wire[0:0] nor_1004_nl;
  wire[0:0] mux_1786_nl;
  wire[0:0] mux_1785_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] mux_1784_nl;
  wire[0:0] mux_1783_nl;
  wire[0:0] mux_1782_nl;
  wire[0:0] nor_1007_nl;
  wire[0:0] mux_1781_nl;
  wire[0:0] nor_1008_nl;
  wire[0:0] nor_1009_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] mux_1780_nl;
  wire[0:0] nor_1011_nl;
  wire[0:0] nor_1012_nl;
  wire[0:0] mux_1842_nl;
  wire[0:0] mux_1841_nl;
  wire[0:0] mux_1840_nl;
  wire[0:0] nor_967_nl;
  wire[0:0] mux_1839_nl;
  wire[0:0] mux_1838_nl;
  wire[0:0] nand_272_nl;
  wire[0:0] or_1832_nl;
  wire[0:0] or_1830_nl;
  wire[0:0] nor_968_nl;
  wire[0:0] mux_1837_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] mux_1836_nl;
  wire[0:0] nor_970_nl;
  wire[0:0] mux_1835_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] nor_972_nl;
  wire[0:0] mux_1834_nl;
  wire[0:0] and_580_nl;
  wire[0:0] mux_1833_nl;
  wire[0:0] nand_274_nl;
  wire[0:0] mux_1832_nl;
  wire[0:0] or_1820_nl;
  wire[0:0] mux_1831_nl;
  wire[0:0] nor_973_nl;
  wire[0:0] mux_1830_nl;
  wire[0:0] nand_398_nl;
  wire[0:0] mux_1829_nl;
  wire[0:0] or_1815_nl;
  wire[0:0] nor_974_nl;
  wire[0:0] mux_1828_nl;
  wire[0:0] mux_1827_nl;
  wire[0:0] mux_1826_nl;
  wire[0:0] nor_975_nl;
  wire[0:0] mux_1825_nl;
  wire[0:0] or_1811_nl;
  wire[0:0] or_1809_nl;
  wire[0:0] nor_976_nl;
  wire[0:0] mux_1824_nl;
  wire[0:0] mux_1823_nl;
  wire[0:0] or_1803_nl;
  wire[0:0] nor_977_nl;
  wire[0:0] mux_1822_nl;
  wire[0:0] mux_1821_nl;
  wire[0:0] or_1799_nl;
  wire[0:0] or_1797_nl;
  wire[0:0] mux_1819_nl;
  wire[0:0] nor_978_nl;
  wire[0:0] mux_1818_nl;
  wire[0:0] mux_1817_nl;
  wire[0:0] or_1792_nl;
  wire[0:0] or_1790_nl;
  wire[0:0] mux_1816_nl;
  wire[0:0] nand_277_nl;
  wire[0:0] or_1788_nl;
  wire[0:0] mux_1815_nl;
  wire[0:0] nor_979_nl;
  wire[0:0] mux_1814_nl;
  wire[0:0] nor_980_nl;
  wire[0:0] nor_981_nl;
  wire[0:0] mux_1813_nl;
  wire[0:0] or_1783_nl;
  wire[0:0] or_1781_nl;
  wire[0:0] mux_1875_nl;
  wire[0:0] and_575_nl;
  wire[0:0] mux_1874_nl;
  wire[0:0] nor_938_nl;
  wire[0:0] mux_1873_nl;
  wire[0:0] or_1889_nl;
  wire[0:0] or_1888_nl;
  wire[0:0] mux_1872_nl;
  wire[0:0] nor_939_nl;
  wire[0:0] mux_1871_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] nor_941_nl;
  wire[0:0] mux_1870_nl;
  wire[0:0] mux_1869_nl;
  wire[0:0] mux_1868_nl;
  wire[0:0] nor_942_nl;
  wire[0:0] mux_1867_nl;
  wire[0:0] mux_1866_nl;
  wire[0:0] nor_944_nl;
  wire[0:0] nor_945_nl;
  wire[0:0] nand_265_nl;
  wire[0:0] mux_1865_nl;
  wire[0:0] nor_946_nl;
  wire[0:0] mux_1864_nl;
  wire[0:0] nor_947_nl;
  wire[0:0] nor_948_nl;
  wire[0:0] mux_1863_nl;
  wire[0:0] mux_1862_nl;
  wire[0:0] nor_949_nl;
  wire[0:0] nor_950_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] mux_1860_nl;
  wire[0:0] mux_1859_nl;
  wire[0:0] mux_1858_nl;
  wire[0:0] mux_1857_nl;
  wire[0:0] and_576_nl;
  wire[0:0] mux_1856_nl;
  wire[0:0] nor_952_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] and_577_nl;
  wire[0:0] mux_1855_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] nor_955_nl;
  wire[0:0] mux_1854_nl;
  wire[0:0] nor_956_nl;
  wire[0:0] nor_957_nl;
  wire[0:0] mux_1852_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] mux_1851_nl;
  wire[0:0] nor_959_nl;
  wire[0:0] and_578_nl;
  wire[0:0] mux_1850_nl;
  wire[0:0] mux_1849_nl;
  wire[0:0] nor_960_nl;
  wire[0:0] nor_961_nl;
  wire[0:0] mux_1848_nl;
  wire[0:0] mux_1847_nl;
  wire[0:0] mux_1846_nl;
  wire[0:0] nor_962_nl;
  wire[0:0] mux_1845_nl;
  wire[0:0] nor_963_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] nor_965_nl;
  wire[0:0] mux_1844_nl;
  wire[0:0] and_579_nl;
  wire[0:0] nor_966_nl;
  wire[0:0] mux_1906_nl;
  wire[0:0] mux_1905_nl;
  wire[0:0] mux_1904_nl;
  wire[0:0] nor_923_nl;
  wire[0:0] mux_1903_nl;
  wire[0:0] mux_1902_nl;
  wire[0:0] or_1944_nl;
  wire[0:0] or_1943_nl;
  wire[0:0] or_1941_nl;
  wire[0:0] nor_924_nl;
  wire[0:0] mux_1901_nl;
  wire[0:0] nor_925_nl;
  wire[0:0] mux_1900_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] mux_1899_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] nor_928_nl;
  wire[0:0] mux_1898_nl;
  wire[0:0] and_574_nl;
  wire[0:0] mux_1897_nl;
  wire[0:0] nand_261_nl;
  wire[0:0] mux_1896_nl;
  wire[0:0] or_1931_nl;
  wire[0:0] mux_1895_nl;
  wire[0:0] nor_929_nl;
  wire[0:0] mux_1894_nl;
  wire[0:0] or_1928_nl;
  wire[0:0] mux_1893_nl;
  wire[0:0] or_1926_nl;
  wire[0:0] nor_930_nl;
  wire[0:0] mux_1892_nl;
  wire[0:0] mux_1891_nl;
  wire[0:0] mux_1890_nl;
  wire[0:0] nor_931_nl;
  wire[0:0] mux_1889_nl;
  wire[0:0] or_1922_nl;
  wire[0:0] or_1920_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] mux_1888_nl;
  wire[0:0] mux_1887_nl;
  wire[0:0] or_1916_nl;
  wire[0:0] nor_933_nl;
  wire[0:0] mux_1886_nl;
  wire[0:0] mux_1885_nl;
  wire[0:0] or_1909_nl;
  wire[0:0] or_1907_nl;
  wire[0:0] mux_1883_nl;
  wire[0:0] nor_934_nl;
  wire[0:0] mux_1882_nl;
  wire[0:0] mux_1881_nl;
  wire[0:0] or_1902_nl;
  wire[0:0] or_1900_nl;
  wire[0:0] mux_1880_nl;
  wire[0:0] or_1899_nl;
  wire[0:0] or_1898_nl;
  wire[0:0] mux_1879_nl;
  wire[0:0] nor_935_nl;
  wire[0:0] mux_1878_nl;
  wire[0:0] nor_936_nl;
  wire[0:0] nor_937_nl;
  wire[0:0] mux_1877_nl;
  wire[0:0] or_1893_nl;
  wire[0:0] or_1891_nl;
  wire[0:0] mux_1939_nl;
  wire[0:0] and_571_nl;
  wire[0:0] mux_1938_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] mux_1937_nl;
  wire[0:0] or_2000_nl;
  wire[0:0] or_1999_nl;
  wire[0:0] mux_1936_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] mux_1935_nl;
  wire[0:0] nor_894_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] mux_1934_nl;
  wire[0:0] mux_1933_nl;
  wire[0:0] mux_1932_nl;
  wire[0:0] nor_896_nl;
  wire[0:0] mux_1931_nl;
  wire[0:0] mux_1930_nl;
  wire[0:0] nor_898_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] or_1986_nl;
  wire[0:0] mux_1929_nl;
  wire[0:0] nor_900_nl;
  wire[0:0] mux_1928_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] mux_1927_nl;
  wire[0:0] mux_1926_nl;
  wire[0:0] nor_903_nl;
  wire[0:0] nor_904_nl;
  wire[0:0] nor_905_nl;
  wire[0:0] mux_1924_nl;
  wire[0:0] mux_1923_nl;
  wire[0:0] mux_1922_nl;
  wire[0:0] mux_1921_nl;
  wire[0:0] and_572_nl;
  wire[0:0] mux_1920_nl;
  wire[0:0] nor_906_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] and_573_nl;
  wire[0:0] mux_1919_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] mux_1918_nl;
  wire[0:0] nor_910_nl;
  wire[0:0] nor_911_nl;
  wire[0:0] mux_1916_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] mux_1915_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] nor_914_nl;
  wire[0:0] mux_1914_nl;
  wire[0:0] mux_1913_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] mux_1912_nl;
  wire[0:0] mux_1911_nl;
  wire[0:0] mux_1910_nl;
  wire[0:0] nor_917_nl;
  wire[0:0] mux_1909_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] mux_1908_nl;
  wire[0:0] nor_921_nl;
  wire[0:0] nor_922_nl;
  wire[0:0] mux_1970_nl;
  wire[0:0] mux_1969_nl;
  wire[0:0] mux_1968_nl;
  wire[0:0] nor_877_nl;
  wire[0:0] mux_1967_nl;
  wire[0:0] mux_1966_nl;
  wire[0:0] nand_250_nl;
  wire[0:0] or_2054_nl;
  wire[0:0] or_2052_nl;
  wire[0:0] nor_878_nl;
  wire[0:0] mux_1965_nl;
  wire[0:0] nor_879_nl;
  wire[0:0] mux_1964_nl;
  wire[0:0] nor_880_nl;
  wire[0:0] mux_1963_nl;
  wire[0:0] nor_881_nl;
  wire[0:0] nor_882_nl;
  wire[0:0] mux_1962_nl;
  wire[0:0] and_570_nl;
  wire[0:0] mux_1961_nl;
  wire[0:0] nand_252_nl;
  wire[0:0] mux_1960_nl;
  wire[0:0] or_2042_nl;
  wire[0:0] mux_1959_nl;
  wire[0:0] nor_883_nl;
  wire[0:0] mux_1958_nl;
  wire[0:0] nand_397_nl;
  wire[0:0] mux_1957_nl;
  wire[0:0] or_2037_nl;
  wire[0:0] nor_884_nl;
  wire[0:0] mux_1956_nl;
  wire[0:0] mux_1955_nl;
  wire[0:0] mux_1954_nl;
  wire[0:0] nor_885_nl;
  wire[0:0] mux_1953_nl;
  wire[0:0] or_2033_nl;
  wire[0:0] or_2031_nl;
  wire[0:0] nor_886_nl;
  wire[0:0] mux_1952_nl;
  wire[0:0] mux_1951_nl;
  wire[0:0] or_2027_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] mux_1950_nl;
  wire[0:0] mux_1949_nl;
  wire[0:0] or_2020_nl;
  wire[0:0] or_2018_nl;
  wire[0:0] mux_1947_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_1946_nl;
  wire[0:0] mux_1945_nl;
  wire[0:0] or_2013_nl;
  wire[0:0] or_2011_nl;
  wire[0:0] mux_1944_nl;
  wire[0:0] nand_255_nl;
  wire[0:0] or_2009_nl;
  wire[0:0] mux_1943_nl;
  wire[0:0] nor_889_nl;
  wire[0:0] mux_1942_nl;
  wire[0:0] nor_890_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] mux_1941_nl;
  wire[0:0] or_2004_nl;
  wire[0:0] or_2002_nl;
  wire[0:0] mux_2003_nl;
  wire[0:0] and_565_nl;
  wire[0:0] mux_2002_nl;
  wire[0:0] nor_848_nl;
  wire[0:0] mux_2001_nl;
  wire[0:0] or_2111_nl;
  wire[0:0] or_2110_nl;
  wire[0:0] mux_2000_nl;
  wire[0:0] nor_849_nl;
  wire[0:0] mux_1999_nl;
  wire[0:0] nor_850_nl;
  wire[0:0] nor_851_nl;
  wire[0:0] mux_1998_nl;
  wire[0:0] mux_1997_nl;
  wire[0:0] mux_1996_nl;
  wire[0:0] nor_852_nl;
  wire[0:0] mux_1995_nl;
  wire[0:0] mux_1994_nl;
  wire[0:0] nor_854_nl;
  wire[0:0] nor_855_nl;
  wire[0:0] nand_243_nl;
  wire[0:0] mux_1993_nl;
  wire[0:0] nor_856_nl;
  wire[0:0] mux_1992_nl;
  wire[0:0] nor_857_nl;
  wire[0:0] nor_858_nl;
  wire[0:0] mux_1991_nl;
  wire[0:0] mux_1990_nl;
  wire[0:0] nor_859_nl;
  wire[0:0] nor_860_nl;
  wire[0:0] nor_861_nl;
  wire[0:0] mux_1988_nl;
  wire[0:0] mux_1987_nl;
  wire[0:0] mux_1986_nl;
  wire[0:0] mux_1985_nl;
  wire[0:0] and_566_nl;
  wire[0:0] mux_1984_nl;
  wire[0:0] nor_862_nl;
  wire[0:0] nor_863_nl;
  wire[0:0] and_567_nl;
  wire[0:0] mux_1983_nl;
  wire[0:0] nor_864_nl;
  wire[0:0] nor_865_nl;
  wire[0:0] mux_1982_nl;
  wire[0:0] nor_866_nl;
  wire[0:0] nor_867_nl;
  wire[0:0] mux_1980_nl;
  wire[0:0] nor_868_nl;
  wire[0:0] mux_1979_nl;
  wire[0:0] nor_869_nl;
  wire[0:0] and_568_nl;
  wire[0:0] mux_1978_nl;
  wire[0:0] mux_1977_nl;
  wire[0:0] nor_870_nl;
  wire[0:0] nor_871_nl;
  wire[0:0] mux_1976_nl;
  wire[0:0] mux_1975_nl;
  wire[0:0] mux_1974_nl;
  wire[0:0] nor_872_nl;
  wire[0:0] mux_1973_nl;
  wire[0:0] nor_873_nl;
  wire[0:0] nor_874_nl;
  wire[0:0] nor_875_nl;
  wire[0:0] mux_1972_nl;
  wire[0:0] and_569_nl;
  wire[0:0] nor_876_nl;
  wire[0:0] mux_2034_nl;
  wire[0:0] mux_2033_nl;
  wire[0:0] mux_2032_nl;
  wire[0:0] nor_833_nl;
  wire[0:0] mux_2031_nl;
  wire[0:0] mux_2030_nl;
  wire[0:0] nand_235_nl;
  wire[0:0] or_2164_nl;
  wire[0:0] or_2162_nl;
  wire[0:0] nor_834_nl;
  wire[0:0] mux_2029_nl;
  wire[0:0] nor_835_nl;
  wire[0:0] mux_2028_nl;
  wire[0:0] nor_836_nl;
  wire[0:0] mux_2027_nl;
  wire[0:0] nor_837_nl;
  wire[0:0] nor_838_nl;
  wire[0:0] mux_2026_nl;
  wire[0:0] and_563_nl;
  wire[0:0] mux_2025_nl;
  wire[0:0] nand_236_nl;
  wire[0:0] mux_2024_nl;
  wire[0:0] or_2152_nl;
  wire[0:0] mux_2023_nl;
  wire[0:0] nor_839_nl;
  wire[0:0] mux_2022_nl;
  wire[0:0] nand_396_nl;
  wire[0:0] mux_2021_nl;
  wire[0:0] or_2147_nl;
  wire[0:0] nor_840_nl;
  wire[0:0] mux_2020_nl;
  wire[0:0] mux_2019_nl;
  wire[0:0] mux_2018_nl;
  wire[0:0] nor_841_nl;
  wire[0:0] mux_2017_nl;
  wire[0:0] or_2143_nl;
  wire[0:0] or_2141_nl;
  wire[0:0] nor_842_nl;
  wire[0:0] mux_2016_nl;
  wire[0:0] mux_2015_nl;
  wire[0:0] or_2135_nl;
  wire[0:0] nor_843_nl;
  wire[0:0] mux_2014_nl;
  wire[0:0] mux_2013_nl;
  wire[0:0] or_2131_nl;
  wire[0:0] or_2129_nl;
  wire[0:0] mux_2011_nl;
  wire[0:0] nor_844_nl;
  wire[0:0] mux_2010_nl;
  wire[0:0] mux_2009_nl;
  wire[0:0] or_2124_nl;
  wire[0:0] or_2122_nl;
  wire[0:0] mux_2008_nl;
  wire[0:0] nand_239_nl;
  wire[0:0] or_2120_nl;
  wire[0:0] mux_2007_nl;
  wire[0:0] nor_845_nl;
  wire[0:0] mux_2006_nl;
  wire[0:0] nor_846_nl;
  wire[0:0] nor_847_nl;
  wire[0:0] mux_2005_nl;
  wire[0:0] or_2115_nl;
  wire[0:0] or_2113_nl;
  wire[0:0] mux_2067_nl;
  wire[0:0] and_558_nl;
  wire[0:0] mux_2066_nl;
  wire[0:0] nor_804_nl;
  wire[0:0] mux_2065_nl;
  wire[0:0] or_2221_nl;
  wire[0:0] or_2220_nl;
  wire[0:0] mux_2064_nl;
  wire[0:0] nor_805_nl;
  wire[0:0] mux_2063_nl;
  wire[0:0] nor_806_nl;
  wire[0:0] nor_807_nl;
  wire[0:0] mux_2062_nl;
  wire[0:0] mux_2061_nl;
  wire[0:0] mux_2060_nl;
  wire[0:0] nor_808_nl;
  wire[0:0] mux_2059_nl;
  wire[0:0] mux_2058_nl;
  wire[0:0] nor_810_nl;
  wire[0:0] nor_811_nl;
  wire[0:0] nand_228_nl;
  wire[0:0] mux_2057_nl;
  wire[0:0] nor_812_nl;
  wire[0:0] mux_2056_nl;
  wire[0:0] nor_813_nl;
  wire[0:0] nor_814_nl;
  wire[0:0] mux_2055_nl;
  wire[0:0] mux_2054_nl;
  wire[0:0] nor_815_nl;
  wire[0:0] nor_816_nl;
  wire[0:0] nor_817_nl;
  wire[0:0] mux_2052_nl;
  wire[0:0] mux_2051_nl;
  wire[0:0] mux_2050_nl;
  wire[0:0] mux_2049_nl;
  wire[0:0] and_559_nl;
  wire[0:0] mux_2048_nl;
  wire[0:0] nor_818_nl;
  wire[0:0] nor_819_nl;
  wire[0:0] and_560_nl;
  wire[0:0] mux_2047_nl;
  wire[0:0] nor_820_nl;
  wire[0:0] nor_821_nl;
  wire[0:0] mux_2046_nl;
  wire[0:0] nor_822_nl;
  wire[0:0] nor_823_nl;
  wire[0:0] mux_2044_nl;
  wire[0:0] nor_824_nl;
  wire[0:0] mux_2043_nl;
  wire[0:0] nor_825_nl;
  wire[0:0] and_561_nl;
  wire[0:0] mux_2042_nl;
  wire[0:0] mux_2041_nl;
  wire[0:0] nor_826_nl;
  wire[0:0] nor_827_nl;
  wire[0:0] mux_2040_nl;
  wire[0:0] mux_2039_nl;
  wire[0:0] mux_2038_nl;
  wire[0:0] nor_828_nl;
  wire[0:0] mux_2037_nl;
  wire[0:0] nor_829_nl;
  wire[0:0] nor_830_nl;
  wire[0:0] nor_831_nl;
  wire[0:0] mux_2036_nl;
  wire[0:0] and_562_nl;
  wire[0:0] nor_832_nl;
  wire[0:0] mux_2098_nl;
  wire[0:0] mux_2097_nl;
  wire[0:0] mux_2096_nl;
  wire[0:0] nor_789_nl;
  wire[0:0] mux_2095_nl;
  wire[0:0] mux_2094_nl;
  wire[0:0] and_554_nl;
  wire[0:0] or_2271_nl;
  wire[0:0] nor_790_nl;
  wire[0:0] mux_2093_nl;
  wire[0:0] nor_791_nl;
  wire[0:0] mux_2092_nl;
  wire[0:0] nor_792_nl;
  wire[0:0] mux_2091_nl;
  wire[0:0] nor_793_nl;
  wire[0:0] nor_794_nl;
  wire[0:0] mux_2090_nl;
  wire[0:0] and_555_nl;
  wire[0:0] mux_2089_nl;
  wire[0:0] nand_215_nl;
  wire[0:0] mux_2088_nl;
  wire[0:0] or_2261_nl;
  wire[0:0] mux_2087_nl;
  wire[0:0] nor_795_nl;
  wire[0:0] mux_2086_nl;
  wire[0:0] nand_395_nl;
  wire[0:0] mux_2085_nl;
  wire[0:0] or_2256_nl;
  wire[0:0] nor_796_nl;
  wire[0:0] mux_2084_nl;
  wire[0:0] mux_2083_nl;
  wire[0:0] mux_2082_nl;
  wire[0:0] nor_797_nl;
  wire[0:0] mux_2081_nl;
  wire[0:0] or_2253_nl;
  wire[0:0] or_2251_nl;
  wire[0:0] nor_798_nl;
  wire[0:0] mux_2080_nl;
  wire[0:0] mux_2079_nl;
  wire[0:0] or_2245_nl;
  wire[0:0] nor_799_nl;
  wire[0:0] mux_2078_nl;
  wire[0:0] mux_2077_nl;
  wire[0:0] or_2241_nl;
  wire[0:0] nand_219_nl;
  wire[0:0] mux_2075_nl;
  wire[0:0] nor_800_nl;
  wire[0:0] mux_2074_nl;
  wire[0:0] mux_2073_nl;
  wire[0:0] or_2234_nl;
  wire[0:0] or_2232_nl;
  wire[0:0] mux_2072_nl;
  wire[0:0] nand_220_nl;
  wire[0:0] nand_221_nl;
  wire[0:0] mux_2071_nl;
  wire[0:0] nor_801_nl;
  wire[0:0] mux_2070_nl;
  wire[0:0] nor_802_nl;
  wire[0:0] nor_803_nl;
  wire[0:0] mux_2069_nl;
  wire[0:0] or_2225_nl;
  wire[0:0] nand_223_nl;
  wire[0:0] mux_2131_nl;
  wire[0:0] and_546_nl;
  wire[0:0] mux_2130_nl;
  wire[0:0] nor_763_nl;
  wire[0:0] mux_2129_nl;
  wire[0:0] nand_199_nl;
  wire[0:0] or_2327_nl;
  wire[0:0] mux_2128_nl;
  wire[0:0] nor_764_nl;
  wire[0:0] mux_2127_nl;
  wire[0:0] nor_765_nl;
  wire[0:0] nor_766_nl;
  wire[0:0] mux_2126_nl;
  wire[0:0] mux_2125_nl;
  wire[0:0] mux_2124_nl;
  wire[0:0] nor_767_nl;
  wire[0:0] mux_2123_nl;
  wire[0:0] mux_2122_nl;
  wire[0:0] nor_769_nl;
  wire[0:0] nor_770_nl;
  wire[0:0] nand_203_nl;
  wire[0:0] mux_2121_nl;
  wire[0:0] nor_771_nl;
  wire[0:0] mux_2120_nl;
  wire[0:0] and_547_nl;
  wire[0:0] nor_772_nl;
  wire[0:0] mux_2119_nl;
  wire[0:0] mux_2118_nl;
  wire[0:0] nor_773_nl;
  wire[0:0] nor_774_nl;
  wire[0:0] nor_775_nl;
  wire[0:0] mux_2116_nl;
  wire[0:0] mux_2115_nl;
  wire[0:0] mux_2114_nl;
  wire[0:0] mux_2113_nl;
  wire[0:0] and_548_nl;
  wire[0:0] mux_2112_nl;
  wire[0:0] nor_776_nl;
  wire[0:0] nor_777_nl;
  wire[0:0] and_549_nl;
  wire[0:0] mux_2111_nl;
  wire[0:0] nor_778_nl;
  wire[0:0] and_759_nl;
  wire[0:0] mux_2110_nl;
  wire[0:0] nor_780_nl;
  wire[0:0] nor_781_nl;
  wire[0:0] mux_2108_nl;
  wire[0:0] nor_782_nl;
  wire[0:0] mux_2107_nl;
  wire[0:0] and_550_nl;
  wire[0:0] and_551_nl;
  wire[0:0] mux_2106_nl;
  wire[0:0] mux_2105_nl;
  wire[0:0] nor_783_nl;
  wire[0:0] nor_784_nl;
  wire[0:0] mux_2104_nl;
  wire[0:0] mux_2103_nl;
  wire[0:0] mux_2102_nl;
  wire[0:0] nor_785_nl;
  wire[0:0] mux_2101_nl;
  wire[0:0] nor_786_nl;
  wire[0:0] nor_787_nl;
  wire[0:0] and_552_nl;
  wire[0:0] mux_2100_nl;
  wire[0:0] and_553_nl;
  wire[0:0] nor_788_nl;
  wire[0:0] mux_3811_nl;
  wire[0:0] nor_1648_nl;
  wire[0:0] mux_3810_nl;
  wire[0:0] mux_3809_nl;
  wire[0:0] or_3467_nl;
  wire[0:0] or_3466_nl;
  wire[0:0] or_3465_nl;
  wire[0:0] mux_3808_nl;
  wire[0:0] nor_1649_nl;
  wire[0:0] mux_3807_nl;
  wire[0:0] mux_3806_nl;
  wire[0:0] mux_3805_nl;
  wire[0:0] nor_1650_nl;
  wire[0:0] nor_1651_nl;
  wire[0:0] nor_1652_nl;
  wire[0:0] and_nl;
  wire[0:0] mux_3804_nl;
  wire[0:0] or_3456_nl;
  wire[0:0] mux_3803_nl;
  wire[0:0] mux_3802_nl;
  wire[0:0] and_1158_nl;
  wire[0:0] mux_3801_nl;
  wire[0:0] nor_1653_nl;
  wire[0:0] nor_1654_nl;
  wire[0:0] mux_3800_nl;
  wire[0:0] nor_1655_nl;
  wire[0:0] nor_1656_nl;
  wire[0:0] mux_3828_nl;
  wire[0:0] or_3448_nl;
  wire[0:0] mux_3821_nl;
  wire[0:0] mux_3829_nl;
  wire[0:0] or_3510_nl;
  wire[0:0] mux_3842_nl;
  wire[0:0] or_3520_nl;
  wire[0:0] or_3527_nl;
  wire[0:0] mux_3849_nl;
  wire[0:0] mux_3893_nl;
  wire[0:0] or_3564_nl;
  wire[0:0] mux_3904_nl;
  wire[0:0] or_3586_nl;
  wire[0:0] or_3585_nl;
  wire[0:0] mux_3907_nl;
  wire[0:0] or_3584_nl;
  wire[0:0] or_3583_nl;
  wire[11:0] operator_64_false_1_mux_2_nl;
  wire[9:0] operator_64_false_1_mux_3_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_72_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_73_nl;
  wire[62:0] COMP_LOOP_mux1h_575_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_and_938_nl;
  wire[0:0] COMP_LOOP_nor_695_nl;
  wire[12:0] COMP_LOOP_acc_105_nl;
  wire[13:0] nl_COMP_LOOP_acc_105_nl;
  wire[6:0] COMP_LOOP_mux1h_576_nl;
  wire[2:0] COMP_LOOP_mux1h_577_nl;
  wire[0:0] COMP_LOOP_or_69_nl;
  wire[10:0] acc_3_nl;
  wire[11:0] nl_acc_3_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_74_nl;
  wire[8:0] COMP_LOOP_COMP_LOOP_mux_18_nl;
  wire[0:0] COMP_LOOP_or_70_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_mux_19_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_75_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_76_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_78_nl;
  wire[9:0] COMP_LOOP_mux_82_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_mux_20_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_79_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_80_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_81_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_82_nl;
  wire[3:0] COMP_LOOP_or_71_nl;
  wire[3:0] COMP_LOOP_mux1h_578_nl;
  wire[0:0] and_1178_nl;
  wire[0:0] and_1179_nl;
  wire[0:0] and_1180_nl;
  wire[0:0] and_1181_nl;
  wire[0:0] and_1182_nl;
  wire[0:0] and_1183_nl;
  wire[0:0] and_1184_nl;
  wire[0:0] and_1185_nl;
  wire[65:0] acc_6_nl;
  wire[66:0] nl_acc_6_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_83_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_84_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_85_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_86_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_87_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_88_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_89_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_90_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_91_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_92_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_93_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_94_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_95_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_96_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_97_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_98_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_99_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_100_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_101_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_102_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_103_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_104_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_105_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_106_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_107_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_108_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_109_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_110_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_111_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_112_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_113_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_114_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_115_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_116_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_117_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_118_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_119_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_120_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_121_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_122_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_123_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_124_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_125_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_126_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_127_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_128_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_129_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_130_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_131_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_132_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_133_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_134_nl;
  wire[3:0] COMP_LOOP_COMP_LOOP_or_135_nl;
  wire[3:0] COMP_LOOP_and_398_nl;
  wire[3:0] COMP_LOOP_mux_83_nl;
  wire[0:0] COMP_LOOP_or_72_nl;
  wire[0:0] COMP_LOOP_or_73_nl;
  wire[0:0] COMP_LOOP_mux1h_579_nl;
  wire[6:0] COMP_LOOP_mux1h_580_nl;
  wire[0:0] COMP_LOOP_or_74_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_136_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_137_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_138_nl;
  wire[2:0] COMP_LOOP_or_75_nl;
  wire[2:0] COMP_LOOP_and_401_nl;
  wire[2:0] COMP_LOOP_COMP_LOOP_mux_21_nl;
  wire[0:0] COMP_LOOP_nor_706_nl;
  wire[1:0] COMP_LOOP_COMP_LOOP_or_139_nl;
  wire[1:0] COMP_LOOP_and_402_nl;
  wire[0:0] COMP_LOOP_nor_707_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_140_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_141_nl;
  wire[7:0] acc_7_nl;
  wire[8:0] nl_acc_7_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_142_nl;
  wire[5:0] COMP_LOOP_mux1h_581_nl;
  wire[0:0] COMP_LOOP_or_76_nl;
  wire[4:0] COMP_LOOP_COMP_LOOP_mux_22_nl;
  wire[0:0] COMP_LOOP_or_77_nl;
  wire[0:0] COMP_LOOP_COMP_LOOP_or_143_nl;
  wire[63:0] modExp_while_if_mux_1_nl;
  wire[0:0] mux_3947_nl;
  wire[0:0] mux_3948_nl;
  wire[0:0] nor_1711_nl;
  wire[0:0] mux_3949_nl;
  wire[0:0] or_3639_nl;
  wire[0:0] mux_3950_nl;
  wire[0:0] or_3640_nl;
  wire[0:0] mux_3951_nl;
  wire[0:0] and_1186_nl;
  wire[0:0] mux_3952_nl;
  wire[0:0] mux_3953_nl;
  wire[0:0] nor_1712_nl;
  wire[0:0] mux_3954_nl;
  wire[0:0] or_3641_nl;
  wire[0:0] or_3642_nl;
  wire[0:0] nor_1713_nl;
  wire[0:0] mux_3955_nl;
  wire[0:0] nand_428_nl;
  wire[0:0] or_3643_nl;
  wire[0:0] mux_3956_nl;
  wire[0:0] mux_3957_nl;
  wire[0:0] and_1187_nl;
  wire[0:0] mux_3958_nl;
  wire[0:0] and_1188_nl;
  wire[0:0] mux_3959_nl;
  wire[0:0] or_3644_nl;
  wire[0:0] nor_1714_nl;
  wire[0:0] mux_3960_nl;
  wire[0:0] or_3645_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [10:0] nl_operator_66_true_div_cmp_b;
  assign nl_operator_66_true_div_cmp_b = {1'b0, operator_66_true_div_cmp_b_9_0};
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0 = ~ (z_out_1[64]);
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0 = ~ COMP_LOOP_nor_11_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_512_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_512_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_576_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_576_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_640_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_640_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_704_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_704_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_768_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_768_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_832_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_832_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_896_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_896_tr0 = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_960_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_960_tr0 = ~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0
      = ~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm;
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0 = z_out[12];
  wire [0:0] nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0;
  assign nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0 = ~ STAGE_LOOP_acc_itm_2_1;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd64)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd64)) r_rsci (
      .dat(r_rsc_dat),
      .idat(r_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_15_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_14_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_13_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_12_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_11_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_10_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_9_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_8_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_7_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_6_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_5_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_4_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_3_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_2_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_1_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) vec_rsc_triosy_0_0_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(vec_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_vec_rsc_triosy_0_15_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_rem #(.width_a(32'sd64),
  .width_b(32'sd64),
  .signd(32'sd1)) modulo_result_rem_cmp (
      .a(modulo_result_rem_cmp_a),
      .b(modulo_result_rem_cmp_b),
      .z(modulo_result_rem_cmp_z)
    );
  mgc_div #(.width_a(32'sd65),
  .width_b(32'sd11),
  .signd(32'sd1)) operator_66_true_div_cmp (
      .a(operator_66_true_div_cmp_a),
      .b(nl_operator_66_true_div_cmp_b[10:0]),
      .z(operator_66_true_div_cmp_z)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd10)) STAGE_LOOP_lshift_rg (
      .a(1'b1),
      .s(STAGE_LOOP_i_3_0_sva),
      .z(STAGE_LOOP_lshift_psp_sva_mx0w0)
    );
  inPlaceNTT_DIT_core_core_fsm inPlaceNTT_DIT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .STAGE_LOOP_C_8_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_8_tr0[0:0]),
      .modExp_while_C_38_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_1_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_1_tr0[0:0]),
      .COMP_LOOP_1_modExp_1_while_C_38_tr0(COMP_LOOP_COMP_LOOP_and_137_itm),
      .COMP_LOOP_C_64_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_64_tr0[0:0]),
      .COMP_LOOP_2_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_2_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_128_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_128_tr0[0:0]),
      .COMP_LOOP_3_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_3_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_192_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_192_tr0[0:0]),
      .COMP_LOOP_4_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_4_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_256_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_256_tr0[0:0]),
      .COMP_LOOP_5_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_5_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_320_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_320_tr0[0:0]),
      .COMP_LOOP_6_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_6_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_384_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_384_tr0[0:0]),
      .COMP_LOOP_7_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_7_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_448_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_448_tr0[0:0]),
      .COMP_LOOP_8_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_8_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_512_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_512_tr0[0:0]),
      .COMP_LOOP_9_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_9_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_576_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_576_tr0[0:0]),
      .COMP_LOOP_10_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_10_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_640_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_640_tr0[0:0]),
      .COMP_LOOP_11_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_11_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_704_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_704_tr0[0:0]),
      .COMP_LOOP_12_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_12_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_768_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_768_tr0[0:0]),
      .COMP_LOOP_13_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_13_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_832_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_832_tr0[0:0]),
      .COMP_LOOP_14_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_14_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_896_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_896_tr0[0:0]),
      .COMP_LOOP_15_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_15_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_960_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_C_960_tr0[0:0]),
      .COMP_LOOP_16_modExp_1_while_C_38_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_COMP_LOOP_16_modExp_1_while_C_38_tr0[0:0]),
      .COMP_LOOP_C_1024_tr0(COMP_LOOP_COMP_LOOP_and_10_itm),
      .VEC_LOOP_C_0_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_VEC_LOOP_C_0_tr0[0:0]),
      .STAGE_LOOP_C_9_tr0(nl_inPlaceNTT_DIT_core_core_fsm_inst_STAGE_LOOP_C_9_tr0[0:0])
    );
  assign nor_1445_cse = ~((fsm_output[7]) | (fsm_output[3]) | (~ (fsm_output[9]))
      | (fsm_output[2]) | (fsm_output[10]));
  assign or_651_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_650_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (VEC_LOOP_j_sva_11_0[2]) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign mux_1157_cse = MUX_s_1_2_2(or_651_nl, or_650_nl, fsm_output[5]);
  assign or_638_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_637_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1149_cse = MUX_s_1_2_2(or_638_nl, or_637_nl, fsm_output[5]);
  assign nand_332_cse = ~((VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign or_859_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_858_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1277_cse = MUX_s_1_2_2(or_859_nl, or_858_nl, fsm_output[5]);
  assign nand_324_cse = ~((~ (fsm_output[1])) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign or_1093_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1092_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]);
  assign mux_1413_cse = MUX_s_1_2_2(or_1093_nl, or_1092_nl, fsm_output[5]);
  assign or_1080_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_1079_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1405_cse = MUX_s_1_2_2(or_1080_nl, or_1079_nl, fsm_output[5]);
  assign or_1301_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_1300_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1533_cse = MUX_s_1_2_2(or_1301_nl, or_1300_nl, fsm_output[5]);
  assign or_1535_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1534_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]);
  assign mux_1669_cse = MUX_s_1_2_2(or_1535_nl, or_1534_nl, fsm_output[5]);
  assign or_1522_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_1521_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1661_cse = MUX_s_1_2_2(or_1522_nl, or_1521_nl, fsm_output[5]);
  assign or_1743_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_1742_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1789_cse = MUX_s_1_2_2(or_1743_nl, or_1742_nl, fsm_output[5]);
  assign nand_259_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) & (fsm_output[7])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10])));
  assign or_1976_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]);
  assign mux_1925_cse = MUX_s_1_2_2(nand_259_nl, or_1976_nl, fsm_output[5]);
  assign or_1964_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]);
  assign or_1963_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_1917_cse = MUX_s_1_2_2(or_1964_nl, or_1963_nl, fsm_output[5]);
  assign nand_231_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (~ (fsm_output[10])));
  assign or_2184_nl = (fsm_output[7]) | (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) |
      (fsm_output[3]) | (fsm_output[9]) | not_tmp_253;
  assign mux_2045_cse = MUX_s_1_2_2(nand_231_nl, or_2184_nl, fsm_output[5]);
  assign or_3388_cse = (fsm_output[1:0]!=2'b00);
  assign and_527_cse = or_3388_cse & (fsm_output[2]);
  assign and_526_cse = (fsm_output[1:0]==2'b11);
  assign or_2377_cse = and_526_cse | (fsm_output[2]);
  assign or_2368_cse = (fsm_output[2:1]!=2'b00);
  assign and_529_cse = (fsm_output[2:1]==2'b11);
  assign nor_758_cse = ~((fsm_output[2:1]!=2'b00));
  assign nand_196_cse = ~((fsm_output[2:1]==2'b11));
  assign or_2419_cse = (~ (fsm_output[1])) | (fsm_output[9]);
  assign nor_297_cse = ~((fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[9])));
  assign nor_303_cse = ~((fsm_output[1]) | (~ (fsm_output[9])));
  assign nor_1584_nl = ~((fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6])
      | (~ (fsm_output[10])));
  assign and_739_nl = (fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]) & (~ (fsm_output[10]));
  assign mux_125_cse = MUX_s_1_2_2(nor_1584_nl, and_739_nl, fsm_output[7]);
  assign and_536_cse = (fsm_output[2:0]==3'b111);
  assign nor_753_cse = ~((fsm_output[1:0]!=2'b00));
  assign or_2387_cse = (fsm_output[10:8]!=3'b110);
  assign or_2414_cse = (fsm_output[10:9]!=2'b00);
  assign or_2407_cse = (fsm_output[10:8]!=3'b010);
  assign mux_2171_cse = MUX_s_1_2_2((fsm_output[7]), or_tmp_2276, fsm_output[9]);
  assign mux_2203_cse = MUX_s_1_2_2(or_tmp_2281, (fsm_output[7]), fsm_output[9]);
  assign or_2400_cse = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[9]);
  assign and_521_cse = (~((fsm_output[1:0]==2'b11))) & (fsm_output[9]);
  assign or_2421_cse = nor_753_cse | (fsm_output[9]);
  assign nand_356_cse = ~((fsm_output[5]) & (fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]));
  assign or_491_cse = (fsm_output[4:2]!=3'b000);
  assign nand_357_cse = ~((fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]));
  assign nand_358_cse = ~((fsm_output[10:9]==2'b11));
  assign or_2921_cse = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign or_2918_cse = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_2912_cse = (fsm_output[1]) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[6]) | (~ (fsm_output[10]));
  assign or_2905_cse = (~ (fsm_output[1])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign nor_697_cse = ~(and_526_cse | (fsm_output[2]));
  assign mux_3254_cse = MUX_s_1_2_2(or_2947_cse, or_2921_cse, fsm_output[0]);
  assign mux_3245_cse = MUX_s_1_2_2(mux_3281_cse, or_2905_cse, fsm_output[0]);
  assign or_2914_cse = (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[2]) |
      (fsm_output[6]) | (~ (fsm_output[10]));
  assign or_2920_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_3255_nl = MUX_s_1_2_2(mux_3254_cse, or_2920_nl, fsm_output[3]);
  assign nor_640_nl = ~((fsm_output[4]) | (~ (fsm_output[8])) | mux_3255_nl);
  assign mux_3252_nl = MUX_s_1_2_2(or_2918_cse, mux_3281_cse, fsm_output[0]);
  assign and_421_nl = (fsm_output[8]) & (fsm_output[3]) & (~ mux_3252_nl);
  assign nor_642_nl = ~((fsm_output[2]) | (fsm_output[6]) | (fsm_output[10]));
  assign nor_643_nl = ~((~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_3250_nl = MUX_s_1_2_2(nor_642_nl, nor_643_nl, fsm_output[9]);
  assign nand_85_nl = ~((fsm_output[1:0]==2'b11) & mux_3250_nl);
  assign mux_3249_nl = MUX_s_1_2_2(or_2914_cse, or_2912_cse, fsm_output[0]);
  assign mux_3251_nl = MUX_s_1_2_2(nand_85_nl, mux_3249_nl, fsm_output[3]);
  assign nor_641_nl = ~((fsm_output[8]) | mux_3251_nl);
  assign mux_3253_nl = MUX_s_1_2_2(and_421_nl, nor_641_nl, fsm_output[4]);
  assign mux_3256_nl = MUX_s_1_2_2(nor_640_nl, mux_3253_nl, fsm_output[5]);
  assign or_2910_nl = (~ (fsm_output[1])) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign mux_3246_nl = MUX_s_1_2_2(or_2910_nl, or_2947_cse, fsm_output[0]);
  assign and_423_nl = (fsm_output[3]) & (~ mux_3246_nl);
  assign nor_644_nl = ~((fsm_output[3]) | mux_3245_cse);
  assign mux_3247_nl = MUX_s_1_2_2(and_423_nl, nor_644_nl, fsm_output[8]);
  assign and_422_nl = (fsm_output[4]) & mux_3247_nl;
  assign nor_645_nl = ~((fsm_output[4]) | (fsm_output[8]) | (fsm_output[3]) | (~
      (fsm_output[0])) | (fsm_output[1]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[6])
      | (~ (fsm_output[10])));
  assign mux_3248_nl = MUX_s_1_2_2(and_422_nl, nor_645_nl, fsm_output[5]);
  assign mux_3257_nl = MUX_s_1_2_2(mux_3256_nl, mux_3248_nl, fsm_output[7]);
  assign and_323_nl = mux_3257_nl & COMP_LOOP_nor_11_itm;
  assign modExp_while_if_and_nl = modExp_while_and_3 & not_tmp_557;
  assign modExp_while_if_and_1_nl = modExp_while_and_5 & not_tmp_557;
  assign modExp_while_if_mux1h_nl = MUX1HOT_v_64_6_2(z_out_8, 64'b0000000000000000000000000000000000000000000000000000000000000001,
      COMP_LOOP_1_modExp_1_while_if_mul_mut_1, modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w6,
      COMP_LOOP_1_acc_5_mut_mx0w5, {and_dcpl_237 , (~ mux_2757_itm) , and_323_nl
      , modExp_while_if_and_nl , modExp_while_if_and_1_nl , not_tmp_441});
  assign and_261_nl = and_dcpl_93 & and_dcpl_127;
  assign or_2578_nl = (fsm_output[2:0]!=3'b000) | (~ nor_tmp_324);
  assign mux_2540_nl = MUX_s_1_2_2(or_2578_nl, or_2541_cse, fsm_output[9]);
  assign mux_2629_nl = MUX_s_1_2_2((~ or_tmp_2393), (fsm_output[5]), or_2368_cse);
  assign mux_2628_nl = MUX_s_1_2_2((~ or_tmp_2393), (fsm_output[5]), and_527_cse);
  assign mux_2630_nl = MUX_s_1_2_2(mux_2629_nl, mux_2628_nl, fsm_output[9]);
  assign mux_2541_nl = MUX_s_1_2_2(mux_2540_nl, mux_2630_nl, fsm_output[6]);
  assign or_2624_nl = (~(and_526_cse | (fsm_output[2]) | (fsm_output[5]))) | (fsm_output[10]);
  assign mux_2609_nl = MUX_s_1_2_2((~ or_2534_cse), or_2624_nl, fsm_output[9]);
  assign mux_2607_nl = MUX_s_1_2_2(mux_2494_cse, mux_2516_cse, and_526_cse);
  assign or_2622_nl = (~((fsm_output[2:0]!=3'b000))) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_2608_nl = MUX_s_1_2_2(mux_2607_nl, or_2622_nl, fsm_output[9]);
  assign mux_2610_nl = MUX_s_1_2_2(mux_2609_nl, mux_2608_nl, fsm_output[6]);
  assign mux_2542_nl = MUX_s_1_2_2(mux_2541_nl, mux_2610_nl, fsm_output[8]);
  assign mux_2615_nl = MUX_s_1_2_2(nor_tmp_324, mux_2486_cse, and_527_cse);
  assign mux_2616_nl = MUX_s_1_2_2((~ or_2528_cse), mux_2615_nl, fsm_output[9]);
  assign nor_696_nl = ~(nor_697_cse | (fsm_output[5]) | (fsm_output[10]));
  assign or_2627_nl = (~((~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[5])))
      | (fsm_output[10]);
  assign mux_2614_nl = MUX_s_1_2_2(nor_696_nl, or_2627_nl, fsm_output[9]);
  assign mux_2617_nl = MUX_s_1_2_2(mux_2616_nl, mux_2614_nl, fsm_output[6]);
  assign mux_2598_nl = MUX_s_1_2_2((fsm_output[5]), nor_tmp_324, and_527_cse);
  assign mux_2599_nl = MUX_s_1_2_2(mux_2598_nl, or_tmp_2474, fsm_output[9]);
  assign mux_2600_nl = MUX_s_1_2_2(mux_2599_nl, mux_2465_cse, fsm_output[6]);
  assign mux_2532_nl = MUX_s_1_2_2(mux_2617_nl, mux_2600_nl, fsm_output[8]);
  assign mux_2543_nl = MUX_s_1_2_2(mux_2542_nl, mux_2532_nl, fsm_output[7]);
  assign mux_2520_nl = MUX_s_1_2_2((fsm_output[5]), nor_tmp_324, or_2368_cse);
  assign mux_2623_nl = MUX_s_1_2_2(mux_2494_cse, mux_2515_cse, fsm_output[1]);
  assign mux_2622_nl = MUX_s_1_2_2(mux_2516_cse, mux_2515_cse, fsm_output[1]);
  assign mux_2624_nl = MUX_s_1_2_2(mux_2623_nl, mux_2622_nl, fsm_output[0]);
  assign mux_2521_nl = MUX_s_1_2_2(mux_2520_nl, mux_2624_nl, fsm_output[9]);
  assign mux_2619_nl = MUX_s_1_2_2((fsm_output[5]), nor_tmp_324, or_2377_cse);
  assign mux_2620_nl = MUX_s_1_2_2((~ nand_173_cse), mux_2619_nl, fsm_output[9]);
  assign mux_2522_nl = MUX_s_1_2_2(mux_2521_nl, mux_2620_nl, fsm_output[6]);
  assign mux_2603_nl = MUX_s_1_2_2((fsm_output[5]), or_tmp_2474, fsm_output[9]);
  assign mux_2586_nl = MUX_s_1_2_2(or_tmp_2474, (fsm_output[5]), and_529_cse);
  assign or_2620_nl = (~(nor_697_cse | (fsm_output[5]))) | (fsm_output[10]);
  assign mux_2602_nl = MUX_s_1_2_2((~ mux_2586_nl), or_2620_nl, fsm_output[9]);
  assign mux_2604_nl = MUX_s_1_2_2(mux_2603_nl, mux_2602_nl, fsm_output[6]);
  assign mux_2523_nl = MUX_s_1_2_2(mux_2522_nl, mux_2604_nl, fsm_output[8]);
  assign or_2625_nl = (fsm_output[9]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_2613_nl = MUX_s_1_2_2(mux_2465_cse, or_2625_nl, fsm_output[6]);
  assign mux_2594_nl = MUX_s_1_2_2(or_tmp_2474, nor_tmp_324, and_529_cse);
  assign mux_2595_nl = MUX_s_1_2_2(or_2528_cse, mux_2594_nl, fsm_output[0]);
  assign or_2616_nl = (~((~ (fsm_output[2])) | (fsm_output[5]))) | (fsm_output[10]);
  assign mux_2596_nl = MUX_s_1_2_2((~ mux_2595_nl), or_2616_nl, fsm_output[9]);
  assign nor_704_nl = ~((fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[10])));
  assign or_2612_nl = (~((fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[5])))
      | (fsm_output[10]);
  assign mux_2593_nl = MUX_s_1_2_2(nor_704_nl, or_2612_nl, fsm_output[9]);
  assign mux_2597_nl = MUX_s_1_2_2(mux_2596_nl, mux_2593_nl, fsm_output[6]);
  assign mux_2508_nl = MUX_s_1_2_2(mux_2613_nl, mux_2597_nl, fsm_output[8]);
  assign mux_2524_nl = MUX_s_1_2_2(mux_2523_nl, mux_2508_nl, fsm_output[7]);
  assign mux_2544_nl = MUX_s_1_2_2(mux_2543_nl, mux_2524_nl, fsm_output[4]);
  assign mux_2495_nl = MUX_s_1_2_2(or_2540_cse, mux_2494_cse, fsm_output[1]);
  assign mux_2496_nl = MUX_s_1_2_2(or_2528_cse, mux_2495_nl, fsm_output[0]);
  assign mux_2497_nl = MUX_s_1_2_2(mux_2496_nl, or_2540_cse, fsm_output[9]);
  assign mux_2498_nl = MUX_s_1_2_2(mux_2497_nl, (fsm_output[5]), fsm_output[6]);
  assign nor_707_nl = ~(nor_758_cse | (~ (fsm_output[5])) | (fsm_output[10]));
  assign or_2591_nl = (or_3388_cse & (fsm_output[2]) & (fsm_output[5])) | (fsm_output[10]);
  assign mux_2560_nl = MUX_s_1_2_2(nor_707_nl, or_2591_nl, fsm_output[9]);
  assign or_2589_nl = (~((fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[5]))))
      | (fsm_output[10]);
  assign mux_2559_nl = MUX_s_1_2_2((~ nand_386_cse), or_2589_nl, fsm_output[9]);
  assign mux_2561_nl = MUX_s_1_2_2(mux_2560_nl, mux_2559_nl, fsm_output[6]);
  assign mux_2499_nl = MUX_s_1_2_2(mux_2498_nl, mux_2561_nl, fsm_output[8]);
  assign mux_2574_nl = MUX_s_1_2_2(mux_2486_cse, or_tmp_2393, or_2377_cse);
  assign mux_2575_nl = MUX_s_1_2_2((~ (fsm_output[5])), mux_2574_nl, fsm_output[9]);
  assign mux_2570_nl = MUX_s_1_2_2(or_tmp_2474, nor_tmp_324, or_2368_cse);
  assign mux_2571_nl = MUX_s_1_2_2((~ mux_2570_nl), nand_173_cse, fsm_output[0]);
  assign or_2602_nl = (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign mux_2572_nl = MUX_s_1_2_2(mux_2571_nl, or_2602_nl, fsm_output[9]);
  assign mux_2576_nl = MUX_s_1_2_2(mux_2575_nl, mux_2572_nl, fsm_output[6]);
  assign nor_709_nl = ~(and_526_cse | (fsm_output[2]) | (~ nor_tmp_324));
  assign mux_2552_nl = MUX_s_1_2_2(nor_709_nl, (fsm_output[10]), fsm_output[9]);
  assign mux_2550_nl = MUX_s_1_2_2((fsm_output[5]), or_tmp_2394, and_529_cse);
  assign mux_2551_nl = MUX_s_1_2_2((~ mux_2550_nl), or_tmp_2393, fsm_output[9]);
  assign mux_2553_nl = MUX_s_1_2_2(mux_2552_nl, mux_2551_nl, fsm_output[6]);
  assign mux_2490_nl = MUX_s_1_2_2(mux_2576_nl, mux_2553_nl, fsm_output[8]);
  assign mux_2500_nl = MUX_s_1_2_2(mux_2499_nl, mux_2490_nl, fsm_output[7]);
  assign mux_2581_nl = MUX_s_1_2_2((~ nor_tmp_324), or_tmp_2474, fsm_output[2]);
  assign mux_2582_nl = MUX_s_1_2_2(or_2541_cse, mux_2581_nl, fsm_output[1]);
  assign mux_2580_nl = MUX_s_1_2_2(or_2541_cse, or_2540_cse, fsm_output[1]);
  assign mux_2583_nl = MUX_s_1_2_2(mux_2582_nl, mux_2580_nl, fsm_output[0]);
  assign mux_2584_nl = MUX_s_1_2_2(or_2540_cse, mux_2583_nl, fsm_output[9]);
  assign or_2608_nl = (fsm_output[2:1]!=2'b00) | (~ nor_tmp_324);
  assign or_2606_nl = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[5])
      | (fsm_output[10]);
  assign mux_2578_nl = MUX_s_1_2_2(or_2608_nl, or_2606_nl, fsm_output[0]);
  assign mux_2579_nl = MUX_s_1_2_2(or_2540_cse, mux_2578_nl, fsm_output[9]);
  assign mux_2585_nl = MUX_s_1_2_2(mux_2584_nl, mux_2579_nl, fsm_output[6]);
  assign mux_2556_nl = MUX_s_1_2_2((fsm_output[5]), nor_tmp_324, and_529_cse);
  assign mux_2557_nl = MUX_s_1_2_2(mux_2556_nl, or_tmp_2474, fsm_output[9]);
  assign mux_2558_nl = MUX_s_1_2_2(mux_2557_nl, mux_2465_cse, fsm_output[6]);
  assign mux_2477_nl = MUX_s_1_2_2((~ mux_2585_nl), mux_2558_nl, fsm_output[8]);
  assign mux_2566_nl = MUX_s_1_2_2((fsm_output[5]), or_tmp_2394, or_2368_cse);
  assign mux_2567_nl = MUX_s_1_2_2(mux_2566_nl, or_2534_cse, fsm_output[0]);
  assign or_2598_nl = (~((fsm_output[2]) | (fsm_output[5]))) | (fsm_output[10]);
  assign mux_2568_nl = MUX_s_1_2_2((~ mux_2567_nl), or_2598_nl, fsm_output[9]);
  assign mux_2564_nl = MUX_s_1_2_2(or_tmp_2474, (fsm_output[5]), and_527_cse);
  assign mux_2565_nl = MUX_s_1_2_2(mux_2564_nl, or_2528_cse, fsm_output[9]);
  assign mux_2569_nl = MUX_s_1_2_2(mux_2568_nl, mux_2565_nl, fsm_output[6]);
  assign or_2582_nl = (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign mux_2548_nl = MUX_s_1_2_2(nand_386_cse, or_2582_nl, fsm_output[9]);
  assign mux_2546_nl = MUX_s_1_2_2((~ or_tmp_2393), (fsm_output[5]), and_529_cse);
  assign or_2580_nl = (or_2377_cse & (fsm_output[5])) | (fsm_output[10]);
  assign mux_2547_nl = MUX_s_1_2_2(mux_2546_nl, or_2580_nl, fsm_output[9]);
  assign mux_2549_nl = MUX_s_1_2_2(mux_2548_nl, mux_2547_nl, fsm_output[6]);
  assign mux_2464_nl = MUX_s_1_2_2(mux_2569_nl, mux_2549_nl, fsm_output[8]);
  assign mux_2478_nl = MUX_s_1_2_2(mux_2477_nl, mux_2464_nl, fsm_output[7]);
  assign mux_2501_nl = MUX_s_1_2_2(mux_2500_nl, mux_2478_nl, fsm_output[4]);
  assign mux_2545_nl = MUX_s_1_2_2(mux_2544_nl, mux_2501_nl, fsm_output[3]);
  assign operator_64_false_mux1h_2_rgt = MUX1HOT_v_65_3_2(z_out_6, ({2'b00 , operator_64_false_slc_modExp_exp_63_1_3}),
      ({1'b0 , modExp_while_if_mux1h_nl}), {and_261_nl , and_dcpl_247 , (~ mux_2545_nl)});
  assign or_3532_cse = (fsm_output[6]) | and_757_cse;
  assign or_3609_nl = (~ (fsm_output[10])) | (fsm_output[6]) | (~ (fsm_output[2]))
      | (fsm_output[9]);
  assign mux_3935_cse = MUX_s_1_2_2(or_2965_cse, or_3609_nl, fsm_output[1]);
  assign mux_554_cse = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[6]);
  assign or_181_cse = (fsm_output[5]) | (fsm_output[3]);
  assign or_2644_cse = (fsm_output[3:2]!=2'b00);
  assign mux_544_cse = MUX_s_1_2_2((~ or_tmp_167), (fsm_output[10]), fsm_output[9]);
  assign mux_2643_cse = MUX_s_1_2_2(mux_tmp_2640, and_756_cse, fsm_output[6]);
  assign and_273_m1c = and_dcpl_147 & and_dcpl_90 & and_dcpl_107;
  assign and_756_cse = (fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]);
  assign and_757_cse = (fsm_output[10:9]==2'b11);
  assign modExp_result_and_rgt = (~ modExp_while_and_5) & and_273_m1c;
  assign modExp_result_and_1_rgt = modExp_while_and_5 & and_273_m1c;
  assign and_458_cse = (fsm_output[7]) & (fsm_output[9]);
  assign and_459_cse = (fsm_output[3:1]==3'b111);
  assign nand_166_nl = ~((fsm_output[2]) & (fsm_output[9]) & (fsm_output[1]) & (fsm_output[6])
      & (~ (fsm_output[10])));
  assign mux_2769_nl = MUX_s_1_2_2(nand_166_nl, or_tmp_2651, fsm_output[0]);
  assign nor_678_nl = ~((~ (fsm_output[4])) | (fsm_output[8]) | (~ (fsm_output[3]))
      | mux_2769_nl);
  assign or_2716_nl = (~ (fsm_output[2])) | (~ (fsm_output[9])) | (fsm_output[1])
      | not_tmp_49;
  assign or_2714_nl = (fsm_output[2]) | (fsm_output[9]) | (fsm_output[1]) | not_tmp_49;
  assign mux_2767_nl = MUX_s_1_2_2(or_2716_nl, or_2714_nl, fsm_output[0]);
  assign or_2717_nl = (fsm_output[3]) | mux_2767_nl;
  assign mux_2766_nl = MUX_s_1_2_2(or_2921_cse, mux_tmp_2760, fsm_output[0]);
  assign nand_58_nl = ~((fsm_output[3]) & (~ mux_2766_nl));
  assign mux_2768_nl = MUX_s_1_2_2(or_2717_nl, nand_58_nl, fsm_output[8]);
  assign nor_679_nl = ~((fsm_output[4]) | mux_2768_nl);
  assign mux_2770_nl = MUX_s_1_2_2(nor_678_nl, nor_679_nl, fsm_output[5]);
  assign mux_2762_nl = MUX_s_1_2_2(or_tmp_2651, or_2918_cse, fsm_output[0]);
  assign or_2708_nl = (fsm_output[0]) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[1])
      | not_tmp_49;
  assign mux_2763_nl = MUX_s_1_2_2(mux_2762_nl, or_2708_nl, fsm_output[3]);
  assign nor_680_nl = ~((fsm_output[8]) | mux_2763_nl);
  assign or_2702_nl = (fsm_output[2]) | (~ (fsm_output[9])) | (~ (fsm_output[1]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2761_nl = MUX_s_1_2_2(mux_tmp_2760, or_2702_nl, fsm_output[0]);
  assign nor_681_nl = ~((~ (fsm_output[8])) | (fsm_output[3]) | mux_2761_nl);
  assign mux_2764_nl = MUX_s_1_2_2(nor_680_nl, nor_681_nl, fsm_output[4]);
  assign nor_682_nl = ~((~ (fsm_output[0])) | (~ (fsm_output[2])) | (fsm_output[9])
      | (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign nor_683_nl = ~((fsm_output[2]) | (~ (fsm_output[9])) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (fsm_output[10]));
  assign nor_684_nl = ~((~ (fsm_output[2])) | (fsm_output[9]) | (fsm_output[1]) |
      not_tmp_49);
  assign mux_2758_nl = MUX_s_1_2_2(nor_683_nl, nor_684_nl, fsm_output[0]);
  assign mux_2759_nl = MUX_s_1_2_2(nor_682_nl, mux_2758_nl, fsm_output[3]);
  assign and_451_nl = (fsm_output[4]) & (fsm_output[8]) & mux_2759_nl;
  assign mux_2765_nl = MUX_s_1_2_2(mux_2764_nl, and_451_nl, fsm_output[5]);
  assign mux_2771_m1c = MUX_s_1_2_2(mux_2770_nl, mux_2765_nl, fsm_output[7]);
  assign or_470_cse = (fsm_output[9:8]!=2'b00);
  assign or_469_cse = (fsm_output[10:8]!=3'b100);
  assign mux_2926_cse = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[7]);
  assign mux_1036_cse = MUX_s_1_2_2((~ or_tmp_93), or_tmp_88, fsm_output[9]);
  assign mux_981_cse = MUX_s_1_2_2(or_tmp_94, or_tmp_93, fsm_output[9]);
  assign nor_685_nl = ~((fsm_output[6]) | (~ (fsm_output[5])) | (fsm_output[3]));
  assign nor_686_nl = ~((~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[3])));
  assign mux_2743_nl = MUX_s_1_2_2(nor_685_nl, nor_686_nl, fsm_output[0]);
  assign and_317_m1c = mux_2743_nl & and_dcpl_245 & (~ (fsm_output[8])) & (fsm_output[4])
      & (~ (fsm_output[1])) & nor_609_cse;
  assign or_80_cse = (fsm_output[9]) | (fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign nand_159_cse = ~((fsm_output[3]) & (fsm_output[10]));
  assign nor_657_cse = ~((~ (fsm_output[9])) | (fsm_output[2]));
  assign nor_653_cse = ~((~((~ (fsm_output[0])) | (fsm_output[9]))) | (fsm_output[2]));
  assign mux_498_cse = MUX_s_1_2_2(mux_tmp_165, or_2991_cse, fsm_output[4]);
  assign COMP_LOOP_or_32_cse = and_dcpl_117 | and_dcpl_130 | and_dcpl_140 | and_dcpl_149
      | and_dcpl_155 | and_dcpl_164 | and_dcpl_171 | and_dcpl_178 | and_dcpl_185
      | and_dcpl_189 | and_dcpl_197 | and_dcpl_202 | and_dcpl_211 | and_dcpl_219
      | and_dcpl_226 | and_dcpl_231;
  assign or_2855_cse = (~ (fsm_output[9])) | (fsm_output[2]);
  assign or_2991_cse = (fsm_output[10:8]!=3'b001);
  assign or_2998_cse = (fsm_output[10:8]!=3'b000);
  assign or_2947_cse = (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[2]) |
      (fsm_output[6]) | (fsm_output[10]);
  assign or_3008_cse = (fsm_output[9]) | nand_138_cse;
  assign or_2962_nl = (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_2961_nl = (fsm_output[9]) | nand_367_cse;
  assign mux_3281_cse = MUX_s_1_2_2(or_2962_nl, or_2961_nl, fsm_output[1]);
  assign or_2965_cse = (fsm_output[9]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[10]);
  assign nand_367_cse = ~((fsm_output[2]) & (fsm_output[6]) & (fsm_output[10]));
  assign and_407_cse = (fsm_output[5:4]==2'b11);
  assign or_3039_cse = (fsm_output[3:1]!=3'b000);
  assign or_3427_cse = (fsm_output[7]) | (fsm_output[5]);
  assign and_404_cse = (fsm_output[8:7]==2'b11);
  assign or_259_cse = (fsm_output[9:8]!=2'b01);
  assign and_676_cse = (fsm_output[5]) & (fsm_output[2]);
  assign and_672_cse = ((fsm_output[9]) | (fsm_output[6])) & (fsm_output[10]);
  assign and_395_cse = (fsm_output[7]) & (fsm_output[10]);
  assign or_3063_cse = (fsm_output[5:4]!=2'b00);
  assign or_352_cse = (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_3417_cse = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[6]);
  assign or_361_cse = (fsm_output[10:9]!=2'b01);
  assign or_3079_cse = (fsm_output[8:6]!=3'b000);
  assign or_3074_cse = (fsm_output[8:5]!=4'b0000);
  assign nor_609_cse = ~((fsm_output[10:9]!=2'b00));
  assign nand_142_cse = ~((fsm_output[8]) & (fsm_output[6]) & (fsm_output[10]));
  assign and_366_cse = (fsm_output[2]) & (fsm_output[4]);
  assign nand_138_cse = ~((fsm_output[8]) & (fsm_output[10]));
  assign mux_3555_cse = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), fsm_output[9]);
  assign and_350_cse = (fsm_output[7]) & (fsm_output[5]);
  assign nl_STAGE_LOOP_i_3_0_sva_2 = STAGE_LOOP_i_3_0_sva + 4'b0001;
  assign STAGE_LOOP_i_3_0_sva_2 = nl_STAGE_LOOP_i_3_0_sva_2[3:0];
  assign nl_COMP_LOOP_acc_psp_sva_1 = (VEC_LOOP_j_sva_11_0[11:4]) + conv_u2u_5_8(COMP_LOOP_k_9_4_sva_4_0);
  assign COMP_LOOP_acc_psp_sva_1 = nl_COMP_LOOP_acc_psp_sva_1[7:0];
  assign nl_COMP_LOOP_1_acc_5_mut_mx0w5 = tmp_10_lpi_4_dfm + COMP_LOOP_10_mul_mut;
  assign COMP_LOOP_1_acc_5_mut_mx0w5 = nl_COMP_LOOP_1_acc_5_mut_mx0w5[63:0];
  assign nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1 = $signed(operator_64_false_acc_mut_63_0)
      * $signed(COMP_LOOP_10_mul_mut);
  assign COMP_LOOP_1_modExp_1_while_if_mul_mut_1 = nl_COMP_LOOP_1_modExp_1_while_if_mul_mut_1[63:0];
  assign operator_64_false_slc_modExp_exp_63_1_3 = MUX_v_63_2_2((operator_66_true_div_cmp_z[63:1]),
      (tmp_10_lpi_4_dfm[63:1]), and_dcpl_256);
  assign nl_modulo_qr_sva_1_mx0w6 = modulo_result_rem_cmp_z + p_sva;
  assign modulo_qr_sva_1_mx0w6 = nl_modulo_qr_sva_1_mx0w6[63:0];
  assign or_70_cse = (fsm_output[2]) | (fsm_output[6]) | (~ (fsm_output[1])) | (~
      (fsm_output[8])) | (fsm_output[4]) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign or_56_cse = (fsm_output[2]) | (~ (fsm_output[6])) | (fsm_output[1]) | (~
      (fsm_output[8])) | (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign mux_340_cse = MUX_s_1_2_2(mux_tmp_141, or_tmp_94, fsm_output[4]);
  assign mux_375_cse = MUX_s_1_2_2(mux_tmp_130, or_2998_cse, fsm_output[4]);
  assign nl_COMP_LOOP_acc_1_cse_6_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0101});
  assign COMP_LOOP_acc_1_cse_6_sva_1 = nl_COMP_LOOP_acc_1_cse_6_sva_1[11:0];
  assign nl_COMP_LOOP_acc_1_cse_2_sva_1 = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0001});
  assign COMP_LOOP_acc_1_cse_2_sva_1 = nl_COMP_LOOP_acc_1_cse_2_sva_1[11:0];
  assign modExp_while_and_3 = (~ (modulo_result_rem_cmp_z[63])) & COMP_LOOP_nor_11_itm;
  assign modExp_while_and_5 = (modulo_result_rem_cmp_z[63]) & COMP_LOOP_nor_11_itm;
  assign nor_tmp_4 = (fsm_output[3]) & (fsm_output[5]);
  assign or_18_nl = (fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]);
  assign mux_tmp_14 = MUX_s_1_2_2((fsm_output[5]), or_18_nl, fsm_output[7]);
  assign not_tmp_39 = ~((fsm_output[4]) & (fsm_output[10]));
  assign or_tmp_68 = (fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3])) | (fsm_output[8])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign not_tmp_49 = ~((fsm_output[6]) & (fsm_output[10]));
  assign or_84_nl = (fsm_output[8]) | not_tmp_49;
  assign or_83_nl = (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_tmp_119 = MUX_s_1_2_2(or_84_nl, or_83_nl, fsm_output[3]);
  assign or_tmp_88 = (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_tmp_130 = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_88, fsm_output[9]);
  assign mux_tmp_131 = MUX_s_1_2_2(or_2991_cse, mux_tmp_130, fsm_output[4]);
  assign or_tmp_93 = (fsm_output[8]) | (~ (fsm_output[10]));
  assign nand_tmp_4 = ~((fsm_output[4]) & (~ mux_tmp_130));
  assign or_tmp_94 = (fsm_output[8]) | (fsm_output[10]);
  assign mux_tmp_139 = MUX_s_1_2_2((fsm_output[8]), or_tmp_94, fsm_output[9]);
  assign mux_tmp_141 = MUX_s_1_2_2(nand_138_cse, or_tmp_88, fsm_output[9]);
  assign or_tmp_96 = (fsm_output[4]) | mux_tmp_130;
  assign or_108_nl = (~ (fsm_output[4])) | (fsm_output[9]);
  assign mux_155_cse = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_88, or_108_nl);
  assign mux_161_cse = MUX_s_1_2_2(mux_tmp_130, or_3008_cse, fsm_output[4]);
  assign mux_tmp_165 = MUX_s_1_2_2(or_tmp_93, or_tmp_94, fsm_output[9]);
  assign mux_171_cse = MUX_s_1_2_2(or_469_cse, or_tmp_88, fsm_output[4]);
  assign or_tmp_104 = (fsm_output[10:9]!=2'b10);
  assign mux_tmp_214 = MUX_s_1_2_2(and_757_cse, or_tmp_104, fsm_output[5]);
  assign mux_tmp_215 = MUX_s_1_2_2(or_2414_cse, and_757_cse, fsm_output[5]);
  assign nand_tmp_7 = ~((fsm_output[5]) & (~ and_757_cse));
  assign mux_tmp_227 = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[9]);
  assign nor_tmp_23 = ((~ (fsm_output[5])) | (fsm_output[9])) & (fsm_output[10]);
  assign mux_tmp_228 = MUX_s_1_2_2(or_tmp_104, and_757_cse, fsm_output[5]);
  assign mux_tmp_231 = MUX_s_1_2_2(and_757_cse, or_2414_cse, fsm_output[5]);
  assign mux_tmp_236 = MUX_s_1_2_2(and_757_cse, mux_tmp_227, fsm_output[5]);
  assign or_tmp_114 = (fsm_output[5]) | and_757_cse;
  assign mux_259_cse = MUX_s_1_2_2((fsm_output[9]), and_757_cse, fsm_output[5]);
  assign or_163_cse = (~ (fsm_output[4])) | (fsm_output[8]);
  assign and_dcpl_1 = (~ (fsm_output[4])) & (fsm_output[1]);
  assign and_dcpl_2 = and_dcpl_1 & (fsm_output[0]);
  assign and_dcpl_4 = (fsm_output[8:7]==2'b01);
  assign and_dcpl_5 = and_dcpl_4 & (fsm_output[6]);
  assign and_dcpl_6 = nor_tmp_4 & (~ (fsm_output[2]));
  assign nor_1580_cse = ~((fsm_output[5]) | (fsm_output[7]));
  assign not_tmp_90 = ~((fsm_output[7:6]!=2'b00));
  assign or_tmp_167 = (fsm_output[6]) | (fsm_output[10]);
  assign nor_tmp_48 = (fsm_output[6]) & (fsm_output[10]);
  assign and_707_cse = (fsm_output[5]) & (fsm_output[8]);
  assign mux_648_cse = MUX_s_1_2_2((~ (fsm_output[8])), and_707_cse, fsm_output[6]);
  assign or_tmp_222 = (fsm_output[5]) | (fsm_output[8]);
  assign not_tmp_133 = ~((fsm_output[8:7]!=2'b00));
  assign nor_tmp_82 = (fsm_output[9:8]==2'b11);
  assign or_tmp_258 = (fsm_output[7]) | (fsm_output[9]);
  assign and_dcpl_19 = (fsm_output[4]) & (fsm_output[1]);
  assign and_dcpl_26 = (fsm_output[4]) & (~ (fsm_output[1]));
  assign and_dcpl_27 = and_dcpl_26 & (fsm_output[0]);
  assign and_dcpl_33 = (fsm_output[10:9]==2'b01);
  assign and_dcpl_34 = ~((fsm_output[4]) | (fsm_output[1]));
  assign and_dcpl_39 = (fsm_output[5]) & (~ (fsm_output[3]));
  assign and_dcpl_40 = and_dcpl_39 & (~ (fsm_output[2]));
  assign and_dcpl_44 = and_dcpl_4 & (~ (fsm_output[6]));
  assign and_dcpl_48 = and_dcpl_1 & (~ (fsm_output[0]));
  assign and_dcpl_55 = and_dcpl_26 & (~ (fsm_output[0]));
  assign and_dcpl_59 = (fsm_output[10:9]==2'b10);
  assign or_3394_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[9]) | (fsm_output[10]);
  assign mux_1077_nl = MUX_s_1_2_2(or_3394_nl, nand_356_cse, or_491_cse);
  assign mux_1078_nl = MUX_s_1_2_2(mux_1077_nl, nand_357_cse, fsm_output[6]);
  assign not_tmp_208 = MUX_s_1_2_2(mux_1078_nl, nand_358_cse, fsm_output[8]);
  assign and_dcpl_87 = and_dcpl_34 & (~ (fsm_output[0]));
  assign and_dcpl_88 = and_dcpl_87 & nor_609_cse;
  assign and_dcpl_90 = not_tmp_133 & (~ (fsm_output[6]));
  assign and_dcpl_91 = ~((fsm_output[3]) | (fsm_output[5]));
  assign and_dcpl_92 = and_dcpl_91 & (~ (fsm_output[2]));
  assign and_dcpl_93 = and_dcpl_92 & and_dcpl_90;
  assign and_dcpl_98 = and_dcpl_2 & and_757_cse;
  assign and_dcpl_103 = and_dcpl_40 & and_dcpl_44;
  assign and_dcpl_107 = and_dcpl_27 & nor_609_cse;
  assign and_dcpl_108 = and_dcpl_40 & and_dcpl_90;
  assign and_dcpl_109 = and_dcpl_108 & and_dcpl_107;
  assign and_dcpl_111 = and_dcpl_19 & (~ (fsm_output[0]));
  assign and_dcpl_112 = and_dcpl_111 & nor_609_cse;
  assign and_dcpl_113 = not_tmp_133 & (fsm_output[6]);
  assign and_dcpl_114 = (fsm_output[3]) & (~ (fsm_output[5]));
  assign and_dcpl_115 = and_dcpl_114 & (~ (fsm_output[2]));
  assign and_dcpl_117 = and_dcpl_115 & and_dcpl_113 & and_dcpl_112;
  assign and_dcpl_118 = and_dcpl_91 & (fsm_output[2]);
  assign or_tmp_453 = (fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[4]) | (~
      (fsm_output[8])) | (fsm_output[10]);
  assign or_510_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[10]);
  assign or_508_nl = (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[4])) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_1081_nl = MUX_s_1_2_2(or_tmp_453, or_508_nl, fsm_output[0]);
  assign mux_tmp_1082 = MUX_s_1_2_2(or_510_nl, mux_1081_nl, fsm_output[3]);
  assign and_dcpl_126 = and_dcpl_34 & (fsm_output[0]);
  assign and_dcpl_127 = and_dcpl_126 & nor_609_cse;
  assign and_dcpl_130 = and_dcpl_92 & and_dcpl_5 & and_dcpl_127;
  assign and_dcpl_135 = (fsm_output[8:7]==2'b10);
  assign and_dcpl_136 = and_dcpl_135 & (~ (fsm_output[6]));
  assign and_dcpl_139 = and_dcpl_6 & and_dcpl_136;
  assign and_dcpl_140 = and_dcpl_139 & and_dcpl_88;
  assign and_dcpl_144 = and_dcpl_2 & nor_609_cse;
  assign and_dcpl_146 = and_404_cse & (~ (fsm_output[6]));
  assign and_dcpl_147 = and_dcpl_114 & (fsm_output[2]);
  assign and_dcpl_149 = and_dcpl_147 & and_dcpl_146 & and_dcpl_144;
  assign and_dcpl_152 = and_404_cse & (fsm_output[6]);
  assign and_dcpl_153 = and_dcpl_39 & (fsm_output[2]);
  assign and_dcpl_155 = and_dcpl_153 & and_dcpl_152 & and_dcpl_112;
  assign and_dcpl_162 = and_dcpl_27 & and_dcpl_33;
  assign and_dcpl_164 = and_dcpl_147 & and_dcpl_113 & and_dcpl_162;
  assign and_dcpl_170 = and_dcpl_118 & and_dcpl_5;
  assign and_dcpl_171 = and_dcpl_170 & and_dcpl_87 & and_dcpl_33;
  assign and_dcpl_177 = and_dcpl_2 & and_dcpl_33;
  assign and_dcpl_178 = and_dcpl_139 & and_dcpl_177;
  assign and_dcpl_185 = and_dcpl_92 & and_dcpl_146 & and_dcpl_111 & and_dcpl_33;
  assign and_dcpl_189 = and_dcpl_6 & and_dcpl_152 & and_dcpl_162;
  assign and_dcpl_191 = ~((fsm_output[8]) | (fsm_output[6]));
  assign and_dcpl_196 = and_dcpl_40 & and_dcpl_113;
  assign and_dcpl_197 = and_dcpl_196 & and_dcpl_87 & and_dcpl_59;
  assign and_dcpl_202 = and_dcpl_170 & and_dcpl_2 & and_dcpl_59;
  assign and_dcpl_208 = and_dcpl_48 & and_dcpl_59;
  assign and_dcpl_209 = nor_tmp_4 & (fsm_output[2]);
  assign and_dcpl_211 = and_dcpl_209 & and_dcpl_136 & and_dcpl_208;
  assign and_dcpl_219 = and_dcpl_118 & and_dcpl_146 & and_dcpl_27 & and_dcpl_59;
  assign and_dcpl_224 = and_dcpl_55 & and_dcpl_59;
  assign and_dcpl_226 = and_dcpl_209 & and_dcpl_152 & and_dcpl_224;
  assign and_dcpl_231 = and_dcpl_196 & and_dcpl_98;
  assign not_tmp_248 = ~((fsm_output[5]) & (fsm_output[10]));
  assign or_580_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (fsm_output[10]);
  assign or_579_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (fsm_output[10]);
  assign mux_tmp_1116 = MUX_s_1_2_2(or_580_nl, or_579_nl, fsm_output[2]);
  assign or_tmp_532 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (~ (fsm_output[10]));
  assign or_586_cse = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000);
  assign or_591_cse = (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (fsm_output[10]);
  assign nand_337_cse = ~((fsm_output[9]) & (fsm_output[5]) & (fsm_output[10]));
  assign not_tmp_253 = ~((fsm_output[2]) & (fsm_output[10]));
  assign or_691_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (fsm_output[10]);
  assign or_690_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (fsm_output[10]);
  assign mux_tmp_1180 = MUX_s_1_2_2(or_691_nl, or_690_nl, fsm_output[2]);
  assign or_tmp_643 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (~ (fsm_output[10]));
  assign nand_334_cse = ~((VEC_LOOP_j_sva_11_0[0]) & (fsm_output[9]) & (fsm_output[5])
      & (fsm_output[10]));
  assign or_702_cse = (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (fsm_output[10]);
  assign or_802_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (fsm_output[10]);
  assign or_801_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010)
      | (fsm_output[10]);
  assign mux_tmp_1244 = MUX_s_1_2_2(or_802_nl, or_801_nl, fsm_output[2]);
  assign or_tmp_756 = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010)
      | (~ (fsm_output[10]));
  assign nor_209_cse = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001));
  assign or_912_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (fsm_output[10]);
  assign or_911_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011)
      | (fsm_output[10]);
  assign mux_tmp_1308 = MUX_s_1_2_2(or_912_nl, or_911_nl, fsm_output[2]);
  assign or_tmp_866 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011)
      | (~ (fsm_output[10]));
  assign or_1022_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (fsm_output[10]);
  assign or_1021_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (fsm_output[10]);
  assign mux_tmp_1372 = MUX_s_1_2_2(or_1022_nl, or_1021_nl, fsm_output[2]);
  assign or_tmp_974 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (~ (fsm_output[10]));
  assign or_1028_cse = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010);
  assign or_1133_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (fsm_output[10]);
  assign or_1132_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101)
      | (fsm_output[10]);
  assign mux_tmp_1436 = MUX_s_1_2_2(or_1133_nl, or_1132_nl, fsm_output[2]);
  assign or_tmp_1085 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (~ (fsm_output[10]));
  assign or_1244_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (fsm_output[10]);
  assign or_1243_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110)
      | (fsm_output[10]);
  assign mux_tmp_1500 = MUX_s_1_2_2(or_1244_nl, or_1243_nl, fsm_output[2]);
  assign or_tmp_1198 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (~ (fsm_output[10]));
  assign nor_223_cse = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011));
  assign or_1354_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (fsm_output[10]);
  assign or_1353_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111)
      | (fsm_output[10]);
  assign mux_tmp_1564 = MUX_s_1_2_2(or_1354_nl, or_1353_nl, fsm_output[2]);
  assign or_tmp_1308 = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (~ (fsm_output[10]));
  assign not_tmp_318 = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3]) & (fsm_output[10]));
  assign or_1464_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000) | (fsm_output[10]);
  assign or_1463_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000)
      | (fsm_output[10]);
  assign mux_tmp_1628 = MUX_s_1_2_2(or_1464_nl, or_1463_nl, fsm_output[2]);
  assign or_tmp_1416 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000) | not_tmp_318;
  assign or_1470_cse = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100);
  assign or_1575_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001) | (fsm_output[10]);
  assign or_1574_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001)
      | (fsm_output[10]);
  assign mux_tmp_1692 = MUX_s_1_2_2(or_1575_nl, or_1574_nl, fsm_output[2]);
  assign or_tmp_1527 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001) | not_tmp_318;
  assign or_1686_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010) | (fsm_output[10]);
  assign or_1685_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010)
      | (fsm_output[10]);
  assign mux_tmp_1756 = MUX_s_1_2_2(or_1686_nl, or_1685_nl, fsm_output[2]);
  assign or_tmp_1640 = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010) | not_tmp_318;
  assign nor_239_cse = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101));
  assign or_1796_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011) | (fsm_output[10]);
  assign or_1795_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011)
      | (fsm_output[10]);
  assign mux_tmp_1820 = MUX_s_1_2_2(or_1796_nl, or_1795_nl, fsm_output[2]);
  assign or_tmp_1750 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011) | not_tmp_318;
  assign not_tmp_357 = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:2]==2'b11) & (fsm_output[10]));
  assign or_1906_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100) | (fsm_output[10]);
  assign or_1905_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100)
      | (fsm_output[10]);
  assign mux_tmp_1884 = MUX_s_1_2_2(or_1906_nl, or_1905_nl, fsm_output[2]);
  assign or_tmp_1858 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | not_tmp_357;
  assign or_1912_cse = (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110);
  assign or_2017_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101) | (fsm_output[10]);
  assign or_2016_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101)
      | (fsm_output[10]);
  assign mux_tmp_1948 = MUX_s_1_2_2(or_2017_nl, or_2016_nl, fsm_output[2]);
  assign or_tmp_1969 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | not_tmp_357;
  assign not_tmp_377 = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:1]==3'b111) & (fsm_output[10]));
  assign or_2128_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110) | (fsm_output[10]);
  assign or_2127_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110)
      | (fsm_output[10]);
  assign mux_tmp_2012 = MUX_s_1_2_2(or_2128_nl, or_2127_nl, fsm_output[2]);
  assign or_tmp_2082 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) | not_tmp_377;
  assign and_564_cse = (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111);
  assign not_tmp_387 = ~((fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111)
      & (fsm_output[10]));
  assign nand_225_nl = ~((~ (fsm_output[7])) & (fsm_output[9]) & (fsm_output[5])
      & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111) & (~ (fsm_output[10])));
  assign or_2237_nl = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1111)
      | (fsm_output[10]);
  assign mux_tmp_2076 = MUX_s_1_2_2(nand_225_nl, or_2237_nl, fsm_output[2]);
  assign not_tmp_390 = ~((COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111) & (fsm_output[10]));
  assign or_tmp_2192 = (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[5]) |
      not_tmp_390;
  assign nor_tmp_265 = (fsm_output[9]) & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111)
      & (fsm_output[10]);
  assign and_dcpl_235 = and_dcpl_48 & nor_609_cse;
  assign and_dcpl_236 = and_dcpl_115 & and_dcpl_90;
  assign and_dcpl_237 = and_dcpl_236 & and_dcpl_235;
  assign or_tmp_2274 = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (fsm_output[7])
      | (fsm_output[10]);
  assign or_tmp_2276 = (fsm_output[7]) | (fsm_output[10]);
  assign or_tmp_2277 = and_526_cse | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[10]);
  assign or_tmp_2280 = (~ (fsm_output[7])) | (fsm_output[10]);
  assign or_tmp_2281 = (fsm_output[7]) | (~ (fsm_output[10]));
  assign mux_tmp_2159 = MUX_s_1_2_2((~ (fsm_output[7])), or_tmp_2280, fsm_output[9]);
  assign or_tmp_2294 = nor_753_cse | (~ (fsm_output[2])) | (~ (fsm_output[7])) |
      (fsm_output[10]);
  assign mux_tmp_2172 = MUX_s_1_2_2((fsm_output[7]), and_395_cse, and_529_cse);
  assign or_tmp_2297 = nor_758_cse | (fsm_output[7]) | (fsm_output[10]);
  assign mux_2175_nl = MUX_s_1_2_2(or_tmp_2276, (fsm_output[7]), and_529_cse);
  assign mux_tmp_2176 = MUX_s_1_2_2(or_tmp_2297, mux_2175_nl, fsm_output[0]);
  assign mux_tmp_2178 = MUX_s_1_2_2((~ and_395_cse), or_tmp_2276, fsm_output[2]);
  assign or_tmp_2302 = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[10]);
  assign mux_2234_nl = MUX_s_1_2_2(mux_tmp_139, mux_tmp_165, or_3388_cse);
  assign mux_tmp_2235 = MUX_s_1_2_2(mux_tmp_139, mux_2234_nl, fsm_output[3]);
  assign mux_2239_nl = MUX_s_1_2_2(mux_tmp_141, or_3008_cse, fsm_output[1]);
  assign mux_tmp_2241 = MUX_s_1_2_2(mux_tmp_130, mux_2239_nl, fsm_output[3]);
  assign or_tmp_2340 = nor_303_cse | (fsm_output[8]) | (fsm_output[10]);
  assign or_tmp_2341 = (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[8]) |
      (fsm_output[10]);
  assign mux_tmp_2262 = MUX_s_1_2_2(mux_tmp_141, or_3008_cse, and_526_cse);
  assign and_524_cse = (fsm_output[3]) & (fsm_output[0]) & (fsm_output[1]);
  assign mux_tmp_2287 = MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, and_524_cse);
  assign mux_tmp_2289 = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), nor_303_cse);
  assign mux_tmp_2293 = MUX_s_1_2_2(or_259_cse, or_2991_cse, fsm_output[1]);
  assign or_tmp_2360 = (fsm_output[1]) | (fsm_output[9]) | nand_138_cse;
  assign mux_tmp_2311 = MUX_s_1_2_2(or_3008_cse, or_2991_cse, fsm_output[1]);
  assign or_tmp_2376 = (fsm_output[4]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_tmp_2389 = (~ (fsm_output[8])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign nand_188_nl = ~((fsm_output[8]) & (fsm_output[5]));
  assign mux_tmp_2347 = MUX_s_1_2_2(nand_188_nl, or_tmp_2389, fsm_output[9]);
  assign or_tmp_2390 = (~ (fsm_output[8])) | (fsm_output[5]) | (fsm_output[10]);
  assign or_2447_nl = (~ (fsm_output[8])) | (fsm_output[5]);
  assign mux_tmp_2348 = MUX_s_1_2_2(or_2447_nl, or_tmp_2390, fsm_output[9]);
  assign mux_tmp_2350 = MUX_s_1_2_2(mux_tmp_2348, or_tmp_2389, fsm_output[6]);
  assign not_tmp_431 = ~((fsm_output[8]) & (fsm_output[5]) & (fsm_output[10]));
  assign mux_2352_nl = MUX_s_1_2_2(not_tmp_431, or_tmp_2389, fsm_output[9]);
  assign or_2448_nl = (fsm_output[9]) | (fsm_output[8]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_tmp_2353 = MUX_s_1_2_2(mux_2352_nl, or_2448_nl, fsm_output[6]);
  assign or_tmp_2393 = (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_tmp_2394 = (fsm_output[5]) | (~ (fsm_output[10]));
  assign mux_tmp_2355 = MUX_s_1_2_2(or_tmp_2394, or_tmp_2393, fsm_output[8]);
  assign or_2451_nl = (fsm_output[9]) | mux_tmp_2355;
  assign mux_tmp_2356 = MUX_s_1_2_2(mux_tmp_2348, or_2451_nl, fsm_output[6]);
  assign or_tmp_2396 = (fsm_output[6]) | mux_tmp_2347;
  assign or_tmp_2397 = (fsm_output[8]) | (fsm_output[5]) | (fsm_output[10]);
  assign or_tmp_2399 = (fsm_output[8]) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign mux_tmp_2359 = MUX_s_1_2_2(or_tmp_2399, or_tmp_2397, fsm_output[9]);
  assign or_2457_nl = (fsm_output[9:8]!=2'b10) | not_tmp_248;
  assign mux_tmp_2361 = MUX_s_1_2_2(mux_tmp_2347, or_2457_nl, fsm_output[6]);
  assign mux_tmp_2363 = MUX_s_1_2_2(or_tmp_222, or_tmp_2397, fsm_output[9]);
  assign or_2459_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_tmp_2364 = MUX_s_1_2_2(or_2459_nl, mux_tmp_2363, fsm_output[6]);
  assign or_tmp_2404 = (fsm_output[8]) | not_tmp_248;
  assign mux_tmp_2365 = MUX_s_1_2_2(mux_tmp_2347, or_tmp_2404, fsm_output[6]);
  assign nand_tmp_54 = ~((fsm_output[6]) & (~ mux_tmp_2363));
  assign or_tmp_2405 = (fsm_output[8]) | (~ (fsm_output[5]));
  assign mux_tmp_2369 = MUX_s_1_2_2(or_tmp_2404, or_tmp_2405, fsm_output[9]);
  assign mux_tmp_2370 = MUX_s_1_2_2(or_tmp_2389, mux_tmp_2355, fsm_output[9]);
  assign mux_tmp_2371 = MUX_s_1_2_2(mux_tmp_2370, mux_tmp_2369, fsm_output[6]);
  assign mux_2375_nl = MUX_s_1_2_2(mux_tmp_2355, or_tmp_2399, fsm_output[9]);
  assign mux_tmp_2376 = MUX_s_1_2_2(mux_2375_nl, or_tmp_2405, fsm_output[6]);
  assign mux_tmp_2377 = MUX_s_1_2_2(or_tmp_2399, or_tmp_222, fsm_output[9]);
  assign mux_tmp_2378 = MUX_s_1_2_2(mux_tmp_2377, or_tmp_2405, fsm_output[6]);
  assign or_2462_nl = (fsm_output[9]) | not_tmp_431;
  assign mux_tmp_2382 = MUX_s_1_2_2(or_2462_nl, or_tmp_2397, fsm_output[6]);
  assign or_tmp_2407 = (fsm_output[8]) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign mux_2385_nl = MUX_s_1_2_2(or_tmp_2405, or_tmp_2407, fsm_output[9]);
  assign mux_tmp_2386 = MUX_s_1_2_2(mux_tmp_2377, mux_2385_nl, fsm_output[6]);
  assign mux_2387_nl = MUX_s_1_2_2(or_tmp_2393, or_tmp_2394, fsm_output[8]);
  assign mux_2388_nl = MUX_s_1_2_2(mux_2387_nl, or_tmp_2407, fsm_output[9]);
  assign mux_tmp_2389 = MUX_s_1_2_2(mux_tmp_2377, mux_2388_nl, fsm_output[6]);
  assign or_2475_nl = (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_2474_nl = (fsm_output[1]) | not_tmp_49;
  assign mux_tmp_2424 = MUX_s_1_2_2(or_2475_nl, or_2474_nl, fsm_output[3]);
  assign nand_183_cse = ~((fsm_output[1]) & (fsm_output[6]) & (fsm_output[10]));
  assign or_2488_nl = (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[10]);
  assign or_2487_nl = (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[7]) | (~
      (fsm_output[3])) | (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_2430_nl = MUX_s_1_2_2(or_2488_nl, or_2487_nl, fsm_output[0]);
  assign nor_741_nl = ~((fsm_output[5]) | mux_2430_nl);
  assign or_2484_nl = (fsm_output[3]) | (~ (fsm_output[1])) | (fsm_output[6]) | (~
      (fsm_output[10]));
  assign nand_182_nl = ~((fsm_output[3]) & (fsm_output[1]) & (fsm_output[6]) & (~
      (fsm_output[10])));
  assign mux_2427_nl = MUX_s_1_2_2(or_2484_nl, nand_182_nl, fsm_output[7]);
  assign nor_742_nl = ~((~ (fsm_output[9])) | (fsm_output[2]) | mux_2427_nl);
  assign nor_743_nl = ~((fsm_output[9]) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | mux_tmp_2424);
  assign mux_2428_nl = MUX_s_1_2_2(nor_742_nl, nor_743_nl, fsm_output[0]);
  assign or_2479_nl = (fsm_output[7]) | (fsm_output[3]) | (fsm_output[1]) | (~ (fsm_output[6]))
      | (fsm_output[10]);
  assign or_2478_nl = (fsm_output[7]) | (fsm_output[3]) | nand_183_cse;
  assign mux_2425_nl = MUX_s_1_2_2(or_2479_nl, or_2478_nl, fsm_output[2]);
  assign nor_744_nl = ~((fsm_output[9]) | mux_2425_nl);
  assign nor_745_nl = ~((~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[7]) |
      mux_tmp_2424);
  assign mux_2426_nl = MUX_s_1_2_2(nor_744_nl, nor_745_nl, fsm_output[0]);
  assign mux_2429_nl = MUX_s_1_2_2(mux_2428_nl, mux_2426_nl, fsm_output[5]);
  assign mux_2431_nl = MUX_s_1_2_2(nor_741_nl, mux_2429_nl, fsm_output[4]);
  assign nor_746_nl = ~((fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[7]) |
      (fsm_output[3]) | (fsm_output[1]) | not_tmp_49);
  assign nor_747_nl = ~((~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[7]) |
      (fsm_output[3]) | (fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign mux_2421_nl = MUX_s_1_2_2(nor_746_nl, nor_747_nl, fsm_output[0]);
  assign nor_748_nl = ~((~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[10]));
  assign nand_388_nl = ~((fsm_output[7]) & (fsm_output[3]) & (fsm_output[1]) & (~
      (fsm_output[6])) & (fsm_output[10]));
  assign or_2465_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[10]);
  assign mux_2419_nl = MUX_s_1_2_2(nand_388_nl, or_2465_nl, fsm_output[2]);
  assign nor_749_nl = ~((fsm_output[9]) | mux_2419_nl);
  assign mux_2420_nl = MUX_s_1_2_2(nor_748_nl, nor_749_nl, fsm_output[0]);
  assign mux_2422_nl = MUX_s_1_2_2(mux_2421_nl, mux_2420_nl, fsm_output[5]);
  assign nor_750_nl = ~((~ (fsm_output[5])) | (fsm_output[0]) | (fsm_output[9]) |
      (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[1]))
      | (fsm_output[6]) | (fsm_output[10]));
  assign mux_2423_nl = MUX_s_1_2_2(mux_2422_nl, nor_750_nl, fsm_output[4]);
  assign not_tmp_441 = MUX_s_1_2_2(mux_2431_nl, mux_2423_nl, fsm_output[8]);
  assign or_tmp_2436 = ~((fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]) & (~
      (fsm_output[10])));
  assign or_2512_nl = (fsm_output[3]) | (fsm_output[8]) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_2442_nl = MUX_s_1_2_2(or_tmp_2436, or_2512_nl, fsm_output[7]);
  assign nor_729_nl = ~((fsm_output[2]) | (~ (fsm_output[5])) | mux_2442_nl);
  assign nor_730_nl = ~((~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[7]) |
      (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_2443_nl = MUX_s_1_2_2(nor_729_nl, nor_730_nl, fsm_output[9]);
  assign nor_1628_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (~ (fsm_output[3])) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[7])
      | (~ (fsm_output[10])));
  assign mux_2444_nl = MUX_s_1_2_2(mux_2443_nl, nor_1628_nl, fsm_output[4]);
  assign nor_732_nl = ~((fsm_output[9]) | (~ (fsm_output[2])) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (~((fsm_output[3]) & (fsm_output[8]) & (fsm_output[6])
      & (fsm_output[10]))));
  assign nor_733_nl = ~((fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[7])) |
      (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]));
  assign nor_734_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign nor_735_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[3]) |
      (fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_2439_nl = MUX_s_1_2_2(nor_734_nl, nor_735_nl, fsm_output[2]);
  assign mux_2440_nl = MUX_s_1_2_2(nor_733_nl, mux_2439_nl, fsm_output[9]);
  assign mux_2441_nl = MUX_s_1_2_2(nor_732_nl, mux_2440_nl, fsm_output[4]);
  assign mux_2445_nl = MUX_s_1_2_2(mux_2444_nl, mux_2441_nl, fsm_output[1]);
  assign nor_736_nl = ~((fsm_output[9]) | (fsm_output[2]) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]));
  assign nor_737_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (fsm_output[8]) | (fsm_output[6]) | (~ (fsm_output[10])));
  assign nor_738_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      nand_142_cse);
  assign mux_2435_nl = MUX_s_1_2_2(nor_737_nl, nor_738_nl, fsm_output[2]);
  assign nor_739_nl = ~((~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_2436_nl = MUX_s_1_2_2(mux_2435_nl, nor_739_nl, fsm_output[9]);
  assign mux_2437_nl = MUX_s_1_2_2(nor_736_nl, mux_2436_nl, fsm_output[4]);
  assign or_2494_nl = (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) | (~
      (fsm_output[10]));
  assign mux_2433_nl = MUX_s_1_2_2(or_2494_nl, or_tmp_2436, fsm_output[7]);
  assign or_2495_nl = (~ (fsm_output[2])) | (fsm_output[5]) | mux_2433_nl;
  assign or_2490_nl = (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[7]) | (~
      (fsm_output[3])) | (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_2434_nl = MUX_s_1_2_2(or_2495_nl, or_2490_nl, fsm_output[9]);
  assign nor_740_nl = ~((fsm_output[4]) | mux_2434_nl);
  assign mux_2438_nl = MUX_s_1_2_2(mux_2437_nl, nor_740_nl, fsm_output[1]);
  assign not_tmp_446 = MUX_s_1_2_2(mux_2445_nl, mux_2438_nl, fsm_output[0]);
  assign mux_2447_nl = MUX_s_1_2_2((fsm_output[3]), (~ (fsm_output[3])), or_2368_cse);
  assign nor_1612_nl = ~(nor_758_cse | (fsm_output[3]));
  assign mux_2448_nl = MUX_s_1_2_2(mux_2447_nl, nor_1612_nl, fsm_output[0]);
  assign and_dcpl_241 = mux_2448_nl & nor_1580_cse & and_dcpl_191 & (~ (fsm_output[4]))
      & nor_609_cse;
  assign and_dcpl_245 = ~((fsm_output[2]) | (fsm_output[7]));
  assign nor_726_nl = ~((fsm_output[5:3]!=3'b110));
  assign nor_727_nl = ~((fsm_output[5:3]!=3'b001));
  assign mux_2453_nl = MUX_s_1_2_2(nor_726_nl, nor_727_nl, fsm_output[0]);
  assign and_dcpl_247 = mux_2453_nl & and_dcpl_245 & and_dcpl_191 & (~ (fsm_output[1]))
      & nor_609_cse;
  assign nor_tmp_324 = (fsm_output[5]) & (fsm_output[10]);
  assign nand_386_cse = ~((~(or_3388_cse & (fsm_output[2]))) & nor_tmp_324);
  assign or_2528_cse = nor_758_cse | (fsm_output[5]) | (fsm_output[10]);
  assign or_tmp_2474 = (fsm_output[5]) | (fsm_output[10]);
  assign or_2534_cse = and_529_cse | (fsm_output[5]) | (~ (fsm_output[10]));
  assign mux_2465_cse = MUX_s_1_2_2((~ (fsm_output[5])), or_tmp_2393, fsm_output[9]);
  assign or_2540_cse = (~ (fsm_output[2])) | (fsm_output[5]) | (fsm_output[10]);
  assign or_2541_cse = (fsm_output[2]) | (~ nor_tmp_324);
  assign nand_173_cse = ~(nand_196_cse & nor_tmp_324);
  assign mux_2486_cse = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), fsm_output[5]);
  assign mux_2494_cse = MUX_s_1_2_2(or_tmp_2474, (fsm_output[5]), fsm_output[2]);
  assign mux_2515_cse = MUX_s_1_2_2((fsm_output[5]), nor_tmp_324, fsm_output[2]);
  assign mux_2516_cse = MUX_s_1_2_2(or_tmp_2474, nor_tmp_324, fsm_output[2]);
  assign mux_tmp_2640 = MUX_s_1_2_2(nor_609_cse, and_757_cse, fsm_output[7]);
  assign nor_694_cse = ~((fsm_output[7]) | (fsm_output[9]) | (fsm_output[10]));
  assign and_465_cse = (fsm_output[5]) & (fsm_output[7]) & (fsm_output[9]) & (fsm_output[10]);
  assign mux_tmp_2659 = MUX_s_1_2_2(nor_694_cse, and_756_cse, fsm_output[5]);
  assign and_dcpl_256 = and_dcpl_108 & and_dcpl_55 & nor_609_cse;
  assign mux_tmp_2669 = MUX_s_1_2_2((~ (fsm_output[6])), or_352_cse, fsm_output[9]);
  assign mux_tmp_2672 = MUX_s_1_2_2(and_757_cse, mux_tmp_2669, fsm_output[7]);
  assign mux_tmp_2675 = MUX_s_1_2_2((fsm_output[6]), or_tmp_167, fsm_output[9]);
  assign not_tmp_500 = MUX_s_1_2_2(or_tmp_167, (~ mux_554_cse), fsm_output[9]);
  assign mux_2681_nl = MUX_s_1_2_2(mux_554_cse, nor_tmp_48, fsm_output[9]);
  assign mux_tmp_2682 = MUX_s_1_2_2((~ mux_2681_nl), mux_tmp_2675, fsm_output[7]);
  assign mux_tmp_2690 = MUX_s_1_2_2(mux_tmp_2675, and_757_cse, fsm_output[7]);
  assign mux_tmp_2691 = MUX_s_1_2_2(mux_tmp_2675, and_672_cse, fsm_output[7]);
  assign mux_tmp_2693 = MUX_s_1_2_2(nor_tmp_48, or_tmp_167, fsm_output[9]);
  assign or_tmp_2603 = (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_2698_itm = MUX_s_1_2_2(or_tmp_2603, (fsm_output[6]), fsm_output[9]);
  assign or_tmp_2604 = (fsm_output[9]) | (~ mux_554_cse);
  assign mux_tmp_2700 = MUX_s_1_2_2((~ mux_2698_itm), or_tmp_2604, fsm_output[7]);
  assign mux_tmp_2702 = MUX_s_1_2_2((~ nor_tmp_48), or_352_cse, fsm_output[9]);
  assign mux_tmp_2703 = MUX_s_1_2_2((~ mux_2698_itm), mux_tmp_2702, fsm_output[7]);
  assign mux_tmp_2706 = MUX_s_1_2_2((~ mux_2698_itm), mux_tmp_2669, fsm_output[7]);
  assign mux_2708_nl = MUX_s_1_2_2(or_tmp_2603, or_tmp_167, fsm_output[9]);
  assign mux_tmp_2709 = MUX_s_1_2_2((~ mux_2708_nl), mux_tmp_2669, fsm_output[7]);
  assign mux_tmp_2715 = MUX_s_1_2_2(and_672_cse, mux_tmp_2669, fsm_output[7]);
  assign nor_1575_nl = ~((fsm_output[9]) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_tmp_2736 = MUX_s_1_2_2(nor_1575_nl, mux_tmp_2669, fsm_output[7]);
  assign and_dcpl_257 = and_dcpl_108 & and_dcpl_112;
  assign and_dcpl_260 = and_dcpl_92 & and_dcpl_136;
  assign and_dcpl_262 = and_dcpl_135 & (fsm_output[6]);
  assign and_dcpl_270 = and_dcpl_147 & and_dcpl_44;
  assign and_dcpl_278 = and_dcpl_6 & and_dcpl_90;
  assign and_dcpl_280 = and_dcpl_19 & (fsm_output[0]);
  assign or_2678_nl = (~ (fsm_output[1])) | (~ (fsm_output[2])) | (~ (fsm_output[6]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign or_2677_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[8])
      | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_tmp_2745 = MUX_s_1_2_2(or_2678_nl, or_2677_nl, fsm_output[9]);
  assign or_2694_nl = (fsm_output[2]) | (fsm_output[6]) | (~ (fsm_output[8])) | (fsm_output[4])
      | (fsm_output[10]);
  assign or_2693_nl = (~ (fsm_output[2])) | (fsm_output[6]) | (~ (fsm_output[8]))
      | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_2754_nl = MUX_s_1_2_2(or_2694_nl, or_2693_nl, fsm_output[1]);
  assign or_2695_nl = (fsm_output[9]) | mux_2754_nl;
  assign mux_2755_nl = MUX_s_1_2_2(or_2695_nl, or_70_cse, fsm_output[0]);
  assign or_2696_nl = (fsm_output[3]) | mux_2755_nl;
  assign or_2690_nl = (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[6])
      | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_2752_nl = MUX_s_1_2_2(or_2690_nl, mux_tmp_2745, fsm_output[0]);
  assign or_2689_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[8])
      | not_tmp_39;
  assign or_2687_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (~ (fsm_output[6]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_2750_nl = MUX_s_1_2_2(or_2689_nl, or_2687_nl, fsm_output[9]);
  assign or_2686_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[6]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (~ (fsm_output[10]));
  assign or_2684_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[8])
      | not_tmp_39;
  assign mux_2749_nl = MUX_s_1_2_2(or_2686_nl, or_2684_nl, fsm_output[9]);
  assign mux_2751_nl = MUX_s_1_2_2(mux_2750_nl, mux_2749_nl, fsm_output[0]);
  assign mux_2753_nl = MUX_s_1_2_2(mux_2752_nl, mux_2751_nl, fsm_output[3]);
  assign mux_2756_nl = MUX_s_1_2_2(or_2696_nl, mux_2753_nl, fsm_output[5]);
  assign or_2681_nl = (fsm_output[9]) | (fsm_output[1]) | (~((fsm_output[2]) & (fsm_output[6])
      & (fsm_output[8]) & (fsm_output[4]) & (fsm_output[10])));
  assign mux_2747_nl = MUX_s_1_2_2(or_2681_nl, or_56_cse, fsm_output[0]);
  assign or_2675_nl = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[4]))
      | (fsm_output[10]);
  assign or_2674_nl = (~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[8]) | not_tmp_39;
  assign mux_2744_nl = MUX_s_1_2_2(or_2675_nl, or_2674_nl, fsm_output[1]);
  assign or_2676_nl = (fsm_output[9]) | mux_2744_nl;
  assign mux_2746_nl = MUX_s_1_2_2(mux_tmp_2745, or_2676_nl, fsm_output[0]);
  assign mux_2748_nl = MUX_s_1_2_2(mux_2747_nl, mux_2746_nl, fsm_output[3]);
  assign or_2682_nl = (fsm_output[5]) | mux_2748_nl;
  assign mux_2757_itm = MUX_s_1_2_2(mux_2756_nl, or_2682_nl, fsm_output[7]);
  assign or_2705_nl = (fsm_output[9]) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[10]);
  assign or_2704_nl = (fsm_output[9]) | (~ (fsm_output[1])) | (fsm_output[6]) | (~
      (fsm_output[10]));
  assign mux_tmp_2760 = MUX_s_1_2_2(or_2705_nl, or_2704_nl, fsm_output[2]);
  assign or_tmp_2651 = (fsm_output[2]) | (fsm_output[9]) | (~ (fsm_output[1])) |
      (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_tmp_2682 = (fsm_output[10:7]!=4'b0110);
  assign or_tmp_2683 = ~((fsm_output[10:7]==4'b0111));
  assign or_tmp_2690 = (fsm_output[7]) | (fsm_output[9]) | nand_138_cse;
  assign or_tmp_2693 = (fsm_output[10:7]!=4'b0010);
  assign or_tmp_2696 = (fsm_output[10:7]!=4'b0011);
  assign or_tmp_2697 = (fsm_output[10:7]!=4'b0100);
  assign mux_tmp_2796 = MUX_s_1_2_2(or_3008_cse, or_2998_cse, fsm_output[7]);
  assign or_tmp_2701 = (fsm_output[10:7]!=4'b0001);
  assign or_tmp_2703 = (fsm_output[10:7]!=4'b1000);
  assign or_tmp_2704 = (fsm_output[10:7]!=4'b0101);
  assign or_tmp_2706 = (fsm_output[10:7]!=4'b1100);
  assign or_tmp_2709 = (fsm_output[10:7]!=4'b1001);
  assign or_tmp_2714 = (~ (fsm_output[7])) | (fsm_output[9]) | nand_138_cse;
  assign or_2785_nl = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[7]) | (~ (fsm_output[9]))
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign or_2784_nl = (~((fsm_output[3]) & (fsm_output[6]) & (fsm_output[7]) & (~
      (fsm_output[9])))) | nand_138_cse;
  assign mux_2834_nl = MUX_s_1_2_2(or_tmp_2704, or_tmp_2709, fsm_output[6]);
  assign mux_2832_nl = MUX_s_1_2_2(or_2387_cse, or_2991_cse, fsm_output[7]);
  assign mux_2833_nl = MUX_s_1_2_2(mux_2832_nl, or_tmp_2706, fsm_output[6]);
  assign mux_2835_nl = MUX_s_1_2_2(mux_2834_nl, mux_2833_nl, fsm_output[3]);
  assign mux_2836_nl = MUX_s_1_2_2(or_2784_nl, mux_2835_nl, fsm_output[4]);
  assign mux_2837_nl = MUX_s_1_2_2(or_2785_nl, mux_2836_nl, fsm_output[5]);
  assign nand_394_nl = ~((fsm_output[10:7]==4'b1101));
  assign mux_2829_nl = MUX_s_1_2_2(nand_394_nl, or_tmp_2703, fsm_output[6]);
  assign nand_65_nl = ~((fsm_output[3]) & (~ mux_2829_nl));
  assign mux_2827_nl = MUX_s_1_2_2(or_tmp_2693, or_tmp_2682, fsm_output[6]);
  assign mux_2828_nl = MUX_s_1_2_2(mux_2827_nl, or_tmp_2709, fsm_output[3]);
  assign mux_2830_nl = MUX_s_1_2_2(nand_65_nl, mux_2828_nl, fsm_output[4]);
  assign mux_2826_nl = MUX_s_1_2_2(or_tmp_2696, or_tmp_2693, fsm_output[6]);
  assign or_2780_nl = (fsm_output[4:3]!=2'b00) | mux_2826_nl;
  assign mux_2831_nl = MUX_s_1_2_2(mux_2830_nl, or_2780_nl, fsm_output[5]);
  assign mux_2838_nl = MUX_s_1_2_2(mux_2837_nl, mux_2831_nl, fsm_output[2]);
  assign or_2778_nl = (~ (fsm_output[4])) | (~ (fsm_output[3])) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[9]) | nand_138_cse;
  assign mux_2821_nl = MUX_s_1_2_2(or_tmp_2703, or_tmp_2696, fsm_output[6]);
  assign mux_2820_nl = MUX_s_1_2_2(or_tmp_2714, mux_tmp_2796, fsm_output[6]);
  assign mux_2822_nl = MUX_s_1_2_2(mux_2821_nl, mux_2820_nl, fsm_output[3]);
  assign or_2776_nl = (fsm_output[3]) | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_2823_nl = MUX_s_1_2_2(mux_2822_nl, or_2776_nl, fsm_output[4]);
  assign mux_2824_nl = MUX_s_1_2_2(or_2778_nl, mux_2823_nl, fsm_output[5]);
  assign or_2775_nl = (fsm_output[10:6]!=5'b01010);
  assign mux_2816_nl = MUX_s_1_2_2(or_tmp_2703, or_tmp_2683, fsm_output[6]);
  assign mux_2817_nl = MUX_s_1_2_2(or_2775_nl, mux_2816_nl, fsm_output[3]);
  assign or_2774_nl = (fsm_output[3]) | (~ (fsm_output[7])) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[10]);
  assign mux_2818_nl = MUX_s_1_2_2(mux_2817_nl, or_2774_nl, fsm_output[4]);
  assign mux_2815_nl = MUX_s_1_2_2(or_tmp_2714, or_tmp_2682, fsm_output[6]);
  assign nand_64_nl = ~((fsm_output[4:3]==2'b11) & (~ mux_2815_nl));
  assign mux_2819_nl = MUX_s_1_2_2(mux_2818_nl, nand_64_nl, fsm_output[5]);
  assign mux_2825_nl = MUX_s_1_2_2(mux_2824_nl, mux_2819_nl, fsm_output[2]);
  assign mux_2839_nl = MUX_s_1_2_2(mux_2838_nl, mux_2825_nl, fsm_output[1]);
  assign or_2770_nl = (fsm_output[6]) | (~ (fsm_output[7])) | (fsm_output[9]) | nand_138_cse;
  assign mux_2810_nl = MUX_s_1_2_2(or_tmp_2709, or_tmp_2697, fsm_output[6]);
  assign mux_2811_nl = MUX_s_1_2_2(or_2770_nl, mux_2810_nl, fsm_output[3]);
  assign mux_2807_nl = MUX_s_1_2_2(or_2991_cse, or_3008_cse, fsm_output[7]);
  assign mux_2808_nl = MUX_s_1_2_2(or_tmp_2706, mux_2807_nl, fsm_output[6]);
  assign mux_2809_nl = MUX_s_1_2_2(mux_2808_nl, or_tmp_2704, fsm_output[3]);
  assign mux_2812_nl = MUX_s_1_2_2(mux_2811_nl, mux_2809_nl, fsm_output[4]);
  assign or_2771_nl = (fsm_output[5]) | mux_2812_nl;
  assign mux_2804_nl = MUX_s_1_2_2(or_tmp_2706, or_tmp_2683, fsm_output[6]);
  assign mux_2803_nl = MUX_s_1_2_2(or_tmp_2701, or_tmp_2704, fsm_output[6]);
  assign mux_2805_nl = MUX_s_1_2_2(mux_2804_nl, mux_2803_nl, fsm_output[3]);
  assign mux_2801_nl = MUX_s_1_2_2(or_tmp_2693, or_tmp_2701, fsm_output[6]);
  assign mux_2802_nl = MUX_s_1_2_2(or_tmp_2703, mux_2801_nl, fsm_output[3]);
  assign mux_2806_nl = MUX_s_1_2_2(mux_2805_nl, mux_2802_nl, fsm_output[4]);
  assign nand_63_nl = ~((fsm_output[5]) & (~ mux_2806_nl));
  assign mux_2813_nl = MUX_s_1_2_2(or_2771_nl, nand_63_nl, fsm_output[2]);
  assign mux_2797_nl = MUX_s_1_2_2(mux_tmp_2796, or_tmp_2690, fsm_output[6]);
  assign mux_2795_nl = MUX_s_1_2_2(or_tmp_2697, or_tmp_2696, fsm_output[6]);
  assign mux_2798_nl = MUX_s_1_2_2(mux_2797_nl, mux_2795_nl, fsm_output[3]);
  assign or_2759_nl = (fsm_output[4]) | mux_2798_nl;
  assign or_2754_nl = (fsm_output[10:6]!=5'b10010);
  assign mux_2793_nl = MUX_s_1_2_2(or_tmp_2683, or_tmp_2693, fsm_output[6]);
  assign mux_2794_nl = MUX_s_1_2_2(or_2754_nl, mux_2793_nl, fsm_output[3]);
  assign nand_62_nl = ~((fsm_output[4]) & (~ mux_2794_nl));
  assign mux_2799_nl = MUX_s_1_2_2(or_2759_nl, nand_62_nl, fsm_output[5]);
  assign or_2751_nl = (~ (fsm_output[3])) | (~ (fsm_output[6])) | (fsm_output[7])
      | (~ (fsm_output[9])) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_2789_nl = MUX_s_1_2_2(or_tmp_2682, or_tmp_2690, fsm_output[6]);
  assign mux_2788_nl = MUX_s_1_2_2(or_2407_cse, or_2387_cse, fsm_output[7]);
  assign or_2747_nl = (fsm_output[6]) | mux_2788_nl;
  assign mux_2790_nl = MUX_s_1_2_2(mux_2789_nl, or_2747_nl, fsm_output[3]);
  assign mux_2791_nl = MUX_s_1_2_2(or_2751_nl, mux_2790_nl, fsm_output[4]);
  assign mux_2786_nl = MUX_s_1_2_2(or_tmp_2683, or_tmp_2682, fsm_output[6]);
  assign or_2740_nl = (fsm_output[10:6]!=5'b00001);
  assign mux_2787_nl = MUX_s_1_2_2(mux_2786_nl, or_2740_nl, fsm_output[3]);
  assign or_2743_nl = (fsm_output[4]) | mux_2787_nl;
  assign mux_2792_nl = MUX_s_1_2_2(mux_2791_nl, or_2743_nl, fsm_output[5]);
  assign mux_2800_nl = MUX_s_1_2_2(mux_2799_nl, mux_2792_nl, fsm_output[2]);
  assign mux_2814_nl = MUX_s_1_2_2(mux_2813_nl, mux_2800_nl, fsm_output[1]);
  assign mux_2840_itm = MUX_s_1_2_2(mux_2839_nl, mux_2814_nl, fsm_output[0]);
  assign mux_tmp_2841 = MUX_s_1_2_2((~ or_tmp_2281), (fsm_output[10]), fsm_output[9]);
  assign or_tmp_2729 = (fsm_output[9]) | (fsm_output[7]) | (~ (fsm_output[10]));
  assign or_tmp_2731 = (~((~ (fsm_output[9])) | (fsm_output[7]))) | (fsm_output[10]);
  assign mux_tmp_2843 = MUX_s_1_2_2(or_tmp_2281, or_tmp_2276, fsm_output[9]);
  assign mux_tmp_2844 = MUX_s_1_2_2(mux_tmp_2843, or_tmp_2731, fsm_output[6]);
  assign or_tmp_2734 = (fsm_output[6]) | mux_tmp_2159;
  assign mux_tmp_2848 = MUX_s_1_2_2((~ and_395_cse), or_tmp_2280, fsm_output[9]);
  assign mux_tmp_2850 = MUX_s_1_2_2(mux_2171_cse, mux_tmp_2848, fsm_output[6]);
  assign or_tmp_2736 = (~ (fsm_output[9])) | (fsm_output[7]) | (~ (fsm_output[10]));
  assign mux_tmp_2851 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[10]), fsm_output[9]);
  assign mux_tmp_2856 = MUX_s_1_2_2((fsm_output[7]), or_tmp_2281, fsm_output[9]);
  assign mux_2858_nl = MUX_s_1_2_2((fsm_output[10]), (~ and_395_cse), fsm_output[9]);
  assign nand_tmp_67 = ~((fsm_output[6]) & mux_2858_nl);
  assign mux_tmp_2862 = MUX_s_1_2_2(or_tmp_2276, mux_tmp_2159, fsm_output[6]);
  assign mux_tmp_2863 = MUX_s_1_2_2((~ or_tmp_2276), or_tmp_2280, fsm_output[9]);
  assign or_tmp_2739 = (fsm_output[9]) | (~ (fsm_output[7])) | (fsm_output[10]);
  assign mux_tmp_2867 = MUX_s_1_2_2(or_tmp_2739, mux_2203_cse, fsm_output[6]);
  assign or_tmp_2740 = (fsm_output[7:6]!=2'b01);
  assign mux_2875_nl = MUX_s_1_2_2((~ or_tmp_2276), (fsm_output[10]), fsm_output[9]);
  assign mux_tmp_2876 = MUX_s_1_2_2(or_tmp_2736, mux_2875_nl, fsm_output[6]);
  assign or_2800_nl = (fsm_output[6]) | mux_tmp_2863;
  assign mux_tmp_2878 = MUX_s_1_2_2(or_tmp_2734, or_2800_nl, fsm_output[0]);
  assign mux_tmp_2879 = MUX_s_1_2_2(mux_2203_cse, or_tmp_2280, fsm_output[6]);
  assign or_tmp_2742 = (fsm_output[9]) | (~ (fsm_output[7]));
  assign mux_tmp_2880 = MUX_s_1_2_2(mux_2203_cse, or_tmp_2742, fsm_output[6]);
  assign mux_tmp_2886 = MUX_s_1_2_2(mux_2171_cse, or_tmp_2742, fsm_output[6]);
  assign mux_tmp_2888 = MUX_s_1_2_2(mux_2171_cse, mux_tmp_2159, fsm_output[6]);
  assign mux_tmp_2890 = MUX_s_1_2_2(or_tmp_2280, or_tmp_2281, fsm_output[6]);
  assign or_tmp_2743 = (fsm_output[6]) | mux_tmp_2841;
  assign nand_tmp_68 = ~((fsm_output[6]) & (~ mux_2203_cse));
  assign mux_tmp_2895 = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[7]), fsm_output[9]);
  assign or_tmp_2745 = (fsm_output[6]) | (fsm_output[9]) | (~ (fsm_output[7]));
  assign or_tmp_2746 = (~ (fsm_output[9])) | (~ (fsm_output[7])) | (fsm_output[10]);
  assign mux_2901_nl = MUX_s_1_2_2(or_tmp_2276, (~ and_395_cse), fsm_output[9]);
  assign nand_tmp_69 = ~((fsm_output[6]) & mux_2901_nl);
  assign mux_tmp_2906 = MUX_s_1_2_2(mux_tmp_2843, mux_tmp_2159, fsm_output[6]);
  assign mux_2909_nl = MUX_s_1_2_2((~ or_tmp_2280), (fsm_output[10]), fsm_output[9]);
  assign mux_tmp_2910 = MUX_s_1_2_2(mux_2909_nl, or_tmp_2739, fsm_output[6]);
  assign nand_tmp_70 = ~((fsm_output[6]) & (~ mux_2171_cse));
  assign mux_tmp_2912 = MUX_s_1_2_2(or_tmp_2276, (fsm_output[7]), fsm_output[9]);
  assign nand_tmp_71 = ~((fsm_output[6]) & (~ mux_tmp_2912));
  assign mux_tmp_2916 = MUX_s_1_2_2(or_tmp_2281, mux_tmp_2851, fsm_output[6]);
  assign mux_tmp_2920 = MUX_s_1_2_2(mux_2203_cse, mux_tmp_2848, fsm_output[6]);
  assign or_tmp_2749 = (fsm_output[9]) | (~ and_395_cse);
  assign or_tmp_2774 = (~ (fsm_output[1])) | (~ (fsm_output[8])) | (fsm_output[6])
      | (fsm_output[10]);
  assign or_2835_cse = (~ (fsm_output[1])) | (fsm_output[8]) | not_tmp_49;
  assign mux_tmp_2996 = MUX_s_1_2_2(or_2835_cse, or_tmp_2774, fsm_output[3]);
  assign nor_667_cse = ~((~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[1])
      | (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign or_2840_nl = (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[6]) | (~
      (fsm_output[10]));
  assign mux_2998_cse = MUX_s_1_2_2(or_tmp_2774, or_2840_nl, fsm_output[3]);
  assign nor_661_nl = ~((fsm_output[0]) | (fsm_output[5]) | (~ (fsm_output[7])) |
      (fsm_output[3]) | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[6])) |
      (fsm_output[10]));
  assign or_2842_nl = (fsm_output[3]) | (~ (fsm_output[1])) | (fsm_output[8]) | (~
      (fsm_output[6])) | (fsm_output[10]);
  assign mux_2999_nl = MUX_s_1_2_2(or_2842_nl, mux_tmp_2996, fsm_output[7]);
  assign nor_662_nl = ~((fsm_output[5]) | mux_2999_nl);
  assign nor_663_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | mux_2998_cse);
  assign mux_3000_nl = MUX_s_1_2_2(nor_662_nl, nor_663_nl, fsm_output[0]);
  assign mux_3001_nl = MUX_s_1_2_2(nor_661_nl, mux_3000_nl, fsm_output[2]);
  assign or_2836_nl = (~ (fsm_output[5])) | (fsm_output[7]) | mux_tmp_2996;
  assign or_2831_nl = (fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) | (~
      (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_2997_nl = MUX_s_1_2_2(or_2836_nl, or_2831_nl, fsm_output[0]);
  assign nor_664_nl = ~((fsm_output[2]) | mux_2997_nl);
  assign mux_3002_nl = MUX_s_1_2_2(mux_3001_nl, nor_664_nl, fsm_output[9]);
  assign and_445_nl = (fsm_output[0]) & (fsm_output[5]) & (fsm_output[7]) & (fsm_output[3])
      & (fsm_output[1]) & (fsm_output[8]) & (fsm_output[6]) & (fsm_output[10]);
  assign nor_665_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[6]) | (~ (fsm_output[10])));
  assign nor_666_nl = ~((fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[1]))
      | (fsm_output[8]) | not_tmp_49);
  assign mux_2992_nl = MUX_s_1_2_2(nor_666_nl, nor_667_cse, fsm_output[5]);
  assign mux_2993_nl = MUX_s_1_2_2(nor_665_nl, mux_2992_nl, fsm_output[0]);
  assign mux_2994_nl = MUX_s_1_2_2(and_445_nl, mux_2993_nl, fsm_output[2]);
  assign and_446_nl = (fsm_output[5]) & (fsm_output[7]) & (fsm_output[3]) & (~ (fsm_output[1]))
      & (fsm_output[8]) & (fsm_output[6]) & (~ (fsm_output[10]));
  assign nor_668_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_2990_nl = MUX_s_1_2_2(and_446_nl, nor_668_nl, fsm_output[0]);
  assign nor_669_nl = ~((fsm_output[0]) | (fsm_output[5]) | (fsm_output[7]) | (~
      (fsm_output[3])) | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[6]))
      | (fsm_output[10]));
  assign mux_2991_nl = MUX_s_1_2_2(mux_2990_nl, nor_669_nl, fsm_output[2]);
  assign mux_2995_nl = MUX_s_1_2_2(mux_2994_nl, mux_2991_nl, fsm_output[9]);
  assign not_tmp_557 = MUX_s_1_2_2(mux_3002_nl, mux_2995_nl, fsm_output[4]);
  assign nor_tmp_405 = (fsm_output[8]) & (fsm_output[10]);
  assign mux_3799_nl = MUX_s_1_2_2(or_tmp_88, (~ (fsm_output[8])), fsm_output[2]);
  assign mux_tmp_3007 = MUX_s_1_2_2(mux_3799_nl, or_tmp_88, fsm_output[9]);
  assign mux_3006_nl = MUX_s_1_2_2(or_tmp_88, (~ (fsm_output[8])), fsm_output[2]);
  assign or_2848_nl = (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_tmp_3008 = MUX_s_1_2_2(mux_3006_nl, or_2848_nl, fsm_output[9]);
  assign or_tmp_2791 = nor_657_cse | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_tmp_3014 = MUX_s_1_2_2((fsm_output[8]), or_tmp_93, fsm_output[2]);
  assign or_tmp_2795 = (fsm_output[2]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign or_tmp_2802 = (fsm_output[9]) | (fsm_output[2]) | (~ nor_tmp_405);
  assign or_tmp_2803 = (fsm_output[2]) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign or_2863_nl = (fsm_output[2]) | (~ nor_tmp_405);
  assign mux_tmp_3024 = MUX_s_1_2_2(or_2863_nl, or_tmp_2803, fsm_output[9]);
  assign mux_3031_nl = MUX_s_1_2_2((fsm_output[8]), nor_tmp_405, fsm_output[2]);
  assign mux_tmp_3032 = MUX_s_1_2_2((~ mux_3031_nl), or_tmp_88, fsm_output[9]);
  assign mux_tmp_3049 = MUX_s_1_2_2(or_tmp_2791, mux_tmp_3008, fsm_output[0]);
  assign or_tmp_2814 = (fsm_output[2]) | (fsm_output[8]) | (fsm_output[10]);
  assign nor_tmp_410 = (fsm_output[1]) & (fsm_output[4]) & (fsm_output[3]) & (fsm_output[10]);
  assign and_dcpl_304 = and_dcpl_108 & and_dcpl_280 & nor_609_cse;
  assign or_3025_nl = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[3]) | (fsm_output[6])
      | (fsm_output[7]) | (fsm_output[8]);
  assign mux_3321_nl = MUX_s_1_2_2(or_3079_cse, or_3025_nl, and_407_cse);
  assign or_3367_nl = (fsm_output[10]) | mux_3321_nl;
  assign or_3023_nl = and_524_cse | (fsm_output[8:6]!=3'b000);
  assign or_3022_nl = (fsm_output[3]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8]);
  assign mux_3319_nl = MUX_s_1_2_2(or_3023_nl, or_3022_nl, fsm_output[2]);
  assign mux_3320_nl = MUX_s_1_2_2(or_3079_cse, mux_3319_nl, and_407_cse);
  assign nand_149_nl = ~((fsm_output[10]) & mux_3320_nl);
  assign not_tmp_619 = MUX_s_1_2_2(or_3367_nl, nand_149_nl, fsm_output[9]);
  assign mux_tmp_3329 = MUX_s_1_2_2(nor_694_cse, and_757_cse, fsm_output[6]);
  assign nor_tmp_457 = (fsm_output[7:6]==2'b11);
  assign mux_tmp_3341 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), fsm_output[6]);
  assign mux_3342_nl = MUX_s_1_2_2(not_tmp_90, mux_tmp_3341, fsm_output[3]);
  assign mux_tmp_3343 = MUX_s_1_2_2(mux_3342_nl, nor_tmp_457, fsm_output[4]);
  assign mux_tmp_3361 = MUX_s_1_2_2(nor_tmp_4, (fsm_output[5]), fsm_output[2]);
  assign or_tmp_2988 = (~((fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[9]))) | (fsm_output[10]);
  assign or_3061_nl = (fsm_output[9:6]!=4'b0000);
  assign mux_tmp_3378 = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), or_3061_nl);
  assign not_tmp_647 = ~((fsm_output[6]) | (fsm_output[7]) | (fsm_output[10]));
  assign or_3087_nl = (fsm_output[8:7]!=2'b00) | (~ and_dcpl_209);
  assign or_12_nl = (fsm_output[8]) | (fsm_output[7]) | (fsm_output[5]);
  assign mux_tmp_3410 = MUX_s_1_2_2(or_3087_nl, or_12_nl, fsm_output[6]);
  assign mux_tmp_3414 = MUX_s_1_2_2((~ (fsm_output[3])), (fsm_output[3]), fsm_output[5]);
  assign mux_tmp_3415 = MUX_s_1_2_2(mux_tmp_3414, nor_tmp_4, fsm_output[2]);
  assign mux_tmp_3417 = MUX_s_1_2_2((fsm_output[5]), or_181_cse, fsm_output[2]);
  assign or_tmp_3023 = (fsm_output[7]) | mux_tmp_3417;
  assign mux_3416_nl = MUX_s_1_2_2((~ (fsm_output[5])), mux_tmp_3415, fsm_output[7]);
  assign mux_tmp_3418 = MUX_s_1_2_2(or_tmp_3023, mux_3416_nl, fsm_output[8]);
  assign mux_tmp_3420 = MUX_s_1_2_2(nor_tmp_4, (fsm_output[5]), fsm_output[7]);
  assign mux_tmp_3421 = MUX_s_1_2_2((~ mux_tmp_3420), mux_tmp_14, fsm_output[8]);
  assign mux_tmp_3423 = MUX_s_1_2_2(and_dcpl_209, (fsm_output[5]), fsm_output[7]);
  assign mux_tmp_3424 = MUX_s_1_2_2((~ mux_tmp_14), mux_tmp_3423, fsm_output[8]);
  assign mux_tmp_3425 = MUX_s_1_2_2(and_dcpl_91, nor_tmp_4, fsm_output[2]);
  assign mux_3426_nl = MUX_s_1_2_2(mux_tmp_3425, (fsm_output[5]), fsm_output[7]);
  assign mux_3427_nl = MUX_s_1_2_2((~ and_350_cse), mux_3426_nl, fsm_output[8]);
  assign not_tmp_663 = MUX_s_1_2_2(mux_3427_nl, (~ mux_tmp_3424), fsm_output[6]);
  assign mux_3422_nl = MUX_s_1_2_2(mux_tmp_3421, mux_tmp_3418, fsm_output[6]);
  assign mux_tmp_3429 = MUX_s_1_2_2(not_tmp_663, mux_3422_nl, fsm_output[4]);
  assign mux_3430_nl = MUX_s_1_2_2((~ (fsm_output[5])), mux_tmp_3425, fsm_output[7]);
  assign mux_3431_nl = MUX_s_1_2_2(or_3427_cse, mux_3430_nl, fsm_output[8]);
  assign mux_tmp_3432 = MUX_s_1_2_2(mux_tmp_3421, mux_3431_nl, fsm_output[6]);
  assign mux_3433_nl = MUX_s_1_2_2((fsm_output[5]), or_181_cse, fsm_output[7]);
  assign mux_tmp_3434 = MUX_s_1_2_2((~ mux_3433_nl), and_350_cse, fsm_output[8]);
  assign mux_tmp_3435 = MUX_s_1_2_2(and_dcpl_91, mux_tmp_3414, fsm_output[2]);
  assign mux_3436_nl = MUX_s_1_2_2(mux_tmp_3435, (fsm_output[5]), fsm_output[7]);
  assign not_tmp_665 = MUX_s_1_2_2(and_350_cse, (~ mux_3436_nl), fsm_output[8]);
  assign mux_3447_nl = MUX_s_1_2_2(and_dcpl_91, (fsm_output[5]), fsm_output[7]);
  assign mux_3448_nl = MUX_s_1_2_2(and_350_cse, (~ mux_3447_nl), fsm_output[8]);
  assign mux_3449_nl = MUX_s_1_2_2(mux_3448_nl, mux_tmp_3434, fsm_output[6]);
  assign mux_3445_nl = MUX_s_1_2_2((~ mux_tmp_3423), mux_tmp_14, fsm_output[8]);
  assign mux_3443_nl = MUX_s_1_2_2((~ (fsm_output[5])), mux_tmp_3435, fsm_output[7]);
  assign mux_3444_nl = MUX_s_1_2_2(or_3427_cse, mux_3443_nl, fsm_output[8]);
  assign mux_3446_nl = MUX_s_1_2_2(mux_3445_nl, mux_3444_nl, fsm_output[6]);
  assign mux_3450_nl = MUX_s_1_2_2((~ mux_3449_nl), mux_3446_nl, fsm_output[4]);
  assign mux_3441_nl = MUX_s_1_2_2(not_tmp_665, mux_tmp_3424, fsm_output[6]);
  assign mux_3442_nl = MUX_s_1_2_2((~ mux_3441_nl), mux_tmp_3432, fsm_output[4]);
  assign mux_3451_nl = MUX_s_1_2_2(mux_3450_nl, mux_3442_nl, fsm_output[1]);
  assign mux_3438_nl = MUX_s_1_2_2(not_tmp_665, mux_tmp_3434, fsm_output[6]);
  assign mux_3439_nl = MUX_s_1_2_2((~ mux_3438_nl), mux_tmp_3432, fsm_output[4]);
  assign mux_3440_nl = MUX_s_1_2_2(mux_3439_nl, mux_tmp_3429, fsm_output[1]);
  assign mux_3452_nl = MUX_s_1_2_2(mux_3451_nl, mux_3440_nl, fsm_output[0]);
  assign or_3090_nl = (fsm_output[8:6]!=3'b001) | mux_tmp_3361;
  assign mux_3412_nl = MUX_s_1_2_2(or_3090_nl, mux_tmp_3410, fsm_output[4]);
  assign or_3088_nl = (fsm_output[8:5]!=4'b0010);
  assign mux_3411_nl = MUX_s_1_2_2(or_3088_nl, mux_tmp_3410, fsm_output[4]);
  assign mux_3413_nl = MUX_s_1_2_2(mux_3412_nl, mux_3411_nl, fsm_output[1]);
  assign mux_tmp_3453 = MUX_s_1_2_2(mux_3452_nl, mux_3413_nl, fsm_output[9]);
  assign mux_tmp_3456 = MUX_s_1_2_2(mux_tmp_3361, mux_tmp_3417, fsm_output[7]);
  assign mux_tmp_3457 = MUX_s_1_2_2((~ mux_tmp_3456), or_3427_cse, fsm_output[8]);
  assign mux_3454_nl = MUX_s_1_2_2((~ (fsm_output[5])), nor_tmp_4, fsm_output[7]);
  assign mux_3455_nl = MUX_s_1_2_2(or_tmp_3023, mux_3454_nl, fsm_output[8]);
  assign mux_tmp_3458 = MUX_s_1_2_2(mux_tmp_3457, mux_3455_nl, fsm_output[6]);
  assign mux_tmp_3459 = MUX_s_1_2_2(nor_1580_cse, mux_tmp_3420, fsm_output[8]);
  assign mux_3460_nl = MUX_s_1_2_2(mux_tmp_3415, (fsm_output[5]), fsm_output[7]);
  assign not_tmp_672 = MUX_s_1_2_2(and_350_cse, (~ mux_3460_nl), fsm_output[8]);
  assign mux_3462_nl = MUX_s_1_2_2(not_tmp_672, mux_tmp_3459, fsm_output[6]);
  assign mux_tmp_3463 = MUX_s_1_2_2((~ mux_3462_nl), mux_tmp_3458, fsm_output[4]);
  assign mux_tmp_3464 = MUX_s_1_2_2(nor_tmp_4, mux_tmp_3417, fsm_output[7]);
  assign mux_3469_nl = MUX_s_1_2_2(not_tmp_672, mux_tmp_3424, fsm_output[6]);
  assign mux_3470_nl = MUX_s_1_2_2((~ mux_3469_nl), mux_tmp_3458, fsm_output[4]);
  assign mux_3471_nl = MUX_s_1_2_2(mux_tmp_3429, mux_3470_nl, fsm_output[1]);
  assign mux_3465_nl = MUX_s_1_2_2((~ mux_tmp_3464), or_3427_cse, fsm_output[8]);
  assign mux_3466_nl = MUX_s_1_2_2(mux_3465_nl, mux_tmp_3418, fsm_output[6]);
  assign mux_3467_nl = MUX_s_1_2_2(not_tmp_663, mux_3466_nl, fsm_output[4]);
  assign mux_3468_nl = MUX_s_1_2_2(mux_3467_nl, mux_tmp_3463, fsm_output[1]);
  assign mux_tmp_3472 = MUX_s_1_2_2(mux_3471_nl, mux_3468_nl, fsm_output[0]);
  assign mux_tmp_3473 = MUX_s_1_2_2((~ (fsm_output[5])), mux_tmp_3361, fsm_output[7]);
  assign or_3095_nl = (fsm_output[7]) | (fsm_output[5]) | (fsm_output[3]);
  assign mux_tmp_3474 = MUX_s_1_2_2(or_3095_nl, mux_tmp_3473, fsm_output[8]);
  assign mux_3475_nl = MUX_s_1_2_2(mux_tmp_3361, or_181_cse, fsm_output[7]);
  assign mux_3476_nl = MUX_s_1_2_2((~ mux_3475_nl), or_3427_cse, fsm_output[8]);
  assign mux_tmp_3477 = MUX_s_1_2_2(mux_3476_nl, mux_tmp_3474, fsm_output[6]);
  assign mux_3479_nl = MUX_s_1_2_2(and_350_cse, (~ mux_tmp_3456), fsm_output[8]);
  assign mux_3478_nl = MUX_s_1_2_2(nor_1580_cse, mux_tmp_3464, fsm_output[8]);
  assign mux_3480_nl = MUX_s_1_2_2(mux_3479_nl, mux_3478_nl, fsm_output[6]);
  assign mux_tmp_3481 = MUX_s_1_2_2((~ mux_3480_nl), mux_tmp_3477, fsm_output[4]);
  assign mux_3484_nl = MUX_s_1_2_2(and_350_cse, (~ mux_tmp_3420), fsm_output[8]);
  assign mux_3485_itm = MUX_s_1_2_2(mux_3484_nl, mux_tmp_3459, fsm_output[6]);
  assign mux_3488_nl = MUX_s_1_2_2(and_350_cse, (~ mux_tmp_3464), fsm_output[8]);
  assign mux_3489_nl = MUX_s_1_2_2(mux_3488_nl, mux_tmp_3459, fsm_output[6]);
  assign mux_3490_nl = MUX_s_1_2_2((~ mux_3489_nl), mux_tmp_3477, fsm_output[4]);
  assign mux_tmp_3491 = MUX_s_1_2_2(mux_tmp_3463, mux_3490_nl, fsm_output[1]);
  assign mux_3482_nl = MUX_s_1_2_2(or_tmp_3023, mux_tmp_3473, fsm_output[8]);
  assign mux_3483_nl = MUX_s_1_2_2(mux_tmp_3457, mux_3482_nl, fsm_output[6]);
  assign mux_3486_nl = MUX_s_1_2_2((~ mux_3485_itm), mux_3483_nl, fsm_output[4]);
  assign mux_3487_nl = MUX_s_1_2_2(mux_3486_nl, mux_tmp_3481, fsm_output[1]);
  assign mux_3492_nl = MUX_s_1_2_2(mux_tmp_3491, mux_3487_nl, fsm_output[0]);
  assign mux_3493_nl = MUX_s_1_2_2(mux_3492_nl, mux_tmp_3472, fsm_output[9]);
  assign mux_3494_itm = MUX_s_1_2_2(mux_3493_nl, mux_tmp_3453, fsm_output[10]);
  assign or_3116_nl = (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[8])) | (fsm_output[4])
      | (fsm_output[10]);
  assign or_3115_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[8]))
      | (fsm_output[4]) | (~ (fsm_output[10]));
  assign mux_3504_nl = MUX_s_1_2_2(or_3116_nl, or_3115_nl, fsm_output[2]);
  assign or_3117_nl = (fsm_output[9]) | mux_3504_nl;
  assign mux_3505_nl = MUX_s_1_2_2(or_3117_nl, or_70_cse, fsm_output[0]);
  assign nor_603_nl = ~((fsm_output[3]) | mux_3505_nl);
  assign and_376_nl = (fsm_output[0]) & (~ mux_tmp_2745);
  assign nor_604_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[8])
      | not_tmp_39);
  assign nor_605_nl = ~((fsm_output[2]) | (~ (fsm_output[1])) | (~ (fsm_output[6]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]));
  assign mux_3501_nl = MUX_s_1_2_2(nor_604_nl, nor_605_nl, fsm_output[9]);
  assign nor_606_nl = ~((~ (fsm_output[2])) | (fsm_output[1]) | (~ (fsm_output[6]))
      | (~ (fsm_output[8])) | (fsm_output[4]) | (~ (fsm_output[10])));
  assign nor_607_nl = ~((fsm_output[2]) | (~ (fsm_output[1])) | (fsm_output[6]) |
      (fsm_output[8]) | not_tmp_39);
  assign mux_3500_nl = MUX_s_1_2_2(nor_606_nl, nor_607_nl, fsm_output[9]);
  assign mux_3502_nl = MUX_s_1_2_2(mux_3501_nl, mux_3500_nl, fsm_output[0]);
  assign mux_3503_nl = MUX_s_1_2_2(and_376_nl, mux_3502_nl, fsm_output[3]);
  assign mux_3506_nl = MUX_s_1_2_2(nor_603_nl, mux_3503_nl, fsm_output[5]);
  assign or_3104_nl = (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[1]) | (~((fsm_output[6])
      & (fsm_output[8]) & (fsm_output[4]) & (fsm_output[10])));
  assign mux_3498_nl = MUX_s_1_2_2(or_3104_nl, or_56_cse, fsm_output[0]);
  assign or_3098_nl = (fsm_output[1]) | (fsm_output[6]) | (fsm_output[8]) | (~ (fsm_output[4]))
      | (fsm_output[10]);
  assign or_3097_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[8]) | not_tmp_39;
  assign mux_3495_nl = MUX_s_1_2_2(or_3098_nl, or_3097_nl, fsm_output[2]);
  assign or_3099_nl = (fsm_output[9]) | mux_3495_nl;
  assign mux_3497_nl = MUX_s_1_2_2(mux_tmp_2745, or_3099_nl, fsm_output[0]);
  assign mux_3499_nl = MUX_s_1_2_2(mux_3498_nl, mux_3497_nl, fsm_output[3]);
  assign nor_608_nl = ~((fsm_output[5]) | mux_3499_nl);
  assign not_tmp_688 = MUX_s_1_2_2(mux_3506_nl, nor_608_nl, fsm_output[7]);
  assign or_tmp_3053 = (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[2])) |
      (fsm_output[8]) | not_tmp_49;
  assign or_3154_nl = (fsm_output[8]) | nand_183_cse;
  assign mux_tmp_3529 = MUX_s_1_2_2(or_3154_nl, or_tmp_2774, fsm_output[3]);
  assign nor_584_nl = ~((fsm_output[5]) | (fsm_output[4]) | (~ (fsm_output[7])) |
      (fsm_output[3]) | (fsm_output[8]) | (fsm_output[1]) | (~ (fsm_output[6])) |
      (fsm_output[10]));
  assign nand_103_nl = ~((fsm_output[7]) & (~ mux_tmp_3529));
  assign or_3157_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[8]))
      | (fsm_output[1]) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_3532_nl = MUX_s_1_2_2(nand_103_nl, or_3157_nl, fsm_output[4]);
  assign nor_585_nl = ~((fsm_output[5]) | mux_3532_nl);
  assign mux_3533_nl = MUX_s_1_2_2(nor_584_nl, nor_585_nl, fsm_output[2]);
  assign nor_586_nl = ~((fsm_output[7]) | mux_tmp_3529);
  assign nor_587_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[8]))
      | (fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign mux_3530_nl = MUX_s_1_2_2(nor_586_nl, nor_587_nl, fsm_output[4]);
  assign and_371_nl = (fsm_output[5]) & mux_3530_nl;
  assign nor_588_nl = ~((fsm_output[5]) | (~ (fsm_output[4])) | (fsm_output[7]) |
      (~ (fsm_output[3])) | (fsm_output[8]) | (fsm_output[1]) | (~ (fsm_output[6]))
      | (fsm_output[10]));
  assign mux_3531_nl = MUX_s_1_2_2(and_371_nl, nor_588_nl, fsm_output[2]);
  assign mux_3534_nl = MUX_s_1_2_2(mux_3533_nl, mux_3531_nl, fsm_output[9]);
  assign nor_589_nl = ~((fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[1])) |
      (fsm_output[6]) | (fsm_output[10]));
  assign and_373_nl = (fsm_output[3]) & (fsm_output[8]) & (fsm_output[1]) & (fsm_output[6])
      & (fsm_output[10]);
  assign mux_3526_nl = MUX_s_1_2_2(nor_589_nl, and_373_nl, fsm_output[7]);
  assign and_372_nl = (fsm_output[5:4]==2'b11) & mux_3526_nl;
  assign nor_590_nl = ~((~ (fsm_output[4])) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (fsm_output[8]) | nand_183_cse);
  assign nor_591_nl = ~((fsm_output[7]) | mux_2998_cse);
  assign mux_3524_nl = MUX_s_1_2_2(nor_591_nl, nor_667_cse, fsm_output[4]);
  assign mux_3525_nl = MUX_s_1_2_2(nor_590_nl, mux_3524_nl, fsm_output[5]);
  assign mux_3527_nl = MUX_s_1_2_2(and_372_nl, mux_3525_nl, fsm_output[2]);
  assign or_3142_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[8]) | (~
      (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_3141_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[8]))
      | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_3522_nl = MUX_s_1_2_2(or_3142_nl, or_3141_nl, fsm_output[4]);
  assign nor_593_nl = ~((fsm_output[2]) | (fsm_output[5]) | mux_3522_nl);
  assign mux_3528_nl = MUX_s_1_2_2(mux_3527_nl, nor_593_nl, fsm_output[9]);
  assign not_tmp_701 = MUX_s_1_2_2(mux_3534_nl, mux_3528_nl, fsm_output[0]);
  assign or_tmp_3095 = (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[6]) |
      (fsm_output[8]) | (fsm_output[10]);
  assign or_3178_nl = (fsm_output[2]) | (fsm_output[4]);
  assign mux_tmp_3547 = MUX_s_1_2_2(or_2991_cse, mux_tmp_130, or_3178_nl);
  assign mux_tmp_3551 = MUX_s_1_2_2(mux_tmp_131, mux_155_cse, fsm_output[2]);
  assign mux_tmp_3574 = MUX_s_1_2_2(mux_375_cse, mux_340_cse, fsm_output[2]);
  assign mux_460_nl = MUX_s_1_2_2(mux_tmp_130, or_tmp_94, fsm_output[4]);
  assign mux_tmp_3576 = MUX_s_1_2_2(or_tmp_96, mux_460_nl, fsm_output[2]);
  assign mux_tmp_3577 = MUX_s_1_2_2(or_tmp_96, mux_375_cse, fsm_output[2]);
  assign or_3199_nl = (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_tmp_3618 = MUX_s_1_2_2(or_3199_nl, or_2835_cse, fsm_output[2]);
  assign or_tmp_3135 = (~ (fsm_output[2])) | (~ (fsm_output[1])) | (~ (fsm_output[8]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign or_3222_nl = (fsm_output[7]) | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[4])
      | (fsm_output[10]);
  assign or_3221_nl = (fsm_output[7]) | (~ (fsm_output[3])) | (fsm_output[8]) | not_tmp_39;
  assign mux_tmp_3632 = MUX_s_1_2_2(or_3222_nl, or_3221_nl, fsm_output[5]);
  assign or_tmp_3176 = (~ (fsm_output[4])) | (fsm_output[8]) | (~ (fsm_output[9]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign or_tmp_3190 = (fsm_output[1]) | (~ (fsm_output[2])) | (fsm_output[6]) |
      (~ (fsm_output[9]));
  assign mux_tmp_3673 = MUX_s_1_2_2(mux_tmp_215, mux_tmp_214, fsm_output[7]);
  assign mux_tmp_3674 = MUX_s_1_2_2(mux_tmp_215, or_tmp_114, fsm_output[7]);
  assign or_127_nl = (~((fsm_output[5]) | (~ (fsm_output[9])))) | (fsm_output[10]);
  assign mux_tmp_3679 = MUX_s_1_2_2(or_127_nl, nand_tmp_7, fsm_output[7]);
  assign mux_tmp_3681 = MUX_s_1_2_2(or_2414_cse, nand_tmp_7, fsm_output[7]);
  assign and_tmp_28 = (fsm_output[5]) & or_tmp_104;
  assign mux_tmp_3691 = MUX_s_1_2_2(and_tmp_28, or_361_cse, fsm_output[7]);
  assign or_tmp_3224 = (fsm_output[7]) | mux_tmp_231;
  assign or_134_nl = (fsm_output[5]) | mux_tmp_227;
  assign mux_tmp_3698 = MUX_s_1_2_2(mux_tmp_231, or_134_nl, fsm_output[7]);
  assign mux_262_nl = MUX_s_1_2_2(and_757_cse, (fsm_output[9]), fsm_output[5]);
  assign mux_tmp_3701 = MUX_s_1_2_2(mux_262_nl, or_tmp_114, fsm_output[7]);
  assign mux_tmp_3705 = MUX_s_1_2_2(mux_tmp_236, or_tmp_114, fsm_output[7]);
  assign mux_tmp_3720 = MUX_s_1_2_2((~ mux_tmp_214), mux_tmp_228, fsm_output[7]);
  assign mux_tmp_3724 = MUX_s_1_2_2((~ and_757_cse), mux_tmp_228, fsm_output[7]);
  assign mux_tmp_3736 = MUX_s_1_2_2(mux_tmp_227, or_361_cse, fsm_output[5]);
  assign mux_tmp_3737 = MUX_s_1_2_2(and_tmp_28, mux_tmp_3736, fsm_output[7]);
  assign mux_3738_nl = MUX_s_1_2_2(or_tmp_104, or_361_cse, fsm_output[5]);
  assign mux_tmp_3739 = MUX_s_1_2_2(and_tmp_28, mux_3738_nl, fsm_output[7]);
  assign mux_tmp_3753 = MUX_s_1_2_2(nor_tmp_23, or_tmp_114, fsm_output[7]);
  assign STAGE_LOOP_i_3_0_sva_mx0c1 = and_dcpl_103 & and_dcpl_98;
  assign VEC_LOOP_j_sva_11_0_mx0c1 = and_dcpl_103 & and_dcpl_48 & and_757_cse;
  assign nor_693_nl = ~((fsm_output[2]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[9])
      | (fsm_output[10]));
  assign mux_2654_nl = MUX_s_1_2_2(nor_694_cse, nor_693_nl, fsm_output[3]);
  assign and_467_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[7]) & (fsm_output[9])
      & (fsm_output[10]);
  assign mux_2653_nl = MUX_s_1_2_2(and_467_nl, and_756_cse, or_2644_cse);
  assign mux_2655_nl = MUX_s_1_2_2(mux_2654_nl, mux_2653_nl, fsm_output[5]);
  assign mux_2656_nl = MUX_s_1_2_2(mux_2655_nl, and_465_cse, fsm_output[4]);
  assign mux_2657_nl = MUX_s_1_2_2(mux_2656_nl, and_756_cse, fsm_output[6]);
  assign modExp_result_sva_mx0c0 = MUX_s_1_2_2(mux_2657_nl, and_757_cse, fsm_output[8]);
  assign nl_STAGE_LOOP_acc_nl = (STAGE_LOOP_i_3_0_sva_2[3:1]) + 3'b011;
  assign STAGE_LOOP_acc_nl = nl_STAGE_LOOP_acc_nl[2:0];
  assign STAGE_LOOP_acc_itm_2_1 = readslicef_3_1_2(STAGE_LOOP_acc_nl);
  assign and_279_m1c = and_dcpl_115 & and_dcpl_44 & and_dcpl_107;
  assign and_281_m1c = and_dcpl_260 & and_dcpl_88;
  assign and_284_m1c = and_dcpl_153 & and_dcpl_262 & and_dcpl_144;
  assign and_286_m1c = and_dcpl_147 & and_dcpl_152 & and_dcpl_235;
  assign and_288_m1c = and_dcpl_153 & and_dcpl_90 & and_dcpl_162;
  assign and_291_m1c = and_dcpl_270 & and_dcpl_55 & and_dcpl_33;
  assign and_292_m1c = and_dcpl_260 & and_dcpl_177;
  assign and_295_m1c = and_dcpl_6 & and_dcpl_262 & and_dcpl_48 & and_dcpl_33;
  assign and_297_m1c = and_dcpl_92 & and_dcpl_152 & and_dcpl_162;
  assign and_299_m1c = and_dcpl_278 & and_dcpl_224;
  assign and_302_m1c = and_dcpl_270 & and_dcpl_280 & and_dcpl_59;
  assign and_304_m1c = and_dcpl_118 & and_dcpl_136 & and_dcpl_208;
  assign and_307_m1c = and_dcpl_209 & and_dcpl_262 & and_dcpl_126 & and_dcpl_59;
  assign and_309_m1c = and_dcpl_118 & and_dcpl_152 & and_dcpl_224;
  assign and_311_m1c = and_dcpl_278 & and_dcpl_280 & and_757_cse;
  assign and_139_nl = and_dcpl_118 & and_dcpl_44 & and_dcpl_88;
  assign or_522_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[0]) | (~((fsm_output[1])
      & (fsm_output[6]) & (fsm_output[4]) & (fsm_output[8]) & (fsm_output[10])));
  assign or_520_nl = (fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[0]))
      | (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[4]) | nand_138_cse;
  assign mux_1091_nl = MUX_s_1_2_2(or_522_nl, or_520_nl, fsm_output[5]);
  assign or_518_nl = (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[4]) | nand_138_cse;
  assign mux_1089_nl = MUX_s_1_2_2(or_518_nl, mux_tmp_1082, fsm_output[7]);
  assign or_515_nl = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[4]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1087_nl = MUX_s_1_2_2(or_515_nl, or_tmp_453, fsm_output[0]);
  assign or_516_nl = (fsm_output[3]) | mux_1087_nl;
  assign or_513_nl = (~ (fsm_output[3])) | (fsm_output[0]) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1088_nl = MUX_s_1_2_2(or_516_nl, or_513_nl, fsm_output[7]);
  assign mux_1090_nl = MUX_s_1_2_2(mux_1089_nl, mux_1088_nl, fsm_output[5]);
  assign mux_1092_nl = MUX_s_1_2_2(mux_1091_nl, mux_1090_nl, fsm_output[2]);
  assign or_512_nl = (fsm_output[3]) | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[4]) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign or_511_nl = (~ (fsm_output[3])) | (fsm_output[0]) | (~ (fsm_output[1]))
      | (fsm_output[6]) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[10]);
  assign mux_1084_nl = MUX_s_1_2_2(or_512_nl, or_511_nl, fsm_output[7]);
  assign or_506_nl = (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6])
      | (fsm_output[4]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_1083_nl = MUX_s_1_2_2(mux_tmp_1082, or_506_nl, fsm_output[7]);
  assign mux_1085_nl = MUX_s_1_2_2(mux_1084_nl, mux_1083_nl, fsm_output[5]);
  assign or_504_nl = (fsm_output[5]) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (~ (fsm_output[0])) | (~ (fsm_output[1])) | (~ (fsm_output[6])) | (fsm_output[4])
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_1086_nl = MUX_s_1_2_2(mux_1085_nl, or_504_nl, fsm_output[2]);
  assign mux_1093_nl = MUX_s_1_2_2(mux_1092_nl, mux_1086_nl, fsm_output[9]);
  assign nor_1513_nl = ~((fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (fsm_output[5]));
  assign nor_1514_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (~((fsm_output[6:5]==2'b11))));
  assign mux_1094_nl = MUX_s_1_2_2(nor_1513_nl, nor_1514_nl, fsm_output[0]);
  assign and_144_nl = mux_1094_nl & (fsm_output[3]) & (~ (fsm_output[2])) & (fsm_output[7])
      & (~ (fsm_output[8])) & nor_609_cse;
  assign nor_1511_nl = ~((~ (fsm_output[8])) | (fsm_output[7]) | (fsm_output[2])
      | (fsm_output[5]) | (fsm_output[3]));
  assign nor_1512_nl = ~((fsm_output[8]) | (~((fsm_output[7]) & (fsm_output[2]) &
      (fsm_output[5]) & (fsm_output[3]))));
  assign mux_1095_nl = MUX_s_1_2_2(nor_1511_nl, nor_1512_nl, fsm_output[0]);
  assign and_153_nl = mux_1095_nl & (fsm_output[6]) & (fsm_output[4]) & (fsm_output[1])
      & nor_609_cse;
  assign nor_1509_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (~ (fsm_output[6]))
      | (fsm_output[7]) | (~ (fsm_output[2])) | (fsm_output[3]));
  assign nor_1510_nl = ~((fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[6])
      | (~ (fsm_output[7])) | (fsm_output[2]) | (~ (fsm_output[3])));
  assign mux_1096_nl = MUX_s_1_2_2(nor_1509_nl, nor_1510_nl, fsm_output[0]);
  assign and_162_nl = mux_1096_nl & and_707_cse & nor_609_cse;
  assign and_758_nl = (fsm_output[0]) & (fsm_output[6]) & (fsm_output[8]) & (fsm_output[7])
      & (fsm_output[2]) & (~ (fsm_output[5])) & (fsm_output[3]);
  assign nor_1508_nl = ~((fsm_output[0]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[7])
      | (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[3]));
  assign mux_1097_nl = MUX_s_1_2_2(and_758_nl, nor_1508_nl, fsm_output[9]);
  assign and_170_nl = mux_1097_nl & and_dcpl_34 & (~ (fsm_output[10]));
  assign nor_1505_nl = ~((fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[7])
      | (~ (fsm_output[5])));
  assign nor_1506_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (~ (fsm_output[7]))
      | (fsm_output[5]));
  assign mux_1098_nl = MUX_s_1_2_2(nor_1505_nl, nor_1506_nl, fsm_output[0]);
  assign and_180_nl = mux_1098_nl & (~ (fsm_output[3])) & (fsm_output[2]) & (~ (fsm_output[8]))
      & (~ (fsm_output[6])) & and_dcpl_33;
  assign nor_1503_nl = ~((fsm_output[4]) | (~((fsm_output[6]) & (fsm_output[2]) &
      (fsm_output[5]))));
  assign nor_1504_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | (fsm_output[2])
      | (fsm_output[5]));
  assign mux_1099_nl = MUX_s_1_2_2(nor_1503_nl, nor_1504_nl, fsm_output[0]);
  assign and_187_nl = mux_1099_nl & (fsm_output[3]) & and_dcpl_4 & (fsm_output[1])
      & and_dcpl_33;
  assign nor_1501_nl = ~((~ (fsm_output[1])) | (fsm_output[4]) | (fsm_output[6])
      | (fsm_output[2]));
  assign nor_1502_nl = ~((fsm_output[1]) | (~((fsm_output[4]) & (fsm_output[6]) &
      (fsm_output[2]))));
  assign mux_1100_nl = MUX_s_1_2_2(nor_1501_nl, nor_1502_nl, fsm_output[0]);
  assign and_195_nl = mux_1100_nl & (~ (fsm_output[3])) & nor_1580_cse & (fsm_output[8])
      & and_dcpl_33;
  assign nor_1499_nl = ~((~ (fsm_output[4])) | (fsm_output[6]) | (~((fsm_output[7])
      & (fsm_output[2]))));
  assign nor_1500_nl = ~((fsm_output[4]) | (~ (fsm_output[6])) | (fsm_output[7])
      | (fsm_output[2]));
  assign mux_1101_nl = MUX_s_1_2_2(nor_1499_nl, nor_1500_nl, fsm_output[0]);
  assign and_201_nl = mux_1101_nl & (fsm_output[3]) & and_707_cse & (~ (fsm_output[1]))
      & and_dcpl_33;
  assign or_3445_nl = (~ (fsm_output[9])) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[4])) | (~ (fsm_output[6])) | (~ (fsm_output[8])) | (~ (fsm_output[7]))
      | (fsm_output[5]);
  assign or_3446_nl = (fsm_output[9]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8]) | (fsm_output[7]) | (~
      (fsm_output[5]));
  assign mux_1102_nl = MUX_s_1_2_2(or_3445_nl, or_3446_nl, fsm_output[10]);
  assign nor_1625_nl = ~(mux_1102_nl | (fsm_output[3:2]!=2'b00));
  assign nor_1495_nl = ~((fsm_output[4]) | (~ (fsm_output[7])) | (fsm_output[2])
      | (fsm_output[5]) | (~ (fsm_output[3])));
  assign nor_1496_nl = ~((~ (fsm_output[4])) | (fsm_output[7]) | (~ (fsm_output[2]))
      | (~ (fsm_output[5])) | (fsm_output[3]));
  assign mux_1103_nl = MUX_s_1_2_2(nor_1495_nl, nor_1496_nl, fsm_output[0]);
  assign and_213_nl = mux_1103_nl & and_dcpl_191 & (fsm_output[1]) & and_dcpl_59;
  assign nor_1493_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[2]))
      | (fsm_output[5]) | (~ (fsm_output[3])));
  assign nor_1494_nl = ~((fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[2])
      | (~ (fsm_output[5])) | (fsm_output[3]));
  assign mux_1104_nl = MUX_s_1_2_2(nor_1493_nl, nor_1494_nl, fsm_output[0]);
  assign and_219_nl = mux_1104_nl & and_dcpl_4 & (fsm_output[4]) & and_dcpl_59;
  assign and_760_nl = (fsm_output[4]) & (fsm_output[6]) & (~ (fsm_output[2])) & (fsm_output[3]);
  assign nor_1492_nl = ~((fsm_output[4]) | (fsm_output[6]) | (~ (fsm_output[2]))
      | (fsm_output[3]));
  assign mux_1105_nl = MUX_s_1_2_2(and_760_nl, nor_1492_nl, fsm_output[0]);
  assign and_225_nl = mux_1105_nl & (~ (fsm_output[5])) & and_dcpl_135 & (~ (fsm_output[1]))
      & and_dcpl_59;
  assign nor_1489_nl = ~((fsm_output[1]) | (fsm_output[4]) | (~ (fsm_output[6]))
      | (fsm_output[7]));
  assign and_748_nl = (fsm_output[1]) & (fsm_output[4]) & (~ (fsm_output[6])) & (fsm_output[7]);
  assign mux_1106_nl = MUX_s_1_2_2(nor_1489_nl, and_748_nl, fsm_output[0]);
  assign and_235_nl = mux_1106_nl & (fsm_output[3]) & and_676_cse & (fsm_output[8])
      & and_dcpl_59;
  assign and_627_nl = (fsm_output[0]) & (fsm_output[4]) & (fsm_output[6]) & (fsm_output[8])
      & (fsm_output[7]) & (~ (fsm_output[2])) & (~ (fsm_output[5]));
  assign nor_1488_nl = ~((fsm_output[0]) | (fsm_output[4]) | (fsm_output[6]) | (fsm_output[8])
      | (fsm_output[7]) | (~ and_676_cse));
  assign mux_1107_nl = MUX_s_1_2_2(and_627_nl, nor_1488_nl, fsm_output[9]);
  assign and_241_nl = mux_1107_nl & (~ (fsm_output[3])) & (fsm_output[1]) & (fsm_output[10]);
  assign nor_1486_nl = ~((~ (fsm_output[1])) | (~ (fsm_output[4])) | (fsm_output[7])
      | (fsm_output[2]) | (~ (fsm_output[5])));
  assign nor_1487_nl = ~((fsm_output[1]) | (fsm_output[4]) | (~ (fsm_output[7]))
      | (~ (fsm_output[2])) | (fsm_output[5]));
  assign mux_1108_nl = MUX_s_1_2_2(nor_1486_nl, nor_1487_nl, fsm_output[0]);
  assign and_249_nl = mux_1108_nl & (fsm_output[3]) & (~ (fsm_output[8])) & (~ (fsm_output[6]))
      & and_757_cse;
  assign vec_rsc_0_0_i_adra_d_pff = MUX1HOT_v_8_19_2(COMP_LOOP_acc_psp_sva_1, (z_out_2_12_1[11:4]),
      COMP_LOOP_acc_psp_sva, (COMP_LOOP_acc_10_cse_12_1_1_sva[11:4]), (COMP_LOOP_acc_1_cse_2_sva[11:4]),
      (COMP_LOOP_acc_11_psp_sva[10:3]), (COMP_LOOP_acc_1_cse_4_sva[11:4]), (COMP_LOOP_acc_13_psp_sva[9:2]),
      (COMP_LOOP_acc_1_cse_6_sva[11:4]), (COMP_LOOP_acc_14_psp_sva[10:3]), (COMP_LOOP_acc_1_cse_8_sva[11:4]),
      (COMP_LOOP_acc_16_psp_sva[8:1]), (COMP_LOOP_acc_1_cse_10_sva[11:4]), (COMP_LOOP_acc_17_psp_sva[10:3]),
      (COMP_LOOP_acc_1_cse_12_sva[11:4]), (COMP_LOOP_acc_19_psp_sva[9:2]), (COMP_LOOP_acc_1_cse_14_sva[11:4]),
      (COMP_LOOP_acc_20_psp_sva[10:3]), (COMP_LOOP_acc_1_cse_sva[11:4]), {and_dcpl_109
      , COMP_LOOP_or_32_cse , and_139_nl , (~ mux_1093_nl) , and_144_nl , and_153_nl
      , and_162_nl , and_170_nl , and_180_nl , and_187_nl , and_195_nl , and_201_nl
      , nor_1625_nl , and_213_nl , and_219_nl , and_225_nl , and_235_nl , and_241_nl
      , and_249_nl});
  assign vec_rsc_0_0_i_da_d_pff = COMP_LOOP_10_mul_mut;
  assign or_618_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_617_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (~ (fsm_output[10]));
  assign mux_1134_nl = MUX_s_1_2_2(or_618_nl, or_617_nl, fsm_output[7]);
  assign or_615_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b00) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1135_nl = MUX_s_1_2_2(mux_1134_nl, or_615_nl, fsm_output[2]);
  assign nor_1471_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1135_nl);
  assign nor_1472_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (~ (fsm_output[10])));
  assign mux_1136_nl = MUX_s_1_2_2(nor_1471_nl, nor_1472_nl, fsm_output[8]);
  assign nor_1473_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1474_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (fsm_output[10]));
  assign nor_1475_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (fsm_output[10]));
  assign nor_1476_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1131_nl = MUX_s_1_2_2(nor_1475_nl, nor_1476_nl, fsm_output[4]);
  assign mux_1132_nl = MUX_s_1_2_2(nor_1474_nl, mux_1131_nl, fsm_output[6]);
  assign mux_1133_nl = MUX_s_1_2_2(nor_1473_nl, mux_1132_nl, fsm_output[8]);
  assign mux_1137_nl = MUX_s_1_2_2(mux_1136_nl, mux_1133_nl, fsm_output[0]);
  assign or_606_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (VEC_LOOP_j_sva_11_0[2]) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_605_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[2]) | (fsm_output[7])
      | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[9]) | (fsm_output[5]) | (~
      (fsm_output[10]));
  assign mux_1128_nl = MUX_s_1_2_2(mux_tmp_1116, or_605_nl, fsm_output[4]);
  assign mux_1129_nl = MUX_s_1_2_2(or_606_nl, mux_1128_nl, fsm_output[6]);
  assign and_626_nl = (fsm_output[8]) & (~ mux_1129_nl);
  assign or_602_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_600_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (~ (fsm_output[10]));
  assign mux_1125_nl = MUX_s_1_2_2(or_600_nl, or_tmp_532, fsm_output[2]);
  assign mux_1126_nl = MUX_s_1_2_2(or_602_nl, mux_1125_nl, fsm_output[4]);
  assign nor_1477_nl = ~((fsm_output[6]) | mux_1126_nl);
  assign nor_1478_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1127_nl = MUX_s_1_2_2(nor_1477_nl, nor_1478_nl, fsm_output[8]);
  assign mux_1130_nl = MUX_s_1_2_2(and_626_nl, mux_1127_nl, fsm_output[0]);
  assign mux_1138_nl = MUX_s_1_2_2(mux_1137_nl, mux_1130_nl, fsm_output[3]);
  assign or_596_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[0]) | nand_337_cse;
  assign or_594_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (~ (fsm_output[10]));
  assign mux_1121_nl = MUX_s_1_2_2(or_596_nl, or_594_nl, fsm_output[4]);
  assign nor_1479_nl = ~((fsm_output[6]) | mux_1121_nl);
  assign or_590_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (~ (fsm_output[10]));
  assign mux_1119_nl = MUX_s_1_2_2(or_591_cse, or_590_nl, fsm_output[7]);
  assign mux_1120_nl = MUX_s_1_2_2(mux_1119_nl, or_tmp_532, or_586_cse);
  assign nor_1480_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1120_nl);
  assign mux_1122_nl = MUX_s_1_2_2(nor_1479_nl, nor_1480_nl, fsm_output[8]);
  assign or_583_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_581_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1117_nl = MUX_s_1_2_2(or_583_nl, or_581_nl, fsm_output[2]);
  assign mux_1118_nl = MUX_s_1_2_2(mux_1117_nl, mux_tmp_1116, fsm_output[4]);
  assign nor_1481_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1118_nl);
  assign mux_1123_nl = MUX_s_1_2_2(mux_1122_nl, nor_1481_nl, fsm_output[0]);
  assign or_576_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_574_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (fsm_output[10]);
  assign mux_1113_nl = MUX_s_1_2_2(or_576_nl, or_574_nl, fsm_output[4]);
  assign or_573_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9])) | (~
      (fsm_output[5])) | (fsm_output[10]);
  assign or_572_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (fsm_output[10]);
  assign mux_1112_nl = MUX_s_1_2_2(or_573_nl, or_572_nl, fsm_output[4]);
  assign mux_1114_nl = MUX_s_1_2_2(mux_1113_nl, mux_1112_nl, fsm_output[6]);
  assign nor_1482_nl = ~((fsm_output[8]) | mux_1114_nl);
  assign nor_1483_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1484_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (fsm_output[9]) | not_tmp_248);
  assign or_567_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000)
      | (~ (fsm_output[10]));
  assign or_565_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0000) | (fsm_output[10]);
  assign mux_1109_nl = MUX_s_1_2_2(or_567_nl, or_565_nl, fsm_output[2]);
  assign nor_1485_nl = ~((fsm_output[4]) | mux_1109_nl);
  assign mux_1110_nl = MUX_s_1_2_2(nor_1484_nl, nor_1485_nl, fsm_output[6]);
  assign mux_1111_nl = MUX_s_1_2_2(nor_1483_nl, mux_1110_nl, fsm_output[8]);
  assign mux_1115_nl = MUX_s_1_2_2(nor_1482_nl, mux_1111_nl, fsm_output[0]);
  assign mux_1124_nl = MUX_s_1_2_2(mux_1123_nl, mux_1115_nl, fsm_output[3]);
  assign vec_rsc_0_0_i_wea_d_pff = MUX_s_1_2_2(mux_1138_nl, mux_1124_nl, fsm_output[1]);
  assign or_674_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0000) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_673_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0000) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1169_nl = MUX_s_1_2_2(or_674_nl, or_673_nl, fsm_output[5]);
  assign nor_1440_nl = ~((fsm_output[1]) | mux_1169_nl);
  assign nor_1441_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0000)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1442_nl = ~((z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1443_nl = ~((z_out_2_12_1[3:0]!=4'b0000) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1167_nl = MUX_s_1_2_2(nor_1442_nl, nor_1443_nl, fsm_output[5]);
  assign mux_1168_nl = MUX_s_1_2_2(nor_1441_nl, mux_1167_nl, fsm_output[1]);
  assign mux_1170_nl = MUX_s_1_2_2(nor_1440_nl, mux_1168_nl, fsm_output[0]);
  assign and_623_nl = (fsm_output[6]) & mux_1170_nl;
  assign nor_1444_nl = ~((z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1446_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1162_nl = MUX_s_1_2_2(nor_1445_cse, nor_1446_nl, fsm_output[5]);
  assign nor_1447_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_660_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1163_nl = MUX_s_1_2_2(mux_1162_nl, nor_1447_nl, or_660_nl);
  assign mux_1164_nl = MUX_s_1_2_2(nor_1444_nl, mux_1163_nl, fsm_output[1]);
  assign nor_1448_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1449_nl = ~((z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1450_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1160_nl = MUX_s_1_2_2(nor_1449_nl, nor_1450_nl, fsm_output[5]);
  assign mux_1161_nl = MUX_s_1_2_2(nor_1448_nl, mux_1160_nl, fsm_output[1]);
  assign mux_1165_nl = MUX_s_1_2_2(mux_1164_nl, mux_1161_nl, fsm_output[0]);
  assign nor_1451_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0000) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1452_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0000) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1158_nl = MUX_s_1_2_2(nor_1451_nl, nor_1452_nl, fsm_output[1]);
  assign nor_1453_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1157_cse);
  assign mux_1159_nl = MUX_s_1_2_2(mux_1158_nl, nor_1453_nl, fsm_output[0]);
  assign mux_1166_nl = MUX_s_1_2_2(mux_1165_nl, mux_1159_nl, fsm_output[6]);
  assign mux_1171_nl = MUX_s_1_2_2(and_623_nl, mux_1166_nl, fsm_output[8]);
  assign nor_1454_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0000) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1455_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0000) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1152_nl = MUX_s_1_2_2(nor_1454_nl, nor_1455_nl, fsm_output[5]);
  assign and_624_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1152_nl;
  assign nor_1456_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1457_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0000) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1151_nl = MUX_s_1_2_2(nor_1456_nl, nor_1457_nl, fsm_output[5]);
  assign and_625_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1151_nl;
  assign mux_1153_nl = MUX_s_1_2_2(and_624_nl, and_625_nl, fsm_output[1]);
  assign nor_1458_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (VEC_LOOP_j_sva_11_0[1]) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2]) | (fsm_output[7]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1459_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1149_cse);
  assign mux_1150_nl = MUX_s_1_2_2(nor_1458_nl, nor_1459_nl, fsm_output[1]);
  assign mux_1154_nl = MUX_s_1_2_2(mux_1153_nl, mux_1150_nl, fsm_output[0]);
  assign nor_1460_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1461_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1462_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1147_nl = MUX_s_1_2_2(nor_1461_nl, nor_1462_nl, fsm_output[1]);
  assign mux_1148_nl = MUX_s_1_2_2(nor_1460_nl, mux_1147_nl, fsm_output[0]);
  assign mux_1155_nl = MUX_s_1_2_2(mux_1154_nl, mux_1148_nl, fsm_output[6]);
  assign nor_1463_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0000) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1464_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0000)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1145_nl = MUX_s_1_2_2(nor_1463_nl, nor_1464_nl, fsm_output[0]);
  assign nor_1465_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1466_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0000)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1467_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0000) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1141_nl = MUX_s_1_2_2(nor_1466_nl, nor_1467_nl, fsm_output[5]);
  assign mux_1142_nl = MUX_s_1_2_2(nor_1465_nl, mux_1141_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1468_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0000)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1143_nl = MUX_s_1_2_2(mux_1142_nl, nor_1468_nl, fsm_output[1]);
  assign nor_1469_nl = ~((z_out_2_12_1[3:0]!=4'b0000) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1470_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1140_nl = MUX_s_1_2_2(nor_1469_nl, nor_1470_nl, fsm_output[1]);
  assign mux_1144_nl = MUX_s_1_2_2(mux_1143_nl, mux_1140_nl, fsm_output[0]);
  assign mux_1146_nl = MUX_s_1_2_2(mux_1145_nl, mux_1144_nl, fsm_output[6]);
  assign mux_1156_nl = MUX_s_1_2_2(mux_1155_nl, mux_1146_nl, fsm_output[8]);
  assign vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1171_nl,
      mux_1156_nl, fsm_output[4]);
  assign or_729_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_728_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (~ (fsm_output[10]));
  assign mux_1198_nl = MUX_s_1_2_2(or_729_nl, or_728_nl, fsm_output[7]);
  assign or_726_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b00) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1199_nl = MUX_s_1_2_2(mux_1198_nl, or_726_nl, fsm_output[2]);
  assign nor_1425_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1199_nl);
  assign nor_1426_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (~ (fsm_output[10])));
  assign mux_1200_nl = MUX_s_1_2_2(nor_1425_nl, nor_1426_nl, fsm_output[8]);
  assign nor_1427_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1428_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (fsm_output[10]));
  assign nor_1429_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (fsm_output[10]));
  assign nor_1430_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1195_nl = MUX_s_1_2_2(nor_1429_nl, nor_1430_nl, fsm_output[4]);
  assign mux_1196_nl = MUX_s_1_2_2(nor_1428_nl, mux_1195_nl, fsm_output[6]);
  assign mux_1197_nl = MUX_s_1_2_2(nor_1427_nl, mux_1196_nl, fsm_output[8]);
  assign mux_1201_nl = MUX_s_1_2_2(mux_1200_nl, mux_1197_nl, fsm_output[0]);
  assign or_717_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (VEC_LOOP_j_sva_11_0[2]) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_716_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[2]) | (fsm_output[7])
      | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[9]) | (fsm_output[5]) | (~
      (fsm_output[10]));
  assign mux_1192_nl = MUX_s_1_2_2(mux_tmp_1180, or_716_nl, fsm_output[4]);
  assign mux_1193_nl = MUX_s_1_2_2(or_717_nl, mux_1192_nl, fsm_output[6]);
  assign and_622_nl = (fsm_output[8]) & (~ mux_1193_nl);
  assign or_713_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_711_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (~ (fsm_output[10]));
  assign mux_1189_nl = MUX_s_1_2_2(or_711_nl, or_tmp_643, fsm_output[2]);
  assign mux_1190_nl = MUX_s_1_2_2(or_713_nl, mux_1189_nl, fsm_output[4]);
  assign nor_1431_nl = ~((fsm_output[6]) | mux_1190_nl);
  assign nor_1432_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1191_nl = MUX_s_1_2_2(nor_1431_nl, nor_1432_nl, fsm_output[8]);
  assign mux_1194_nl = MUX_s_1_2_2(and_622_nl, mux_1191_nl, fsm_output[0]);
  assign mux_1202_nl = MUX_s_1_2_2(mux_1201_nl, mux_1194_nl, fsm_output[3]);
  assign or_707_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_705_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (~ (fsm_output[10]));
  assign mux_1185_nl = MUX_s_1_2_2(or_707_nl, or_705_nl, fsm_output[4]);
  assign nor_1433_nl = ~((fsm_output[6]) | mux_1185_nl);
  assign or_701_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (~ (fsm_output[10]));
  assign mux_1183_nl = MUX_s_1_2_2(or_702_cse, or_701_nl, fsm_output[7]);
  assign mux_1184_nl = MUX_s_1_2_2(mux_1183_nl, or_tmp_643, or_586_cse);
  assign nor_1434_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1184_nl);
  assign mux_1186_nl = MUX_s_1_2_2(nor_1433_nl, nor_1434_nl, fsm_output[8]);
  assign or_694_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_692_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1181_nl = MUX_s_1_2_2(or_694_nl, or_692_nl, fsm_output[2]);
  assign mux_1182_nl = MUX_s_1_2_2(mux_1181_nl, mux_tmp_1180, fsm_output[4]);
  assign nor_1435_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1182_nl);
  assign mux_1187_nl = MUX_s_1_2_2(mux_1186_nl, nor_1435_nl, fsm_output[0]);
  assign or_687_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b000) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_685_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (fsm_output[10]);
  assign mux_1177_nl = MUX_s_1_2_2(or_687_nl, or_685_nl, fsm_output[4]);
  assign or_684_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b000) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_683_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (fsm_output[10]);
  assign mux_1176_nl = MUX_s_1_2_2(or_684_nl, or_683_nl, fsm_output[4]);
  assign mux_1178_nl = MUX_s_1_2_2(mux_1177_nl, mux_1176_nl, fsm_output[6]);
  assign nor_1436_nl = ~((fsm_output[8]) | mux_1178_nl);
  assign nor_1437_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1438_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (fsm_output[9]) | not_tmp_248);
  assign or_678_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001)
      | (~ (fsm_output[10]));
  assign or_676_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0001) | (fsm_output[10]);
  assign mux_1173_nl = MUX_s_1_2_2(or_678_nl, or_676_nl, fsm_output[2]);
  assign nor_1439_nl = ~((fsm_output[4]) | mux_1173_nl);
  assign mux_1174_nl = MUX_s_1_2_2(nor_1438_nl, nor_1439_nl, fsm_output[6]);
  assign mux_1175_nl = MUX_s_1_2_2(nor_1437_nl, mux_1174_nl, fsm_output[8]);
  assign mux_1179_nl = MUX_s_1_2_2(nor_1436_nl, mux_1175_nl, fsm_output[0]);
  assign mux_1188_nl = MUX_s_1_2_2(mux_1187_nl, mux_1179_nl, fsm_output[3]);
  assign vec_rsc_0_1_i_wea_d_pff = MUX_s_1_2_2(mux_1202_nl, mux_1188_nl, fsm_output[1]);
  assign or_785_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0001) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_784_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0001) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1233_nl = MUX_s_1_2_2(or_785_nl, or_784_nl, fsm_output[5]);
  assign nor_1394_nl = ~((fsm_output[1]) | mux_1233_nl);
  assign nor_1395_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0001)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1396_nl = ~((z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1397_nl = ~((z_out_2_12_1[3:0]!=4'b0001) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1231_nl = MUX_s_1_2_2(nor_1396_nl, nor_1397_nl, fsm_output[5]);
  assign mux_1232_nl = MUX_s_1_2_2(nor_1395_nl, mux_1231_nl, fsm_output[1]);
  assign mux_1234_nl = MUX_s_1_2_2(nor_1394_nl, mux_1232_nl, fsm_output[0]);
  assign and_619_nl = (fsm_output[6]) & mux_1234_nl;
  assign nor_1398_nl = ~((z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1400_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1226_nl = MUX_s_1_2_2(nor_1445_cse, nor_1400_nl, fsm_output[5]);
  assign nor_1401_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_771_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1227_nl = MUX_s_1_2_2(mux_1226_nl, nor_1401_nl, or_771_nl);
  assign mux_1228_nl = MUX_s_1_2_2(nor_1398_nl, mux_1227_nl, fsm_output[1]);
  assign nor_1402_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1403_nl = ~((z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1404_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1224_nl = MUX_s_1_2_2(nor_1403_nl, nor_1404_nl, fsm_output[5]);
  assign mux_1225_nl = MUX_s_1_2_2(nor_1402_nl, mux_1224_nl, fsm_output[1]);
  assign mux_1229_nl = MUX_s_1_2_2(mux_1228_nl, mux_1225_nl, fsm_output[0]);
  assign nor_1405_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0001) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1406_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0001) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1222_nl = MUX_s_1_2_2(nor_1405_nl, nor_1406_nl, fsm_output[1]);
  assign nor_1407_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1157_cse);
  assign mux_1223_nl = MUX_s_1_2_2(mux_1222_nl, nor_1407_nl, fsm_output[0]);
  assign mux_1230_nl = MUX_s_1_2_2(mux_1229_nl, mux_1223_nl, fsm_output[6]);
  assign mux_1235_nl = MUX_s_1_2_2(and_619_nl, mux_1230_nl, fsm_output[8]);
  assign nor_1408_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0001) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1409_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0001) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1216_nl = MUX_s_1_2_2(nor_1408_nl, nor_1409_nl, fsm_output[5]);
  assign and_620_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1216_nl;
  assign nor_1410_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1411_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0001) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1215_nl = MUX_s_1_2_2(nor_1410_nl, nor_1411_nl, fsm_output[5]);
  assign and_621_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1215_nl;
  assign mux_1217_nl = MUX_s_1_2_2(and_620_nl, and_621_nl, fsm_output[1]);
  assign nor_1412_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (VEC_LOOP_j_sva_11_0[1]) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1413_nl = ~(nand_332_cse | mux_1149_cse);
  assign mux_1214_nl = MUX_s_1_2_2(nor_1412_nl, nor_1413_nl, fsm_output[1]);
  assign mux_1218_nl = MUX_s_1_2_2(mux_1217_nl, mux_1214_nl, fsm_output[0]);
  assign nor_1414_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1415_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1416_nl = ~((~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b000) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1211_nl = MUX_s_1_2_2(nor_1415_nl, nor_1416_nl, fsm_output[1]);
  assign mux_1212_nl = MUX_s_1_2_2(nor_1414_nl, mux_1211_nl, fsm_output[0]);
  assign mux_1219_nl = MUX_s_1_2_2(mux_1218_nl, mux_1212_nl, fsm_output[6]);
  assign nor_1417_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0001) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1418_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0001)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1209_nl = MUX_s_1_2_2(nor_1417_nl, nor_1418_nl, fsm_output[0]);
  assign nor_1419_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1420_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0001)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1421_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0001) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1205_nl = MUX_s_1_2_2(nor_1420_nl, nor_1421_nl, fsm_output[5]);
  assign mux_1206_nl = MUX_s_1_2_2(nor_1419_nl, mux_1205_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1422_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0001)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1207_nl = MUX_s_1_2_2(mux_1206_nl, nor_1422_nl, fsm_output[1]);
  assign nor_1423_nl = ~((z_out_2_12_1[3:0]!=4'b0001) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1424_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b000) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1204_nl = MUX_s_1_2_2(nor_1423_nl, nor_1424_nl, fsm_output[1]);
  assign mux_1208_nl = MUX_s_1_2_2(mux_1207_nl, mux_1204_nl, fsm_output[0]);
  assign mux_1210_nl = MUX_s_1_2_2(mux_1209_nl, mux_1208_nl, fsm_output[6]);
  assign mux_1220_nl = MUX_s_1_2_2(mux_1219_nl, mux_1210_nl, fsm_output[8]);
  assign vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1235_nl,
      mux_1220_nl, fsm_output[4]);
  assign or_839_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b01);
  assign or_838_nl = (~ (fsm_output[5])) | (~ (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010)
      | (~ (fsm_output[10]));
  assign mux_1262_nl = MUX_s_1_2_2(or_839_nl, or_838_nl, fsm_output[7]);
  assign or_836_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b00) | (~ (fsm_output[7])) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[5]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b00);
  assign mux_1263_nl = MUX_s_1_2_2(mux_1262_nl, or_836_nl, fsm_output[2]);
  assign nor_1379_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1263_nl);
  assign nor_1380_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010)
      | (~ (fsm_output[10])));
  assign mux_1264_nl = MUX_s_1_2_2(nor_1379_nl, nor_1380_nl, fsm_output[8]);
  assign nor_1381_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (~ (fsm_output[10])));
  assign nor_1382_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[5])
      | (~ (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (fsm_output[10]));
  assign nor_1383_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (fsm_output[10]));
  assign nor_1384_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[10]));
  assign mux_1259_nl = MUX_s_1_2_2(nor_1383_nl, nor_1384_nl, fsm_output[4]);
  assign mux_1260_nl = MUX_s_1_2_2(nor_1382_nl, mux_1259_nl, fsm_output[6]);
  assign mux_1261_nl = MUX_s_1_2_2(nor_1381_nl, mux_1260_nl, fsm_output[8]);
  assign mux_1265_nl = MUX_s_1_2_2(mux_1264_nl, mux_1261_nl, fsm_output[0]);
  assign or_827_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (VEC_LOOP_j_sva_11_0[2]) | (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b01);
  assign or_826_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[2]) | (fsm_output[7])
      | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[5]) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[10:9]!=2'b10);
  assign mux_1256_nl = MUX_s_1_2_2(mux_tmp_1244, or_826_nl, fsm_output[4]);
  assign mux_1257_nl = MUX_s_1_2_2(or_827_nl, mux_1256_nl, fsm_output[6]);
  assign and_618_nl = (fsm_output[8]) & (~ mux_1257_nl);
  assign or_823_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[5]) | nand_358_cse;
  assign or_821_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (~ (fsm_output[10]));
  assign mux_1253_nl = MUX_s_1_2_2(or_821_nl, or_tmp_756, fsm_output[2]);
  assign mux_1254_nl = MUX_s_1_2_2(or_823_nl, mux_1253_nl, fsm_output[4]);
  assign nor_1385_nl = ~((fsm_output[6]) | mux_1254_nl);
  assign nor_1386_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[10]));
  assign mux_1255_nl = MUX_s_1_2_2(nor_1385_nl, nor_1386_nl, fsm_output[8]);
  assign mux_1258_nl = MUX_s_1_2_2(and_618_nl, mux_1255_nl, fsm_output[0]);
  assign mux_1266_nl = MUX_s_1_2_2(mux_1265_nl, mux_1258_nl, fsm_output[3]);
  assign or_817_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | nand_358_cse;
  assign or_815_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (~ (fsm_output[10]));
  assign mux_1249_nl = MUX_s_1_2_2(or_817_nl, or_815_nl, fsm_output[4]);
  assign nor_1387_nl = ~((fsm_output[6]) | mux_1249_nl);
  assign or_809_nl = (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010)
      | (~ (fsm_output[10]));
  assign mux_1247_nl = MUX_s_1_2_2(or_591_cse, or_809_nl, fsm_output[7]);
  assign mux_1248_nl = MUX_s_1_2_2(or_tmp_756, mux_1247_nl, nor_209_cse);
  assign nor_1388_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1248_nl);
  assign mux_1250_nl = MUX_s_1_2_2(nor_1387_nl, nor_1388_nl, fsm_output[8]);
  assign or_805_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010) | (fsm_output[7])
      | (~ (fsm_output[5])) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign or_803_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (~ (fsm_output[7]))
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign mux_1245_nl = MUX_s_1_2_2(or_805_nl, or_803_nl, fsm_output[2]);
  assign mux_1246_nl = MUX_s_1_2_2(mux_1245_nl, mux_tmp_1244, fsm_output[4]);
  assign nor_1389_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1246_nl);
  assign mux_1251_nl = MUX_s_1_2_2(mux_1250_nl, nor_1389_nl, fsm_output[0]);
  assign or_798_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (fsm_output[5]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b10);
  assign or_796_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[5]) | (~
      (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (fsm_output[10]);
  assign mux_1241_nl = MUX_s_1_2_2(or_798_nl, or_796_nl, fsm_output[4]);
  assign or_795_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b01);
  assign or_794_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (fsm_output[10]);
  assign mux_1240_nl = MUX_s_1_2_2(or_795_nl, or_794_nl, fsm_output[4]);
  assign mux_1242_nl = MUX_s_1_2_2(mux_1241_nl, mux_1240_nl, fsm_output[6]);
  assign nor_1390_nl = ~((fsm_output[8]) | mux_1242_nl);
  assign nor_1391_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[10]));
  assign nor_1392_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (~ (fsm_output[5])) | (fsm_output[9])
      | (~ (fsm_output[10])));
  assign or_789_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010)
      | (~ (fsm_output[10]));
  assign or_787_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0010) | (fsm_output[10]);
  assign mux_1237_nl = MUX_s_1_2_2(or_789_nl, or_787_nl, fsm_output[2]);
  assign nor_1393_nl = ~((fsm_output[4]) | mux_1237_nl);
  assign mux_1238_nl = MUX_s_1_2_2(nor_1392_nl, nor_1393_nl, fsm_output[6]);
  assign mux_1239_nl = MUX_s_1_2_2(nor_1391_nl, mux_1238_nl, fsm_output[8]);
  assign mux_1243_nl = MUX_s_1_2_2(nor_1390_nl, mux_1239_nl, fsm_output[0]);
  assign mux_1252_nl = MUX_s_1_2_2(mux_1251_nl, mux_1243_nl, fsm_output[3]);
  assign vec_rsc_0_2_i_wea_d_pff = MUX_s_1_2_2(mux_1266_nl, mux_1252_nl, fsm_output[1]);
  assign or_895_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0010) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_894_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0010) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1297_nl = MUX_s_1_2_2(or_895_nl, or_894_nl, fsm_output[5]);
  assign nor_1348_nl = ~((fsm_output[1]) | mux_1297_nl);
  assign nor_1349_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0010)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1350_nl = ~((z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1351_nl = ~((z_out_2_12_1[3:0]!=4'b0010) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1295_nl = MUX_s_1_2_2(nor_1350_nl, nor_1351_nl, fsm_output[5]);
  assign mux_1296_nl = MUX_s_1_2_2(nor_1349_nl, mux_1295_nl, fsm_output[1]);
  assign mux_1298_nl = MUX_s_1_2_2(nor_1348_nl, mux_1296_nl, fsm_output[0]);
  assign and_615_nl = (fsm_output[6]) & mux_1298_nl;
  assign nor_1352_nl = ~((z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1354_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1290_nl = MUX_s_1_2_2(nor_1445_cse, nor_1354_nl, fsm_output[5]);
  assign nor_1355_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_881_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1291_nl = MUX_s_1_2_2(mux_1290_nl, nor_1355_nl, or_881_nl);
  assign mux_1292_nl = MUX_s_1_2_2(nor_1352_nl, mux_1291_nl, fsm_output[1]);
  assign nor_1356_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1357_nl = ~((z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1358_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1288_nl = MUX_s_1_2_2(nor_1357_nl, nor_1358_nl, fsm_output[5]);
  assign mux_1289_nl = MUX_s_1_2_2(nor_1356_nl, mux_1288_nl, fsm_output[1]);
  assign mux_1293_nl = MUX_s_1_2_2(mux_1292_nl, mux_1289_nl, fsm_output[0]);
  assign nor_1359_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0010) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1360_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0010) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1286_nl = MUX_s_1_2_2(nor_1359_nl, nor_1360_nl, fsm_output[1]);
  assign nor_1361_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1157_cse);
  assign mux_1287_nl = MUX_s_1_2_2(mux_1286_nl, nor_1361_nl, fsm_output[0]);
  assign mux_1294_nl = MUX_s_1_2_2(mux_1293_nl, mux_1287_nl, fsm_output[6]);
  assign mux_1299_nl = MUX_s_1_2_2(and_615_nl, mux_1294_nl, fsm_output[8]);
  assign nor_1362_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0010) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1363_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0010) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1280_nl = MUX_s_1_2_2(nor_1362_nl, nor_1363_nl, fsm_output[5]);
  assign and_616_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1280_nl;
  assign nor_1364_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1365_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0010) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1279_nl = MUX_s_1_2_2(nor_1364_nl, nor_1365_nl, fsm_output[5]);
  assign and_617_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1279_nl;
  assign mux_1281_nl = MUX_s_1_2_2(and_616_nl, and_617_nl, fsm_output[1]);
  assign nor_1366_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1367_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1277_cse);
  assign mux_1278_nl = MUX_s_1_2_2(nor_1366_nl, nor_1367_nl, fsm_output[1]);
  assign mux_1282_nl = MUX_s_1_2_2(mux_1281_nl, mux_1278_nl, fsm_output[0]);
  assign nor_1368_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1369_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1370_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1275_nl = MUX_s_1_2_2(nor_1369_nl, nor_1370_nl, fsm_output[1]);
  assign mux_1276_nl = MUX_s_1_2_2(nor_1368_nl, mux_1275_nl, fsm_output[0]);
  assign mux_1283_nl = MUX_s_1_2_2(mux_1282_nl, mux_1276_nl, fsm_output[6]);
  assign nor_1371_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0010) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1372_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0010)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1273_nl = MUX_s_1_2_2(nor_1371_nl, nor_1372_nl, fsm_output[0]);
  assign nor_1373_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1374_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0010)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1375_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0010) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1269_nl = MUX_s_1_2_2(nor_1374_nl, nor_1375_nl, fsm_output[5]);
  assign mux_1270_nl = MUX_s_1_2_2(nor_1373_nl, mux_1269_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1376_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0010)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1271_nl = MUX_s_1_2_2(mux_1270_nl, nor_1376_nl, fsm_output[1]);
  assign nor_1377_nl = ~((z_out_2_12_1[3:0]!=4'b0010) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1378_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1268_nl = MUX_s_1_2_2(nor_1377_nl, nor_1378_nl, fsm_output[1]);
  assign mux_1272_nl = MUX_s_1_2_2(mux_1271_nl, mux_1268_nl, fsm_output[0]);
  assign mux_1274_nl = MUX_s_1_2_2(mux_1273_nl, mux_1272_nl, fsm_output[6]);
  assign mux_1284_nl = MUX_s_1_2_2(mux_1283_nl, mux_1274_nl, fsm_output[8]);
  assign vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1299_nl,
      mux_1284_nl, fsm_output[4]);
  assign or_949_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign nand_404_nl = ~((fsm_output[9]) & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b0011)
      & (fsm_output[10]));
  assign mux_1326_nl = MUX_s_1_2_2(or_949_nl, nand_404_nl, fsm_output[7]);
  assign or_946_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b00) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1327_nl = MUX_s_1_2_2(mux_1326_nl, or_946_nl, fsm_output[2]);
  assign nor_1333_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1327_nl);
  assign nor_1334_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011)
      | (~ (fsm_output[10])));
  assign mux_1328_nl = MUX_s_1_2_2(nor_1333_nl, nor_1334_nl, fsm_output[8]);
  assign nor_1335_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1336_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011)
      | (fsm_output[10]));
  assign nor_1337_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (fsm_output[10]));
  assign nor_1338_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1323_nl = MUX_s_1_2_2(nor_1337_nl, nor_1338_nl, fsm_output[4]);
  assign mux_1324_nl = MUX_s_1_2_2(nor_1336_nl, mux_1323_nl, fsm_output[6]);
  assign mux_1325_nl = MUX_s_1_2_2(nor_1335_nl, mux_1324_nl, fsm_output[8]);
  assign mux_1329_nl = MUX_s_1_2_2(mux_1328_nl, mux_1325_nl, fsm_output[0]);
  assign nand_327_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) & (fsm_output[4]) & (fsm_output[2])
      & (~ (VEC_LOOP_j_sva_11_0[2])) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_936_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (fsm_output[2]) | (fsm_output[7])
      | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[9]) | (fsm_output[5]) | (~
      (fsm_output[10]));
  assign mux_1320_nl = MUX_s_1_2_2(mux_tmp_1308, or_936_nl, fsm_output[4]);
  assign mux_1321_nl = MUX_s_1_2_2(nand_327_nl, mux_1320_nl, fsm_output[6]);
  assign and_614_nl = (fsm_output[8]) & (~ mux_1321_nl);
  assign or_933_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0011) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_931_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (~ (fsm_output[10]));
  assign mux_1317_nl = MUX_s_1_2_2(or_931_nl, or_tmp_866, fsm_output[2]);
  assign mux_1318_nl = MUX_s_1_2_2(or_933_nl, mux_1317_nl, fsm_output[4]);
  assign nor_1339_nl = ~((fsm_output[6]) | mux_1318_nl);
  assign nor_1340_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1319_nl = MUX_s_1_2_2(nor_1339_nl, nor_1340_nl, fsm_output[8]);
  assign mux_1322_nl = MUX_s_1_2_2(and_614_nl, mux_1319_nl, fsm_output[0]);
  assign mux_1330_nl = MUX_s_1_2_2(mux_1329_nl, mux_1322_nl, fsm_output[3]);
  assign or_927_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_925_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (~ (fsm_output[10]));
  assign mux_1313_nl = MUX_s_1_2_2(or_927_nl, or_925_nl, fsm_output[4]);
  assign nor_1341_nl = ~((fsm_output[6]) | mux_1313_nl);
  assign or_919_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011)
      | (~ (fsm_output[10]));
  assign mux_1311_nl = MUX_s_1_2_2(or_702_cse, or_919_nl, fsm_output[7]);
  assign mux_1312_nl = MUX_s_1_2_2(or_tmp_866, mux_1311_nl, nor_209_cse);
  assign nor_1342_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1312_nl);
  assign mux_1314_nl = MUX_s_1_2_2(nor_1341_nl, nor_1342_nl, fsm_output[8]);
  assign or_915_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_913_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1309_nl = MUX_s_1_2_2(or_915_nl, or_913_nl, fsm_output[2]);
  assign mux_1310_nl = MUX_s_1_2_2(mux_1309_nl, mux_tmp_1308, fsm_output[4]);
  assign nor_1343_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1310_nl);
  assign mux_1315_nl = MUX_s_1_2_2(mux_1314_nl, nor_1343_nl, fsm_output[0]);
  assign or_908_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b001) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_906_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (fsm_output[10]);
  assign mux_1305_nl = MUX_s_1_2_2(or_908_nl, or_906_nl, fsm_output[4]);
  assign or_905_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_904_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (fsm_output[10]);
  assign mux_1304_nl = MUX_s_1_2_2(or_905_nl, or_904_nl, fsm_output[4]);
  assign mux_1306_nl = MUX_s_1_2_2(mux_1305_nl, mux_1304_nl, fsm_output[6]);
  assign nor_1344_nl = ~((fsm_output[8]) | mux_1306_nl);
  assign nor_1345_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1346_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (fsm_output[9]) | not_tmp_248);
  assign or_899_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011)
      | (~ (fsm_output[10]));
  assign or_897_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0011) | (fsm_output[10]);
  assign mux_1301_nl = MUX_s_1_2_2(or_899_nl, or_897_nl, fsm_output[2]);
  assign nor_1347_nl = ~((fsm_output[4]) | mux_1301_nl);
  assign mux_1302_nl = MUX_s_1_2_2(nor_1346_nl, nor_1347_nl, fsm_output[6]);
  assign mux_1303_nl = MUX_s_1_2_2(nor_1345_nl, mux_1302_nl, fsm_output[8]);
  assign mux_1307_nl = MUX_s_1_2_2(nor_1344_nl, mux_1303_nl, fsm_output[0]);
  assign mux_1316_nl = MUX_s_1_2_2(mux_1315_nl, mux_1307_nl, fsm_output[3]);
  assign vec_rsc_0_3_i_wea_d_pff = MUX_s_1_2_2(mux_1330_nl, mux_1316_nl, fsm_output[1]);
  assign or_1005_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0011) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1004_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0011) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1361_nl = MUX_s_1_2_2(or_1005_nl, or_1004_nl, fsm_output[5]);
  assign nor_1302_nl = ~((fsm_output[1]) | mux_1361_nl);
  assign nor_1303_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0011)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1304_nl = ~((z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1305_nl = ~((z_out_2_12_1[3:0]!=4'b0011) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1359_nl = MUX_s_1_2_2(nor_1304_nl, nor_1305_nl, fsm_output[5]);
  assign mux_1360_nl = MUX_s_1_2_2(nor_1303_nl, mux_1359_nl, fsm_output[1]);
  assign mux_1362_nl = MUX_s_1_2_2(nor_1302_nl, mux_1360_nl, fsm_output[0]);
  assign and_611_nl = (fsm_output[6]) & mux_1362_nl;
  assign nor_1306_nl = ~((z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1308_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1354_nl = MUX_s_1_2_2(nor_1445_cse, nor_1308_nl, fsm_output[5]);
  assign nor_1309_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0011)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_991_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0011) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1355_nl = MUX_s_1_2_2(mux_1354_nl, nor_1309_nl, or_991_nl);
  assign mux_1356_nl = MUX_s_1_2_2(nor_1306_nl, mux_1355_nl, fsm_output[1]);
  assign nor_1310_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b00) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1311_nl = ~((z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1312_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1352_nl = MUX_s_1_2_2(nor_1311_nl, nor_1312_nl, fsm_output[5]);
  assign mux_1353_nl = MUX_s_1_2_2(nor_1310_nl, mux_1352_nl, fsm_output[1]);
  assign mux_1357_nl = MUX_s_1_2_2(mux_1356_nl, mux_1353_nl, fsm_output[0]);
  assign nor_1313_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0011) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1314_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0011) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1350_nl = MUX_s_1_2_2(nor_1313_nl, nor_1314_nl, fsm_output[1]);
  assign nor_1315_nl = ~(nand_324_cse | mux_1157_cse);
  assign mux_1351_nl = MUX_s_1_2_2(mux_1350_nl, nor_1315_nl, fsm_output[0]);
  assign mux_1358_nl = MUX_s_1_2_2(mux_1357_nl, mux_1351_nl, fsm_output[6]);
  assign mux_1363_nl = MUX_s_1_2_2(and_611_nl, mux_1358_nl, fsm_output[8]);
  assign nor_1316_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0011) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1317_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0011) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1344_nl = MUX_s_1_2_2(nor_1316_nl, nor_1317_nl, fsm_output[5]);
  assign and_612_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1344_nl;
  assign nor_1318_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0011)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1319_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0011) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1343_nl = MUX_s_1_2_2(nor_1318_nl, nor_1319_nl, fsm_output[5]);
  assign and_613_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1343_nl;
  assign mux_1345_nl = MUX_s_1_2_2(and_612_nl, and_613_nl, fsm_output[1]);
  assign nor_1320_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1321_nl = ~(nand_332_cse | mux_1277_cse);
  assign mux_1342_nl = MUX_s_1_2_2(nor_1320_nl, nor_1321_nl, fsm_output[1]);
  assign mux_1346_nl = MUX_s_1_2_2(mux_1345_nl, mux_1342_nl, fsm_output[0]);
  assign nor_1322_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1323_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1324_nl = ~((~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b001) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1339_nl = MUX_s_1_2_2(nor_1323_nl, nor_1324_nl, fsm_output[1]);
  assign mux_1340_nl = MUX_s_1_2_2(nor_1322_nl, mux_1339_nl, fsm_output[0]);
  assign mux_1347_nl = MUX_s_1_2_2(mux_1346_nl, mux_1340_nl, fsm_output[6]);
  assign nor_1325_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0011) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1326_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0011)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1337_nl = MUX_s_1_2_2(nor_1325_nl, nor_1326_nl, fsm_output[0]);
  assign nor_1327_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0011)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1328_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0011)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1329_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0011) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1333_nl = MUX_s_1_2_2(nor_1328_nl, nor_1329_nl, fsm_output[5]);
  assign mux_1334_nl = MUX_s_1_2_2(nor_1327_nl, mux_1333_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1330_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0011)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1335_nl = MUX_s_1_2_2(mux_1334_nl, nor_1330_nl, fsm_output[1]);
  assign nor_1331_nl = ~((z_out_2_12_1[3:0]!=4'b0011) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1332_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b001) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1332_nl = MUX_s_1_2_2(nor_1331_nl, nor_1332_nl, fsm_output[1]);
  assign mux_1336_nl = MUX_s_1_2_2(mux_1335_nl, mux_1332_nl, fsm_output[0]);
  assign mux_1338_nl = MUX_s_1_2_2(mux_1337_nl, mux_1336_nl, fsm_output[6]);
  assign mux_1348_nl = MUX_s_1_2_2(mux_1347_nl, mux_1338_nl, fsm_output[8]);
  assign vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1363_nl,
      mux_1348_nl, fsm_output[4]);
  assign or_1060_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1059_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (~ (fsm_output[10]));
  assign mux_1390_nl = MUX_s_1_2_2(or_1060_nl, or_1059_nl, fsm_output[7]);
  assign or_1057_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b01) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1391_nl = MUX_s_1_2_2(mux_1390_nl, or_1057_nl, fsm_output[2]);
  assign nor_1287_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1391_nl);
  assign nor_1288_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (~ (fsm_output[10])));
  assign mux_1392_nl = MUX_s_1_2_2(nor_1287_nl, nor_1288_nl, fsm_output[8]);
  assign nor_1289_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1290_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (fsm_output[10]));
  assign nor_1291_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (fsm_output[10]));
  assign nor_1292_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1387_nl = MUX_s_1_2_2(nor_1291_nl, nor_1292_nl, fsm_output[4]);
  assign mux_1388_nl = MUX_s_1_2_2(nor_1290_nl, mux_1387_nl, fsm_output[6]);
  assign mux_1389_nl = MUX_s_1_2_2(nor_1289_nl, mux_1388_nl, fsm_output[8]);
  assign mux_1393_nl = MUX_s_1_2_2(mux_1392_nl, mux_1389_nl, fsm_output[0]);
  assign or_1048_nl = (COMP_LOOP_acc_16_psp_sva[0]) | (~ (fsm_output[4])) | (~ (fsm_output[2]))
      | (~ (VEC_LOOP_j_sva_11_0[2])) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1047_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1384_nl = MUX_s_1_2_2(mux_tmp_1372, or_1047_nl, fsm_output[4]);
  assign mux_1385_nl = MUX_s_1_2_2(or_1048_nl, mux_1384_nl, fsm_output[6]);
  assign and_610_nl = (fsm_output[8]) & (~ mux_1385_nl);
  assign or_1044_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_1042_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (~ (fsm_output[10]));
  assign mux_1381_nl = MUX_s_1_2_2(or_1042_nl, or_tmp_974, fsm_output[2]);
  assign mux_1382_nl = MUX_s_1_2_2(or_1044_nl, mux_1381_nl, fsm_output[4]);
  assign nor_1293_nl = ~((fsm_output[6]) | mux_1382_nl);
  assign nor_1294_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1383_nl = MUX_s_1_2_2(nor_1293_nl, nor_1294_nl, fsm_output[8]);
  assign mux_1386_nl = MUX_s_1_2_2(and_610_nl, mux_1383_nl, fsm_output[0]);
  assign mux_1394_nl = MUX_s_1_2_2(mux_1393_nl, mux_1386_nl, fsm_output[3]);
  assign or_1038_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[0]) | nand_337_cse;
  assign or_1036_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (~ (fsm_output[10]));
  assign mux_1377_nl = MUX_s_1_2_2(or_1038_nl, or_1036_nl, fsm_output[4]);
  assign nor_1295_nl = ~((fsm_output[6]) | mux_1377_nl);
  assign or_1032_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (~ (fsm_output[10]));
  assign mux_1375_nl = MUX_s_1_2_2(or_591_cse, or_1032_nl, fsm_output[7]);
  assign mux_1376_nl = MUX_s_1_2_2(mux_1375_nl, or_tmp_974, or_1028_cse);
  assign nor_1296_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1376_nl);
  assign mux_1378_nl = MUX_s_1_2_2(nor_1295_nl, nor_1296_nl, fsm_output[8]);
  assign or_1025_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1023_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1373_nl = MUX_s_1_2_2(or_1025_nl, or_1023_nl, fsm_output[2]);
  assign mux_1374_nl = MUX_s_1_2_2(mux_1373_nl, mux_tmp_1372, fsm_output[4]);
  assign nor_1297_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1374_nl);
  assign mux_1379_nl = MUX_s_1_2_2(mux_1378_nl, nor_1297_nl, fsm_output[0]);
  assign or_1018_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1016_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (fsm_output[10]);
  assign mux_1369_nl = MUX_s_1_2_2(or_1018_nl, or_1016_nl, fsm_output[4]);
  assign or_1015_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9])) | (~
      (fsm_output[5])) | (fsm_output[10]);
  assign or_1014_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (fsm_output[10]);
  assign mux_1368_nl = MUX_s_1_2_2(or_1015_nl, or_1014_nl, fsm_output[4]);
  assign mux_1370_nl = MUX_s_1_2_2(mux_1369_nl, mux_1368_nl, fsm_output[6]);
  assign nor_1298_nl = ~((fsm_output[8]) | mux_1370_nl);
  assign nor_1299_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1300_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (fsm_output[9]) | not_tmp_248);
  assign or_1009_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100)
      | (~ (fsm_output[10]));
  assign or_1007_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0100) | (fsm_output[10]);
  assign mux_1365_nl = MUX_s_1_2_2(or_1009_nl, or_1007_nl, fsm_output[2]);
  assign nor_1301_nl = ~((fsm_output[4]) | mux_1365_nl);
  assign mux_1366_nl = MUX_s_1_2_2(nor_1300_nl, nor_1301_nl, fsm_output[6]);
  assign mux_1367_nl = MUX_s_1_2_2(nor_1299_nl, mux_1366_nl, fsm_output[8]);
  assign mux_1371_nl = MUX_s_1_2_2(nor_1298_nl, mux_1367_nl, fsm_output[0]);
  assign mux_1380_nl = MUX_s_1_2_2(mux_1379_nl, mux_1371_nl, fsm_output[3]);
  assign vec_rsc_0_4_i_wea_d_pff = MUX_s_1_2_2(mux_1394_nl, mux_1380_nl, fsm_output[1]);
  assign or_1116_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0100) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1115_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0100) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1425_nl = MUX_s_1_2_2(or_1116_nl, or_1115_nl, fsm_output[5]);
  assign nor_1256_nl = ~((fsm_output[1]) | mux_1425_nl);
  assign nor_1257_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0100)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1258_nl = ~((z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1259_nl = ~((z_out_2_12_1[3:0]!=4'b0100) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1423_nl = MUX_s_1_2_2(nor_1258_nl, nor_1259_nl, fsm_output[5]);
  assign mux_1424_nl = MUX_s_1_2_2(nor_1257_nl, mux_1423_nl, fsm_output[1]);
  assign mux_1426_nl = MUX_s_1_2_2(nor_1256_nl, mux_1424_nl, fsm_output[0]);
  assign and_607_nl = (fsm_output[6]) & mux_1426_nl;
  assign nor_1260_nl = ~((z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1262_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1418_nl = MUX_s_1_2_2(nor_1445_cse, nor_1262_nl, fsm_output[5]);
  assign nor_1263_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1102_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1419_nl = MUX_s_1_2_2(mux_1418_nl, nor_1263_nl, or_1102_nl);
  assign mux_1420_nl = MUX_s_1_2_2(nor_1260_nl, mux_1419_nl, fsm_output[1]);
  assign nor_1264_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1265_nl = ~((z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1266_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1416_nl = MUX_s_1_2_2(nor_1265_nl, nor_1266_nl, fsm_output[5]);
  assign mux_1417_nl = MUX_s_1_2_2(nor_1264_nl, mux_1416_nl, fsm_output[1]);
  assign mux_1421_nl = MUX_s_1_2_2(mux_1420_nl, mux_1417_nl, fsm_output[0]);
  assign nor_1267_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1268_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0100) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1414_nl = MUX_s_1_2_2(nor_1267_nl, nor_1268_nl, fsm_output[1]);
  assign nor_1269_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1413_cse);
  assign mux_1415_nl = MUX_s_1_2_2(mux_1414_nl, nor_1269_nl, fsm_output[0]);
  assign mux_1422_nl = MUX_s_1_2_2(mux_1421_nl, mux_1415_nl, fsm_output[6]);
  assign mux_1427_nl = MUX_s_1_2_2(and_607_nl, mux_1422_nl, fsm_output[8]);
  assign nor_1270_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0100) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1271_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0100) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1408_nl = MUX_s_1_2_2(nor_1270_nl, nor_1271_nl, fsm_output[5]);
  assign and_608_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1408_nl;
  assign nor_1272_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1273_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0100) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1407_nl = MUX_s_1_2_2(nor_1272_nl, nor_1273_nl, fsm_output[5]);
  assign and_609_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1407_nl;
  assign mux_1409_nl = MUX_s_1_2_2(and_608_nl, and_609_nl, fsm_output[1]);
  assign nor_1274_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (VEC_LOOP_j_sva_11_0[1]) | (VEC_LOOP_j_sva_11_0[0])
      | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2])) | (fsm_output[7]) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1275_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1405_cse);
  assign mux_1406_nl = MUX_s_1_2_2(nor_1274_nl, nor_1275_nl, fsm_output[1]);
  assign mux_1410_nl = MUX_s_1_2_2(mux_1409_nl, mux_1406_nl, fsm_output[0]);
  assign nor_1276_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1277_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1278_nl = ~((COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1403_nl = MUX_s_1_2_2(nor_1277_nl, nor_1278_nl, fsm_output[1]);
  assign mux_1404_nl = MUX_s_1_2_2(nor_1276_nl, mux_1403_nl, fsm_output[0]);
  assign mux_1411_nl = MUX_s_1_2_2(mux_1410_nl, mux_1404_nl, fsm_output[6]);
  assign nor_1279_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0100) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1280_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0100)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1401_nl = MUX_s_1_2_2(nor_1279_nl, nor_1280_nl, fsm_output[0]);
  assign nor_1281_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1282_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0100)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1283_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0100) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1397_nl = MUX_s_1_2_2(nor_1282_nl, nor_1283_nl, fsm_output[5]);
  assign mux_1398_nl = MUX_s_1_2_2(nor_1281_nl, mux_1397_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1284_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0100)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1399_nl = MUX_s_1_2_2(mux_1398_nl, nor_1284_nl, fsm_output[1]);
  assign nor_1285_nl = ~((z_out_2_12_1[3:0]!=4'b0100) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1286_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1396_nl = MUX_s_1_2_2(nor_1285_nl, nor_1286_nl, fsm_output[1]);
  assign mux_1400_nl = MUX_s_1_2_2(mux_1399_nl, mux_1396_nl, fsm_output[0]);
  assign mux_1402_nl = MUX_s_1_2_2(mux_1401_nl, mux_1400_nl, fsm_output[6]);
  assign mux_1412_nl = MUX_s_1_2_2(mux_1411_nl, mux_1402_nl, fsm_output[8]);
  assign vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1427_nl,
      mux_1412_nl, fsm_output[4]);
  assign or_1171_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign nand_403_nl = ~((fsm_output[9]) & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b0101)
      & (fsm_output[10]));
  assign mux_1454_nl = MUX_s_1_2_2(or_1171_nl, nand_403_nl, fsm_output[7]);
  assign or_1168_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b01) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1455_nl = MUX_s_1_2_2(mux_1454_nl, or_1168_nl, fsm_output[2]);
  assign nor_1241_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1455_nl);
  assign nor_1242_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101)
      | (~ (fsm_output[10])));
  assign mux_1456_nl = MUX_s_1_2_2(nor_1241_nl, nor_1242_nl, fsm_output[8]);
  assign nor_1243_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1244_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101)
      | (fsm_output[10]));
  assign nor_1245_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (fsm_output[10]));
  assign nor_1246_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1451_nl = MUX_s_1_2_2(nor_1245_nl, nor_1246_nl, fsm_output[4]);
  assign mux_1452_nl = MUX_s_1_2_2(nor_1244_nl, mux_1451_nl, fsm_output[6]);
  assign mux_1453_nl = MUX_s_1_2_2(nor_1243_nl, mux_1452_nl, fsm_output[8]);
  assign mux_1457_nl = MUX_s_1_2_2(mux_1456_nl, mux_1453_nl, fsm_output[0]);
  assign nand_318_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b01)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_1158_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1448_nl = MUX_s_1_2_2(mux_tmp_1436, or_1158_nl, fsm_output[4]);
  assign mux_1449_nl = MUX_s_1_2_2(nand_318_nl, mux_1448_nl, fsm_output[6]);
  assign and_606_nl = (fsm_output[8]) & (~ mux_1449_nl);
  assign or_1155_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0101) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_1153_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (~ (fsm_output[10]));
  assign mux_1445_nl = MUX_s_1_2_2(or_1153_nl, or_tmp_1085, fsm_output[2]);
  assign mux_1446_nl = MUX_s_1_2_2(or_1155_nl, mux_1445_nl, fsm_output[4]);
  assign nor_1247_nl = ~((fsm_output[6]) | mux_1446_nl);
  assign nor_1248_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1447_nl = MUX_s_1_2_2(nor_1247_nl, nor_1248_nl, fsm_output[8]);
  assign mux_1450_nl = MUX_s_1_2_2(and_606_nl, mux_1447_nl, fsm_output[0]);
  assign mux_1458_nl = MUX_s_1_2_2(mux_1457_nl, mux_1450_nl, fsm_output[3]);
  assign or_1149_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_1147_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (~ (fsm_output[10]));
  assign mux_1441_nl = MUX_s_1_2_2(or_1149_nl, or_1147_nl, fsm_output[4]);
  assign nor_1249_nl = ~((fsm_output[6]) | mux_1441_nl);
  assign or_1143_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101)
      | (~ (fsm_output[10]));
  assign mux_1439_nl = MUX_s_1_2_2(or_702_cse, or_1143_nl, fsm_output[7]);
  assign mux_1440_nl = MUX_s_1_2_2(mux_1439_nl, or_tmp_1085, or_1028_cse);
  assign nor_1250_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1440_nl);
  assign mux_1442_nl = MUX_s_1_2_2(nor_1249_nl, nor_1250_nl, fsm_output[8]);
  assign or_1136_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1134_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1437_nl = MUX_s_1_2_2(or_1136_nl, or_1134_nl, fsm_output[2]);
  assign mux_1438_nl = MUX_s_1_2_2(mux_1437_nl, mux_tmp_1436, fsm_output[4]);
  assign nor_1251_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1438_nl);
  assign mux_1443_nl = MUX_s_1_2_2(mux_1442_nl, nor_1251_nl, fsm_output[0]);
  assign or_1129_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b010) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1127_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (fsm_output[10]);
  assign mux_1433_nl = MUX_s_1_2_2(or_1129_nl, or_1127_nl, fsm_output[4]);
  assign or_1126_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b010) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1125_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (fsm_output[10]);
  assign mux_1432_nl = MUX_s_1_2_2(or_1126_nl, or_1125_nl, fsm_output[4]);
  assign mux_1434_nl = MUX_s_1_2_2(mux_1433_nl, mux_1432_nl, fsm_output[6]);
  assign nor_1252_nl = ~((fsm_output[8]) | mux_1434_nl);
  assign nor_1253_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1254_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (fsm_output[9]) | not_tmp_248);
  assign or_1120_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101)
      | (~ (fsm_output[10]));
  assign or_1118_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0101) | (fsm_output[10]);
  assign mux_1429_nl = MUX_s_1_2_2(or_1120_nl, or_1118_nl, fsm_output[2]);
  assign nor_1255_nl = ~((fsm_output[4]) | mux_1429_nl);
  assign mux_1430_nl = MUX_s_1_2_2(nor_1254_nl, nor_1255_nl, fsm_output[6]);
  assign mux_1431_nl = MUX_s_1_2_2(nor_1253_nl, mux_1430_nl, fsm_output[8]);
  assign mux_1435_nl = MUX_s_1_2_2(nor_1252_nl, mux_1431_nl, fsm_output[0]);
  assign mux_1444_nl = MUX_s_1_2_2(mux_1443_nl, mux_1435_nl, fsm_output[3]);
  assign vec_rsc_0_5_i_wea_d_pff = MUX_s_1_2_2(mux_1458_nl, mux_1444_nl, fsm_output[1]);
  assign or_1227_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0101) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1226_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0101) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1489_nl = MUX_s_1_2_2(or_1227_nl, or_1226_nl, fsm_output[5]);
  assign nor_1210_nl = ~((fsm_output[1]) | mux_1489_nl);
  assign nor_1211_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0101)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1212_nl = ~((z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1213_nl = ~((z_out_2_12_1[3:0]!=4'b0101) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1487_nl = MUX_s_1_2_2(nor_1212_nl, nor_1213_nl, fsm_output[5]);
  assign mux_1488_nl = MUX_s_1_2_2(nor_1211_nl, mux_1487_nl, fsm_output[1]);
  assign mux_1490_nl = MUX_s_1_2_2(nor_1210_nl, mux_1488_nl, fsm_output[0]);
  assign and_603_nl = (fsm_output[6]) & mux_1490_nl;
  assign nor_1214_nl = ~((z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1216_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1482_nl = MUX_s_1_2_2(nor_1445_cse, nor_1216_nl, fsm_output[5]);
  assign nor_1217_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0101)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1213_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0101) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1483_nl = MUX_s_1_2_2(mux_1482_nl, nor_1217_nl, or_1213_nl);
  assign mux_1484_nl = MUX_s_1_2_2(nor_1214_nl, mux_1483_nl, fsm_output[1]);
  assign nor_1218_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1219_nl = ~((z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1220_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1480_nl = MUX_s_1_2_2(nor_1219_nl, nor_1220_nl, fsm_output[5]);
  assign mux_1481_nl = MUX_s_1_2_2(nor_1218_nl, mux_1480_nl, fsm_output[1]);
  assign mux_1485_nl = MUX_s_1_2_2(mux_1484_nl, mux_1481_nl, fsm_output[0]);
  assign nor_1221_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0101) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1222_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0101) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1478_nl = MUX_s_1_2_2(nor_1221_nl, nor_1222_nl, fsm_output[1]);
  assign nor_1223_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1413_cse);
  assign mux_1479_nl = MUX_s_1_2_2(mux_1478_nl, nor_1223_nl, fsm_output[0]);
  assign mux_1486_nl = MUX_s_1_2_2(mux_1485_nl, mux_1479_nl, fsm_output[6]);
  assign mux_1491_nl = MUX_s_1_2_2(and_603_nl, mux_1486_nl, fsm_output[8]);
  assign nor_1224_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0101) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1225_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0101) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1472_nl = MUX_s_1_2_2(nor_1224_nl, nor_1225_nl, fsm_output[5]);
  assign and_604_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1472_nl;
  assign nor_1226_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0101)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1227_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0101) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1471_nl = MUX_s_1_2_2(nor_1226_nl, nor_1227_nl, fsm_output[5]);
  assign and_605_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1471_nl;
  assign mux_1473_nl = MUX_s_1_2_2(and_604_nl, and_605_nl, fsm_output[1]);
  assign nor_1228_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (VEC_LOOP_j_sva_11_0[1]) | (~
      (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1229_nl = ~(nand_332_cse | mux_1405_cse);
  assign mux_1470_nl = MUX_s_1_2_2(nor_1228_nl, nor_1229_nl, fsm_output[1]);
  assign mux_1474_nl = MUX_s_1_2_2(mux_1473_nl, mux_1470_nl, fsm_output[0]);
  assign nor_1230_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1231_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1232_nl = ~((~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b010) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1467_nl = MUX_s_1_2_2(nor_1231_nl, nor_1232_nl, fsm_output[1]);
  assign mux_1468_nl = MUX_s_1_2_2(nor_1230_nl, mux_1467_nl, fsm_output[0]);
  assign mux_1475_nl = MUX_s_1_2_2(mux_1474_nl, mux_1468_nl, fsm_output[6]);
  assign nor_1233_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0101) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1234_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0101)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1465_nl = MUX_s_1_2_2(nor_1233_nl, nor_1234_nl, fsm_output[0]);
  assign nor_1235_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0101)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1236_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0101)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1237_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0101) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1461_nl = MUX_s_1_2_2(nor_1236_nl, nor_1237_nl, fsm_output[5]);
  assign mux_1462_nl = MUX_s_1_2_2(nor_1235_nl, mux_1461_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1238_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0101)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1463_nl = MUX_s_1_2_2(mux_1462_nl, nor_1238_nl, fsm_output[1]);
  assign nor_1239_nl = ~((z_out_2_12_1[3:0]!=4'b0101) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1240_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b010) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1460_nl = MUX_s_1_2_2(nor_1239_nl, nor_1240_nl, fsm_output[1]);
  assign mux_1464_nl = MUX_s_1_2_2(mux_1463_nl, mux_1460_nl, fsm_output[0]);
  assign mux_1466_nl = MUX_s_1_2_2(mux_1465_nl, mux_1464_nl, fsm_output[6]);
  assign mux_1476_nl = MUX_s_1_2_2(mux_1475_nl, mux_1466_nl, fsm_output[8]);
  assign vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1491_nl,
      mux_1476_nl, fsm_output[4]);
  assign or_1281_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign nand_402_nl = ~((fsm_output[9]) & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b0110)
      & (fsm_output[10]));
  assign mux_1518_nl = MUX_s_1_2_2(or_1281_nl, nand_402_nl, fsm_output[7]);
  assign or_1278_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b01) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1519_nl = MUX_s_1_2_2(mux_1518_nl, or_1278_nl, fsm_output[2]);
  assign nor_1195_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1519_nl);
  assign nor_1196_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110)
      | (~ (fsm_output[10])));
  assign mux_1520_nl = MUX_s_1_2_2(nor_1195_nl, nor_1196_nl, fsm_output[8]);
  assign nor_1197_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1198_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110)
      | (fsm_output[10]));
  assign nor_1199_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (fsm_output[10]));
  assign nor_1200_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1515_nl = MUX_s_1_2_2(nor_1199_nl, nor_1200_nl, fsm_output[4]);
  assign mux_1516_nl = MUX_s_1_2_2(nor_1198_nl, mux_1515_nl, fsm_output[6]);
  assign mux_1517_nl = MUX_s_1_2_2(nor_1197_nl, mux_1516_nl, fsm_output[8]);
  assign mux_1521_nl = MUX_s_1_2_2(mux_1520_nl, mux_1517_nl, fsm_output[0]);
  assign nand_313_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b10)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_1268_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1512_nl = MUX_s_1_2_2(mux_tmp_1500, or_1268_nl, fsm_output[4]);
  assign mux_1513_nl = MUX_s_1_2_2(nand_313_nl, mux_1512_nl, fsm_output[6]);
  assign and_602_nl = (fsm_output[8]) & (~ mux_1513_nl);
  assign or_1265_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_1263_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (~ (fsm_output[10]));
  assign mux_1509_nl = MUX_s_1_2_2(or_1263_nl, or_tmp_1198, fsm_output[2]);
  assign mux_1510_nl = MUX_s_1_2_2(or_1265_nl, mux_1509_nl, fsm_output[4]);
  assign nor_1201_nl = ~((fsm_output[6]) | mux_1510_nl);
  assign nor_1202_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1511_nl = MUX_s_1_2_2(nor_1201_nl, nor_1202_nl, fsm_output[8]);
  assign mux_1514_nl = MUX_s_1_2_2(and_602_nl, mux_1511_nl, fsm_output[0]);
  assign mux_1522_nl = MUX_s_1_2_2(mux_1521_nl, mux_1514_nl, fsm_output[3]);
  assign or_1259_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[0]) | nand_337_cse;
  assign or_1257_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (~ (fsm_output[10]));
  assign mux_1505_nl = MUX_s_1_2_2(or_1259_nl, or_1257_nl, fsm_output[4]);
  assign nor_1203_nl = ~((fsm_output[6]) | mux_1505_nl);
  assign or_1251_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110)
      | (~ (fsm_output[10]));
  assign mux_1503_nl = MUX_s_1_2_2(or_591_cse, or_1251_nl, fsm_output[7]);
  assign mux_1504_nl = MUX_s_1_2_2(or_tmp_1198, mux_1503_nl, nor_223_cse);
  assign nor_1204_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1504_nl);
  assign mux_1506_nl = MUX_s_1_2_2(nor_1203_nl, nor_1204_nl, fsm_output[8]);
  assign or_1247_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1245_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1501_nl = MUX_s_1_2_2(or_1247_nl, or_1245_nl, fsm_output[2]);
  assign mux_1502_nl = MUX_s_1_2_2(mux_1501_nl, mux_tmp_1500, fsm_output[4]);
  assign nor_1205_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1502_nl);
  assign mux_1507_nl = MUX_s_1_2_2(mux_1506_nl, nor_1205_nl, fsm_output[0]);
  assign or_1240_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1238_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (fsm_output[10]);
  assign mux_1497_nl = MUX_s_1_2_2(or_1240_nl, or_1238_nl, fsm_output[4]);
  assign or_1237_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b011) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9])) | (~
      (fsm_output[5])) | (fsm_output[10]);
  assign or_1236_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (fsm_output[10]);
  assign mux_1496_nl = MUX_s_1_2_2(or_1237_nl, or_1236_nl, fsm_output[4]);
  assign mux_1498_nl = MUX_s_1_2_2(mux_1497_nl, mux_1496_nl, fsm_output[6]);
  assign nor_1206_nl = ~((fsm_output[8]) | mux_1498_nl);
  assign nor_1207_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1208_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (fsm_output[9]) | not_tmp_248);
  assign or_1231_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110)
      | (~ (fsm_output[10]));
  assign or_1229_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0110) | (fsm_output[10]);
  assign mux_1493_nl = MUX_s_1_2_2(or_1231_nl, or_1229_nl, fsm_output[2]);
  assign nor_1209_nl = ~((fsm_output[4]) | mux_1493_nl);
  assign mux_1494_nl = MUX_s_1_2_2(nor_1208_nl, nor_1209_nl, fsm_output[6]);
  assign mux_1495_nl = MUX_s_1_2_2(nor_1207_nl, mux_1494_nl, fsm_output[8]);
  assign mux_1499_nl = MUX_s_1_2_2(nor_1206_nl, mux_1495_nl, fsm_output[0]);
  assign mux_1508_nl = MUX_s_1_2_2(mux_1507_nl, mux_1499_nl, fsm_output[3]);
  assign vec_rsc_0_6_i_wea_d_pff = MUX_s_1_2_2(mux_1522_nl, mux_1508_nl, fsm_output[1]);
  assign or_1337_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0110) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1336_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0110) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1553_nl = MUX_s_1_2_2(or_1337_nl, or_1336_nl, fsm_output[5]);
  assign nor_1164_nl = ~((fsm_output[1]) | mux_1553_nl);
  assign nor_1165_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0110)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1166_nl = ~((z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1167_nl = ~((z_out_2_12_1[3:0]!=4'b0110) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1551_nl = MUX_s_1_2_2(nor_1166_nl, nor_1167_nl, fsm_output[5]);
  assign mux_1552_nl = MUX_s_1_2_2(nor_1165_nl, mux_1551_nl, fsm_output[1]);
  assign mux_1554_nl = MUX_s_1_2_2(nor_1164_nl, mux_1552_nl, fsm_output[0]);
  assign and_599_nl = (fsm_output[6]) & mux_1554_nl;
  assign nor_1168_nl = ~((z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1170_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1546_nl = MUX_s_1_2_2(nor_1445_cse, nor_1170_nl, fsm_output[5]);
  assign nor_1171_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0110)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1323_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0110) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1547_nl = MUX_s_1_2_2(mux_1546_nl, nor_1171_nl, or_1323_nl);
  assign mux_1548_nl = MUX_s_1_2_2(nor_1168_nl, mux_1547_nl, fsm_output[1]);
  assign nor_1172_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1173_nl = ~((z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1174_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1544_nl = MUX_s_1_2_2(nor_1173_nl, nor_1174_nl, fsm_output[5]);
  assign mux_1545_nl = MUX_s_1_2_2(nor_1172_nl, mux_1544_nl, fsm_output[1]);
  assign mux_1549_nl = MUX_s_1_2_2(mux_1548_nl, mux_1545_nl, fsm_output[0]);
  assign nor_1175_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0110) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1176_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0110) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1542_nl = MUX_s_1_2_2(nor_1175_nl, nor_1176_nl, fsm_output[1]);
  assign nor_1177_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1413_cse);
  assign mux_1543_nl = MUX_s_1_2_2(mux_1542_nl, nor_1177_nl, fsm_output[0]);
  assign mux_1550_nl = MUX_s_1_2_2(mux_1549_nl, mux_1543_nl, fsm_output[6]);
  assign mux_1555_nl = MUX_s_1_2_2(and_599_nl, mux_1550_nl, fsm_output[8]);
  assign nor_1178_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0110) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1179_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0110) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1536_nl = MUX_s_1_2_2(nor_1178_nl, nor_1179_nl, fsm_output[5]);
  assign and_600_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1536_nl;
  assign nor_1180_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b0110)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1181_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0110) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1535_nl = MUX_s_1_2_2(nor_1180_nl, nor_1181_nl, fsm_output[5]);
  assign and_601_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1535_nl;
  assign mux_1537_nl = MUX_s_1_2_2(and_600_nl, and_601_nl, fsm_output[1]);
  assign nor_1182_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1183_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1533_cse);
  assign mux_1534_nl = MUX_s_1_2_2(nor_1182_nl, nor_1183_nl, fsm_output[1]);
  assign mux_1538_nl = MUX_s_1_2_2(mux_1537_nl, mux_1534_nl, fsm_output[0]);
  assign nor_1184_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1185_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1186_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b011) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1531_nl = MUX_s_1_2_2(nor_1185_nl, nor_1186_nl, fsm_output[1]);
  assign mux_1532_nl = MUX_s_1_2_2(nor_1184_nl, mux_1531_nl, fsm_output[0]);
  assign mux_1539_nl = MUX_s_1_2_2(mux_1538_nl, mux_1532_nl, fsm_output[6]);
  assign nor_1187_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0110) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1188_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0110)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1529_nl = MUX_s_1_2_2(nor_1187_nl, nor_1188_nl, fsm_output[0]);
  assign nor_1189_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0110)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1190_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0110)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1191_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0110) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1525_nl = MUX_s_1_2_2(nor_1190_nl, nor_1191_nl, fsm_output[5]);
  assign mux_1526_nl = MUX_s_1_2_2(nor_1189_nl, mux_1525_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1192_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0110)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1527_nl = MUX_s_1_2_2(mux_1526_nl, nor_1192_nl, fsm_output[1]);
  assign nor_1193_nl = ~((z_out_2_12_1[3:0]!=4'b0110) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1194_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1524_nl = MUX_s_1_2_2(nor_1193_nl, nor_1194_nl, fsm_output[1]);
  assign mux_1528_nl = MUX_s_1_2_2(mux_1527_nl, mux_1524_nl, fsm_output[0]);
  assign mux_1530_nl = MUX_s_1_2_2(mux_1529_nl, mux_1528_nl, fsm_output[6]);
  assign mux_1540_nl = MUX_s_1_2_2(mux_1539_nl, mux_1530_nl, fsm_output[8]);
  assign vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1555_nl,
      mux_1540_nl, fsm_output[4]);
  assign nand_302_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b01) & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[5]) & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[10:9]==2'b01));
  assign nand_401_nl = ~((fsm_output[5]) & (fsm_output[9]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b0111)
      & (fsm_output[10]));
  assign mux_1582_nl = MUX_s_1_2_2(nand_302_nl, nand_401_nl, fsm_output[7]);
  assign or_1388_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b01) | (~ (fsm_output[7])) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[5]) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (fsm_output[10:9]!=2'b00);
  assign mux_1583_nl = MUX_s_1_2_2(mux_1582_nl, or_1388_nl, fsm_output[2]);
  assign nor_1149_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1583_nl);
  assign nor_1150_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111)
      | (~ (fsm_output[10])));
  assign mux_1584_nl = MUX_s_1_2_2(nor_1149_nl, nor_1150_nl, fsm_output[8]);
  assign and_762_nl = (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b0111) & (fsm_output[6])
      & (fsm_output[4]) & (~ (fsm_output[2])) & (fsm_output[7]) & (fsm_output[5])
      & (~ (fsm_output[9])) & (fsm_output[10]);
  assign nor_1152_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[5])
      | (~ (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (fsm_output[10]));
  assign nor_1153_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (fsm_output[10]));
  assign nor_1154_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b0111) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[10]));
  assign mux_1579_nl = MUX_s_1_2_2(nor_1153_nl, nor_1154_nl, fsm_output[4]);
  assign mux_1580_nl = MUX_s_1_2_2(nor_1152_nl, mux_1579_nl, fsm_output[6]);
  assign mux_1581_nl = MUX_s_1_2_2(and_762_nl, mux_1580_nl, fsm_output[8]);
  assign mux_1585_nl = MUX_s_1_2_2(mux_1584_nl, mux_1581_nl, fsm_output[0]);
  assign nand_305_nl = ~((~ (COMP_LOOP_acc_16_psp_sva[0])) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1]) & (fsm_output[5])
      & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[10:9]==2'b01));
  assign or_1378_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (fsm_output[2]) |
      (fsm_output[7]) | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[5]) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (fsm_output[10:9]!=2'b10);
  assign mux_1576_nl = MUX_s_1_2_2(mux_tmp_1564, or_1378_nl, fsm_output[4]);
  assign mux_1577_nl = MUX_s_1_2_2(nand_305_nl, mux_1576_nl, fsm_output[6]);
  assign and_598_nl = (fsm_output[8]) & (~ mux_1577_nl);
  assign or_1375_nl = (~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b0111) & (fsm_output[2])
      & (fsm_output[7]) & (~ (fsm_output[5])))) | nand_358_cse;
  assign nand_400_nl = ~((~ (fsm_output[7])) & (fsm_output[5]) & (fsm_output[9])
      & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b0111) & (fsm_output[10]));
  assign mux_1573_nl = MUX_s_1_2_2(nand_400_nl, or_tmp_1308, fsm_output[2]);
  assign mux_1574_nl = MUX_s_1_2_2(or_1375_nl, mux_1573_nl, fsm_output[4]);
  assign nor_1155_nl = ~((fsm_output[6]) | mux_1574_nl);
  assign nor_1156_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[10]));
  assign mux_1575_nl = MUX_s_1_2_2(nor_1155_nl, nor_1156_nl, fsm_output[8]);
  assign mux_1578_nl = MUX_s_1_2_2(and_598_nl, mux_1575_nl, fsm_output[0]);
  assign mux_1586_nl = MUX_s_1_2_2(mux_1585_nl, mux_1578_nl, fsm_output[3]);
  assign or_1369_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_1367_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (~ (fsm_output[10]));
  assign mux_1569_nl = MUX_s_1_2_2(or_1369_nl, or_1367_nl, fsm_output[4]);
  assign nor_1157_nl = ~((fsm_output[6]) | mux_1569_nl);
  assign or_1361_nl = (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111)
      | (~ (fsm_output[10]));
  assign mux_1567_nl = MUX_s_1_2_2(or_702_cse, or_1361_nl, fsm_output[7]);
  assign mux_1568_nl = MUX_s_1_2_2(or_tmp_1308, mux_1567_nl, nor_223_cse);
  assign nor_1158_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1568_nl);
  assign mux_1570_nl = MUX_s_1_2_2(nor_1157_nl, nor_1158_nl, fsm_output[8]);
  assign or_1357_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0111) | (fsm_output[7])
      | (~ (fsm_output[5])) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign or_1355_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0111) | (~ (fsm_output[7]))
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign mux_1565_nl = MUX_s_1_2_2(or_1357_nl, or_1355_nl, fsm_output[2]);
  assign mux_1566_nl = MUX_s_1_2_2(mux_1565_nl, mux_tmp_1564, fsm_output[4]);
  assign nor_1159_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1566_nl);
  assign mux_1571_nl = MUX_s_1_2_2(mux_1570_nl, nor_1159_nl, fsm_output[0]);
  assign or_1350_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b011) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (fsm_output[5]) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[10:9]!=2'b10);
  assign or_1348_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[5]) | (~
      (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (fsm_output[10]);
  assign mux_1561_nl = MUX_s_1_2_2(or_1350_nl, or_1348_nl, fsm_output[4]);
  assign nand_310_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b011) & (fsm_output[2])
      & (fsm_output[7]) & (fsm_output[5]) & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[10:9]==2'b01));
  assign or_1346_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (fsm_output[10]);
  assign mux_1560_nl = MUX_s_1_2_2(nand_310_nl, or_1346_nl, fsm_output[4]);
  assign mux_1562_nl = MUX_s_1_2_2(mux_1561_nl, mux_1560_nl, fsm_output[6]);
  assign nor_1160_nl = ~((fsm_output[8]) | mux_1562_nl);
  assign nor_1161_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[10]));
  assign and_763_nl = (fsm_output[4]) & (fsm_output[2]) & (fsm_output[7]) & (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b0111)
      & (fsm_output[5]) & (~ (fsm_output[9])) & (fsm_output[10]);
  assign or_1341_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111)
      | (~ (fsm_output[10]));
  assign or_1339_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b0111) | (fsm_output[10]);
  assign mux_1557_nl = MUX_s_1_2_2(or_1341_nl, or_1339_nl, fsm_output[2]);
  assign nor_1163_nl = ~((fsm_output[4]) | mux_1557_nl);
  assign mux_1558_nl = MUX_s_1_2_2(and_763_nl, nor_1163_nl, fsm_output[6]);
  assign mux_1559_nl = MUX_s_1_2_2(nor_1161_nl, mux_1558_nl, fsm_output[8]);
  assign mux_1563_nl = MUX_s_1_2_2(nor_1160_nl, mux_1559_nl, fsm_output[0]);
  assign mux_1572_nl = MUX_s_1_2_2(mux_1571_nl, mux_1563_nl, fsm_output[3]);
  assign vec_rsc_0_7_i_wea_d_pff = MUX_s_1_2_2(mux_1586_nl, mux_1572_nl, fsm_output[1]);
  assign or_1447_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0111) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1446_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0111) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1617_nl = MUX_s_1_2_2(or_1447_nl, or_1446_nl, fsm_output[5]);
  assign nor_1120_nl = ~((fsm_output[1]) | mux_1617_nl);
  assign nor_1121_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0111)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1122_nl = ~((z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1123_nl = ~((z_out_2_12_1[3:0]!=4'b0111) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1615_nl = MUX_s_1_2_2(nor_1122_nl, nor_1123_nl, fsm_output[5]);
  assign mux_1616_nl = MUX_s_1_2_2(nor_1121_nl, mux_1615_nl, fsm_output[1]);
  assign mux_1618_nl = MUX_s_1_2_2(nor_1120_nl, mux_1616_nl, fsm_output[0]);
  assign and_593_nl = (fsm_output[6]) & mux_1618_nl;
  assign nor_1124_nl = ~((z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1126_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1610_nl = MUX_s_1_2_2(nor_1445_cse, nor_1126_nl, fsm_output[5]);
  assign nor_1127_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0111)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nand_295_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b0111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1611_nl = MUX_s_1_2_2(mux_1610_nl, nor_1127_nl, nand_295_nl);
  assign mux_1612_nl = MUX_s_1_2_2(nor_1124_nl, mux_1611_nl, fsm_output[1]);
  assign nor_1128_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b01) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1129_nl = ~((z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1130_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1608_nl = MUX_s_1_2_2(nor_1129_nl, nor_1130_nl, fsm_output[5]);
  assign mux_1609_nl = MUX_s_1_2_2(nor_1128_nl, mux_1608_nl, fsm_output[1]);
  assign mux_1613_nl = MUX_s_1_2_2(mux_1612_nl, mux_1609_nl, fsm_output[0]);
  assign nor_1131_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b0111) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1132_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b0111) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1606_nl = MUX_s_1_2_2(nor_1131_nl, nor_1132_nl, fsm_output[1]);
  assign nor_1133_nl = ~(nand_324_cse | mux_1413_cse);
  assign mux_1607_nl = MUX_s_1_2_2(mux_1606_nl, nor_1133_nl, fsm_output[0]);
  assign mux_1614_nl = MUX_s_1_2_2(mux_1613_nl, mux_1607_nl, fsm_output[6]);
  assign mux_1619_nl = MUX_s_1_2_2(and_593_nl, mux_1614_nl, fsm_output[8]);
  assign nor_1134_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b0111) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1135_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b0111) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1600_nl = MUX_s_1_2_2(nor_1134_nl, nor_1135_nl, fsm_output[5]);
  assign and_594_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1600_nl;
  assign nor_1136_nl = ~((~((fsm_output[7]) & (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b0111)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_1137_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b0111) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1599_nl = MUX_s_1_2_2(nor_1136_nl, nor_1137_nl, fsm_output[5]);
  assign and_595_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1599_nl;
  assign mux_1601_nl = MUX_s_1_2_2(and_594_nl, and_595_nl, fsm_output[1]);
  assign nor_1138_nl = ~((VEC_LOOP_j_sva_11_0[3]) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1139_nl = ~(nand_332_cse | mux_1533_cse);
  assign mux_1598_nl = MUX_s_1_2_2(nor_1138_nl, nor_1139_nl, fsm_output[1]);
  assign mux_1602_nl = MUX_s_1_2_2(mux_1601_nl, mux_1598_nl, fsm_output[0]);
  assign nor_1140_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1141_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b0111) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign and_596_nl = (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b011) & (fsm_output[7])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign mux_1595_nl = MUX_s_1_2_2(nor_1141_nl, and_596_nl, fsm_output[1]);
  assign mux_1596_nl = MUX_s_1_2_2(nor_1140_nl, mux_1595_nl, fsm_output[0]);
  assign mux_1603_nl = MUX_s_1_2_2(mux_1602_nl, mux_1596_nl, fsm_output[6]);
  assign nor_1142_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b0111) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1143_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b0111)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1593_nl = MUX_s_1_2_2(nor_1142_nl, nor_1143_nl, fsm_output[0]);
  assign nor_1144_nl = ~((~((fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b0111)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_1145_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b0111)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1146_nl = ~((~((fsm_output[7]) & (z_out_2_12_1[3:0]==4'b0111) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign mux_1589_nl = MUX_s_1_2_2(nor_1145_nl, nor_1146_nl, fsm_output[5]);
  assign mux_1590_nl = MUX_s_1_2_2(nor_1144_nl, mux_1589_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1147_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b0111)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1591_nl = MUX_s_1_2_2(mux_1590_nl, nor_1147_nl, fsm_output[1]);
  assign and_597_nl = (z_out_2_12_1[3:0]==4'b0111) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (~ (fsm_output[10]));
  assign nor_1148_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b011) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1588_nl = MUX_s_1_2_2(and_597_nl, nor_1148_nl, fsm_output[1]);
  assign mux_1592_nl = MUX_s_1_2_2(mux_1591_nl, mux_1588_nl, fsm_output[0]);
  assign mux_1594_nl = MUX_s_1_2_2(mux_1593_nl, mux_1592_nl, fsm_output[6]);
  assign mux_1604_nl = MUX_s_1_2_2(mux_1603_nl, mux_1594_nl, fsm_output[8]);
  assign vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1619_nl,
      mux_1604_nl, fsm_output[4]);
  assign or_1502_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1501_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000)
      | not_tmp_318;
  assign mux_1646_nl = MUX_s_1_2_2(or_1502_nl, or_1501_nl, fsm_output[7]);
  assign or_1499_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b10) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1647_nl = MUX_s_1_2_2(mux_1646_nl, or_1499_nl, fsm_output[2]);
  assign nor_1105_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1647_nl);
  assign nor_1106_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000)
      | not_tmp_318);
  assign mux_1648_nl = MUX_s_1_2_2(nor_1105_nl, nor_1106_nl, fsm_output[8]);
  assign nor_1107_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1108_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000)
      | (fsm_output[10]));
  assign nor_1109_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000) | (fsm_output[10]));
  assign nor_1110_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1643_nl = MUX_s_1_2_2(nor_1109_nl, nor_1110_nl, fsm_output[4]);
  assign mux_1644_nl = MUX_s_1_2_2(nor_1108_nl, mux_1643_nl, fsm_output[6]);
  assign mux_1645_nl = MUX_s_1_2_2(nor_1107_nl, mux_1644_nl, fsm_output[8]);
  assign mux_1649_nl = MUX_s_1_2_2(mux_1648_nl, mux_1645_nl, fsm_output[0]);
  assign or_1490_nl = (~ (COMP_LOOP_acc_16_psp_sva[0])) | (~ (fsm_output[4])) | (~
      (fsm_output[2])) | (VEC_LOOP_j_sva_11_0[2]) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1489_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1640_nl = MUX_s_1_2_2(mux_tmp_1628, or_1489_nl, fsm_output[4]);
  assign mux_1641_nl = MUX_s_1_2_2(or_1490_nl, mux_1640_nl, fsm_output[6]);
  assign and_592_nl = (fsm_output[8]) & (~ mux_1641_nl);
  assign or_1486_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_1484_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000) | not_tmp_318;
  assign mux_1637_nl = MUX_s_1_2_2(or_1484_nl, or_tmp_1416, fsm_output[2]);
  assign mux_1638_nl = MUX_s_1_2_2(or_1486_nl, mux_1637_nl, fsm_output[4]);
  assign nor_1111_nl = ~((fsm_output[6]) | mux_1638_nl);
  assign nor_1112_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1639_nl = MUX_s_1_2_2(nor_1111_nl, nor_1112_nl, fsm_output[8]);
  assign mux_1642_nl = MUX_s_1_2_2(and_592_nl, mux_1639_nl, fsm_output[0]);
  assign mux_1650_nl = MUX_s_1_2_2(mux_1649_nl, mux_1642_nl, fsm_output[3]);
  assign or_1480_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[0]) | nand_337_cse;
  assign or_1478_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000) | not_tmp_318;
  assign mux_1633_nl = MUX_s_1_2_2(or_1480_nl, or_1478_nl, fsm_output[4]);
  assign nor_1113_nl = ~((fsm_output[6]) | mux_1633_nl);
  assign or_1474_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000)
      | not_tmp_318;
  assign mux_1631_nl = MUX_s_1_2_2(or_591_cse, or_1474_nl, fsm_output[7]);
  assign mux_1632_nl = MUX_s_1_2_2(mux_1631_nl, or_tmp_1416, or_1470_cse);
  assign nor_1114_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1632_nl);
  assign mux_1634_nl = MUX_s_1_2_2(nor_1113_nl, nor_1114_nl, fsm_output[8]);
  assign or_1467_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1465_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1629_nl = MUX_s_1_2_2(or_1467_nl, or_1465_nl, fsm_output[2]);
  assign mux_1630_nl = MUX_s_1_2_2(mux_1629_nl, mux_tmp_1628, fsm_output[4]);
  assign nor_1115_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1630_nl);
  assign mux_1635_nl = MUX_s_1_2_2(mux_1634_nl, nor_1115_nl, fsm_output[0]);
  assign or_1460_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1458_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000) | (fsm_output[10]);
  assign mux_1625_nl = MUX_s_1_2_2(or_1460_nl, or_1458_nl, fsm_output[4]);
  assign or_1457_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9])) | (~
      (fsm_output[5])) | (fsm_output[10]);
  assign or_1456_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000) | (fsm_output[10]);
  assign mux_1624_nl = MUX_s_1_2_2(or_1457_nl, or_1456_nl, fsm_output[4]);
  assign mux_1626_nl = MUX_s_1_2_2(mux_1625_nl, mux_1624_nl, fsm_output[6]);
  assign nor_1116_nl = ~((fsm_output[8]) | mux_1626_nl);
  assign nor_1117_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1118_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (fsm_output[9]) | not_tmp_248);
  assign or_1451_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b000)
      | not_tmp_318;
  assign or_1449_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1000) | (fsm_output[10]);
  assign mux_1621_nl = MUX_s_1_2_2(or_1451_nl, or_1449_nl, fsm_output[2]);
  assign nor_1119_nl = ~((fsm_output[4]) | mux_1621_nl);
  assign mux_1622_nl = MUX_s_1_2_2(nor_1118_nl, nor_1119_nl, fsm_output[6]);
  assign mux_1623_nl = MUX_s_1_2_2(nor_1117_nl, mux_1622_nl, fsm_output[8]);
  assign mux_1627_nl = MUX_s_1_2_2(nor_1116_nl, mux_1623_nl, fsm_output[0]);
  assign mux_1636_nl = MUX_s_1_2_2(mux_1635_nl, mux_1627_nl, fsm_output[3]);
  assign vec_rsc_0_8_i_wea_d_pff = MUX_s_1_2_2(mux_1650_nl, mux_1636_nl, fsm_output[1]);
  assign or_1558_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1000) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1557_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1000) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1681_nl = MUX_s_1_2_2(or_1558_nl, or_1557_nl, fsm_output[5]);
  assign nor_1074_nl = ~((fsm_output[1]) | mux_1681_nl);
  assign nor_1075_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1000)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1076_nl = ~((z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1077_nl = ~((z_out_2_12_1[3:0]!=4'b1000) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1679_nl = MUX_s_1_2_2(nor_1076_nl, nor_1077_nl, fsm_output[5]);
  assign mux_1680_nl = MUX_s_1_2_2(nor_1075_nl, mux_1679_nl, fsm_output[1]);
  assign mux_1682_nl = MUX_s_1_2_2(nor_1074_nl, mux_1680_nl, fsm_output[0]);
  assign and_589_nl = (fsm_output[6]) & mux_1682_nl;
  assign nor_1078_nl = ~((z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1080_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1674_nl = MUX_s_1_2_2(nor_1445_cse, nor_1080_nl, fsm_output[5]);
  assign nor_1081_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1544_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1000) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1675_nl = MUX_s_1_2_2(mux_1674_nl, nor_1081_nl, or_1544_nl);
  assign mux_1676_nl = MUX_s_1_2_2(nor_1078_nl, mux_1675_nl, fsm_output[1]);
  assign nor_1082_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1083_nl = ~((z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1084_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1672_nl = MUX_s_1_2_2(nor_1083_nl, nor_1084_nl, fsm_output[5]);
  assign mux_1673_nl = MUX_s_1_2_2(nor_1082_nl, mux_1672_nl, fsm_output[1]);
  assign mux_1677_nl = MUX_s_1_2_2(mux_1676_nl, mux_1673_nl, fsm_output[0]);
  assign nor_1085_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1000) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1086_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1000) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1670_nl = MUX_s_1_2_2(nor_1085_nl, nor_1086_nl, fsm_output[1]);
  assign nor_1087_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1669_cse);
  assign mux_1671_nl = MUX_s_1_2_2(mux_1670_nl, nor_1087_nl, fsm_output[0]);
  assign mux_1678_nl = MUX_s_1_2_2(mux_1677_nl, mux_1671_nl, fsm_output[6]);
  assign mux_1683_nl = MUX_s_1_2_2(and_589_nl, mux_1678_nl, fsm_output[8]);
  assign nor_1088_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1000) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1089_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1000) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1664_nl = MUX_s_1_2_2(nor_1088_nl, nor_1089_nl, fsm_output[5]);
  assign and_590_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1664_nl;
  assign nor_1090_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1091_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1000) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1663_nl = MUX_s_1_2_2(nor_1090_nl, nor_1091_nl, fsm_output[5]);
  assign and_591_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1663_nl;
  assign mux_1665_nl = MUX_s_1_2_2(and_590_nl, and_591_nl, fsm_output[1]);
  assign nor_1092_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (VEC_LOOP_j_sva_11_0[1])
      | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1093_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1661_cse);
  assign mux_1662_nl = MUX_s_1_2_2(nor_1092_nl, nor_1093_nl, fsm_output[1]);
  assign mux_1666_nl = MUX_s_1_2_2(mux_1665_nl, mux_1662_nl, fsm_output[0]);
  assign nor_1094_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1095_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1096_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1659_nl = MUX_s_1_2_2(nor_1095_nl, nor_1096_nl, fsm_output[1]);
  assign mux_1660_nl = MUX_s_1_2_2(nor_1094_nl, mux_1659_nl, fsm_output[0]);
  assign mux_1667_nl = MUX_s_1_2_2(mux_1666_nl, mux_1660_nl, fsm_output[6]);
  assign nor_1097_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1000) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1098_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1000)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1657_nl = MUX_s_1_2_2(nor_1097_nl, nor_1098_nl, fsm_output[0]);
  assign nor_1099_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1000)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1100_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1000)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1101_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1000) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1653_nl = MUX_s_1_2_2(nor_1100_nl, nor_1101_nl, fsm_output[5]);
  assign mux_1654_nl = MUX_s_1_2_2(nor_1099_nl, mux_1653_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1102_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1000)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1655_nl = MUX_s_1_2_2(mux_1654_nl, nor_1102_nl, fsm_output[1]);
  assign nor_1103_nl = ~((z_out_2_12_1[3:0]!=4'b1000) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1104_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1652_nl = MUX_s_1_2_2(nor_1103_nl, nor_1104_nl, fsm_output[1]);
  assign mux_1656_nl = MUX_s_1_2_2(mux_1655_nl, mux_1652_nl, fsm_output[0]);
  assign mux_1658_nl = MUX_s_1_2_2(mux_1657_nl, mux_1656_nl, fsm_output[6]);
  assign mux_1668_nl = MUX_s_1_2_2(mux_1667_nl, mux_1658_nl, fsm_output[8]);
  assign vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1683_nl,
      mux_1668_nl, fsm_output[4]);
  assign or_1613_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1612_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001)
      | not_tmp_318;
  assign mux_1710_nl = MUX_s_1_2_2(or_1613_nl, or_1612_nl, fsm_output[7]);
  assign or_1610_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b10) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1711_nl = MUX_s_1_2_2(mux_1710_nl, or_1610_nl, fsm_output[2]);
  assign nor_1059_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1711_nl);
  assign nor_1060_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001)
      | not_tmp_318);
  assign mux_1712_nl = MUX_s_1_2_2(nor_1059_nl, nor_1060_nl, fsm_output[8]);
  assign nor_1061_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_1062_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001)
      | (fsm_output[10]));
  assign nor_1063_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001) | (fsm_output[10]));
  assign nor_1064_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1707_nl = MUX_s_1_2_2(nor_1063_nl, nor_1064_nl, fsm_output[4]);
  assign mux_1708_nl = MUX_s_1_2_2(nor_1062_nl, mux_1707_nl, fsm_output[6]);
  assign mux_1709_nl = MUX_s_1_2_2(nor_1061_nl, mux_1708_nl, fsm_output[8]);
  assign mux_1713_nl = MUX_s_1_2_2(mux_1712_nl, mux_1709_nl, fsm_output[0]);
  assign nand_287_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (~ (VEC_LOOP_j_sva_11_0[2])) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b01)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_1600_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1704_nl = MUX_s_1_2_2(mux_tmp_1692, or_1600_nl, fsm_output[4]);
  assign mux_1705_nl = MUX_s_1_2_2(nand_287_nl, mux_1704_nl, fsm_output[6]);
  assign and_588_nl = (fsm_output[8]) & (~ mux_1705_nl);
  assign or_1597_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1001) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_1595_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001) | not_tmp_318;
  assign mux_1701_nl = MUX_s_1_2_2(or_1595_nl, or_tmp_1527, fsm_output[2]);
  assign mux_1702_nl = MUX_s_1_2_2(or_1597_nl, mux_1701_nl, fsm_output[4]);
  assign nor_1065_nl = ~((fsm_output[6]) | mux_1702_nl);
  assign nor_1066_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1703_nl = MUX_s_1_2_2(nor_1065_nl, nor_1066_nl, fsm_output[8]);
  assign mux_1706_nl = MUX_s_1_2_2(and_588_nl, mux_1703_nl, fsm_output[0]);
  assign mux_1714_nl = MUX_s_1_2_2(mux_1713_nl, mux_1706_nl, fsm_output[3]);
  assign or_1591_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_1589_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001) | not_tmp_318;
  assign mux_1697_nl = MUX_s_1_2_2(or_1591_nl, or_1589_nl, fsm_output[4]);
  assign nor_1067_nl = ~((fsm_output[6]) | mux_1697_nl);
  assign or_1585_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001)
      | not_tmp_318;
  assign mux_1695_nl = MUX_s_1_2_2(or_702_cse, or_1585_nl, fsm_output[7]);
  assign mux_1696_nl = MUX_s_1_2_2(mux_1695_nl, or_tmp_1527, or_1470_cse);
  assign nor_1068_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1696_nl);
  assign mux_1698_nl = MUX_s_1_2_2(nor_1067_nl, nor_1068_nl, fsm_output[8]);
  assign or_1578_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1576_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1693_nl = MUX_s_1_2_2(or_1578_nl, or_1576_nl, fsm_output[2]);
  assign mux_1694_nl = MUX_s_1_2_2(mux_1693_nl, mux_tmp_1692, fsm_output[4]);
  assign nor_1069_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1694_nl);
  assign mux_1699_nl = MUX_s_1_2_2(mux_1698_nl, nor_1069_nl, fsm_output[0]);
  assign or_1571_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b100) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1569_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001) | (fsm_output[10]);
  assign mux_1689_nl = MUX_s_1_2_2(or_1571_nl, or_1569_nl, fsm_output[4]);
  assign or_1568_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b100) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[9]))
      | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1567_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001) | (fsm_output[10]);
  assign mux_1688_nl = MUX_s_1_2_2(or_1568_nl, or_1567_nl, fsm_output[4]);
  assign mux_1690_nl = MUX_s_1_2_2(mux_1689_nl, mux_1688_nl, fsm_output[6]);
  assign nor_1070_nl = ~((fsm_output[8]) | mux_1690_nl);
  assign nor_1071_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_1072_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (fsm_output[9]) | not_tmp_248);
  assign or_1562_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b001)
      | not_tmp_318;
  assign or_1560_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1001) | (fsm_output[10]);
  assign mux_1685_nl = MUX_s_1_2_2(or_1562_nl, or_1560_nl, fsm_output[2]);
  assign nor_1073_nl = ~((fsm_output[4]) | mux_1685_nl);
  assign mux_1686_nl = MUX_s_1_2_2(nor_1072_nl, nor_1073_nl, fsm_output[6]);
  assign mux_1687_nl = MUX_s_1_2_2(nor_1071_nl, mux_1686_nl, fsm_output[8]);
  assign mux_1691_nl = MUX_s_1_2_2(nor_1070_nl, mux_1687_nl, fsm_output[0]);
  assign mux_1700_nl = MUX_s_1_2_2(mux_1699_nl, mux_1691_nl, fsm_output[3]);
  assign vec_rsc_0_9_i_wea_d_pff = MUX_s_1_2_2(mux_1714_nl, mux_1700_nl, fsm_output[1]);
  assign or_1669_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1001) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1668_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1001) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1745_nl = MUX_s_1_2_2(or_1669_nl, or_1668_nl, fsm_output[5]);
  assign nor_1028_nl = ~((fsm_output[1]) | mux_1745_nl);
  assign nor_1029_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1001)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1030_nl = ~((z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1031_nl = ~((z_out_2_12_1[3:0]!=4'b1001) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1743_nl = MUX_s_1_2_2(nor_1030_nl, nor_1031_nl, fsm_output[5]);
  assign mux_1744_nl = MUX_s_1_2_2(nor_1029_nl, mux_1743_nl, fsm_output[1]);
  assign mux_1746_nl = MUX_s_1_2_2(nor_1028_nl, mux_1744_nl, fsm_output[0]);
  assign and_585_nl = (fsm_output[6]) & mux_1746_nl;
  assign nor_1032_nl = ~((z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1034_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1738_nl = MUX_s_1_2_2(nor_1445_cse, nor_1034_nl, fsm_output[5]);
  assign nor_1035_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1655_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1001) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1739_nl = MUX_s_1_2_2(mux_1738_nl, nor_1035_nl, or_1655_nl);
  assign mux_1740_nl = MUX_s_1_2_2(nor_1032_nl, mux_1739_nl, fsm_output[1]);
  assign nor_1036_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_1037_nl = ~((z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_1038_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1736_nl = MUX_s_1_2_2(nor_1037_nl, nor_1038_nl, fsm_output[5]);
  assign mux_1737_nl = MUX_s_1_2_2(nor_1036_nl, mux_1736_nl, fsm_output[1]);
  assign mux_1741_nl = MUX_s_1_2_2(mux_1740_nl, mux_1737_nl, fsm_output[0]);
  assign nor_1039_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1001) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_1040_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1001) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1734_nl = MUX_s_1_2_2(nor_1039_nl, nor_1040_nl, fsm_output[1]);
  assign nor_1041_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1669_cse);
  assign mux_1735_nl = MUX_s_1_2_2(mux_1734_nl, nor_1041_nl, fsm_output[0]);
  assign mux_1742_nl = MUX_s_1_2_2(mux_1741_nl, mux_1735_nl, fsm_output[6]);
  assign mux_1747_nl = MUX_s_1_2_2(and_585_nl, mux_1742_nl, fsm_output[8]);
  assign nor_1042_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1001) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1043_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1001) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1728_nl = MUX_s_1_2_2(nor_1042_nl, nor_1043_nl, fsm_output[5]);
  assign and_586_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1728_nl;
  assign nor_1044_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1045_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1001) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1727_nl = MUX_s_1_2_2(nor_1044_nl, nor_1045_nl, fsm_output[5]);
  assign and_587_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1727_nl;
  assign mux_1729_nl = MUX_s_1_2_2(and_586_nl, and_587_nl, fsm_output[1]);
  assign nor_1046_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (VEC_LOOP_j_sva_11_0[1])
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1047_nl = ~(nand_332_cse | mux_1661_cse);
  assign mux_1726_nl = MUX_s_1_2_2(nor_1046_nl, nor_1047_nl, fsm_output[1]);
  assign mux_1730_nl = MUX_s_1_2_2(mux_1729_nl, mux_1726_nl, fsm_output[0]);
  assign nor_1048_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1049_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1050_nl = ~((~ (VEC_LOOP_j_sva_11_0[0])) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b100) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1723_nl = MUX_s_1_2_2(nor_1049_nl, nor_1050_nl, fsm_output[1]);
  assign mux_1724_nl = MUX_s_1_2_2(nor_1048_nl, mux_1723_nl, fsm_output[0]);
  assign mux_1731_nl = MUX_s_1_2_2(mux_1730_nl, mux_1724_nl, fsm_output[6]);
  assign nor_1051_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1001) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1052_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1001)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1721_nl = MUX_s_1_2_2(nor_1051_nl, nor_1052_nl, fsm_output[0]);
  assign nor_1053_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1001)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1054_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1001)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1055_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1001) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1717_nl = MUX_s_1_2_2(nor_1054_nl, nor_1055_nl, fsm_output[5]);
  assign mux_1718_nl = MUX_s_1_2_2(nor_1053_nl, mux_1717_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1056_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1001)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1719_nl = MUX_s_1_2_2(mux_1718_nl, nor_1056_nl, fsm_output[1]);
  assign nor_1057_nl = ~((z_out_2_12_1[3:0]!=4'b1001) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1058_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b100) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1716_nl = MUX_s_1_2_2(nor_1057_nl, nor_1058_nl, fsm_output[1]);
  assign mux_1720_nl = MUX_s_1_2_2(mux_1719_nl, mux_1716_nl, fsm_output[0]);
  assign mux_1722_nl = MUX_s_1_2_2(mux_1721_nl, mux_1720_nl, fsm_output[6]);
  assign mux_1732_nl = MUX_s_1_2_2(mux_1731_nl, mux_1722_nl, fsm_output[8]);
  assign vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1747_nl,
      mux_1732_nl, fsm_output[4]);
  assign or_1723_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b10) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b01);
  assign or_1722_nl = (~ (fsm_output[5])) | (~ (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010)
      | not_tmp_318;
  assign mux_1774_nl = MUX_s_1_2_2(or_1723_nl, or_1722_nl, fsm_output[7]);
  assign or_1720_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b10) | (~ (fsm_output[7])) | (~
      (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[5]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b00);
  assign mux_1775_nl = MUX_s_1_2_2(mux_1774_nl, or_1720_nl, fsm_output[2]);
  assign nor_1013_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1775_nl);
  assign nor_1014_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010)
      | not_tmp_318);
  assign mux_1776_nl = MUX_s_1_2_2(nor_1013_nl, nor_1014_nl, fsm_output[8]);
  assign nor_1015_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (~ (fsm_output[10])));
  assign nor_1016_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (fsm_output[5])
      | (~ (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010) | (fsm_output[10]));
  assign nor_1017_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010) | (fsm_output[10]));
  assign nor_1018_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[10]));
  assign mux_1771_nl = MUX_s_1_2_2(nor_1017_nl, nor_1018_nl, fsm_output[4]);
  assign mux_1772_nl = MUX_s_1_2_2(nor_1016_nl, mux_1771_nl, fsm_output[6]);
  assign mux_1773_nl = MUX_s_1_2_2(nor_1015_nl, mux_1772_nl, fsm_output[8]);
  assign mux_1777_nl = MUX_s_1_2_2(mux_1776_nl, mux_1773_nl, fsm_output[0]);
  assign nand_282_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (~ (VEC_LOOP_j_sva_11_0[2])) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1])
      & (fsm_output[5]) & (~ (VEC_LOOP_j_sva_11_0[0])) & (fsm_output[10:9]==2'b01));
  assign or_1710_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[2]) |
      (fsm_output[7]) | (~ (VEC_LOOP_j_sva_11_0[1])) | (fsm_output[5]) | (VEC_LOOP_j_sva_11_0[0])
      | (fsm_output[10:9]!=2'b10);
  assign mux_1768_nl = MUX_s_1_2_2(mux_tmp_1756, or_1710_nl, fsm_output[4]);
  assign mux_1769_nl = MUX_s_1_2_2(nand_282_nl, mux_1768_nl, fsm_output[6]);
  assign and_584_nl = (fsm_output[8]) & (~ mux_1769_nl);
  assign or_1707_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (fsm_output[5]) | nand_358_cse;
  assign or_1705_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010) | not_tmp_318;
  assign mux_1765_nl = MUX_s_1_2_2(or_1705_nl, or_tmp_1640, fsm_output[2]);
  assign mux_1766_nl = MUX_s_1_2_2(or_1707_nl, mux_1765_nl, fsm_output[4]);
  assign nor_1019_nl = ~((fsm_output[6]) | mux_1766_nl);
  assign nor_1020_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[10]));
  assign mux_1767_nl = MUX_s_1_2_2(nor_1019_nl, nor_1020_nl, fsm_output[8]);
  assign mux_1770_nl = MUX_s_1_2_2(and_584_nl, mux_1767_nl, fsm_output[0]);
  assign mux_1778_nl = MUX_s_1_2_2(mux_1777_nl, mux_1770_nl, fsm_output[3]);
  assign or_1701_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | nand_358_cse;
  assign or_1699_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010) | not_tmp_318;
  assign mux_1761_nl = MUX_s_1_2_2(or_1701_nl, or_1699_nl, fsm_output[4]);
  assign nor_1021_nl = ~((fsm_output[6]) | mux_1761_nl);
  assign or_1693_nl = (fsm_output[5]) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010)
      | not_tmp_318;
  assign mux_1759_nl = MUX_s_1_2_2(or_591_cse, or_1693_nl, fsm_output[7]);
  assign mux_1760_nl = MUX_s_1_2_2(or_tmp_1640, mux_1759_nl, nor_239_cse);
  assign nor_1022_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1760_nl);
  assign mux_1762_nl = MUX_s_1_2_2(nor_1021_nl, nor_1022_nl, fsm_output[8]);
  assign or_1689_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010) | (fsm_output[7])
      | (~ (fsm_output[5])) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign or_1687_nl = (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (~ (fsm_output[7]))
      | (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[10]);
  assign mux_1757_nl = MUX_s_1_2_2(or_1689_nl, or_1687_nl, fsm_output[2]);
  assign mux_1758_nl = MUX_s_1_2_2(mux_1757_nl, mux_tmp_1756, fsm_output[4]);
  assign nor_1023_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1758_nl);
  assign mux_1763_nl = MUX_s_1_2_2(mux_1762_nl, nor_1023_nl, fsm_output[0]);
  assign or_1682_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (fsm_output[5]) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b10);
  assign or_1680_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[5]) | (~
      (fsm_output[9])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010) | (fsm_output[10]);
  assign mux_1753_nl = MUX_s_1_2_2(or_1682_nl, or_1680_nl, fsm_output[4]);
  assign or_1679_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b101) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[10:9]!=2'b01);
  assign or_1678_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010) | (fsm_output[10]);
  assign mux_1752_nl = MUX_s_1_2_2(or_1679_nl, or_1678_nl, fsm_output[4]);
  assign mux_1754_nl = MUX_s_1_2_2(mux_1753_nl, mux_1752_nl, fsm_output[6]);
  assign nor_1024_nl = ~((fsm_output[8]) | mux_1754_nl);
  assign nor_1025_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (fsm_output[10]));
  assign and_761_nl = (fsm_output[4]) & (fsm_output[2]) & (fsm_output[7]) & (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1010)
      & (fsm_output[5]) & (~ (fsm_output[9])) & (fsm_output[10]);
  assign or_1673_nl = (fsm_output[7]) | (~ (fsm_output[5])) | (fsm_output[9]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b010)
      | not_tmp_318;
  assign or_1671_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (~ (fsm_output[9]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1010) | (fsm_output[10]);
  assign mux_1749_nl = MUX_s_1_2_2(or_1673_nl, or_1671_nl, fsm_output[2]);
  assign nor_1027_nl = ~((fsm_output[4]) | mux_1749_nl);
  assign mux_1750_nl = MUX_s_1_2_2(and_761_nl, nor_1027_nl, fsm_output[6]);
  assign mux_1751_nl = MUX_s_1_2_2(nor_1025_nl, mux_1750_nl, fsm_output[8]);
  assign mux_1755_nl = MUX_s_1_2_2(nor_1024_nl, mux_1751_nl, fsm_output[0]);
  assign mux_1764_nl = MUX_s_1_2_2(mux_1763_nl, mux_1755_nl, fsm_output[3]);
  assign vec_rsc_0_10_i_wea_d_pff = MUX_s_1_2_2(mux_1778_nl, mux_1764_nl, fsm_output[1]);
  assign or_1779_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1010) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1778_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1010) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1809_nl = MUX_s_1_2_2(or_1779_nl, or_1778_nl, fsm_output[5]);
  assign nor_982_nl = ~((fsm_output[1]) | mux_1809_nl);
  assign nor_983_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1010)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_984_nl = ~((z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_985_nl = ~((z_out_2_12_1[3:0]!=4'b1010) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1807_nl = MUX_s_1_2_2(nor_984_nl, nor_985_nl, fsm_output[5]);
  assign mux_1808_nl = MUX_s_1_2_2(nor_983_nl, mux_1807_nl, fsm_output[1]);
  assign mux_1810_nl = MUX_s_1_2_2(nor_982_nl, mux_1808_nl, fsm_output[0]);
  assign and_581_nl = (fsm_output[6]) & mux_1810_nl;
  assign nor_986_nl = ~((z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_988_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1802_nl = MUX_s_1_2_2(nor_1445_cse, nor_988_nl, fsm_output[5]);
  assign nor_989_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1765_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1010) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1803_nl = MUX_s_1_2_2(mux_1802_nl, nor_989_nl, or_1765_nl);
  assign mux_1804_nl = MUX_s_1_2_2(nor_986_nl, mux_1803_nl, fsm_output[1]);
  assign nor_990_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_991_nl = ~((z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_992_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1800_nl = MUX_s_1_2_2(nor_991_nl, nor_992_nl, fsm_output[5]);
  assign mux_1801_nl = MUX_s_1_2_2(nor_990_nl, mux_1800_nl, fsm_output[1]);
  assign mux_1805_nl = MUX_s_1_2_2(mux_1804_nl, mux_1801_nl, fsm_output[0]);
  assign nor_993_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1010) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_994_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1010) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1798_nl = MUX_s_1_2_2(nor_993_nl, nor_994_nl, fsm_output[1]);
  assign nor_995_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1669_cse);
  assign mux_1799_nl = MUX_s_1_2_2(mux_1798_nl, nor_995_nl, fsm_output[0]);
  assign mux_1806_nl = MUX_s_1_2_2(mux_1805_nl, mux_1799_nl, fsm_output[6]);
  assign mux_1811_nl = MUX_s_1_2_2(and_581_nl, mux_1806_nl, fsm_output[8]);
  assign nor_996_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1010) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_997_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1010) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1792_nl = MUX_s_1_2_2(nor_996_nl, nor_997_nl, fsm_output[5]);
  assign and_582_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1792_nl;
  assign nor_998_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_999_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1010) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1791_nl = MUX_s_1_2_2(nor_998_nl, nor_999_nl, fsm_output[5]);
  assign and_583_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1791_nl;
  assign mux_1793_nl = MUX_s_1_2_2(and_582_nl, and_583_nl, fsm_output[1]);
  assign nor_1000_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1001_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1789_cse);
  assign mux_1790_nl = MUX_s_1_2_2(nor_1000_nl, nor_1001_nl, fsm_output[1]);
  assign mux_1794_nl = MUX_s_1_2_2(mux_1793_nl, mux_1790_nl, fsm_output[0]);
  assign nor_1002_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7])
      | (z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1003_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3]))
      | (z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[10]));
  assign nor_1004_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b101) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1787_nl = MUX_s_1_2_2(nor_1003_nl, nor_1004_nl, fsm_output[1]);
  assign mux_1788_nl = MUX_s_1_2_2(nor_1002_nl, mux_1787_nl, fsm_output[0]);
  assign mux_1795_nl = MUX_s_1_2_2(mux_1794_nl, mux_1788_nl, fsm_output[6]);
  assign nor_1005_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1010) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1006_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1010)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1785_nl = MUX_s_1_2_2(nor_1005_nl, nor_1006_nl, fsm_output[0]);
  assign nor_1007_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1010)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_1008_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1010)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_1009_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1010) | (~
      (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign mux_1781_nl = MUX_s_1_2_2(nor_1008_nl, nor_1009_nl, fsm_output[5]);
  assign mux_1782_nl = MUX_s_1_2_2(nor_1007_nl, mux_1781_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_1010_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1010)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1783_nl = MUX_s_1_2_2(mux_1782_nl, nor_1010_nl, fsm_output[1]);
  assign nor_1011_nl = ~((z_out_2_12_1[3:0]!=4'b1010) | (~ (fsm_output[5])) | (~
      (fsm_output[7])) | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_1012_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1780_nl = MUX_s_1_2_2(nor_1011_nl, nor_1012_nl, fsm_output[1]);
  assign mux_1784_nl = MUX_s_1_2_2(mux_1783_nl, mux_1780_nl, fsm_output[0]);
  assign mux_1786_nl = MUX_s_1_2_2(mux_1785_nl, mux_1784_nl, fsm_output[6]);
  assign mux_1796_nl = MUX_s_1_2_2(mux_1795_nl, mux_1786_nl, fsm_output[8]);
  assign vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1811_nl,
      mux_1796_nl, fsm_output[4]);
  assign nand_272_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b10) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_1832_nl = (~((fsm_output[9]) & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]==3'b011)))
      | not_tmp_318;
  assign mux_1838_nl = MUX_s_1_2_2(nand_272_nl, or_1832_nl, fsm_output[7]);
  assign or_1830_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b10) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1839_nl = MUX_s_1_2_2(mux_1838_nl, or_1830_nl, fsm_output[2]);
  assign nor_967_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1839_nl);
  assign nor_968_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2])) |
      (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011)
      | not_tmp_318);
  assign mux_1840_nl = MUX_s_1_2_2(nor_967_nl, nor_968_nl, fsm_output[8]);
  assign nor_969_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1011) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_970_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011)
      | (fsm_output[10]));
  assign nor_971_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) |
      (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011) | (fsm_output[10]));
  assign nor_972_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1011) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1835_nl = MUX_s_1_2_2(nor_971_nl, nor_972_nl, fsm_output[4]);
  assign mux_1836_nl = MUX_s_1_2_2(nor_970_nl, mux_1835_nl, fsm_output[6]);
  assign mux_1837_nl = MUX_s_1_2_2(nor_969_nl, mux_1836_nl, fsm_output[8]);
  assign mux_1841_nl = MUX_s_1_2_2(mux_1840_nl, mux_1837_nl, fsm_output[0]);
  assign nand_274_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (~ (VEC_LOOP_j_sva_11_0[2])) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_1820_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1832_nl = MUX_s_1_2_2(mux_tmp_1820, or_1820_nl, fsm_output[4]);
  assign mux_1833_nl = MUX_s_1_2_2(nand_274_nl, mux_1832_nl, fsm_output[6]);
  assign and_580_nl = (fsm_output[8]) & (~ mux_1833_nl);
  assign nand_398_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1011) & (fsm_output[2])
      & (fsm_output[7]) & (fsm_output[9]) & (~ (fsm_output[5])) & (fsm_output[10]));
  assign or_1815_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011) | not_tmp_318;
  assign mux_1829_nl = MUX_s_1_2_2(or_1815_nl, or_tmp_1750, fsm_output[2]);
  assign mux_1830_nl = MUX_s_1_2_2(nand_398_nl, mux_1829_nl, fsm_output[4]);
  assign nor_973_nl = ~((fsm_output[6]) | mux_1830_nl);
  assign nor_974_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1831_nl = MUX_s_1_2_2(nor_973_nl, nor_974_nl, fsm_output[8]);
  assign mux_1834_nl = MUX_s_1_2_2(and_580_nl, mux_1831_nl, fsm_output[0]);
  assign mux_1842_nl = MUX_s_1_2_2(mux_1841_nl, mux_1834_nl, fsm_output[3]);
  assign or_1811_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_1809_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011) | not_tmp_318;
  assign mux_1825_nl = MUX_s_1_2_2(or_1811_nl, or_1809_nl, fsm_output[4]);
  assign nor_975_nl = ~((fsm_output[6]) | mux_1825_nl);
  assign or_1803_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011)
      | not_tmp_318;
  assign mux_1823_nl = MUX_s_1_2_2(or_702_cse, or_1803_nl, fsm_output[7]);
  assign mux_1824_nl = MUX_s_1_2_2(or_tmp_1750, mux_1823_nl, nor_239_cse);
  assign nor_976_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1824_nl);
  assign mux_1826_nl = MUX_s_1_2_2(nor_975_nl, nor_976_nl, fsm_output[8]);
  assign or_1799_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1011) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1797_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1011)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1821_nl = MUX_s_1_2_2(or_1799_nl, or_1797_nl, fsm_output[2]);
  assign mux_1822_nl = MUX_s_1_2_2(mux_1821_nl, mux_tmp_1820, fsm_output[4]);
  assign nor_977_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1822_nl);
  assign mux_1827_nl = MUX_s_1_2_2(mux_1826_nl, nor_977_nl, fsm_output[0]);
  assign or_1792_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b101) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1790_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011) | (fsm_output[10]);
  assign mux_1817_nl = MUX_s_1_2_2(or_1792_nl, or_1790_nl, fsm_output[4]);
  assign nand_277_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b101) & (fsm_output[2])
      & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[9]) & (fsm_output[5])
      & (~ (fsm_output[10])));
  assign or_1788_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011) | (fsm_output[10]);
  assign mux_1816_nl = MUX_s_1_2_2(nand_277_nl, or_1788_nl, fsm_output[4]);
  assign mux_1818_nl = MUX_s_1_2_2(mux_1817_nl, mux_1816_nl, fsm_output[6]);
  assign nor_978_nl = ~((fsm_output[8]) | mux_1818_nl);
  assign nor_979_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_980_nl = ~((~((fsm_output[4]) & (fsm_output[2]) & (fsm_output[7]) &
      (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1011) & (~ (fsm_output[9])))) | not_tmp_248);
  assign or_1783_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[2:0]!=3'b011)
      | not_tmp_318;
  assign or_1781_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1011) | (fsm_output[10]);
  assign mux_1813_nl = MUX_s_1_2_2(or_1783_nl, or_1781_nl, fsm_output[2]);
  assign nor_981_nl = ~((fsm_output[4]) | mux_1813_nl);
  assign mux_1814_nl = MUX_s_1_2_2(nor_980_nl, nor_981_nl, fsm_output[6]);
  assign mux_1815_nl = MUX_s_1_2_2(nor_979_nl, mux_1814_nl, fsm_output[8]);
  assign mux_1819_nl = MUX_s_1_2_2(nor_978_nl, mux_1815_nl, fsm_output[0]);
  assign mux_1828_nl = MUX_s_1_2_2(mux_1827_nl, mux_1819_nl, fsm_output[3]);
  assign vec_rsc_0_11_i_wea_d_pff = MUX_s_1_2_2(mux_1842_nl, mux_1828_nl, fsm_output[1]);
  assign or_1889_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1011) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1888_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1011) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1873_nl = MUX_s_1_2_2(or_1889_nl, or_1888_nl, fsm_output[5]);
  assign nor_938_nl = ~((fsm_output[1]) | mux_1873_nl);
  assign nor_939_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1011)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_940_nl = ~((z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_941_nl = ~((z_out_2_12_1[3:0]!=4'b1011) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1871_nl = MUX_s_1_2_2(nor_940_nl, nor_941_nl, fsm_output[5]);
  assign mux_1872_nl = MUX_s_1_2_2(nor_939_nl, mux_1871_nl, fsm_output[1]);
  assign mux_1874_nl = MUX_s_1_2_2(nor_938_nl, mux_1872_nl, fsm_output[0]);
  assign and_575_nl = (fsm_output[6]) & mux_1874_nl;
  assign nor_942_nl = ~((z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_944_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1866_nl = MUX_s_1_2_2(nor_1445_cse, nor_944_nl, fsm_output[5]);
  assign nor_945_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1011)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nand_265_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1011) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1867_nl = MUX_s_1_2_2(mux_1866_nl, nor_945_nl, nand_265_nl);
  assign mux_1868_nl = MUX_s_1_2_2(nor_942_nl, mux_1867_nl, fsm_output[1]);
  assign nor_946_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b10) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_947_nl = ~((z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_948_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1864_nl = MUX_s_1_2_2(nor_947_nl, nor_948_nl, fsm_output[5]);
  assign mux_1865_nl = MUX_s_1_2_2(nor_946_nl, mux_1864_nl, fsm_output[1]);
  assign mux_1869_nl = MUX_s_1_2_2(mux_1868_nl, mux_1865_nl, fsm_output[0]);
  assign nor_949_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1011) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_950_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1011) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1862_nl = MUX_s_1_2_2(nor_949_nl, nor_950_nl, fsm_output[1]);
  assign nor_951_nl = ~(nand_324_cse | mux_1669_cse);
  assign mux_1863_nl = MUX_s_1_2_2(mux_1862_nl, nor_951_nl, fsm_output[0]);
  assign mux_1870_nl = MUX_s_1_2_2(mux_1869_nl, mux_1863_nl, fsm_output[6]);
  assign mux_1875_nl = MUX_s_1_2_2(and_575_nl, mux_1870_nl, fsm_output[8]);
  assign nor_952_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1011) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_953_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1011) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1856_nl = MUX_s_1_2_2(nor_952_nl, nor_953_nl, fsm_output[5]);
  assign and_576_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1856_nl;
  assign nor_954_nl = ~((~((fsm_output[7]) & (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1011)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_955_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1011) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1855_nl = MUX_s_1_2_2(nor_954_nl, nor_955_nl, fsm_output[5]);
  assign and_577_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1855_nl;
  assign mux_1857_nl = MUX_s_1_2_2(and_576_nl, and_577_nl, fsm_output[1]);
  assign nor_956_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (VEC_LOOP_j_sva_11_0[2])
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_957_nl = ~(nand_332_cse | mux_1789_cse);
  assign mux_1854_nl = MUX_s_1_2_2(nor_956_nl, nor_957_nl, fsm_output[1]);
  assign mux_1858_nl = MUX_s_1_2_2(mux_1857_nl, mux_1854_nl, fsm_output[0]);
  assign nor_958_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7]) |
      (z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_959_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3])) |
      (z_out_2_12_1[3:0]!=4'b1011) | (~ (fsm_output[9])) | (~ (fsm_output[2])) |
      (fsm_output[10]));
  assign and_578_nl = (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b101) & (fsm_output[7])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign mux_1851_nl = MUX_s_1_2_2(nor_959_nl, and_578_nl, fsm_output[1]);
  assign mux_1852_nl = MUX_s_1_2_2(nor_958_nl, mux_1851_nl, fsm_output[0]);
  assign mux_1859_nl = MUX_s_1_2_2(mux_1858_nl, mux_1852_nl, fsm_output[6]);
  assign nor_960_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1011) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_961_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1011)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1849_nl = MUX_s_1_2_2(nor_960_nl, nor_961_nl, fsm_output[0]);
  assign nor_962_nl = ~((~((fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1011)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_963_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1011)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_964_nl = ~((~((fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1011) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign mux_1845_nl = MUX_s_1_2_2(nor_963_nl, nor_964_nl, fsm_output[5]);
  assign mux_1846_nl = MUX_s_1_2_2(nor_962_nl, mux_1845_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_965_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1011)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1847_nl = MUX_s_1_2_2(mux_1846_nl, nor_965_nl, fsm_output[1]);
  assign and_579_nl = (z_out_2_12_1[3:0]==4'b1011) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (~ (fsm_output[10]));
  assign nor_966_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b101) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1844_nl = MUX_s_1_2_2(and_579_nl, nor_966_nl, fsm_output[1]);
  assign mux_1848_nl = MUX_s_1_2_2(mux_1847_nl, mux_1844_nl, fsm_output[0]);
  assign mux_1850_nl = MUX_s_1_2_2(mux_1849_nl, mux_1848_nl, fsm_output[6]);
  assign mux_1860_nl = MUX_s_1_2_2(mux_1859_nl, mux_1850_nl, fsm_output[8]);
  assign vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1875_nl,
      mux_1860_nl, fsm_output[4]);
  assign or_1944_nl = (COMP_LOOP_acc_13_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ (fsm_output[9])) | (~ (fsm_output[5])) | (fsm_output[10]);
  assign or_1943_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | not_tmp_357;
  assign mux_1902_nl = MUX_s_1_2_2(or_1944_nl, or_1943_nl, fsm_output[7]);
  assign or_1941_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b11) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1903_nl = MUX_s_1_2_2(mux_1902_nl, or_1941_nl, fsm_output[2]);
  assign nor_923_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1903_nl);
  assign nor_924_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2])) |
      (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | not_tmp_357);
  assign mux_1904_nl = MUX_s_1_2_2(nor_923_nl, nor_924_nl, fsm_output[8]);
  assign nor_925_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_926_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100)
      | (fsm_output[10]));
  assign nor_927_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) |
      (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100) | (fsm_output[10]));
  assign nor_928_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1899_nl = MUX_s_1_2_2(nor_927_nl, nor_928_nl, fsm_output[4]);
  assign mux_1900_nl = MUX_s_1_2_2(nor_926_nl, mux_1899_nl, fsm_output[6]);
  assign mux_1901_nl = MUX_s_1_2_2(nor_925_nl, mux_1900_nl, fsm_output[8]);
  assign mux_1905_nl = MUX_s_1_2_2(mux_1904_nl, mux_1901_nl, fsm_output[0]);
  assign nand_261_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b00)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_1931_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1896_nl = MUX_s_1_2_2(mux_tmp_1884, or_1931_nl, fsm_output[4]);
  assign mux_1897_nl = MUX_s_1_2_2(nand_261_nl, mux_1896_nl, fsm_output[6]);
  assign and_574_nl = (fsm_output[8]) & (~ mux_1897_nl);
  assign or_1928_nl = (COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5]) | (~ (fsm_output[10]));
  assign or_1926_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | not_tmp_357;
  assign mux_1893_nl = MUX_s_1_2_2(or_1926_nl, or_tmp_1858, fsm_output[2]);
  assign mux_1894_nl = MUX_s_1_2_2(or_1928_nl, mux_1893_nl, fsm_output[4]);
  assign nor_929_nl = ~((fsm_output[6]) | mux_1894_nl);
  assign nor_930_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1895_nl = MUX_s_1_2_2(nor_929_nl, nor_930_nl, fsm_output[8]);
  assign mux_1898_nl = MUX_s_1_2_2(and_574_nl, mux_1895_nl, fsm_output[0]);
  assign mux_1906_nl = MUX_s_1_2_2(mux_1905_nl, mux_1898_nl, fsm_output[3]);
  assign or_1922_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[0]) | nand_337_cse;
  assign or_1920_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00) | not_tmp_357;
  assign mux_1889_nl = MUX_s_1_2_2(or_1922_nl, or_1920_nl, fsm_output[4]);
  assign nor_931_nl = ~((fsm_output[6]) | mux_1889_nl);
  assign or_1916_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | not_tmp_357;
  assign mux_1887_nl = MUX_s_1_2_2(or_591_cse, or_1916_nl, fsm_output[7]);
  assign mux_1888_nl = MUX_s_1_2_2(mux_1887_nl, or_tmp_1858, or_1912_cse);
  assign nor_932_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1888_nl);
  assign mux_1890_nl = MUX_s_1_2_2(nor_931_nl, nor_932_nl, fsm_output[8]);
  assign or_1909_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_1907_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1885_nl = MUX_s_1_2_2(or_1909_nl, or_1907_nl, fsm_output[2]);
  assign mux_1886_nl = MUX_s_1_2_2(mux_1885_nl, mux_tmp_1884, fsm_output[4]);
  assign nor_933_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1886_nl);
  assign mux_1891_nl = MUX_s_1_2_2(mux_1890_nl, nor_933_nl, fsm_output[0]);
  assign or_1902_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_1900_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100) | (fsm_output[10]);
  assign mux_1881_nl = MUX_s_1_2_2(or_1902_nl, or_1900_nl, fsm_output[4]);
  assign or_1899_nl = (COMP_LOOP_acc_14_psp_sva[2:0]!=3'b110) | (~ (fsm_output[2]))
      | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[9])) | (~
      (fsm_output[5])) | (fsm_output[10]);
  assign or_1898_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100) | (fsm_output[10]);
  assign mux_1880_nl = MUX_s_1_2_2(or_1899_nl, or_1898_nl, fsm_output[4]);
  assign mux_1882_nl = MUX_s_1_2_2(mux_1881_nl, mux_1880_nl, fsm_output[6]);
  assign nor_934_nl = ~((fsm_output[8]) | mux_1882_nl);
  assign nor_935_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_936_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[2])) | (~ (fsm_output[7]))
      | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (fsm_output[9]) | not_tmp_248);
  assign or_1893_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b00)
      | not_tmp_357;
  assign or_1891_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1100) | (fsm_output[10]);
  assign mux_1877_nl = MUX_s_1_2_2(or_1893_nl, or_1891_nl, fsm_output[2]);
  assign nor_937_nl = ~((fsm_output[4]) | mux_1877_nl);
  assign mux_1878_nl = MUX_s_1_2_2(nor_936_nl, nor_937_nl, fsm_output[6]);
  assign mux_1879_nl = MUX_s_1_2_2(nor_935_nl, mux_1878_nl, fsm_output[8]);
  assign mux_1883_nl = MUX_s_1_2_2(nor_934_nl, mux_1879_nl, fsm_output[0]);
  assign mux_1892_nl = MUX_s_1_2_2(mux_1891_nl, mux_1883_nl, fsm_output[3]);
  assign vec_rsc_0_12_i_wea_d_pff = MUX_s_1_2_2(mux_1906_nl, mux_1892_nl, fsm_output[1]);
  assign or_2000_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1100) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_1999_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1100) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_1937_nl = MUX_s_1_2_2(or_2000_nl, or_1999_nl, fsm_output[5]);
  assign nor_892_nl = ~((fsm_output[1]) | mux_1937_nl);
  assign nor_893_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1100)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_894_nl = ~((z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_895_nl = ~((z_out_2_12_1[3:0]!=4'b1100) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1935_nl = MUX_s_1_2_2(nor_894_nl, nor_895_nl, fsm_output[5]);
  assign mux_1936_nl = MUX_s_1_2_2(nor_893_nl, mux_1935_nl, fsm_output[1]);
  assign mux_1938_nl = MUX_s_1_2_2(nor_892_nl, mux_1936_nl, fsm_output[0]);
  assign and_571_nl = (fsm_output[6]) & mux_1938_nl;
  assign nor_896_nl = ~((z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_898_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1930_nl = MUX_s_1_2_2(nor_1445_cse, nor_898_nl, fsm_output[5]);
  assign nor_899_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign or_1986_nl = (COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1100) | (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1931_nl = MUX_s_1_2_2(mux_1930_nl, nor_899_nl, or_1986_nl);
  assign mux_1932_nl = MUX_s_1_2_2(nor_896_nl, mux_1931_nl, fsm_output[1]);
  assign nor_900_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_901_nl = ~((z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_902_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1928_nl = MUX_s_1_2_2(nor_901_nl, nor_902_nl, fsm_output[5]);
  assign mux_1929_nl = MUX_s_1_2_2(nor_900_nl, mux_1928_nl, fsm_output[1]);
  assign mux_1933_nl = MUX_s_1_2_2(mux_1932_nl, mux_1929_nl, fsm_output[0]);
  assign nor_903_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_904_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1100) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1926_nl = MUX_s_1_2_2(nor_903_nl, nor_904_nl, fsm_output[1]);
  assign nor_905_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b00) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1925_cse);
  assign mux_1927_nl = MUX_s_1_2_2(mux_1926_nl, nor_905_nl, fsm_output[0]);
  assign mux_1934_nl = MUX_s_1_2_2(mux_1933_nl, mux_1927_nl, fsm_output[6]);
  assign mux_1939_nl = MUX_s_1_2_2(and_571_nl, mux_1934_nl, fsm_output[8]);
  assign nor_906_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1100) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_907_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1100) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1920_nl = MUX_s_1_2_2(nor_906_nl, nor_907_nl, fsm_output[5]);
  assign and_572_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1920_nl;
  assign nor_908_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_909_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1100) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1919_nl = MUX_s_1_2_2(nor_908_nl, nor_909_nl, fsm_output[5]);
  assign and_573_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1919_nl;
  assign mux_1921_nl = MUX_s_1_2_2(and_572_nl, and_573_nl, fsm_output[1]);
  assign nor_910_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (VEC_LOOP_j_sva_11_0[1]) |
      (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_911_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_1917_cse);
  assign mux_1918_nl = MUX_s_1_2_2(nor_910_nl, nor_911_nl, fsm_output[1]);
  assign mux_1922_nl = MUX_s_1_2_2(mux_1921_nl, mux_1918_nl, fsm_output[0]);
  assign nor_912_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7]) |
      (z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_913_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3])) |
      (z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[9])) | (~ (fsm_output[2])) |
      (fsm_output[10]));
  assign nor_914_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_11_psp_sva[2:0]!=3'b110) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1915_nl = MUX_s_1_2_2(nor_913_nl, nor_914_nl, fsm_output[1]);
  assign mux_1916_nl = MUX_s_1_2_2(nor_912_nl, mux_1915_nl, fsm_output[0]);
  assign mux_1923_nl = MUX_s_1_2_2(mux_1922_nl, mux_1916_nl, fsm_output[6]);
  assign nor_915_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1100) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_916_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1100)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1913_nl = MUX_s_1_2_2(nor_915_nl, nor_916_nl, fsm_output[0]);
  assign nor_917_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1100)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nor_918_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1100)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_919_nl = ~((~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1909_nl = MUX_s_1_2_2(nor_918_nl, nor_919_nl, fsm_output[5]);
  assign mux_1910_nl = MUX_s_1_2_2(nor_917_nl, mux_1909_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_920_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1100)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1911_nl = MUX_s_1_2_2(mux_1910_nl, nor_920_nl, fsm_output[1]);
  assign nor_921_nl = ~((z_out_2_12_1[3:0]!=4'b1100) | (~ (fsm_output[5])) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_922_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1908_nl = MUX_s_1_2_2(nor_921_nl, nor_922_nl, fsm_output[1]);
  assign mux_1912_nl = MUX_s_1_2_2(mux_1911_nl, mux_1908_nl, fsm_output[0]);
  assign mux_1914_nl = MUX_s_1_2_2(mux_1913_nl, mux_1912_nl, fsm_output[6]);
  assign mux_1924_nl = MUX_s_1_2_2(mux_1923_nl, mux_1914_nl, fsm_output[8]);
  assign vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_1939_nl,
      mux_1924_nl, fsm_output[4]);
  assign nand_250_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_11_0[1:0]==2'b01)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_2054_nl = (~((fsm_output[9]) & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]==2'b01)))
      | not_tmp_357;
  assign mux_1966_nl = MUX_s_1_2_2(nand_250_nl, or_2054_nl, fsm_output[7]);
  assign or_2052_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b11) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1967_nl = MUX_s_1_2_2(mux_1966_nl, or_2052_nl, fsm_output[2]);
  assign nor_877_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_1967_nl);
  assign nor_878_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2])) |
      (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01)
      | not_tmp_357);
  assign mux_1968_nl = MUX_s_1_2_2(nor_877_nl, nor_878_nl, fsm_output[8]);
  assign nor_879_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1101) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_880_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101)
      | (fsm_output[10]));
  assign nor_881_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) |
      (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101) | (fsm_output[10]));
  assign nor_882_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1101) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_1963_nl = MUX_s_1_2_2(nor_881_nl, nor_882_nl, fsm_output[4]);
  assign mux_1964_nl = MUX_s_1_2_2(nor_880_nl, mux_1963_nl, fsm_output[6]);
  assign mux_1965_nl = MUX_s_1_2_2(nor_879_nl, mux_1964_nl, fsm_output[8]);
  assign mux_1969_nl = MUX_s_1_2_2(mux_1968_nl, mux_1965_nl, fsm_output[0]);
  assign nand_252_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b01)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_2042_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_1960_nl = MUX_s_1_2_2(mux_tmp_1948, or_2042_nl, fsm_output[4]);
  assign mux_1961_nl = MUX_s_1_2_2(nand_252_nl, mux_1960_nl, fsm_output[6]);
  assign and_570_nl = (fsm_output[8]) & (~ mux_1961_nl);
  assign nand_397_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1101) & (fsm_output[2])
      & (fsm_output[7]) & (fsm_output[9]) & (~ (fsm_output[5])) & (fsm_output[10]));
  assign or_2037_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | not_tmp_357;
  assign mux_1957_nl = MUX_s_1_2_2(or_2037_nl, or_tmp_1969, fsm_output[2]);
  assign mux_1958_nl = MUX_s_1_2_2(nand_397_nl, mux_1957_nl, fsm_output[4]);
  assign nor_883_nl = ~((fsm_output[6]) | mux_1958_nl);
  assign nor_884_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_1959_nl = MUX_s_1_2_2(nor_883_nl, nor_884_nl, fsm_output[8]);
  assign mux_1962_nl = MUX_s_1_2_2(and_570_nl, mux_1959_nl, fsm_output[0]);
  assign mux_1970_nl = MUX_s_1_2_2(mux_1969_nl, mux_1962_nl, fsm_output[3]);
  assign or_2033_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (~ (fsm_output[2]))
      | (fsm_output[7]) | nand_334_cse;
  assign or_2031_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01) | not_tmp_357;
  assign mux_1953_nl = MUX_s_1_2_2(or_2033_nl, or_2031_nl, fsm_output[4]);
  assign nor_885_nl = ~((fsm_output[6]) | mux_1953_nl);
  assign or_2027_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01)
      | not_tmp_357;
  assign mux_1951_nl = MUX_s_1_2_2(or_702_cse, or_2027_nl, fsm_output[7]);
  assign mux_1952_nl = MUX_s_1_2_2(mux_1951_nl, or_tmp_1969, or_1912_cse);
  assign nor_886_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_1952_nl);
  assign mux_1954_nl = MUX_s_1_2_2(nor_885_nl, nor_886_nl, fsm_output[8]);
  assign or_2020_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1101) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_2018_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1101)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_1949_nl = MUX_s_1_2_2(or_2020_nl, or_2018_nl, fsm_output[2]);
  assign mux_1950_nl = MUX_s_1_2_2(mux_1949_nl, mux_tmp_1948, fsm_output[4]);
  assign nor_887_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_1950_nl);
  assign mux_1955_nl = MUX_s_1_2_2(mux_1954_nl, nor_887_nl, fsm_output[0]);
  assign or_2013_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b110) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_2011_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101) | (fsm_output[10]);
  assign mux_1945_nl = MUX_s_1_2_2(or_2013_nl, or_2011_nl, fsm_output[4]);
  assign nand_255_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b110) & (fsm_output[2])
      & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[9]) & (fsm_output[5])
      & (~ (fsm_output[10])));
  assign or_2009_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101) | (fsm_output[10]);
  assign mux_1944_nl = MUX_s_1_2_2(nand_255_nl, or_2009_nl, fsm_output[4]);
  assign mux_1946_nl = MUX_s_1_2_2(mux_1945_nl, mux_1944_nl, fsm_output[6]);
  assign nor_888_nl = ~((fsm_output[8]) | mux_1946_nl);
  assign nor_889_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_890_nl = ~((~((fsm_output[4]) & (fsm_output[2]) & (fsm_output[7]) &
      (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1101) & (~ (fsm_output[9])))) | not_tmp_248);
  assign or_2004_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[1:0]!=2'b01)
      | not_tmp_357;
  assign or_2002_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1101) | (fsm_output[10]);
  assign mux_1941_nl = MUX_s_1_2_2(or_2004_nl, or_2002_nl, fsm_output[2]);
  assign nor_891_nl = ~((fsm_output[4]) | mux_1941_nl);
  assign mux_1942_nl = MUX_s_1_2_2(nor_890_nl, nor_891_nl, fsm_output[6]);
  assign mux_1943_nl = MUX_s_1_2_2(nor_889_nl, mux_1942_nl, fsm_output[8]);
  assign mux_1947_nl = MUX_s_1_2_2(nor_888_nl, mux_1943_nl, fsm_output[0]);
  assign mux_1956_nl = MUX_s_1_2_2(mux_1955_nl, mux_1947_nl, fsm_output[3]);
  assign vec_rsc_0_13_i_wea_d_pff = MUX_s_1_2_2(mux_1970_nl, mux_1956_nl, fsm_output[1]);
  assign or_2111_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1101) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_2110_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1101) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_2001_nl = MUX_s_1_2_2(or_2111_nl, or_2110_nl, fsm_output[5]);
  assign nor_848_nl = ~((fsm_output[1]) | mux_2001_nl);
  assign nor_849_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1101)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_850_nl = ~((z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_851_nl = ~((z_out_2_12_1[3:0]!=4'b1101) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1999_nl = MUX_s_1_2_2(nor_850_nl, nor_851_nl, fsm_output[5]);
  assign mux_2000_nl = MUX_s_1_2_2(nor_849_nl, mux_1999_nl, fsm_output[1]);
  assign mux_2002_nl = MUX_s_1_2_2(nor_848_nl, mux_2000_nl, fsm_output[0]);
  assign and_565_nl = (fsm_output[6]) & mux_2002_nl;
  assign nor_852_nl = ~((z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_854_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_1994_nl = MUX_s_1_2_2(nor_1445_cse, nor_854_nl, fsm_output[5]);
  assign nor_855_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1101)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nand_243_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1101) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_1995_nl = MUX_s_1_2_2(mux_1994_nl, nor_855_nl, nand_243_nl);
  assign mux_1996_nl = MUX_s_1_2_2(nor_852_nl, mux_1995_nl, fsm_output[1]);
  assign nor_856_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_857_nl = ~((z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_858_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_1992_nl = MUX_s_1_2_2(nor_857_nl, nor_858_nl, fsm_output[5]);
  assign mux_1993_nl = MUX_s_1_2_2(nor_856_nl, mux_1992_nl, fsm_output[1]);
  assign mux_1997_nl = MUX_s_1_2_2(mux_1996_nl, mux_1993_nl, fsm_output[0]);
  assign nor_859_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1101) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_860_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1101) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1990_nl = MUX_s_1_2_2(nor_859_nl, nor_860_nl, fsm_output[1]);
  assign nor_861_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b01) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1925_cse);
  assign mux_1991_nl = MUX_s_1_2_2(mux_1990_nl, nor_861_nl, fsm_output[0]);
  assign mux_1998_nl = MUX_s_1_2_2(mux_1997_nl, mux_1991_nl, fsm_output[6]);
  assign mux_2003_nl = MUX_s_1_2_2(and_565_nl, mux_1998_nl, fsm_output[8]);
  assign nor_862_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1101) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_863_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1101) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1984_nl = MUX_s_1_2_2(nor_862_nl, nor_863_nl, fsm_output[5]);
  assign and_566_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_1984_nl;
  assign nor_864_nl = ~((~((fsm_output[7]) & (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1101)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_865_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1101) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1983_nl = MUX_s_1_2_2(nor_864_nl, nor_865_nl, fsm_output[5]);
  assign and_567_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_1983_nl;
  assign mux_1985_nl = MUX_s_1_2_2(and_566_nl, and_567_nl, fsm_output[1]);
  assign nor_866_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (VEC_LOOP_j_sva_11_0[1]) |
      (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_867_nl = ~(nand_332_cse | mux_1917_cse);
  assign mux_1982_nl = MUX_s_1_2_2(nor_866_nl, nor_867_nl, fsm_output[1]);
  assign mux_1986_nl = MUX_s_1_2_2(mux_1985_nl, mux_1982_nl, fsm_output[0]);
  assign nor_868_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7]) |
      (z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_869_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3])) |
      (z_out_2_12_1[3:0]!=4'b1101) | (~ (fsm_output[9])) | (~ (fsm_output[2])) |
      (fsm_output[10]));
  assign and_568_nl = (VEC_LOOP_j_sva_11_0[0]) & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm
      & (fsm_output[5]) & (COMP_LOOP_acc_11_psp_sva[2:0]==3'b110) & (fsm_output[7])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign mux_1979_nl = MUX_s_1_2_2(nor_869_nl, and_568_nl, fsm_output[1]);
  assign mux_1980_nl = MUX_s_1_2_2(nor_868_nl, mux_1979_nl, fsm_output[0]);
  assign mux_1987_nl = MUX_s_1_2_2(mux_1986_nl, mux_1980_nl, fsm_output[6]);
  assign nor_870_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1101) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_871_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1101)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_1977_nl = MUX_s_1_2_2(nor_870_nl, nor_871_nl, fsm_output[0]);
  assign nor_872_nl = ~((~((fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1101)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_873_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1101)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_874_nl = ~((~((fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1101) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign mux_1973_nl = MUX_s_1_2_2(nor_873_nl, nor_874_nl, fsm_output[5]);
  assign mux_1974_nl = MUX_s_1_2_2(nor_872_nl, mux_1973_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_875_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1101)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_1975_nl = MUX_s_1_2_2(mux_1974_nl, nor_875_nl, fsm_output[1]);
  assign and_569_nl = (z_out_2_12_1[3:0]==4'b1101) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (~ (fsm_output[10]));
  assign nor_876_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b110) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_1972_nl = MUX_s_1_2_2(and_569_nl, nor_876_nl, fsm_output[1]);
  assign mux_1976_nl = MUX_s_1_2_2(mux_1975_nl, mux_1972_nl, fsm_output[0]);
  assign mux_1978_nl = MUX_s_1_2_2(mux_1977_nl, mux_1976_nl, fsm_output[6]);
  assign mux_1988_nl = MUX_s_1_2_2(mux_1987_nl, mux_1978_nl, fsm_output[8]);
  assign vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2003_nl,
      mux_1988_nl, fsm_output[4]);
  assign nand_235_nl = ~((COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_11_0[1:0]==2'b10)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_2164_nl = (~ (fsm_output[9])) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | not_tmp_377;
  assign mux_2030_nl = MUX_s_1_2_2(nand_235_nl, or_2164_nl, fsm_output[7]);
  assign or_2162_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b11) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_2031_nl = MUX_s_1_2_2(mux_2030_nl, or_2162_nl, fsm_output[2]);
  assign nor_833_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_2031_nl);
  assign nor_834_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2])) |
      (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | not_tmp_377);
  assign mux_2032_nl = MUX_s_1_2_2(nor_833_nl, nor_834_nl, fsm_output[8]);
  assign nor_835_nl = ~((COMP_LOOP_acc_1_cse_12_sva[3:0]!=4'b1110) | (~ (fsm_output[6]))
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | not_tmp_248);
  assign nor_836_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110)
      | (fsm_output[10]));
  assign nor_837_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) |
      (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110) | (fsm_output[10]));
  assign nor_838_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1110) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_2027_nl = MUX_s_1_2_2(nor_837_nl, nor_838_nl, fsm_output[4]);
  assign mux_2028_nl = MUX_s_1_2_2(nor_836_nl, mux_2027_nl, fsm_output[6]);
  assign mux_2029_nl = MUX_s_1_2_2(nor_835_nl, mux_2028_nl, fsm_output[8]);
  assign mux_2033_nl = MUX_s_1_2_2(mux_2032_nl, mux_2029_nl, fsm_output[0]);
  assign nand_236_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b10)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_2152_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_2024_nl = MUX_s_1_2_2(mux_tmp_2012, or_2152_nl, fsm_output[4]);
  assign mux_2025_nl = MUX_s_1_2_2(nand_236_nl, mux_2024_nl, fsm_output[6]);
  assign and_563_nl = (fsm_output[8]) & (~ mux_2025_nl);
  assign nand_396_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1110) & (fsm_output[2])
      & (fsm_output[7]) & (fsm_output[9]) & (~ (fsm_output[5])) & (fsm_output[10]));
  assign or_2147_nl = (fsm_output[7]) | (~ (fsm_output[9])) | (~ (fsm_output[5]))
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) | not_tmp_377;
  assign mux_2021_nl = MUX_s_1_2_2(or_2147_nl, or_tmp_2082, fsm_output[2]);
  assign mux_2022_nl = MUX_s_1_2_2(nand_396_nl, mux_2021_nl, fsm_output[4]);
  assign nor_839_nl = ~((fsm_output[6]) | mux_2022_nl);
  assign nor_840_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2023_nl = MUX_s_1_2_2(nor_839_nl, nor_840_nl, fsm_output[8]);
  assign mux_2026_nl = MUX_s_1_2_2(and_563_nl, mux_2023_nl, fsm_output[0]);
  assign mux_2034_nl = MUX_s_1_2_2(mux_2033_nl, mux_2026_nl, fsm_output[3]);
  assign or_2143_nl = (COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[0]) | nand_337_cse;
  assign or_2141_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | (~
      (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) | not_tmp_377;
  assign mux_2017_nl = MUX_s_1_2_2(or_2143_nl, or_2141_nl, fsm_output[4]);
  assign nor_841_nl = ~((fsm_output[6]) | mux_2017_nl);
  assign or_2135_nl = (fsm_output[9]) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | not_tmp_377;
  assign mux_2015_nl = MUX_s_1_2_2(or_591_cse, or_2135_nl, fsm_output[7]);
  assign mux_2016_nl = MUX_s_1_2_2(or_tmp_2082, mux_2015_nl, and_564_cse);
  assign nor_842_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_2016_nl);
  assign mux_2018_nl = MUX_s_1_2_2(nor_841_nl, nor_842_nl, fsm_output[8]);
  assign or_2131_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1110) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign or_2129_nl = (~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1110)
      | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_2013_nl = MUX_s_1_2_2(or_2131_nl, or_2129_nl, fsm_output[2]);
  assign mux_2014_nl = MUX_s_1_2_2(mux_2013_nl, mux_tmp_2012, fsm_output[4]);
  assign nor_843_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_2014_nl);
  assign mux_2019_nl = MUX_s_1_2_2(mux_2018_nl, nor_843_nl, fsm_output[0]);
  assign or_2124_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[0]) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_2122_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110) | (fsm_output[10]);
  assign mux_2009_nl = MUX_s_1_2_2(or_2124_nl, or_2122_nl, fsm_output[4]);
  assign nand_239_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[2])
      & (fsm_output[7]) & (~ (VEC_LOOP_j_sva_11_0[0])) & (fsm_output[9]) & (fsm_output[5])
      & (~ (fsm_output[10])));
  assign or_2120_nl = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110) | (fsm_output[10]);
  assign mux_2008_nl = MUX_s_1_2_2(nand_239_nl, or_2120_nl, fsm_output[4]);
  assign mux_2010_nl = MUX_s_1_2_2(mux_2009_nl, mux_2008_nl, fsm_output[6]);
  assign nor_844_nl = ~((fsm_output[8]) | mux_2010_nl);
  assign nor_845_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_846_nl = ~((~((fsm_output[4]) & (fsm_output[2]) & (fsm_output[7]) &
      (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1110) & (~ (fsm_output[9])))) | not_tmp_248);
  assign or_2115_nl = (fsm_output[7]) | (fsm_output[9]) | (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[0])
      | not_tmp_377;
  assign or_2113_nl = (~ (fsm_output[7])) | (~ (fsm_output[9])) | (fsm_output[5])
      | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1110) | (fsm_output[10]);
  assign mux_2005_nl = MUX_s_1_2_2(or_2115_nl, or_2113_nl, fsm_output[2]);
  assign nor_847_nl = ~((fsm_output[4]) | mux_2005_nl);
  assign mux_2006_nl = MUX_s_1_2_2(nor_846_nl, nor_847_nl, fsm_output[6]);
  assign mux_2007_nl = MUX_s_1_2_2(nor_845_nl, mux_2006_nl, fsm_output[8]);
  assign mux_2011_nl = MUX_s_1_2_2(nor_844_nl, mux_2007_nl, fsm_output[0]);
  assign mux_2020_nl = MUX_s_1_2_2(mux_2019_nl, mux_2011_nl, fsm_output[3]);
  assign vec_rsc_0_14_i_wea_d_pff = MUX_s_1_2_2(mux_2034_nl, mux_2020_nl, fsm_output[1]);
  assign or_2221_nl = (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1110) | (fsm_output[3])
      | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]);
  assign or_2220_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1110) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_2065_nl = MUX_s_1_2_2(or_2221_nl, or_2220_nl, fsm_output[5]);
  assign nor_804_nl = ~((fsm_output[1]) | mux_2065_nl);
  assign nor_805_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1110)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_806_nl = ~((z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[7])) | (fsm_output[3])
      | (fsm_output[9]) | not_tmp_253);
  assign nor_807_nl = ~((z_out_2_12_1[3:0]!=4'b1110) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_2063_nl = MUX_s_1_2_2(nor_806_nl, nor_807_nl, fsm_output[5]);
  assign mux_2064_nl = MUX_s_1_2_2(nor_805_nl, mux_2063_nl, fsm_output[1]);
  assign mux_2066_nl = MUX_s_1_2_2(nor_804_nl, mux_2064_nl, fsm_output[0]);
  assign and_558_nl = (fsm_output[6]) & mux_2066_nl;
  assign nor_808_nl = ~((z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_810_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign mux_2058_nl = MUX_s_1_2_2(nor_1445_cse, nor_810_nl, fsm_output[5]);
  assign nor_811_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1110)
      | (~ (fsm_output[3])) | (fsm_output[9]) | not_tmp_253);
  assign nand_228_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1110) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_2059_nl = MUX_s_1_2_2(mux_2058_nl, nor_811_nl, nand_228_nl);
  assign mux_2060_nl = MUX_s_1_2_2(nor_808_nl, mux_2059_nl, fsm_output[1]);
  assign nor_812_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign nor_813_nl = ~((z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign nor_814_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_2056_nl = MUX_s_1_2_2(nor_813_nl, nor_814_nl, fsm_output[5]);
  assign mux_2057_nl = MUX_s_1_2_2(nor_812_nl, mux_2056_nl, fsm_output[1]);
  assign mux_2061_nl = MUX_s_1_2_2(mux_2060_nl, mux_2057_nl, fsm_output[0]);
  assign nor_815_nl = ~((~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_14_sva[3:0]!=4'b1110) | (~ (fsm_output[3]))
      | (fsm_output[9]) | not_tmp_253);
  assign nor_816_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1110) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_2054_nl = MUX_s_1_2_2(nor_815_nl, nor_816_nl, fsm_output[1]);
  assign nor_817_nl = ~((fsm_output[1]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b10) | (~
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | mux_1925_cse);
  assign mux_2055_nl = MUX_s_1_2_2(mux_2054_nl, nor_817_nl, fsm_output[0]);
  assign mux_2062_nl = MUX_s_1_2_2(mux_2061_nl, mux_2055_nl, fsm_output[6]);
  assign mux_2067_nl = MUX_s_1_2_2(and_558_nl, mux_2062_nl, fsm_output[8]);
  assign nor_818_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1110) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_819_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1110) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_2048_nl = MUX_s_1_2_2(nor_818_nl, nor_819_nl, fsm_output[5]);
  assign and_559_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_2048_nl;
  assign nor_820_nl = ~((~((fsm_output[7]) & (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1110)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_821_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]!=4'b1110) | (fsm_output[7])
      | (~ (fsm_output[3])) | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_2047_nl = MUX_s_1_2_2(nor_820_nl, nor_821_nl, fsm_output[5]);
  assign and_560_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_2047_nl;
  assign mux_2049_nl = MUX_s_1_2_2(and_559_nl, and_560_nl, fsm_output[1]);
  assign nor_822_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (VEC_LOOP_j_sva_11_0[0]) | (~ (fsm_output[5])) | (~ (VEC_LOOP_j_sva_11_0[2]))
      | (fsm_output[7]) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_823_nl = ~((VEC_LOOP_j_sva_11_0[0]) | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm)
      | mux_2045_cse);
  assign mux_2046_nl = MUX_s_1_2_2(nor_822_nl, nor_823_nl, fsm_output[1]);
  assign mux_2050_nl = MUX_s_1_2_2(mux_2049_nl, mux_2046_nl, fsm_output[0]);
  assign nor_824_nl = ~((~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[7]) |
      (z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_825_nl = ~((fsm_output[5]) | (fsm_output[7]) | (~ (fsm_output[3])) |
      (z_out_2_12_1[3:0]!=4'b1110) | (~ (fsm_output[9])) | (~ (fsm_output[2])) |
      (fsm_output[10]));
  assign and_561_nl = (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111) & (~ (VEC_LOOP_j_sva_11_0[0]))
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign mux_2043_nl = MUX_s_1_2_2(nor_825_nl, and_561_nl, fsm_output[1]);
  assign mux_2044_nl = MUX_s_1_2_2(nor_824_nl, mux_2043_nl, fsm_output[0]);
  assign mux_2051_nl = MUX_s_1_2_2(mux_2050_nl, mux_2044_nl, fsm_output[6]);
  assign nor_826_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1110) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_827_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1110)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_2041_nl = MUX_s_1_2_2(nor_826_nl, nor_827_nl, fsm_output[0]);
  assign nor_828_nl = ~((~((fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1110)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_829_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1110)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_830_nl = ~((~((fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1110) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign mux_2037_nl = MUX_s_1_2_2(nor_829_nl, nor_830_nl, fsm_output[5]);
  assign mux_2038_nl = MUX_s_1_2_2(nor_828_nl, mux_2037_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign nor_831_nl = ~((~ (fsm_output[5])) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1110)
      | (fsm_output[3]) | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_2039_nl = MUX_s_1_2_2(mux_2038_nl, nor_831_nl, fsm_output[1]);
  assign and_562_nl = (z_out_2_12_1[3:0]==4'b1110) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (~ (fsm_output[10]));
  assign nor_832_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111) | (VEC_LOOP_j_sva_11_0[0])
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_2036_nl = MUX_s_1_2_2(and_562_nl, nor_832_nl, fsm_output[1]);
  assign mux_2040_nl = MUX_s_1_2_2(mux_2039_nl, mux_2036_nl, fsm_output[0]);
  assign mux_2042_nl = MUX_s_1_2_2(mux_2041_nl, mux_2040_nl, fsm_output[6]);
  assign mux_2052_nl = MUX_s_1_2_2(mux_2051_nl, mux_2042_nl, fsm_output[8]);
  assign vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2067_nl,
      mux_2052_nl, fsm_output[4]);
  assign and_554_nl = (COMP_LOOP_acc_13_psp_sva[1:0]==2'b11) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10]));
  assign mux_2094_nl = MUX_s_1_2_2(and_554_nl, nor_tmp_265, fsm_output[7]);
  assign or_2271_nl = (VEC_LOOP_j_sva_11_0[3:2]!=2'b11) | (~ (fsm_output[7])) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (fsm_output[9]) | (fsm_output[5]) | (fsm_output[10]);
  assign mux_2095_nl = MUX_s_1_2_2((~ mux_2094_nl), or_2271_nl, fsm_output[2]);
  assign nor_789_nl = ~((fsm_output[6]) | (fsm_output[4]) | mux_2095_nl);
  assign nor_790_nl = ~((fsm_output[6]) | (fsm_output[4]) | (~ (fsm_output[2])) |
      (fsm_output[7]) | (fsm_output[9]) | (fsm_output[5]) | not_tmp_390);
  assign mux_2096_nl = MUX_s_1_2_2(nor_789_nl, nor_790_nl, fsm_output[8]);
  assign nor_791_nl = ~((~((COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111) & (fsm_output[6])
      & (fsm_output[4]) & (~ (fsm_output[2])) & (fsm_output[7]) & (~ (fsm_output[9]))))
      | not_tmp_248);
  assign nor_792_nl = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]) | (~
      (fsm_output[9])) | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1111)
      | (fsm_output[10]));
  assign nor_793_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) |
      (~ (fsm_output[5])) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1111) | (fsm_output[10]));
  assign nor_794_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]!=4'b1111) | (~ (fsm_output[2]))
      | (fsm_output[7]) | (~ (fsm_output[9])) | (fsm_output[5]) | (fsm_output[10]));
  assign mux_2091_nl = MUX_s_1_2_2(nor_793_nl, nor_794_nl, fsm_output[4]);
  assign mux_2092_nl = MUX_s_1_2_2(nor_792_nl, mux_2091_nl, fsm_output[6]);
  assign mux_2093_nl = MUX_s_1_2_2(nor_791_nl, mux_2092_nl, fsm_output[8]);
  assign mux_2097_nl = MUX_s_1_2_2(mux_2096_nl, mux_2093_nl, fsm_output[0]);
  assign nand_215_nl = ~((COMP_LOOP_acc_16_psp_sva[0]) & (fsm_output[4]) & (fsm_output[2])
      & (VEC_LOOP_j_sva_11_0[2]) & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[1:0]==2'b11)
      & (fsm_output[9]) & (fsm_output[5]) & (~ (fsm_output[10])));
  assign or_2261_nl = (COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (fsm_output[2]) |
      (fsm_output[7]) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign mux_2088_nl = MUX_s_1_2_2(mux_tmp_2076, or_2261_nl, fsm_output[4]);
  assign mux_2089_nl = MUX_s_1_2_2(nand_215_nl, mux_2088_nl, fsm_output[6]);
  assign and_555_nl = (fsm_output[8]) & (~ mux_2089_nl);
  assign nand_395_nl = ~((COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & (fsm_output[2])
      & (fsm_output[7]) & (fsm_output[9]) & (~ (fsm_output[5])) & (fsm_output[10]));
  assign or_2256_nl = (fsm_output[7]) | (~ nor_tmp_265);
  assign mux_2085_nl = MUX_s_1_2_2(or_2256_nl, or_tmp_2192, fsm_output[2]);
  assign mux_2086_nl = MUX_s_1_2_2(nand_395_nl, mux_2085_nl, fsm_output[4]);
  assign nor_795_nl = ~((fsm_output[6]) | mux_2086_nl);
  assign nor_796_nl = ~((COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1111) | (fsm_output[6])
      | (~ (fsm_output[4])) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_2087_nl = MUX_s_1_2_2(nor_795_nl, nor_796_nl, fsm_output[8]);
  assign mux_2090_nl = MUX_s_1_2_2(and_555_nl, mux_2087_nl, fsm_output[0]);
  assign mux_2098_nl = MUX_s_1_2_2(mux_2097_nl, mux_2090_nl, fsm_output[3]);
  assign or_2253_nl = (~((COMP_LOOP_acc_20_psp_sva[2:0]==3'b111) & (fsm_output[2])
      & (~ (fsm_output[7])))) | nand_334_cse;
  assign or_2251_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (fsm_output[9]) | not_tmp_387;
  assign mux_2081_nl = MUX_s_1_2_2(or_2253_nl, or_2251_nl, fsm_output[4]);
  assign nor_797_nl = ~((fsm_output[6]) | mux_2081_nl);
  assign or_2245_nl = (fsm_output[9]) | (fsm_output[5]) | not_tmp_390;
  assign mux_2079_nl = MUX_s_1_2_2(or_702_cse, or_2245_nl, fsm_output[7]);
  assign mux_2080_nl = MUX_s_1_2_2(or_tmp_2192, mux_2079_nl, and_564_cse);
  assign nor_798_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[4])) | (fsm_output[2])
      | mux_2080_nl);
  assign mux_2082_nl = MUX_s_1_2_2(nor_797_nl, nor_798_nl, fsm_output[8]);
  assign or_2241_nl = (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1111) | (fsm_output[7])
      | (fsm_output[9]) | not_tmp_248;
  assign nand_219_nl = ~((fsm_output[7]) & (COMP_LOOP_acc_1_cse_6_sva[3:0]==4'b1111)
      & (fsm_output[9]) & (~ (fsm_output[5])) & (~ (fsm_output[10])));
  assign mux_2077_nl = MUX_s_1_2_2(or_2241_nl, nand_219_nl, fsm_output[2]);
  assign mux_2078_nl = MUX_s_1_2_2(mux_2077_nl, mux_tmp_2076, fsm_output[4]);
  assign nor_799_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_2078_nl);
  assign mux_2083_nl = MUX_s_1_2_2(mux_2082_nl, nor_799_nl, fsm_output[0]);
  assign or_2234_nl = (COMP_LOOP_acc_17_psp_sva[2:0]!=3'b111) | (fsm_output[2]) |
      (~ (fsm_output[7])) | (~ (VEC_LOOP_j_sva_11_0[0])) | (fsm_output[9]) | (fsm_output[5])
      | (~ (fsm_output[10]));
  assign or_2232_nl = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[9]))
      | (fsm_output[5]) | (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]!=4'b1111) | (fsm_output[10]);
  assign mux_2073_nl = MUX_s_1_2_2(or_2234_nl, or_2232_nl, fsm_output[4]);
  assign nand_220_nl = ~((COMP_LOOP_acc_14_psp_sva[2:0]==3'b111) & (fsm_output[2])
      & (fsm_output[7]) & (VEC_LOOP_j_sva_11_0[0]) & (fsm_output[9]) & (fsm_output[5])
      & (~ (fsm_output[10])));
  assign nand_221_nl = ~((fsm_output[2]) & (fsm_output[7]) & (~ (fsm_output[9]))
      & (fsm_output[5]) & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111) & (~ (fsm_output[10])));
  assign mux_2072_nl = MUX_s_1_2_2(nand_220_nl, nand_221_nl, fsm_output[4]);
  assign mux_2074_nl = MUX_s_1_2_2(mux_2073_nl, mux_2072_nl, fsm_output[6]);
  assign nor_800_nl = ~((fsm_output[8]) | mux_2074_nl);
  assign nor_801_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111) | (~ (fsm_output[6]))
      | (fsm_output[4]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[9])
      | (~ (fsm_output[5])) | (fsm_output[10]));
  assign nor_802_nl = ~((~((fsm_output[4]) & (fsm_output[2]) & (fsm_output[7]) &
      (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & (~ (fsm_output[9])))) | not_tmp_248);
  assign or_2225_nl = (fsm_output[7]) | (fsm_output[9]) | not_tmp_387;
  assign nand_223_nl = ~((fsm_output[7]) & (fsm_output[9]) & (~ (fsm_output[5]))
      & (COMP_LOOP_acc_10_cse_12_1_1_sva[3:0]==4'b1111) & (~ (fsm_output[10])));
  assign mux_2069_nl = MUX_s_1_2_2(or_2225_nl, nand_223_nl, fsm_output[2]);
  assign nor_803_nl = ~((fsm_output[4]) | mux_2069_nl);
  assign mux_2070_nl = MUX_s_1_2_2(nor_802_nl, nor_803_nl, fsm_output[6]);
  assign mux_2071_nl = MUX_s_1_2_2(nor_801_nl, mux_2070_nl, fsm_output[8]);
  assign mux_2075_nl = MUX_s_1_2_2(nor_800_nl, mux_2071_nl, fsm_output[0]);
  assign mux_2084_nl = MUX_s_1_2_2(mux_2083_nl, mux_2075_nl, fsm_output[3]);
  assign vec_rsc_0_15_i_wea_d_pff = MUX_s_1_2_2(mux_2098_nl, mux_2084_nl, fsm_output[1]);
  assign nand_199_nl = ~((fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1111) & (~ (fsm_output[3]))
      & (fsm_output[9]) & (fsm_output[2]) & (~ (fsm_output[10])));
  assign or_2327_nl = (fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10]));
  assign mux_2129_nl = MUX_s_1_2_2(nand_199_nl, or_2327_nl, fsm_output[5]);
  assign nor_763_nl = ~((fsm_output[1]) | mux_2129_nl);
  assign nor_764_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (z_out_2_12_1[3:0]!=4'b1111)
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_765_nl = ~((~((z_out_2_12_1[3:0]==4'b1111) & (fsm_output[7]) & (~ (fsm_output[3]))
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_766_nl = ~((z_out_2_12_1[3:0]!=4'b1111) | (fsm_output[7]) | (fsm_output[3])
      | (~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_2127_nl = MUX_s_1_2_2(nor_765_nl, nor_766_nl, fsm_output[5]);
  assign mux_2128_nl = MUX_s_1_2_2(nor_764_nl, mux_2127_nl, fsm_output[1]);
  assign mux_2130_nl = MUX_s_1_2_2(nor_763_nl, mux_2128_nl, fsm_output[0]);
  assign and_546_nl = (fsm_output[6]) & mux_2130_nl;
  assign nor_767_nl = ~((z_out_2_12_1[3:0]!=4'b1111) | (~ (fsm_output[5])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_769_nl = ~((~((~ (fsm_output[7])) & (z_out_2_12_1[3:0]==4'b1111) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign mux_2122_nl = MUX_s_1_2_2(nor_1445_cse, nor_769_nl, fsm_output[5]);
  assign nor_770_nl = ~((~((fsm_output[5]) & (~ (fsm_output[7])) & (z_out_2_12_1[3:0]==4'b1111)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nand_203_nl = ~((COMP_LOOP_acc_1_cse_8_sva[3:0]==4'b1111) & COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm);
  assign mux_2123_nl = MUX_s_1_2_2(mux_2122_nl, nor_770_nl, nand_203_nl);
  assign mux_2124_nl = MUX_s_1_2_2(nor_767_nl, mux_2123_nl, fsm_output[1]);
  assign nor_771_nl = ~((COMP_LOOP_acc_19_psp_sva[1:0]!=2'b11) | (VEC_LOOP_j_sva_11_0[1:0]!=2'b11)
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign and_547_nl = (z_out_2_12_1[3:0]==4'b1111) & (fsm_output[7]) & (fsm_output[3])
      & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign nor_772_nl = ~((fsm_output[7]) | (z_out_2_12_1[3:0]!=4'b1111) | (~ (fsm_output[3]))
      | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign mux_2120_nl = MUX_s_1_2_2(and_547_nl, nor_772_nl, fsm_output[5]);
  assign mux_2121_nl = MUX_s_1_2_2(nor_771_nl, mux_2120_nl, fsm_output[1]);
  assign mux_2125_nl = MUX_s_1_2_2(mux_2124_nl, mux_2121_nl, fsm_output[0]);
  assign nor_773_nl = ~((~(COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5])
      & (~ (fsm_output[7])) & (COMP_LOOP_acc_1_cse_14_sva[3:0]==4'b1111) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_774_nl = ~((~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) | (~ (fsm_output[5]))
      | (fsm_output[7]) | (COMP_LOOP_acc_1_cse_4_sva[3:0]!=4'b1111) | (fsm_output[3])
      | (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_2118_nl = MUX_s_1_2_2(nor_773_nl, nor_774_nl, fsm_output[1]);
  assign nor_775_nl = ~(nand_324_cse | mux_1925_cse);
  assign mux_2119_nl = MUX_s_1_2_2(mux_2118_nl, nor_775_nl, fsm_output[0]);
  assign mux_2126_nl = MUX_s_1_2_2(mux_2125_nl, mux_2119_nl, fsm_output[6]);
  assign mux_2131_nl = MUX_s_1_2_2(and_546_nl, mux_2126_nl, fsm_output[8]);
  assign nor_776_nl = ~((COMP_LOOP_acc_1_cse_2_sva[3:0]!=4'b1111) | (~ (fsm_output[7]))
      | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_777_nl = ~((COMP_LOOP_acc_1_cse_6_sva[3:0]!=4'b1111) | (fsm_output[7])
      | (fsm_output[3]) | (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[10]));
  assign mux_2112_nl = MUX_s_1_2_2(nor_776_nl, nor_777_nl, fsm_output[5]);
  assign and_548_nl = COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & mux_2112_nl;
  assign nor_778_nl = ~((~((fsm_output[7]) & (COMP_LOOP_acc_1_cse_12_sva[3:0]==4'b1111)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign and_759_nl = (COMP_LOOP_acc_1_cse_sva[3:0]==4'b1111) & (~ (fsm_output[7]))
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (fsm_output[10]);
  assign mux_2111_nl = MUX_s_1_2_2(nor_778_nl, and_759_nl, fsm_output[5]);
  assign and_549_nl = COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm & mux_2111_nl;
  assign mux_2113_nl = MUX_s_1_2_2(and_548_nl, and_549_nl, fsm_output[1]);
  assign nor_780_nl = ~((~ (VEC_LOOP_j_sva_11_0[3])) | (~ (VEC_LOOP_j_sva_11_0[1]))
      | (~ (VEC_LOOP_j_sva_11_0[0])) | (~ (fsm_output[5])) | (fsm_output[7]) | (~
      (VEC_LOOP_j_sva_11_0[2])) | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_781_nl = ~(nand_332_cse | mux_2045_cse);
  assign mux_2110_nl = MUX_s_1_2_2(nor_780_nl, nor_781_nl, fsm_output[1]);
  assign mux_2114_nl = MUX_s_1_2_2(mux_2113_nl, mux_2110_nl, fsm_output[0]);
  assign nor_782_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1111) | (fsm_output[5])
      | (fsm_output[7]) | (~ (fsm_output[3])) | (fsm_output[9]) | (fsm_output[2])
      | (fsm_output[10]));
  assign and_550_nl = (~ (fsm_output[5])) & (~ (fsm_output[7])) & (fsm_output[3])
      & (z_out_2_12_1[3:0]==4'b1111) & (fsm_output[9]) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign and_551_nl = (COMP_LOOP_acc_11_psp_sva[2:0]==3'b111) & (VEC_LOOP_j_sva_11_0[0])
      & COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign mux_2107_nl = MUX_s_1_2_2(and_550_nl, and_551_nl, fsm_output[1]);
  assign mux_2108_nl = MUX_s_1_2_2(nor_782_nl, mux_2107_nl, fsm_output[0]);
  assign mux_2115_nl = MUX_s_1_2_2(mux_2114_nl, mux_2108_nl, fsm_output[6]);
  assign nor_783_nl = ~((~ (fsm_output[1])) | (z_out_2_12_1[3:0]!=4'b1111) | (fsm_output[5])
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]));
  assign nor_784_nl = ~((fsm_output[1]) | (fsm_output[5]) | (z_out_2_12_1[3:0]!=4'b1111)
      | (~ (fsm_output[7])) | (fsm_output[3]) | (fsm_output[9]) | not_tmp_253);
  assign mux_2105_nl = MUX_s_1_2_2(nor_783_nl, nor_784_nl, fsm_output[0]);
  assign nor_785_nl = ~((~((fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1111)
      & (fsm_output[3]) & (~ (fsm_output[9])))) | not_tmp_253);
  assign nor_786_nl = ~((~ (fsm_output[7])) | (COMP_LOOP_acc_1_cse_10_sva[3:0]!=4'b1111)
      | (fsm_output[3]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[10]));
  assign nor_787_nl = ~((~((fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1111) & (fsm_output[3])
      & (~ (fsm_output[9])))) | not_tmp_253);
  assign mux_2101_nl = MUX_s_1_2_2(nor_786_nl, nor_787_nl, fsm_output[5]);
  assign mux_2102_nl = MUX_s_1_2_2(nor_785_nl, mux_2101_nl, COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm);
  assign and_552_nl = (fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1111)
      & (~ (fsm_output[3])) & (~ (fsm_output[9])) & (fsm_output[2]) & (~ (fsm_output[10]));
  assign mux_2103_nl = MUX_s_1_2_2(mux_2102_nl, and_552_nl, fsm_output[1]);
  assign and_553_nl = (fsm_output[5]) & (fsm_output[7]) & (z_out_2_12_1[3:0]==4'b1111)
      & (fsm_output[3]) & (fsm_output[9]) & (~ (fsm_output[2])) & (~ (fsm_output[10]));
  assign nor_788_nl = ~((COMP_LOOP_acc_20_psp_sva[2:0]!=3'b111) | (~ (VEC_LOOP_j_sva_11_0[0]))
      | (~ COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (fsm_output[9]) | (fsm_output[2]) | (~ (fsm_output[10])));
  assign mux_2100_nl = MUX_s_1_2_2(and_553_nl, nor_788_nl, fsm_output[1]);
  assign mux_2104_nl = MUX_s_1_2_2(mux_2103_nl, mux_2100_nl, fsm_output[0]);
  assign mux_2106_nl = MUX_s_1_2_2(mux_2105_nl, mux_2104_nl, fsm_output[6]);
  assign mux_2116_nl = MUX_s_1_2_2(mux_2115_nl, mux_2106_nl, fsm_output[8]);
  assign vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = MUX_s_1_2_2(mux_2131_nl,
      mux_2116_nl, fsm_output[4]);
  assign and_dcpl_332 = (fsm_output==11'b11010100010);
  assign and_dcpl_333 = (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_dcpl_338 = (~ (fsm_output[3])) & (fsm_output[5]) & (~ (fsm_output[8]));
  assign and_dcpl_340 = ~((fsm_output[2]) | (fsm_output[9]) | (fsm_output[10]));
  assign and_dcpl_342 = and_dcpl_340 & and_dcpl_338 & (fsm_output[4]) & (~ (fsm_output[7]))
      & (~ (fsm_output[1])) & and_dcpl_333;
  assign and_dcpl_344 = ~((fsm_output[4]) | (fsm_output[7]));
  assign and_dcpl_345 = and_dcpl_344 & (fsm_output[1]);
  assign and_dcpl_349 = and_dcpl_340 & (fsm_output[3]) & (~ (fsm_output[5])) & (~
      (fsm_output[8]));
  assign and_dcpl_350 = and_dcpl_349 & and_dcpl_345 & (~ (fsm_output[6])) & (~ (fsm_output[0]));
  assign and_dcpl_356 = (~ (fsm_output[2])) & (fsm_output[9]) & (fsm_output[10])
      & and_dcpl_338 & and_dcpl_345 & (fsm_output[6]) & (fsm_output[0]);
  assign and_dcpl_359 = and_dcpl_349 & and_dcpl_344 & (~ (fsm_output[1])) & and_dcpl_333;
  assign and_815_cse = (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_816_cse = (fsm_output[4]) & (~ (fsm_output[7]));
  assign and_820_cse = and_dcpl_114 & (~ (fsm_output[8]));
  assign and_dcpl_367 = nor_609_cse & (~ (fsm_output[2]));
  assign and_825_cse = (fsm_output[6]) & (fsm_output[0]);
  assign and_dcpl_371 = (~ (fsm_output[4])) & (fsm_output[7]);
  assign and_827_cse = and_dcpl_371 & (~ (fsm_output[1]));
  assign and_830_cse = and_dcpl_91 & (~ (fsm_output[8]));
  assign nor_1670_cse = ~((fsm_output[6]) | (fsm_output[0]));
  assign and_835_cse = and_dcpl_344 & (~ (fsm_output[1]));
  assign and_dcpl_383 = (fsm_output[3]) & (fsm_output[5]) & (fsm_output[8]);
  assign and_842_cse = and_dcpl_371 & (fsm_output[1]);
  assign and_dcpl_390 = nor_609_cse & (fsm_output[2]);
  assign and_dcpl_393 = (fsm_output[4]) & (fsm_output[7]);
  assign and_849_cse = and_dcpl_393 & (fsm_output[1]);
  assign and_dcpl_403 = and_dcpl_33 & (fsm_output[2]);
  assign and_dcpl_411 = and_dcpl_33 & (~ (fsm_output[2]));
  assign and_dcpl_412 = and_dcpl_411 & and_dcpl_383;
  assign and_870_cse = and_dcpl_91 & (fsm_output[8]);
  assign and_873_cse = and_dcpl_393 & (~ (fsm_output[1]));
  assign and_dcpl_422 = and_dcpl_39 & (~ (fsm_output[8]));
  assign and_dcpl_428 = and_dcpl_59 & (fsm_output[2]);
  assign and_dcpl_432 = and_dcpl_428 & and_dcpl_383;
  assign and_dcpl_446 = and_816_cse & (~ (fsm_output[1]));
  assign and_dcpl_453 = and_dcpl_340 & and_dcpl_39 & (~ (fsm_output[8])) & and_dcpl_446
      & and_dcpl_333;
  assign and_dcpl_460 = and_dcpl_340 & and_820_cse & and_816_cse & (fsm_output[1])
      & and_815_cse;
  assign and_dcpl_468 = and_dcpl_340 & and_830_cse & and_dcpl_371 & (~ (fsm_output[1]))
      & and_825_cse;
  assign and_dcpl_472 = (fsm_output[2]) & (~ (fsm_output[9]));
  assign and_dcpl_473 = and_dcpl_472 & (~ (fsm_output[10]));
  assign and_dcpl_475 = and_dcpl_473 & and_dcpl_114 & (fsm_output[8]) & and_842_cse
      & and_dcpl_333;
  assign and_dcpl_481 = and_dcpl_473 & and_dcpl_39 & (fsm_output[8]) & and_849_cse
      & and_815_cse;
  assign and_dcpl_486 = (fsm_output[2]) & (fsm_output[9]) & (~ (fsm_output[10]))
      & and_820_cse & and_dcpl_446 & and_825_cse;
  assign and_dcpl_488 = (~ (fsm_output[4])) & (~ (fsm_output[7])) & (fsm_output[1]);
  assign and_dcpl_493 = (~ (fsm_output[2])) & (fsm_output[9]) & (~ (fsm_output[10]));
  assign and_dcpl_494 = and_dcpl_493 & and_dcpl_383;
  assign and_dcpl_495 = and_dcpl_494 & and_dcpl_488 & and_dcpl_333;
  assign and_dcpl_500 = and_dcpl_493 & and_870_cse & and_849_cse & nor_1670_cse;
  assign and_dcpl_503 = and_dcpl_494 & and_873_cse & and_825_cse;
  assign and_dcpl_505 = and_dcpl_472 & (fsm_output[10]);
  assign and_dcpl_507 = and_dcpl_505 & and_830_cse & and_842_cse & and_825_cse;
  assign and_dcpl_510 = and_dcpl_505 & and_dcpl_383 & and_dcpl_488 & nor_1670_cse;
  assign and_dcpl_513 = and_dcpl_505 & and_870_cse & and_873_cse & and_dcpl_333;
  assign and_dcpl_531 = nor_609_cse & (fsm_output[2]) & and_dcpl_39 & (fsm_output[8])
      & and_dcpl_393 & (fsm_output[1]) & (fsm_output[6]) & (~ (fsm_output[0]));
  assign and_dcpl_539 = (~ (fsm_output[10])) & (fsm_output[9]) & (~ (fsm_output[2]))
      & and_dcpl_383;
  assign and_dcpl_540 = and_dcpl_539 & and_dcpl_488 & and_dcpl_333;
  assign and_dcpl_544 = and_dcpl_539 & and_873_cse & and_825_cse;
  assign and_dcpl_551 = (fsm_output[10]) & (~ (fsm_output[9])) & (fsm_output[2]);
  assign and_dcpl_553 = and_dcpl_551 & and_dcpl_91 & (~ (fsm_output[8])) & (~ (fsm_output[4]))
      & (fsm_output[7]) & (fsm_output[1]) & and_825_cse;
  assign and_dcpl_557 = and_dcpl_551 & and_dcpl_383 & and_dcpl_488 & (~ (fsm_output[6]))
      & (~ (fsm_output[0]));
  assign and_dcpl_561 = and_dcpl_551 & and_dcpl_91 & (fsm_output[8]) & and_873_cse
      & and_dcpl_333;
  assign and_dcpl_567 = ~((fsm_output[3]) | (fsm_output[5]) | (fsm_output[8]));
  assign and_dcpl_568 = ~((fsm_output[2]) | (fsm_output[9]));
  assign and_dcpl_569 = and_dcpl_568 & (~ (fsm_output[10]));
  assign and_dcpl_594 = (fsm_output[2]) & (fsm_output[9]) & (~ (fsm_output[10]));
  assign and_dcpl_627 = and_dcpl_340 & and_dcpl_338;
  assign and_dcpl_628 = and_dcpl_627 & and_816_cse & (~ (fsm_output[1])) & and_dcpl_333;
  assign and_dcpl_631 = ~((fsm_output[4]) | (fsm_output[7]) | (fsm_output[1]));
  assign and_dcpl_636 = and_dcpl_340 & (fsm_output[3]) & (fsm_output[5]) & (fsm_output[8])
      & and_dcpl_631 & (~ (fsm_output[6])) & (~ (fsm_output[0]));
  assign and_dcpl_642 = (fsm_output[10]) & (~ (fsm_output[9])) & (~ (fsm_output[2]))
      & and_dcpl_338 & and_dcpl_631 & (fsm_output[6]) & (~ (fsm_output[0]));
  assign or_tmp_3282 = (fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[9]))
      | (fsm_output[8]) | (fsm_output[6]);
  assign not_tmp_834 = ~((fsm_output[8]) & (fsm_output[6]));
  assign not_tmp_835 = ~((fsm_output[9]) & (fsm_output[8]) & (fsm_output[6]));
  assign nor_1657_cse = ~((fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[10]))
      | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[6]));
  assign or_3467_nl = (fsm_output[1]) | (~ (fsm_output[2])) | (~ (fsm_output[9]))
      | (~ (fsm_output[8])) | (fsm_output[6]);
  assign or_3466_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]) | (~ (fsm_output[8]))
      | (fsm_output[6]);
  assign mux_3809_nl = MUX_s_1_2_2(or_3467_nl, or_3466_nl, fsm_output[0]);
  assign or_3465_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[6]);
  assign mux_3810_nl = MUX_s_1_2_2(mux_3809_nl, or_3465_nl, fsm_output[10]);
  assign nor_1648_nl = ~((fsm_output[4:3]!=2'b00) | mux_3810_nl);
  assign nor_1649_nl = ~((~ (fsm_output[4])) | (fsm_output[10]) | (fsm_output[0])
      | (~ (fsm_output[1])) | (~ (fsm_output[2])) | (~ (fsm_output[9])) | (fsm_output[8])
      | (fsm_output[6]));
  assign nor_1650_nl = ~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]) | not_tmp_834);
  assign nor_1651_nl = ~((fsm_output[2:1]!=2'b01) | not_tmp_835);
  assign mux_3805_nl = MUX_s_1_2_2(nor_1650_nl, nor_1651_nl, fsm_output[0]);
  assign nor_1652_nl = ~((fsm_output[0]) | (~ (fsm_output[1])) | (~ (fsm_output[2]))
      | (fsm_output[9]) | not_tmp_834);
  assign mux_3806_nl = MUX_s_1_2_2(mux_3805_nl, nor_1652_nl, fsm_output[10]);
  assign or_3456_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[6]);
  assign mux_3804_nl = MUX_s_1_2_2(or_tmp_3282, or_3456_nl, fsm_output[0]);
  assign and_nl = (fsm_output[10]) & (~ mux_3804_nl);
  assign mux_3807_nl = MUX_s_1_2_2(mux_3806_nl, and_nl, fsm_output[4]);
  assign mux_3808_nl = MUX_s_1_2_2(nor_1649_nl, mux_3807_nl, fsm_output[3]);
  assign mux_3811_nl = MUX_s_1_2_2(nor_1648_nl, mux_3808_nl, fsm_output[5]);
  assign nor_1653_nl = ~((fsm_output[2:0]!=3'b010) | not_tmp_835);
  assign nor_1654_nl = ~((~ (fsm_output[0])) | (fsm_output[1]) | (~ (fsm_output[2]))
      | (fsm_output[9]) | not_tmp_834);
  assign mux_3801_nl = MUX_s_1_2_2(nor_1653_nl, nor_1654_nl, fsm_output[10]);
  assign and_1158_nl = (fsm_output[4]) & mux_3801_nl;
  assign nor_1655_nl = ~((fsm_output[10]) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (~ (fsm_output[2])) | (fsm_output[9]) | not_tmp_834);
  assign or_3448_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[9]) | (fsm_output[8])
      | (fsm_output[6]);
  assign mux_3828_nl = MUX_s_1_2_2(or_3448_nl, or_tmp_3282, fsm_output[0]);
  assign nor_1656_nl = ~((fsm_output[10]) | mux_3828_nl);
  assign mux_3800_nl = MUX_s_1_2_2(nor_1655_nl, nor_1656_nl, fsm_output[4]);
  assign mux_3802_nl = MUX_s_1_2_2(and_1158_nl, mux_3800_nl, fsm_output[3]);
  assign mux_3803_nl = MUX_s_1_2_2(mux_3802_nl, nor_1657_cse, fsm_output[5]);
  assign not_tmp_838 = MUX_s_1_2_2(mux_3811_nl, mux_3803_nl, fsm_output[7]);
  assign and_dcpl_647 = and_dcpl_340 & (~ (fsm_output[3])) & (~ (fsm_output[5]))
      & (~ (fsm_output[8])) & and_dcpl_631 & and_dcpl_333;
  assign and_dcpl_650 = and_dcpl_627 & and_816_cse & (fsm_output[1]) & and_dcpl_333;
  assign and_dcpl_660 = (fsm_output[2]) & (fsm_output[9]) & (~ (fsm_output[10]))
      & and_dcpl_91 & (~ (fsm_output[8])) & (~ (fsm_output[4])) & (fsm_output[7])
      & (~ (fsm_output[1])) & and_815_cse;
  assign and_dcpl_669 = (fsm_output[2]) & (~ (fsm_output[9])) & (fsm_output[10])
      & (fsm_output[3]) & (fsm_output[5]) & (fsm_output[8]) & and_dcpl_393 & (~ (fsm_output[1]))
      & and_815_cse;
  assign and_dcpl_678 = (~ (fsm_output[2])) & (~ (fsm_output[9])) & (~ (fsm_output[10]))
      & (fsm_output[3]) & (~ (fsm_output[5])) & (~ (fsm_output[8])) & (fsm_output[4])
      & (~ (fsm_output[7])) & (fsm_output[1]) & and_815_cse;
  assign and_dcpl_686 = (~ (fsm_output[2])) & (fsm_output[9]) & (~ (fsm_output[10]))
      & and_dcpl_91 & (fsm_output[8]) & and_dcpl_393 & (fsm_output[1]) & (~ (fsm_output[6]))
      & (~ (fsm_output[0]));
  assign or_tmp_3307 = (~ (fsm_output[9])) | (fsm_output[10]) | (fsm_output[1]) |
      (~ (fsm_output[2]));
  assign or_tmp_3312 = (~ (fsm_output[9])) | (fsm_output[10]) | (~ (fsm_output[1]))
      | (fsm_output[2]);
  assign mux_3821_nl = MUX_s_1_2_2(nor_758_cse, and_529_cse, fsm_output[10]);
  assign or_tmp_3326 = (fsm_output[9]) | (~ mux_3821_nl);
  assign and_978_ssc = nor_609_cse & (~ (fsm_output[2])) & and_dcpl_39 & (~ (fsm_output[8]))
      & (fsm_output[4]) & (~ (fsm_output[7])) & (~ (fsm_output[1])) & and_dcpl_333;
  assign and_824_ssc = and_dcpl_367 & and_820_cse & and_816_cse & (fsm_output[1])
      & and_815_cse;
  assign COMP_LOOP_or_54_ssc = (and_dcpl_367 & and_830_cse & and_827_cse & and_825_cse)
      | (and_dcpl_367 & and_dcpl_383 & and_835_cse & nor_1670_cse) | (and_dcpl_390
      & and_dcpl_114 & (fsm_output[8]) & and_842_cse & and_dcpl_333) | (and_dcpl_403
      & and_820_cse & and_816_cse & (~ (fsm_output[1])) & and_825_cse) | (and_dcpl_403
      & and_830_cse & and_827_cse & and_815_cse) | (and_dcpl_59 & (~ (fsm_output[2]))
      & and_dcpl_422 & and_835_cse & and_815_cse) | (and_dcpl_432 & and_873_cse &
      and_815_cse) | ((fsm_output[10]) & (fsm_output[9]) & (~ (fsm_output[2])) &
      and_dcpl_422 & and_dcpl_345 & and_825_cse);
  assign COMP_LOOP_or_55_ssc = (and_dcpl_390 & and_dcpl_39 & (fsm_output[8]) & and_849_cse
      & and_815_cse) | (and_dcpl_412 & and_dcpl_345 & and_dcpl_333) | (and_dcpl_412
      & and_873_cse & and_825_cse) | (and_dcpl_428 & and_830_cse & and_842_cse &
      and_825_cse) | (and_dcpl_432 & and_dcpl_345 & nor_1670_cse) | (and_dcpl_428
      & and_870_cse & and_873_cse & and_dcpl_333);
  assign and_872_ssc = and_dcpl_411 & and_870_cse & and_849_cse & nor_1670_cse;
  assign mux_3829_nl = MUX_s_1_2_2(mux_tmp_227, or_tmp_104, and_526_cse);
  assign or_3510_nl = (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign mux_tmp_3828 = MUX_s_1_2_2(mux_3829_nl, or_3510_nl, fsm_output[2]);
  assign mux_tmp_3830 = MUX_s_1_2_2(mux_tmp_227, or_tmp_104, fsm_output[1]);
  assign nor_tmp_549 = or_2400_cse & (fsm_output[10]);
  assign or_tmp_3337 = nor_753_cse | (fsm_output[10:9]!=2'b00);
  assign or_tmp_3339 = nor_297_cse | (fsm_output[10]);
  assign mux_tmp_3839 = MUX_s_1_2_2(or_tmp_3339, and_757_cse, or_2644_cse);
  assign mux_3842_nl = MUX_s_1_2_2(and_757_cse, mux_tmp_227, or_3388_cse);
  assign or_3520_nl = and_526_cse | (fsm_output[10:9]!=2'b10);
  assign mux_tmp_3841 = MUX_s_1_2_2(mux_3842_nl, or_3520_nl, fsm_output[2]);
  assign or_tmp_3344 = (~ (fsm_output[3])) | (~ (fsm_output[2])) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (fsm_output[10]);
  assign nor_tmp_552 = or_2421_cse & (fsm_output[10]);
  assign or_tmp_3347 = nor_303_cse | (fsm_output[10]);
  assign or_3527_nl = (~ (fsm_output[2])) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (fsm_output[10]);
  assign mux_3849_nl = MUX_s_1_2_2(or_tmp_3347, nor_tmp_552, fsm_output[2]);
  assign mux_tmp_3848 = MUX_s_1_2_2(or_3527_nl, mux_3849_nl, fsm_output[3]);
  assign nor_tmp_554 = or_2419_cse & (fsm_output[10]);
  assign or_tmp_3352 = and_521_cse | (fsm_output[10]);
  assign mux_tmp_3856 = MUX_s_1_2_2(or_tmp_3352, nor_tmp_554, fsm_output[2]);
  assign mux_tmp_3864 = MUX_s_1_2_2(or_tmp_3337, nor_tmp_549, fsm_output[2]);
  assign or_tmp_3357 = (fsm_output[2]) | and_526_cse | (~ and_757_cse);
  assign nor_1704_cse = ~(COMP_LOOP_nor_11_itm | (fsm_output[6]));
  assign or_tmp_3381 = (fsm_output[10]) | nor_1704_cse | (fsm_output[2]) | (~ (fsm_output[9]));
  assign or_tmp_3382 = ~((fsm_output[10]) & COMP_LOOP_nor_11_itm & (fsm_output[6])
      & (fsm_output[2]) & (~ (fsm_output[9])));
  assign or_tmp_3384 = nor_1704_cse | (~ (fsm_output[2])) | (fsm_output[9]);
  assign or_3564_nl = (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[6])) | (fsm_output[2])
      | (fsm_output[9]);
  assign mux_3893_nl = MUX_s_1_2_2(or_3564_nl, or_tmp_3384, fsm_output[10]);
  assign mux_tmp_3892 = MUX_s_1_2_2(mux_3893_nl, or_tmp_3382, fsm_output[1]);
  assign not_tmp_882 = ~(COMP_LOOP_nor_11_itm & (fsm_output[6]) & (fsm_output[2])
      & (fsm_output[9]));
  assign not_tmp_883 = ~((fsm_output[2]) & (fsm_output[9]));
  assign or_tmp_3402 = (~ (fsm_output[6])) | (fsm_output[2]) | (~ (fsm_output[9]));
  assign mux_3904_nl = MUX_s_1_2_2(not_tmp_883, or_2855_cse, fsm_output[6]);
  assign mux_tmp_3903 = MUX_s_1_2_2(or_tmp_3402, mux_3904_nl, COMP_LOOP_nor_11_itm);
  assign or_tmp_3403 = (fsm_output[10]) | mux_tmp_3903;
  assign or_3586_nl = (fsm_output[6]) | (fsm_output[2]) | (fsm_output[9]);
  assign or_3585_nl = (~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign mux_tmp_3906 = MUX_s_1_2_2(or_3586_nl, or_3585_nl, fsm_output[10]);
  assign or_3584_nl = (~ COMP_LOOP_nor_11_itm) | (fsm_output[6]) | (fsm_output[2])
      | (fsm_output[9]);
  assign or_3583_nl = (fsm_output[6]) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign mux_3907_nl = MUX_s_1_2_2(or_3584_nl, or_3583_nl, fsm_output[10]);
  assign mux_tmp_3907 = MUX_s_1_2_2(mux_tmp_3906, mux_3907_nl, fsm_output[1]);
  assign or_tmp_3409 = (fsm_output[10]) | (fsm_output[6]) | not_tmp_883;
  assign COMP_LOOP_or_61_itm = and_dcpl_460 | and_dcpl_468 | and_dcpl_475 | and_dcpl_481
      | and_dcpl_486 | and_dcpl_495 | and_dcpl_500 | and_dcpl_503 | and_dcpl_507
      | and_dcpl_510 | and_dcpl_513;
  assign COMP_LOOP_or_24_itm = and_dcpl_531 | and_dcpl_540 | and_dcpl_544 | and_dcpl_553
      | and_dcpl_557 | and_dcpl_561;
  assign COMP_LOOP_nor_633_itm = ~(and_dcpl_628 | and_dcpl_636 | and_dcpl_642);
  assign COMP_LOOP_nor_685_itm = ~(and_dcpl_636 | and_dcpl_642);
  assign COMP_LOOP_or_65_itm = and_dcpl_636 | and_dcpl_642;
  assign COMP_LOOP_nor_687_itm = ~(and_dcpl_636 | and_dcpl_642 | not_tmp_838 | and_dcpl_650);
  always @(posedge clk) begin
    if ( ~ not_tmp_208 ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( (and_dcpl_93 & and_dcpl_88) | STAGE_LOOP_i_3_0_sva_mx0c1 ) begin
      STAGE_LOOP_i_3_0_sva <= MUX_v_4_2_2(4'b0001, STAGE_LOOP_i_3_0_sva_2, STAGE_LOOP_i_3_0_sva_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( ~ not_tmp_208 ) begin
      r_sva <= r_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= 1'b0;
      COMP_LOOP_nor_11_itm <= 1'b0;
      modExp_exp_1_7_1_sva <= 1'b0;
      COMP_LOOP_nor_12_itm <= 1'b0;
      COMP_LOOP_nor_134_itm <= 1'b0;
      COMP_LOOP_nor_137_itm <= 1'b0;
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_nor_1_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_139_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_140_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_141_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_143_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_144_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_145_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_146_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_147_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_148_itm <= 1'b0;
      COMP_LOOP_COMP_LOOP_and_149_itm <= 1'b0;
    end
    else begin
      reg_vec_rsc_triosy_0_15_obj_ld_cse <= and_dcpl_103 & and_dcpl_2 & and_757_cse
          & (~ STAGE_LOOP_acc_itm_2_1);
      COMP_LOOP_nor_11_itm <= (COMP_LOOP_mux1h_428_nl & (mux_2989_nl | (fsm_output[0])))
          | (mux_3077_nl & (fsm_output[0]));
      modExp_exp_1_7_1_sva <= COMP_LOOP_mux1h_464_nl & mux_3521_nl;
      COMP_LOOP_nor_12_itm <= (COMP_LOOP_mux1h_474_nl & mux_3542_nl) | mux_3636_nl;
      COMP_LOOP_nor_134_itm <= (COMP_LOOP_mux1h_477_nl & mux_3649_nl) | mux_3656_nl;
      COMP_LOOP_nor_137_itm <= (COMP_LOOP_mux1h_479_nl & (mux_3663_nl | (fsm_output[10])))
          | mux_3670_nl;
      COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm <= COMP_LOOP_mux1h_480_nl & (~ and_dcpl_257);
      COMP_LOOP_COMP_LOOP_nor_1_itm <= ~((z_out_2_12_1[3:0]!=4'b0000));
      COMP_LOOP_COMP_LOOP_and_139_itm <= (z_out_2_12_1[3:0]==4'b0101);
      COMP_LOOP_COMP_LOOP_and_140_itm <= (z_out_2_12_1[3:0]==4'b0110);
      COMP_LOOP_COMP_LOOP_and_141_itm <= (z_out_2_12_1[3:0]==4'b0111);
      COMP_LOOP_COMP_LOOP_and_143_itm <= (z_out_2_12_1[3:0]==4'b1001);
      COMP_LOOP_COMP_LOOP_and_144_itm <= (z_out_2_12_1[3:0]==4'b1010);
      COMP_LOOP_COMP_LOOP_and_145_itm <= (z_out_2_12_1[3:0]==4'b1011);
      COMP_LOOP_COMP_LOOP_and_146_itm <= (z_out_2_12_1[3:0]==4'b1100);
      COMP_LOOP_COMP_LOOP_and_147_itm <= (z_out_2_12_1[3:0]==4'b1101);
      COMP_LOOP_COMP_LOOP_and_148_itm <= (z_out_2_12_1[3:0]==4'b1110);
      COMP_LOOP_COMP_LOOP_and_149_itm <= (z_out_2_12_1[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    modulo_result_rem_cmp_a <= MUX1HOT_v_64_6_2(z_out_8, operator_64_false_acc_mut_63_0,
        COMP_LOOP_10_acc_8_itm, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, COMP_LOOP_10_mul_mut,
        COMP_LOOP_1_acc_5_mut_mx0w5, {modulo_result_or_nl , (~ mux_2231_nl) , (~
        mux_2331_nl) , (~ mux_2346_nl) , (~ mux_2418_nl) , not_tmp_441});
    modulo_result_rem_cmp_b <= p_sva;
    operator_66_true_div_cmp_a <= MUX_v_65_2_2(z_out_6, ({operator_64_false_acc_mut_64
        , operator_64_false_acc_mut_63_0}), and_dcpl_241);
    operator_66_true_div_cmp_b_9_0 <= MUX_v_10_2_2(STAGE_LOOP_lshift_psp_sva_mx0w0,
        STAGE_LOOP_lshift_psp_sva, and_dcpl_241);
  end
  always @(posedge clk) begin
    if ( ~ mux_2452_nl ) begin
      STAGE_LOOP_lshift_psp_sva <= STAGE_LOOP_lshift_psp_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_3889_nl ) begin
      operator_64_false_acc_mut_64 <= operator_64_false_mux1h_2_rgt[64];
    end
  end
  always @(posedge clk) begin
    if ( ~ mux_3943_nl ) begin
      operator_64_false_acc_mut_63_0 <= operator_64_false_mux1h_2_rgt[63:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      VEC_LOOP_j_sva_11_0 <= 12'b000000000000;
    end
    else if ( and_dcpl_247 | VEC_LOOP_j_sva_11_0_mx0c1 ) begin
      VEC_LOOP_j_sva_11_0 <= MUX_v_12_2_2(12'b000000000000, (z_out[11:0]), VEC_LOOP_j_sva_11_0_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_k_9_4_sva_4_0 <= 5'b00000;
    end
    else if ( mux_3946_nl & (~((fsm_output[8]) | (fsm_output[2]))) ) begin
      COMP_LOOP_k_9_4_sva_4_0 <= MUX_v_5_2_2(5'b00000, (z_out_1[4:0]), or_3508_nl);
    end
  end
  always @(posedge clk) begin
    if ( (modExp_while_and_3 | modExp_while_and_5 | modExp_result_sva_mx0c0 | (~
        mux_2668_nl)) & (modExp_result_sva_mx0c0 | modExp_result_and_rgt | modExp_result_and_1_rgt)
        ) begin
      modExp_result_sva <= MUX1HOT_v_64_3_2(64'b0000000000000000000000000000000000000000000000000000000000000001,
          modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w6, {modExp_result_sva_mx0c0
          , modExp_result_and_rgt , modExp_result_and_1_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      tmp_10_lpi_4_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( MUX_s_1_2_2(mux_2741_nl, mux_2714_nl, fsm_output[4]) ) begin
      tmp_10_lpi_4_dfm <= MUX1HOT_v_64_17_2(({1'b0 , operator_64_false_slc_modExp_exp_63_1_3}),
          vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d, vec_rsc_0_3_i_qa_d,
          vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d, vec_rsc_0_7_i_qa_d,
          vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d, vec_rsc_0_11_i_qa_d,
          vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d, vec_rsc_0_15_i_qa_d,
          {and_dcpl_247 , COMP_LOOP_or_8_nl , COMP_LOOP_or_9_nl , COMP_LOOP_or_10_nl
          , COMP_LOOP_or_11_nl , COMP_LOOP_or_12_nl , COMP_LOOP_or_13_nl , COMP_LOOP_or_14_nl
          , COMP_LOOP_or_15_nl , COMP_LOOP_or_16_nl , COMP_LOOP_or_17_nl , COMP_LOOP_or_18_nl
          , COMP_LOOP_or_19_nl , COMP_LOOP_or_20_nl , COMP_LOOP_or_21_nl , COMP_LOOP_or_22_nl
          , COMP_LOOP_or_23_nl});
    end
  end
  always @(posedge clk) begin
    if ( MUX_s_1_2_2(mux_2981_nl, mux_2925_nl, fsm_output[1]) ) begin
      COMP_LOOP_10_mul_mut <= MUX1HOT_v_64_21_2(r_sva, modulo_result_rem_cmp_z, modulo_qr_sva_1_mx0w6,
          modExp_result_sva, vec_rsc_0_0_i_qa_d, vec_rsc_0_1_i_qa_d, vec_rsc_0_2_i_qa_d,
          vec_rsc_0_3_i_qa_d, vec_rsc_0_4_i_qa_d, vec_rsc_0_5_i_qa_d, vec_rsc_0_6_i_qa_d,
          vec_rsc_0_7_i_qa_d, vec_rsc_0_8_i_qa_d, vec_rsc_0_9_i_qa_d, vec_rsc_0_10_i_qa_d,
          vec_rsc_0_11_i_qa_d, vec_rsc_0_12_i_qa_d, vec_rsc_0_13_i_qa_d, vec_rsc_0_14_i_qa_d,
          vec_rsc_0_15_i_qa_d, COMP_LOOP_1_modExp_1_while_if_mul_mut_1, {and_312_nl
          , COMP_LOOP_or_29_nl , COMP_LOOP_or_30_nl , (~ mux_2757_itm) , COMP_LOOP_and_277_nl
          , COMP_LOOP_COMP_LOOP_and_932_nl , COMP_LOOP_COMP_LOOP_and_934_nl , COMP_LOOP_and_1_nl
          , COMP_LOOP_COMP_LOOP_and_936_nl , COMP_LOOP_and_2_nl , COMP_LOOP_and_3_nl
          , COMP_LOOP_and_4_nl , COMP_LOOP_COMP_LOOP_and_930_nl , COMP_LOOP_and_5_nl
          , COMP_LOOP_and_6_nl , COMP_LOOP_and_7_nl , COMP_LOOP_and_8_nl , COMP_LOOP_and_9_nl
          , COMP_LOOP_and_10_nl , COMP_LOOP_and_11_nl , (~ mux_129_nl)});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= 1'b0;
    end
    else if ( and_dcpl_237 | and_dcpl_304 | and_dcpl_117 | and_dcpl_130 | and_dcpl_140
        | and_dcpl_149 | and_dcpl_155 | and_dcpl_164 | and_dcpl_171 | and_dcpl_178
        | and_dcpl_185 | and_dcpl_189 | and_dcpl_197 | and_dcpl_202 | and_dcpl_211
        | and_dcpl_219 | and_dcpl_226 | and_dcpl_231 ) begin
      COMP_LOOP_COMP_LOOP_and_137_itm <= MUX1HOT_s_1_3_2((~ (z_out_1[63])), (~ (z_out_6[8])),
          COMP_LOOP_COMP_LOOP_and_17_nl, {and_dcpl_237 , and_dcpl_304 , COMP_LOOP_or_32_cse});
    end
  end
  always @(posedge clk) begin
    if ( mux_3288_nl | not_tmp_441 ) begin
      COMP_LOOP_10_acc_8_itm <= MUX_v_64_2_2(z_out_8, COMP_LOOP_1_acc_8_nl, not_tmp_441);
    end
  end
  always @(posedge clk) begin
    if ( ~((fsm_output[3]) | (~ (fsm_output[5])) | (fsm_output[2]) | or_3079_cse
        | (~ (fsm_output[4])) | (fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[9])
        | (fsm_output[10])) ) begin
      COMP_LOOP_acc_psp_sva <= COMP_LOOP_acc_psp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_nor_itm <= ~((VEC_LOOP_j_sva_11_0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_305_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_305_itm <= (COMP_LOOP_acc_1_cse_6_sva_1[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_62_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_62_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_2_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_2_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0011);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_64_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_64_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_4_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_4_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_5_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_5_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_6_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_6_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b0111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_68_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_68_itm <= (COMP_LOOP_acc_1_cse_2_sva_1[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_8_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_8_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1001);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_9_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_9_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1010);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_10_itm <= 1'b0;
    end
    else if ( MUX_s_1_2_2(mux_3334_nl, and_757_cse, fsm_output[8]) ) begin
      COMP_LOOP_COMP_LOOP_and_10_itm <= MUX_s_1_2_2(COMP_LOOP_COMP_LOOP_and_10_nl,
          (~ (readslicef_10_1_9(COMP_LOOP_1_acc_nl))), and_dcpl_231);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_11_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1100);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_12_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_12_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1101);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_13_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_13_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1110);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_COMP_LOOP_and_14_itm <= 1'b0;
    end
    else if ( ~ not_tmp_619 ) begin
      COMP_LOOP_COMP_LOOP_and_14_itm <= (VEC_LOOP_j_sva_11_0[3:0]==4'b1111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_6_sva <= 12'b000000000000;
    end
    else if ( mux_3340_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_1_cse_6_sva <= COMP_LOOP_acc_1_cse_6_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_2_sva <= 12'b000000000000;
    end
    else if ( mux_3350_nl | (fsm_output[10:8]!=3'b000) ) begin
      COMP_LOOP_acc_1_cse_2_sva <= COMP_LOOP_acc_1_cse_2_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_11_psp_sva <= 11'b00000000000;
    end
    else if ( ~((~ mux_3355_nl) & nor_609_cse) ) begin
      COMP_LOOP_acc_11_psp_sva <= nl_COMP_LOOP_acc_11_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_4_sva <= 12'b000000000000;
    end
    else if ( ~((~ mux_3359_nl) & nor_609_cse) ) begin
      COMP_LOOP_acc_1_cse_4_sva <= z_out_6[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_13_psp_sva <= 10'b0000000000;
    end
    else if ( ~(mux_3364_nl & (~ (fsm_output[10]))) ) begin
      COMP_LOOP_acc_13_psp_sva <= z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_14_psp_sva <= 11'b00000000000;
    end
    else if ( mux_3367_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_14_psp_sva <= nl_COMP_LOOP_acc_14_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_8_sva <= 12'b000000000000;
    end
    else if ( mux_3372_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_1_cse_8_sva <= nl_COMP_LOOP_acc_1_cse_8_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_16_psp_sva <= 9'b000000000;
    end
    else if ( mux_3375_nl | (fsm_output[10]) ) begin
      COMP_LOOP_acc_16_psp_sva <= z_out_1[8:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_10_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_tmp_3378, mux_3381_nl, fsm_output[5]) ) begin
      COMP_LOOP_acc_1_cse_10_sva <= nl_COMP_LOOP_acc_1_cse_10_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_17_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(mux_3386_nl, (fsm_output[10]), or_470_cse) ) begin
      COMP_LOOP_acc_17_psp_sva <= nl_COMP_LOOP_acc_17_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_12_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3391_nl, (fsm_output[10]), or_470_cse) ) begin
      COMP_LOOP_acc_1_cse_12_sva <= nl_COMP_LOOP_acc_1_cse_12_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_19_psp_sva <= 10'b0000000000;
    end
    else if ( MUX_s_1_2_2(mux_3396_nl, (fsm_output[10]), fsm_output[9]) ) begin
      COMP_LOOP_acc_19_psp_sva <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_14_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3400_nl, (fsm_output[10]), fsm_output[9]) ) begin
      COMP_LOOP_acc_1_cse_14_sva <= nl_COMP_LOOP_acc_1_cse_14_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_20_psp_sva <= 11'b00000000000;
    end
    else if ( MUX_s_1_2_2(nor_1680_nl, and_1162_nl, fsm_output[9]) ) begin
      COMP_LOOP_acc_20_psp_sva <= nl_COMP_LOOP_acc_20_psp_sva[10:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_1_cse_sva <= 12'b000000000000;
    end
    else if ( MUX_s_1_2_2(mux_3408_nl, and_757_cse, fsm_output[8]) ) begin
      COMP_LOOP_acc_1_cse_sva <= nl_COMP_LOOP_acc_1_cse_sva[11:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      modExp_exp_1_6_1_sva <= 1'b0;
      modExp_exp_1_5_1_sva <= 1'b0;
      modExp_exp_1_4_1_sva <= 1'b0;
    end
    else if ( mux_3494_itm ) begin
      modExp_exp_1_6_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0[2]), modExp_exp_1_7_1_sva,
          (COMP_LOOP_k_9_4_sva_4_0[3]), {and_dcpl_257 , not_tmp_701 , not_tmp_688});
      modExp_exp_1_5_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0[1]), modExp_exp_1_6_1_sva,
          (COMP_LOOP_k_9_4_sva_4_0[2]), {and_dcpl_257 , not_tmp_701 , not_tmp_688});
      modExp_exp_1_4_1_sva <= MUX1HOT_s_1_3_2((COMP_LOOP_k_9_4_sva_4_0[0]), modExp_exp_1_5_1_sva,
          (COMP_LOOP_k_9_4_sva_4_0[1]), {and_dcpl_257 , not_tmp_701 , not_tmp_688});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= 12'b000000000000;
    end
    else if ( COMP_LOOP_or_32_cse ) begin
      COMP_LOOP_acc_10_cse_12_1_1_sva <= z_out_2_12_1;
    end
  end
  always @(posedge clk) begin
    if ( and_dcpl_117 | not_tmp_446 | and_dcpl_130 | and_dcpl_149 | and_dcpl_155
        | and_dcpl_164 | and_dcpl_178 | and_dcpl_185 | and_dcpl_189 | and_dcpl_202
        | and_dcpl_211 | and_dcpl_219 ) begin
      COMP_LOOP_10_slc_COMP_LOOP_acc_9_itm <= MUX_s_1_2_2((z_out_3[9]), (z_out_6[8]),
          not_tmp_446);
    end
  end
  assign modulo_result_or_nl = and_dcpl_237 | not_tmp_446;
  assign mux_2225_nl = MUX_s_1_2_2((fsm_output[7]), and_395_cse, or_2377_cse);
  assign mux_2226_nl = MUX_s_1_2_2(mux_2225_nl, mux_tmp_2172, fsm_output[9]);
  assign nand_195_nl = ~(nand_196_cse & mux_2926_cse);
  assign mux_2224_nl = MUX_s_1_2_2(nand_195_nl, or_tmp_2277, fsm_output[9]);
  assign mux_2227_nl = MUX_s_1_2_2((~ mux_2226_nl), mux_2224_nl, fsm_output[6]);
  assign or_2375_nl = (fsm_output[2:0]!=3'b000);
  assign mux_2221_nl = MUX_s_1_2_2(or_tmp_2280, (~ (fsm_output[7])), or_2375_nl);
  assign mux_2222_nl = MUX_s_1_2_2(mux_2221_nl, or_tmp_2280, fsm_output[9]);
  assign mux_2219_nl = MUX_s_1_2_2(or_tmp_2276, (fsm_output[7]), and_527_cse);
  assign mux_2220_nl = MUX_s_1_2_2(mux_2219_nl, or_tmp_2297, fsm_output[9]);
  assign mux_2223_nl = MUX_s_1_2_2(mux_2222_nl, mux_2220_nl, fsm_output[6]);
  assign mux_2228_nl = MUX_s_1_2_2(mux_2227_nl, mux_2223_nl, fsm_output[8]);
  assign or_2373_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[7]) | (~ (fsm_output[10]));
  assign or_2371_nl = and_527_cse | (fsm_output[7]) | (~ (fsm_output[10]));
  assign mux_2216_nl = MUX_s_1_2_2(or_2373_nl, or_2371_nl, fsm_output[9]);
  assign mux_2214_nl = MUX_s_1_2_2(mux_2926_cse, or_tmp_2280, or_2368_cse);
  assign mux_2215_nl = MUX_s_1_2_2((~ (fsm_output[7])), mux_2214_nl, fsm_output[9]);
  assign mux_2217_nl = MUX_s_1_2_2(mux_2216_nl, mux_2215_nl, fsm_output[6]);
  assign mux_2210_nl = MUX_s_1_2_2((fsm_output[7]), mux_2926_cse, and_529_cse);
  assign mux_2211_nl = MUX_s_1_2_2(mux_tmp_2172, mux_2210_nl, fsm_output[0]);
  assign mux_2212_nl = MUX_s_1_2_2(mux_2211_nl, or_tmp_2276, fsm_output[9]);
  assign or_2367_nl = nor_758_cse | (~ (fsm_output[7])) | (fsm_output[10]);
  assign mux_2209_nl = MUX_s_1_2_2(or_2367_nl, or_tmp_2294, fsm_output[9]);
  assign mux_2213_nl = MUX_s_1_2_2(mux_2212_nl, mux_2209_nl, fsm_output[6]);
  assign mux_2218_nl = MUX_s_1_2_2(mux_2217_nl, mux_2213_nl, fsm_output[8]);
  assign mux_2229_nl = MUX_s_1_2_2(mux_2228_nl, mux_2218_nl, fsm_output[5]);
  assign mux_2204_nl = MUX_s_1_2_2(or_tmp_2276, (fsm_output[7]), or_2377_cse);
  assign mux_2205_nl = MUX_s_1_2_2((fsm_output[7]), mux_2204_nl, fsm_output[9]);
  assign mux_2206_nl = MUX_s_1_2_2(mux_2205_nl, mux_2203_cse, fsm_output[6]);
  assign or_2364_nl = (fsm_output[1]) | (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[10]);
  assign mux_2200_nl = MUX_s_1_2_2(or_2364_nl, or_tmp_2274, fsm_output[0]);
  assign mux_2201_nl = MUX_s_1_2_2(mux_tmp_2178, mux_2200_nl, fsm_output[9]);
  assign mux_2197_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_2281, or_2368_cse);
  assign or_2362_nl = and_529_cse | (fsm_output[7]) | (~ (fsm_output[10]));
  assign mux_2198_nl = MUX_s_1_2_2(mux_2197_nl, or_2362_nl, fsm_output[0]);
  assign or_2360_nl = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[10]);
  assign mux_2199_nl = MUX_s_1_2_2(mux_2198_nl, or_2360_nl, fsm_output[9]);
  assign mux_2202_nl = MUX_s_1_2_2(mux_2201_nl, mux_2199_nl, fsm_output[6]);
  assign mux_2207_nl = MUX_s_1_2_2(mux_2206_nl, mux_2202_nl, fsm_output[8]);
  assign mux_2192_nl = MUX_s_1_2_2((~ or_tmp_2280), or_tmp_2281, fsm_output[2]);
  assign mux_2191_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_2281, fsm_output[2]);
  assign mux_2193_nl = MUX_s_1_2_2(mux_2192_nl, mux_2191_nl, and_526_cse);
  assign mux_2194_nl = MUX_s_1_2_2((~ mux_2193_nl), or_tmp_2280, fsm_output[9]);
  assign mux_2190_nl = MUX_s_1_2_2(mux_tmp_2176, or_tmp_2302, fsm_output[9]);
  assign mux_2195_nl = MUX_s_1_2_2(mux_2194_nl, mux_2190_nl, fsm_output[6]);
  assign mux_2187_nl = MUX_s_1_2_2((fsm_output[7]), and_395_cse, and_527_cse);
  assign mux_2188_nl = MUX_s_1_2_2((~ mux_2187_nl), or_tmp_2280, fsm_output[9]);
  assign mux_2189_nl = MUX_s_1_2_2(mux_tmp_2159, mux_2188_nl, fsm_output[6]);
  assign mux_2196_nl = MUX_s_1_2_2(mux_2195_nl, mux_2189_nl, fsm_output[8]);
  assign mux_2208_nl = MUX_s_1_2_2(mux_2207_nl, mux_2196_nl, fsm_output[5]);
  assign mux_2230_nl = MUX_s_1_2_2(mux_2229_nl, mux_2208_nl, fsm_output[4]);
  assign mux_2180_nl = MUX_s_1_2_2(mux_tmp_2178, or_tmp_2302, fsm_output[1]);
  assign mux_2181_nl = MUX_s_1_2_2(mux_2180_nl, or_tmp_2297, fsm_output[0]);
  assign or_2357_nl = (fsm_output[2]) | (~ and_395_cse);
  assign mux_2179_nl = MUX_s_1_2_2(or_2357_nl, mux_tmp_2178, or_3388_cse);
  assign mux_2182_nl = MUX_s_1_2_2(mux_2181_nl, mux_2179_nl, fsm_output[9]);
  assign or_2355_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[10]));
  assign mux_2177_nl = MUX_s_1_2_2(or_2355_nl, mux_tmp_2176, fsm_output[9]);
  assign mux_2183_nl = MUX_s_1_2_2(mux_2182_nl, mux_2177_nl, fsm_output[6]);
  assign mux_2173_nl = MUX_s_1_2_2((~ mux_tmp_2172), or_tmp_2280, fsm_output[9]);
  assign mux_2174_nl = MUX_s_1_2_2(mux_2173_nl, mux_2171_cse, fsm_output[6]);
  assign mux_2184_nl = MUX_s_1_2_2(mux_2183_nl, mux_2174_nl, fsm_output[8]);
  assign or_2351_nl = (fsm_output[9]) | or_tmp_2294;
  assign mux_2167_nl = MUX_s_1_2_2((fsm_output[7]), and_395_cse, or_2368_cse);
  assign or_2347_nl = and_527_cse | (~ (fsm_output[7])) | (fsm_output[10]);
  assign mux_2168_nl = MUX_s_1_2_2((~ mux_2167_nl), or_2347_nl, fsm_output[9]);
  assign mux_2169_nl = MUX_s_1_2_2(or_2351_nl, mux_2168_nl, fsm_output[6]);
  assign mux_2163_nl = MUX_s_1_2_2((~ mux_2926_cse), or_tmp_2276, fsm_output[2]);
  assign mux_2162_nl = MUX_s_1_2_2((~ mux_2926_cse), (fsm_output[7]), fsm_output[2]);
  assign mux_2164_nl = MUX_s_1_2_2(mux_2163_nl, mux_2162_nl, or_3388_cse);
  assign mux_2160_nl = MUX_s_1_2_2(or_tmp_2276, or_tmp_2280, or_2368_cse);
  assign or_2343_nl = (~(nor_758_cse | (fsm_output[7]))) | (fsm_output[10]);
  assign mux_2161_nl = MUX_s_1_2_2(mux_2160_nl, or_2343_nl, fsm_output[0]);
  assign mux_2165_nl = MUX_s_1_2_2((~ mux_2164_nl), mux_2161_nl, fsm_output[9]);
  assign mux_2166_nl = MUX_s_1_2_2(mux_2165_nl, mux_tmp_2159, fsm_output[6]);
  assign mux_2170_nl = MUX_s_1_2_2(mux_2169_nl, mux_2166_nl, fsm_output[8]);
  assign mux_2185_nl = MUX_s_1_2_2(mux_2184_nl, mux_2170_nl, fsm_output[5]);
  assign mux_2154_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_2281, and_527_cse);
  assign mux_2153_nl = MUX_s_1_2_2((fsm_output[7]), or_tmp_2281, and_536_cse);
  assign mux_2155_nl = MUX_s_1_2_2(mux_2154_nl, mux_2153_nl, fsm_output[9]);
  assign mux_2150_nl = MUX_s_1_2_2((~ mux_2926_cse), or_tmp_2276, and_529_cse);
  assign mux_2149_nl = MUX_s_1_2_2((~ mux_2926_cse), (fsm_output[7]), and_529_cse);
  assign mux_2151_nl = MUX_s_1_2_2(mux_2150_nl, mux_2149_nl, fsm_output[0]);
  assign mux_2147_nl = MUX_s_1_2_2((fsm_output[7]), mux_2926_cse, fsm_output[2]);
  assign mux_2146_nl = MUX_s_1_2_2(and_395_cse, mux_2926_cse, fsm_output[2]);
  assign mux_2148_nl = MUX_s_1_2_2(mux_2147_nl, mux_2146_nl, and_526_cse);
  assign mux_2152_nl = MUX_s_1_2_2((~ mux_2151_nl), mux_2148_nl, fsm_output[9]);
  assign mux_2156_nl = MUX_s_1_2_2(mux_2155_nl, mux_2152_nl, fsm_output[6]);
  assign mux_2143_nl = MUX_s_1_2_2(or_tmp_2276, (fsm_output[7]), or_2368_cse);
  assign mux_2144_nl = MUX_s_1_2_2(mux_2143_nl, or_tmp_2276, fsm_output[9]);
  assign or_2339_nl = (fsm_output[6]) | mux_2144_nl;
  assign mux_2157_nl = MUX_s_1_2_2(mux_2156_nl, or_2339_nl, fsm_output[8]);
  assign mux_2140_nl = MUX_s_1_2_2((~ or_tmp_2281), or_tmp_2280, fsm_output[9]);
  assign or_2335_nl = (~ (fsm_output[9])) | (fsm_output[1]) | (fsm_output[2]);
  assign mux_2139_nl = MUX_s_1_2_2(or_tmp_2276, (fsm_output[7]), or_2335_nl);
  assign mux_2141_nl = MUX_s_1_2_2(mux_2140_nl, mux_2139_nl, fsm_output[6]);
  assign nand_197_nl = ~(nand_196_cse & and_395_cse);
  assign mux_2135_nl = MUX_s_1_2_2((~ and_395_cse), or_tmp_2276, and_529_cse);
  assign mux_2136_nl = MUX_s_1_2_2(nand_197_nl, mux_2135_nl, fsm_output[0]);
  assign mux_2137_nl = MUX_s_1_2_2(mux_2136_nl, or_tmp_2277, fsm_output[9]);
  assign mux_2133_nl = MUX_s_1_2_2((~ and_395_cse), or_tmp_2276, or_2377_cse);
  assign mux_2134_nl = MUX_s_1_2_2(mux_2133_nl, or_tmp_2274, fsm_output[9]);
  assign mux_2138_nl = MUX_s_1_2_2(mux_2137_nl, mux_2134_nl, fsm_output[6]);
  assign mux_2142_nl = MUX_s_1_2_2(mux_2141_nl, mux_2138_nl, fsm_output[8]);
  assign mux_2158_nl = MUX_s_1_2_2(mux_2157_nl, mux_2142_nl, fsm_output[5]);
  assign mux_2186_nl = MUX_s_1_2_2(mux_2185_nl, mux_2158_nl, fsm_output[4]);
  assign mux_2231_nl = MUX_s_1_2_2(mux_2230_nl, mux_2186_nl, fsm_output[3]);
  assign mux_2324_nl = MUX_s_1_2_2(or_3008_cse, or_259_cse, fsm_output[1]);
  assign mux_2325_nl = MUX_s_1_2_2(mux_2324_nl, mux_tmp_2311, fsm_output[0]);
  assign mux_2326_nl = MUX_s_1_2_2(mux_2325_nl, mux_tmp_130, fsm_output[3]);
  assign and_519_nl = or_3388_cse & (fsm_output[9]);
  assign mux_2322_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_93, and_519_nl);
  assign mux_2323_nl = MUX_s_1_2_2(mux_3555_cse, mux_2322_nl, fsm_output[3]);
  assign mux_2327_nl = MUX_s_1_2_2(mux_2326_nl, mux_2323_nl, fsm_output[6]);
  assign mux_2319_nl = MUX_s_1_2_2(or_tmp_2360, or_tmp_2341, fsm_output[0]);
  assign mux_2318_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_94, or_2421_cse);
  assign mux_2320_nl = MUX_s_1_2_2(mux_2319_nl, mux_2318_nl, fsm_output[3]);
  assign mux_2321_nl = MUX_s_1_2_2(mux_2320_nl, mux_tmp_2287, fsm_output[6]);
  assign mux_2328_nl = MUX_s_1_2_2(mux_2327_nl, mux_2321_nl, fsm_output[7]);
  assign mux_2314_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_94, or_2419_cse);
  assign mux_2315_nl = MUX_s_1_2_2(mux_2314_nl, (fsm_output[8]), fsm_output[3]);
  assign mux_2312_nl = MUX_s_1_2_2(mux_tmp_2311, mux_tmp_2293, fsm_output[0]);
  assign mux_2313_nl = MUX_s_1_2_2(mux_tmp_130, mux_2312_nl, fsm_output[3]);
  assign mux_2316_nl = MUX_s_1_2_2(mux_2315_nl, mux_2313_nl, fsm_output[6]);
  assign or_2418_nl = (~((fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]))) |
      (fsm_output[9]);
  assign mux_2309_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_94, or_2418_nl);
  assign mux_2307_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, fsm_output[1]);
  assign mux_2308_nl = MUX_s_1_2_2(mux_2307_nl, or_tmp_2341, fsm_output[3]);
  assign mux_2310_nl = MUX_s_1_2_2(mux_2309_nl, mux_2308_nl, fsm_output[6]);
  assign mux_2317_nl = MUX_s_1_2_2(mux_2316_nl, mux_2310_nl, fsm_output[7]);
  assign mux_2329_nl = MUX_s_1_2_2(mux_2328_nl, mux_2317_nl, fsm_output[5]);
  assign mux_2303_nl = MUX_s_1_2_2(mux_tmp_130, or_tmp_2360, fsm_output[3]);
  assign mux_2301_nl = MUX_s_1_2_2(or_2998_cse, or_2414_cse, or_3388_cse);
  assign mux_2300_nl = MUX_s_1_2_2(mux_1036_cse, mux_tmp_130, or_3388_cse);
  assign mux_2302_nl = MUX_s_1_2_2(mux_2301_nl, mux_2300_nl, fsm_output[3]);
  assign mux_2304_nl = MUX_s_1_2_2(mux_2303_nl, mux_2302_nl, fsm_output[6]);
  assign mux_2296_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_93, or_2419_cse);
  assign mux_2297_nl = MUX_s_1_2_2(mux_tmp_2289, mux_2296_nl, fsm_output[0]);
  assign mux_2298_nl = MUX_s_1_2_2((fsm_output[8]), mux_2297_nl, fsm_output[3]);
  assign or_2408_nl = nor_303_cse | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_2294_nl = MUX_s_1_2_2(mux_tmp_2293, or_2408_nl, fsm_output[0]);
  assign mux_2295_nl = MUX_s_1_2_2(mux_2294_nl, mux_tmp_130, fsm_output[3]);
  assign mux_2299_nl = MUX_s_1_2_2(mux_2298_nl, mux_2295_nl, fsm_output[6]);
  assign mux_2305_nl = MUX_s_1_2_2(mux_2304_nl, mux_2299_nl, fsm_output[7]);
  assign mux_2288_nl = MUX_s_1_2_2(or_2407_cse, mux_tmp_165, fsm_output[1]);
  assign mux_2290_nl = MUX_s_1_2_2(mux_tmp_2289, mux_2288_nl, fsm_output[3]);
  assign mux_2291_nl = MUX_s_1_2_2(mux_2290_nl, mux_tmp_2287, fsm_output[6]);
  assign or_2406_nl = and_526_cse | (fsm_output[10:8]!=3'b100);
  assign or_2404_nl = and_521_cse | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_2285_nl = MUX_s_1_2_2(or_2406_nl, or_2404_nl, fsm_output[3]);
  assign mux_2286_nl = MUX_s_1_2_2(mux_2285_nl, mux_tmp_139, fsm_output[6]);
  assign mux_2292_nl = MUX_s_1_2_2(mux_2291_nl, mux_2286_nl, fsm_output[7]);
  assign mux_2306_nl = MUX_s_1_2_2(mux_2305_nl, mux_2292_nl, fsm_output[5]);
  assign mux_2330_nl = MUX_s_1_2_2(mux_2329_nl, mux_2306_nl, fsm_output[4]);
  assign or_2403_nl = nor_297_cse | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_2280_nl = MUX_s_1_2_2(or_2403_nl, mux_tmp_130, fsm_output[3]);
  assign or_2402_nl = (fsm_output[1]) | (fsm_output[9]);
  assign mux_2278_nl = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), or_2402_nl);
  assign mux_2277_nl = MUX_s_1_2_2(mux_981_cse, or_2998_cse, and_526_cse);
  assign mux_2279_nl = MUX_s_1_2_2(mux_2278_nl, mux_2277_nl, fsm_output[3]);
  assign mux_2281_nl = MUX_s_1_2_2(mux_2280_nl, mux_2279_nl, fsm_output[6]);
  assign mux_2275_nl = MUX_s_1_2_2(or_tmp_2340, (fsm_output[8]), fsm_output[3]);
  assign mux_2276_nl = MUX_s_1_2_2(mux_2275_nl, mux_tmp_2241, fsm_output[6]);
  assign mux_2282_nl = MUX_s_1_2_2(mux_2281_nl, mux_2276_nl, fsm_output[7]);
  assign nor_295_nl = ~((fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]) | (~
      (fsm_output[9])));
  assign mux_2272_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_94, nor_295_nl);
  assign mux_2270_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_88, or_2400_cse);
  assign mux_2271_nl = MUX_s_1_2_2(mux_tmp_2262, mux_2270_nl, fsm_output[3]);
  assign mux_2273_nl = MUX_s_1_2_2(mux_2272_nl, mux_2271_nl, fsm_output[6]);
  assign mux_2267_nl = MUX_s_1_2_2(mux_tmp_141, or_3008_cse, or_3388_cse);
  assign or_2398_nl = nor_297_cse | (fsm_output[8]) | (fsm_output[10]);
  assign mux_2268_nl = MUX_s_1_2_2(mux_2267_nl, or_2398_nl, fsm_output[3]);
  assign mux_2269_nl = MUX_s_1_2_2(mux_tmp_2235, mux_2268_nl, fsm_output[6]);
  assign mux_2274_nl = MUX_s_1_2_2(mux_2273_nl, mux_2269_nl, fsm_output[7]);
  assign mux_2283_nl = MUX_s_1_2_2(mux_2282_nl, mux_2274_nl, fsm_output[5]);
  assign mux_2261_nl = MUX_s_1_2_2(or_tmp_2341, or_tmp_2340, fsm_output[0]);
  assign mux_2263_nl = MUX_s_1_2_2(mux_tmp_2262, mux_2261_nl, fsm_output[3]);
  assign or_2395_nl = (~((fsm_output[9:8]!=2'b10))) | (fsm_output[10]);
  assign mux_2259_nl = MUX_s_1_2_2(or_2395_nl, mux_1036_cse, and_526_cse);
  assign mux_2260_nl = MUX_s_1_2_2(mux_2259_nl, mux_tmp_130, fsm_output[3]);
  assign mux_2264_nl = MUX_s_1_2_2(mux_2263_nl, mux_2260_nl, fsm_output[6]);
  assign mux_2255_nl = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), or_2419_cse);
  assign mux_2251_nl = MUX_s_1_2_2(or_tmp_94, (fsm_output[8]), fsm_output[9]);
  assign mux_2253_nl = MUX_s_1_2_2(mux_981_cse, mux_2251_nl, fsm_output[1]);
  assign mux_2250_nl = MUX_s_1_2_2(or_tmp_94, or_tmp_93, nor_303_cse);
  assign mux_2254_nl = MUX_s_1_2_2(mux_2253_nl, mux_2250_nl, fsm_output[0]);
  assign mux_2256_nl = MUX_s_1_2_2(mux_2255_nl, mux_2254_nl, fsm_output[3]);
  assign or_2392_nl = (~((fsm_output[3]) | (fsm_output[1]))) | (fsm_output[9]);
  assign mux_2249_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_88, or_2392_nl);
  assign mux_2257_nl = MUX_s_1_2_2(mux_2256_nl, mux_2249_nl, fsm_output[6]);
  assign mux_2265_nl = MUX_s_1_2_2(mux_2264_nl, mux_2257_nl, fsm_output[7]);
  assign or_2390_nl = (~((~ (fsm_output[1])) | (fsm_output[9]))) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign or_2385_nl = (fsm_output[9:8]!=2'b10);
  assign mux_2244_nl = MUX_s_1_2_2(or_2387_cse, or_2385_nl, fsm_output[1]);
  assign mux_2245_nl = MUX_s_1_2_2(or_2390_nl, mux_2244_nl, fsm_output[0]);
  assign mux_2243_nl = MUX_s_1_2_2(mux_tmp_165, mux_3555_cse, or_3388_cse);
  assign mux_2246_nl = MUX_s_1_2_2(mux_2245_nl, mux_2243_nl, fsm_output[3]);
  assign mux_2247_nl = MUX_s_1_2_2(mux_2246_nl, mux_tmp_2241, fsm_output[6]);
  assign mux_2236_nl = MUX_s_1_2_2((fsm_output[8]), (~ or_tmp_88), or_2419_cse);
  assign nand_51_nl = ~((fsm_output[3]) & mux_2236_nl);
  assign mux_2237_nl = MUX_s_1_2_2(nand_51_nl, mux_tmp_2235, fsm_output[6]);
  assign mux_2248_nl = MUX_s_1_2_2(mux_2247_nl, mux_2237_nl, fsm_output[7]);
  assign mux_2266_nl = MUX_s_1_2_2(mux_2265_nl, mux_2248_nl, fsm_output[5]);
  assign mux_2284_nl = MUX_s_1_2_2(mux_2283_nl, mux_2266_nl, fsm_output[4]);
  assign mux_2331_nl = MUX_s_1_2_2(mux_2330_nl, mux_2284_nl, fsm_output[2]);
  assign and_517_nl = (fsm_output[4]) & mux_125_cse;
  assign nor_752_nl = ~((fsm_output[4]) | (fsm_output[7]) | mux_tmp_119);
  assign mux_2343_nl = MUX_s_1_2_2(and_517_nl, nor_752_nl, fsm_output[1]);
  assign nand_189_nl = ~((fsm_output[5]) & mux_2343_nl);
  assign or_3386_nl = (fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[7]) | (~
      (fsm_output[3])) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign nand_190_nl = ~((fsm_output[1]) & (fsm_output[4]) & (fsm_output[7]) & (fsm_output[3])
      & (fsm_output[8]) & (fsm_output[6]) & (fsm_output[10]));
  assign mux_2341_nl = MUX_s_1_2_2(or_3386_nl, nand_190_nl, fsm_output[5]);
  assign mux_2344_nl = MUX_s_1_2_2(nand_189_nl, mux_2341_nl, fsm_output[2]);
  assign or_2437_nl = (~ (fsm_output[4])) | (~ (fsm_output[7])) | (fsm_output[3])
      | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2340_nl = MUX_s_1_2_2(or_2437_nl, or_tmp_2376, fsm_output[1]);
  assign or_2438_nl = (~ (fsm_output[2])) | (fsm_output[5]) | mux_2340_nl;
  assign mux_2345_nl = MUX_s_1_2_2(mux_2344_nl, or_2438_nl, fsm_output[9]);
  assign or_2435_nl = (~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[8])
      | not_tmp_49;
  assign or_2433_nl = (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[8]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2335_nl = MUX_s_1_2_2(or_2435_nl, or_2433_nl, fsm_output[4]);
  assign mux_2336_nl = MUX_s_1_2_2(mux_2335_nl, or_tmp_2376, fsm_output[1]);
  assign or_2431_nl = (~ (fsm_output[1])) | (~ (fsm_output[4])) | (fsm_output[7])
      | (fsm_output[3]) | (fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_2337_nl = MUX_s_1_2_2(mux_2336_nl, or_2431_nl, fsm_output[5]);
  assign or_2430_nl = (fsm_output[5]) | (~ (fsm_output[1])) | (~ (fsm_output[4]))
      | (~ (fsm_output[7])) | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6])
      | (~ (fsm_output[10]));
  assign mux_2338_nl = MUX_s_1_2_2(mux_2337_nl, or_2430_nl, fsm_output[2]);
  assign nand_191_nl = ~((fsm_output[5]) & (fsm_output[1]) & (fsm_output[4]) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]) & (~ (fsm_output[10])));
  assign or_2427_nl = (~ (fsm_output[1])) | (~ (fsm_output[4])) | (fsm_output[7])
      | (~ (fsm_output[3])) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_2426_nl = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[7]) | mux_tmp_119;
  assign mux_2333_nl = MUX_s_1_2_2(or_2427_nl, or_2426_nl, fsm_output[5]);
  assign mux_2334_nl = MUX_s_1_2_2(nand_191_nl, mux_2333_nl, fsm_output[2]);
  assign mux_2339_nl = MUX_s_1_2_2(mux_2338_nl, mux_2334_nl, fsm_output[9]);
  assign mux_2346_nl = MUX_s_1_2_2(mux_2345_nl, mux_2339_nl, fsm_output[0]);
  assign mux_2414_nl = MUX_s_1_2_2(mux_tmp_2389, or_tmp_2396, fsm_output[7]);
  assign mux_2413_nl = MUX_s_1_2_2(mux_tmp_2386, mux_tmp_2353, fsm_output[7]);
  assign mux_2415_nl = MUX_s_1_2_2(mux_2414_nl, mux_2413_nl, fsm_output[2]);
  assign mux_2411_nl = MUX_s_1_2_2(mux_tmp_2378, mux_tmp_2382, fsm_output[7]);
  assign mux_2410_nl = MUX_s_1_2_2(mux_tmp_2376, nand_tmp_54, fsm_output[7]);
  assign mux_2412_nl = MUX_s_1_2_2(mux_2411_nl, mux_2410_nl, fsm_output[2]);
  assign mux_2416_nl = MUX_s_1_2_2(mux_2415_nl, mux_2412_nl, fsm_output[3]);
  assign mux_2405_nl = MUX_s_1_2_2(mux_tmp_2347, mux_tmp_2369, fsm_output[6]);
  assign mux_2406_nl = MUX_s_1_2_2(mux_tmp_2371, mux_2405_nl, fsm_output[0]);
  assign mux_2407_nl = MUX_s_1_2_2(mux_2406_nl, nand_tmp_54, fsm_output[7]);
  assign mux_2403_nl = MUX_s_1_2_2(mux_tmp_2365, mux_tmp_2361, fsm_output[0]);
  assign mux_2401_nl = MUX_s_1_2_2(or_tmp_2390, mux_tmp_2363, fsm_output[6]);
  assign mux_2402_nl = MUX_s_1_2_2(mux_tmp_2364, mux_2401_nl, fsm_output[0]);
  assign mux_2404_nl = MUX_s_1_2_2(mux_2403_nl, mux_2402_nl, fsm_output[7]);
  assign mux_2408_nl = MUX_s_1_2_2(mux_2407_nl, mux_2404_nl, fsm_output[2]);
  assign mux_2397_nl = MUX_s_1_2_2(mux_tmp_2348, mux_tmp_2359, fsm_output[6]);
  assign mux_2398_nl = MUX_s_1_2_2(mux_2397_nl, mux_tmp_2356, fsm_output[0]);
  assign mux_2399_nl = MUX_s_1_2_2(or_tmp_2396, mux_2398_nl, fsm_output[7]);
  assign mux_2395_nl = MUX_s_1_2_2(or_tmp_2396, mux_tmp_2353, fsm_output[0]);
  assign mux_2396_nl = MUX_s_1_2_2(mux_2395_nl, mux_tmp_2350, fsm_output[7]);
  assign mux_2400_nl = MUX_s_1_2_2(mux_2399_nl, mux_2396_nl, fsm_output[2]);
  assign mux_2409_nl = MUX_s_1_2_2(mux_2408_nl, mux_2400_nl, fsm_output[3]);
  assign mux_2417_nl = MUX_s_1_2_2(mux_2416_nl, mux_2409_nl, fsm_output[4]);
  assign mux_2390_nl = MUX_s_1_2_2(mux_tmp_2389, mux_tmp_2386, fsm_output[0]);
  assign mux_2391_nl = MUX_s_1_2_2(mux_2390_nl, or_tmp_2396, fsm_output[7]);
  assign mux_2383_nl = MUX_s_1_2_2(mux_tmp_2353, mux_tmp_2382, fsm_output[0]);
  assign mux_2384_nl = MUX_s_1_2_2(mux_tmp_2378, mux_2383_nl, fsm_output[7]);
  assign mux_2392_nl = MUX_s_1_2_2(mux_2391_nl, mux_2384_nl, fsm_output[2]);
  assign mux_2379_nl = MUX_s_1_2_2(mux_tmp_2378, mux_tmp_2376, fsm_output[0]);
  assign mux_2380_nl = MUX_s_1_2_2(mux_2379_nl, nand_tmp_54, fsm_output[7]);
  assign mux_2372_nl = MUX_s_1_2_2(mux_tmp_2370, or_tmp_2405, fsm_output[6]);
  assign mux_2373_nl = MUX_s_1_2_2(mux_2372_nl, mux_tmp_2371, fsm_output[0]);
  assign mux_2374_nl = MUX_s_1_2_2(mux_2373_nl, nand_tmp_54, fsm_output[7]);
  assign mux_2381_nl = MUX_s_1_2_2(mux_2380_nl, mux_2374_nl, fsm_output[2]);
  assign mux_2393_nl = MUX_s_1_2_2(mux_2392_nl, mux_2381_nl, fsm_output[3]);
  assign mux_2366_nl = MUX_s_1_2_2(mux_tmp_2365, mux_tmp_2364, fsm_output[7]);
  assign mux_2360_nl = MUX_s_1_2_2(or_tmp_2390, mux_tmp_2359, fsm_output[6]);
  assign mux_2362_nl = MUX_s_1_2_2(mux_tmp_2361, mux_2360_nl, fsm_output[7]);
  assign mux_2367_nl = MUX_s_1_2_2(mux_2366_nl, mux_2362_nl, fsm_output[2]);
  assign mux_2357_nl = MUX_s_1_2_2(or_tmp_2396, mux_tmp_2356, fsm_output[7]);
  assign mux_2349_nl = MUX_s_1_2_2(mux_tmp_2348, mux_tmp_2347, fsm_output[6]);
  assign mux_2351_nl = MUX_s_1_2_2(mux_tmp_2350, mux_2349_nl, fsm_output[0]);
  assign mux_2354_nl = MUX_s_1_2_2(mux_tmp_2353, mux_2351_nl, fsm_output[7]);
  assign mux_2358_nl = MUX_s_1_2_2(mux_2357_nl, mux_2354_nl, fsm_output[2]);
  assign mux_2368_nl = MUX_s_1_2_2(mux_2367_nl, mux_2358_nl, fsm_output[3]);
  assign mux_2394_nl = MUX_s_1_2_2(mux_2393_nl, mux_2368_nl, fsm_output[4]);
  assign mux_2418_nl = MUX_s_1_2_2(mux_2417_nl, mux_2394_nl, fsm_output[1]);
  assign COMP_LOOP_nor_11_nl = ~((z_out_2_12_1[3:1]!=3'b000));
  assign COMP_LOOP_and_274_nl = (~ and_dcpl_256) & and_dcpl_247;
  assign or_2881_nl = nor_653_cse | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_3065_nl = MUX_s_1_2_2(or_2881_nl, mux_tmp_3049, fsm_output[1]);
  assign mux_3066_nl = MUX_s_1_2_2(mux_3065_nl, mux_1036_cse, fsm_output[4]);
  assign mux_3063_nl = MUX_s_1_2_2(mux_tmp_3024, or_tmp_2802, or_3388_cse);
  assign mux_3064_nl = MUX_s_1_2_2(mux_tmp_130, mux_3063_nl, fsm_output[4]);
  assign mux_3067_nl = MUX_s_1_2_2(mux_3066_nl, mux_3064_nl, fsm_output[7]);
  assign mux_3060_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_3032, and_526_cse);
  assign or_449_nl = (~ (fsm_output[2])) | (fsm_output[9]) | (fsm_output[8]) | (fsm_output[10]);
  assign or_2876_nl = nor_653_cse | (fsm_output[8]) | (fsm_output[10]);
  assign mux_3059_nl = MUX_s_1_2_2(or_449_nl, or_2876_nl, fsm_output[1]);
  assign mux_3061_nl = MUX_s_1_2_2(mux_3060_nl, mux_3059_nl, fsm_output[4]);
  assign mux_3062_nl = MUX_s_1_2_2(mux_3061_nl, mux_tmp_139, fsm_output[7]);
  assign mux_3068_nl = MUX_s_1_2_2(mux_3067_nl, mux_3062_nl, fsm_output[5]);
  assign nor_407_nl = ~((fsm_output[4]) | (~ (fsm_output[1])) | (fsm_output[0]) |
      (fsm_output[9]) | (~ (fsm_output[2])));
  assign mux_3056_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_93, nor_407_nl);
  assign mux_3053_nl = MUX_s_1_2_2(or_tmp_93, or_tmp_2814, fsm_output[9]);
  assign mux_3051_nl = MUX_s_1_2_2(or_tmp_2795, or_tmp_2814, fsm_output[9]);
  assign or_439_nl = (fsm_output[2]) | (fsm_output[9]) | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_3052_nl = MUX_s_1_2_2(mux_3051_nl, or_439_nl, fsm_output[0]);
  assign mux_3054_nl = MUX_s_1_2_2(mux_3053_nl, mux_3052_nl, fsm_output[1]);
  assign mux_3050_nl = MUX_s_1_2_2(mux_tmp_3049, mux_tmp_3007, fsm_output[1]);
  assign mux_3055_nl = MUX_s_1_2_2(mux_3054_nl, mux_3050_nl, fsm_output[4]);
  assign mux_3057_nl = MUX_s_1_2_2(mux_3056_nl, mux_3055_nl, fsm_output[7]);
  assign or_2870_nl = (fsm_output[1]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[8])
      | (~ (fsm_output[10]));
  assign mux_3047_nl = MUX_s_1_2_2(or_2870_nl, mux_tmp_130, fsm_output[4]);
  assign mux_3045_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_3032, or_3388_cse);
  assign mux_3046_nl = MUX_s_1_2_2(mux_tmp_130, mux_3045_nl, fsm_output[4]);
  assign mux_3048_nl = MUX_s_1_2_2(mux_3047_nl, mux_3046_nl, fsm_output[7]);
  assign mux_3058_nl = MUX_s_1_2_2(mux_3057_nl, mux_3048_nl, fsm_output[5]);
  assign mux_3069_nl = MUX_s_1_2_2(mux_3068_nl, mux_3058_nl, fsm_output[6]);
  assign mux_3039_nl = MUX_s_1_2_2((~ mux_tmp_3014), or_tmp_88, fsm_output[9]);
  assign mux_3040_nl = MUX_s_1_2_2(mux_3039_nl, mux_1036_cse, fsm_output[1]);
  assign mux_3035_nl = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), fsm_output[2]);
  assign mux_3036_nl = MUX_s_1_2_2((~ mux_3035_nl), or_tmp_88, fsm_output[9]);
  assign mux_3038_nl = MUX_s_1_2_2(mux_1036_cse, mux_3036_nl, or_3388_cse);
  assign mux_3041_nl = MUX_s_1_2_2(mux_3040_nl, mux_3038_nl, fsm_output[4]);
  assign mux_3033_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_3032, fsm_output[1]);
  assign or_2866_nl = (~((fsm_output[0]) | (~ (fsm_output[9])))) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (fsm_output[10]);
  assign or_2865_nl = nor_657_cse | (fsm_output[8]) | (fsm_output[10]);
  assign mux_3030_nl = MUX_s_1_2_2(or_2866_nl, or_2865_nl, fsm_output[1]);
  assign mux_3034_nl = MUX_s_1_2_2(mux_3033_nl, mux_3030_nl, fsm_output[4]);
  assign mux_3042_nl = MUX_s_1_2_2(mux_3041_nl, mux_3034_nl, fsm_output[7]);
  assign mux_3025_nl = MUX_s_1_2_2((~ nor_tmp_405), or_tmp_2803, fsm_output[9]);
  assign mux_3026_nl = MUX_s_1_2_2(mux_3025_nl, mux_tmp_3024, fsm_output[0]);
  assign mux_3027_nl = MUX_s_1_2_2(mux_3026_nl, or_tmp_2802, fsm_output[1]);
  assign or_2859_nl = (~(nor_753_cse | (fsm_output[9]))) | (fsm_output[2]);
  assign mux_3023_nl = MUX_s_1_2_2(or_tmp_94, (fsm_output[8]), or_2859_nl);
  assign mux_3028_nl = MUX_s_1_2_2(mux_3027_nl, mux_3023_nl, fsm_output[4]);
  assign mux_3029_nl = MUX_s_1_2_2(mux_3028_nl, mux_tmp_139, fsm_output[7]);
  assign mux_3043_nl = MUX_s_1_2_2(mux_3042_nl, mux_3029_nl, fsm_output[5]);
  assign mux_3016_nl = MUX_s_1_2_2((fsm_output[8]), or_tmp_93, or_2855_cse);
  assign mux_3015_nl = MUX_s_1_2_2(or_tmp_2795, mux_tmp_3014, fsm_output[9]);
  assign mux_3017_nl = MUX_s_1_2_2(mux_3016_nl, mux_3015_nl, fsm_output[0]);
  assign mux_3018_nl = MUX_s_1_2_2(mux_tmp_3014, mux_3017_nl, fsm_output[1]);
  assign mux_3019_nl = MUX_s_1_2_2((fsm_output[8]), mux_3018_nl, fsm_output[4]);
  assign or_2851_nl = (~ (fsm_output[1])) | (~ (fsm_output[0])) | (fsm_output[9])
      | (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_3013_nl = MUX_s_1_2_2(or_2851_nl, mux_tmp_130, fsm_output[4]);
  assign mux_3020_nl = MUX_s_1_2_2(mux_3019_nl, mux_3013_nl, fsm_output[7]);
  assign mux_3009_nl = MUX_s_1_2_2(mux_tmp_3008, mux_tmp_3007, fsm_output[0]);
  assign mux_3010_nl = MUX_s_1_2_2(or_tmp_2791, mux_3009_nl, fsm_output[1]);
  assign mux_3011_nl = MUX_s_1_2_2(mux_3010_nl, mux_tmp_130, fsm_output[4]);
  assign or_2846_nl = and_526_cse | (fsm_output[9]) | (fsm_output[2]) | (~ nor_tmp_405);
  assign mux_3005_nl = MUX_s_1_2_2(mux_tmp_130, or_2846_nl, fsm_output[4]);
  assign mux_3012_nl = MUX_s_1_2_2(mux_3011_nl, mux_3005_nl, fsm_output[7]);
  assign mux_3021_nl = MUX_s_1_2_2(mux_3020_nl, mux_3012_nl, fsm_output[5]);
  assign mux_3044_nl = MUX_s_1_2_2(mux_3043_nl, mux_3021_nl, fsm_output[6]);
  assign mux_3070_nl = MUX_s_1_2_2(mux_3069_nl, mux_3044_nl, fsm_output[3]);
  assign COMP_LOOP_mux1h_428_nl = MUX1HOT_s_1_6_2((operator_66_true_div_cmp_z[0]),
      (tmp_10_lpi_4_dfm[0]), (z_out[5]), COMP_LOOP_nor_12_itm, COMP_LOOP_nor_11_itm,
      COMP_LOOP_nor_11_nl, {COMP_LOOP_and_274_nl , and_dcpl_256 , and_dcpl_109 ,
      not_tmp_557 , (~ mux_3070_nl) , COMP_LOOP_or_32_cse});
  assign or_2821_nl = (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[4]) | (fsm_output[1])
      | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[10]);
  assign nor_671_nl = ~((fsm_output[6]) | nand_159_cse);
  assign nor_672_nl = ~((fsm_output[6]) | (fsm_output[3]) | (fsm_output[10]));
  assign mux_2986_nl = MUX_s_1_2_2(nor_671_nl, nor_672_nl, fsm_output[1]);
  assign nand_74_nl = ~((~((fsm_output[8]) | (~ (fsm_output[4])))) & mux_2986_nl);
  assign or_2818_nl = (~ (fsm_output[8])) | (fsm_output[4]) | (~ (fsm_output[1]))
      | (~ (fsm_output[6])) | (~ (fsm_output[3])) | (fsm_output[10]);
  assign mux_2987_nl = MUX_s_1_2_2(nand_74_nl, or_2818_nl, fsm_output[9]);
  assign mux_2988_nl = MUX_s_1_2_2(or_2821_nl, mux_2987_nl, fsm_output[5]);
  assign or_3440_nl = (fsm_output[7]) | mux_2988_nl;
  assign or_3441_nl = (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[8])) | (fsm_output[4])
      | (~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[3]) | (~ (fsm_output[10]));
  assign and_447_nl = (fsm_output[1]) & (fsm_output[6]) & (fsm_output[3]) & (~ (fsm_output[10]));
  assign nor_675_nl = ~((fsm_output[1]) | (~ (fsm_output[6])) | (fsm_output[3]) |
      (~ (fsm_output[10])));
  assign mux_2983_nl = MUX_s_1_2_2(and_447_nl, nor_675_nl, fsm_output[4]);
  assign nand_73_nl = ~((fsm_output[8]) & mux_2983_nl);
  assign or_2811_nl = (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[1]) | (fsm_output[6])
      | (~ (fsm_output[3])) | (fsm_output[10]);
  assign mux_2984_nl = MUX_s_1_2_2(nand_73_nl, or_2811_nl, fsm_output[9]);
  assign or_3442_nl = (fsm_output[5]) | mux_2984_nl;
  assign mux_2985_nl = MUX_s_1_2_2(or_3441_nl, or_3442_nl, fsm_output[7]);
  assign mux_2989_nl = MUX_s_1_2_2(or_3440_nl, mux_2985_nl, fsm_output[2]);
  assign nor_647_nl = ~((fsm_output[1]) | (~ (fsm_output[4])) | (~ (fsm_output[3]))
      | (fsm_output[10]));
  assign mux_3075_nl = MUX_s_1_2_2(nor_647_nl, nor_tmp_410, fsm_output[2]);
  assign nor_646_nl = ~((fsm_output[7:5]!=3'b100) | (~ mux_3075_nl));
  assign nor_648_nl = ~((fsm_output[4]) | nand_159_cse);
  assign nor_649_nl = ~((fsm_output[4]) | (fsm_output[3]) | (fsm_output[10]));
  assign mux_3074_nl = MUX_s_1_2_2(nor_648_nl, nor_649_nl, fsm_output[1]);
  assign and_439_nl = (~ (fsm_output[7])) & (fsm_output[6]) & (fsm_output[5]) & (fsm_output[2])
      & mux_3074_nl;
  assign mux_3076_nl = MUX_s_1_2_2(nor_646_nl, and_439_nl, fsm_output[8]);
  assign nor_650_nl = ~((fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[3]) |
      (fsm_output[10]));
  assign mux_3072_nl = MUX_s_1_2_2(nor_tmp_410, nor_650_nl, fsm_output[2]);
  assign and_440_nl = (~((fsm_output[7:5]!=3'b001))) & mux_3072_nl;
  assign nor_651_nl = ~((fsm_output[6]) | (fsm_output[5]) | (fsm_output[2]) | (~
      (fsm_output[1])) | (fsm_output[4]) | (fsm_output[3]) | (fsm_output[10]));
  assign nor_652_nl = ~((~ (fsm_output[6])) | (fsm_output[5]) | (fsm_output[2]) |
      (fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[3]) | (fsm_output[10]));
  assign mux_3071_nl = MUX_s_1_2_2(nor_651_nl, nor_652_nl, fsm_output[7]);
  assign mux_3073_nl = MUX_s_1_2_2(and_440_nl, mux_3071_nl, fsm_output[8]);
  assign mux_3077_nl = MUX_s_1_2_2(mux_3076_nl, mux_3073_nl, fsm_output[9]);
  assign COMP_LOOP_mux1h_464_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0[3]), COMP_LOOP_nor_134_itm,
      modExp_exp_1_7_1_sva, (COMP_LOOP_k_9_4_sva_4_0[4]), {and_dcpl_257 , and_dcpl_304
      , (~ mux_3494_itm) , not_tmp_688});
  assign or_3501_nl = (~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[9]) | (~
      (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign or_3502_nl = (fsm_output[5]) | (~ (fsm_output[9])) | (~ (fsm_output[2]))
      | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign or_3503_nl = (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_3517_nl = MUX_s_1_2_2(or_3502_nl, or_3503_nl, fsm_output[7]);
  assign mux_3518_nl = MUX_s_1_2_2(or_3501_nl, mux_3517_nl, fsm_output[3]);
  assign mux_3519_nl = MUX_s_1_2_2(or_80_cse, mux_3518_nl, fsm_output[4]);
  assign or_3133_nl = (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[8]) | not_tmp_49;
  assign mux_3515_nl = MUX_s_1_2_2(or_3133_nl, or_tmp_3053, fsm_output[7]);
  assign or_3131_nl = (~ (fsm_output[5])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign or_3130_nl = (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[2])) | (~
      (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_3514_nl = MUX_s_1_2_2(or_3131_nl, or_3130_nl, fsm_output[7]);
  assign mux_3516_nl = MUX_s_1_2_2(mux_3515_nl, mux_3514_nl, fsm_output[3]);
  assign or_3504_nl = (fsm_output[4]) | mux_3516_nl;
  assign mux_3520_nl = MUX_s_1_2_2(mux_3519_nl, or_3504_nl, fsm_output[1]);
  assign or_3505_nl = (~ (fsm_output[3])) | (fsm_output[7]) | (~ (fsm_output[5]))
      | (fsm_output[9]) | (~ (fsm_output[2])) | (~ (fsm_output[8])) | (fsm_output[6])
      | (~ (fsm_output[10]));
  assign nor_600_nl = ~((~ (fsm_output[9])) | (fsm_output[2]) | (~ (fsm_output[8]))
      | (fsm_output[6]) | (fsm_output[10]));
  assign nor_601_nl = ~((fsm_output[9]) | (~ (fsm_output[2])) | (~ (fsm_output[8]))
      | (~ (fsm_output[6])) | (fsm_output[10]));
  assign mux_3511_nl = MUX_s_1_2_2(nor_600_nl, nor_601_nl, fsm_output[5]);
  assign nand_412_nl = ~((~((fsm_output[3]) | (~ (fsm_output[7])))) & mux_3511_nl);
  assign mux_3512_nl = MUX_s_1_2_2(or_3505_nl, nand_412_nl, fsm_output[4]);
  assign or_3124_nl = (~ (fsm_output[5])) | (fsm_output[9]) | (~ (fsm_output[2]))
      | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign or_3123_nl = (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[2]) | (fsm_output[8])
      | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_3509_nl = MUX_s_1_2_2(or_3124_nl, or_3123_nl, fsm_output[7]);
  assign or_3506_nl = (fsm_output[3]) | mux_3509_nl;
  assign or_3120_nl = (~ (fsm_output[5])) | (fsm_output[9]) | (fsm_output[2]) | nand_142_cse;
  assign mux_3508_nl = MUX_s_1_2_2(or_tmp_3053, or_3120_nl, fsm_output[7]);
  assign nand_413_nl = ~((fsm_output[3]) & (~ mux_3508_nl));
  assign mux_3510_nl = MUX_s_1_2_2(or_3506_nl, nand_413_nl, fsm_output[4]);
  assign mux_3513_nl = MUX_s_1_2_2(mux_3512_nl, mux_3510_nl, fsm_output[1]);
  assign mux_3521_nl = MUX_s_1_2_2(mux_3520_nl, mux_3513_nl, fsm_output[0]);
  assign COMP_LOOP_nor_12_nl = ~((z_out_2_12_1[3]) | (z_out_2_12_1[2]) | (z_out_2_12_1[0]));
  assign mux_3610_nl = MUX_s_1_2_2(nand_tmp_4, mux_155_cse, fsm_output[2]);
  assign mux_3611_nl = MUX_s_1_2_2(mux_3610_nl, mux_tmp_3551, fsm_output[0]);
  assign mux_3609_nl = MUX_s_1_2_2(mux_tmp_3551, mux_tmp_3547, fsm_output[0]);
  assign mux_3612_nl = MUX_s_1_2_2(mux_3611_nl, mux_3609_nl, fsm_output[1]);
  assign mux_3606_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, fsm_output[4]);
  assign mux_3607_nl = MUX_s_1_2_2(mux_3606_nl, or_tmp_96, fsm_output[2]);
  assign mux_3605_nl = MUX_s_1_2_2(mux_161_cse, or_tmp_96, fsm_output[2]);
  assign mux_3608_nl = MUX_s_1_2_2(mux_3607_nl, mux_3605_nl, or_3388_cse);
  assign mux_3613_nl = MUX_s_1_2_2(mux_3612_nl, mux_3608_nl, fsm_output[7]);
  assign mux_3602_nl = MUX_s_1_2_2(mux_tmp_3576, mux_tmp_3574, fsm_output[0]);
  assign mux_3603_nl = MUX_s_1_2_2(mux_tmp_3577, mux_3602_nl, fsm_output[1]);
  assign mux_3604_nl = MUX_s_1_2_2(mux_3603_nl, mux_tmp_139, fsm_output[7]);
  assign mux_3614_nl = MUX_s_1_2_2(mux_3613_nl, mux_3604_nl, fsm_output[5]);
  assign or_3192_nl = (~(and_529_cse | (fsm_output[4]))) | (fsm_output[9]);
  assign mux_3599_nl = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), or_3192_nl);
  assign mux_3596_nl = MUX_s_1_2_2(mux_498_cse, mux_171_cse, fsm_output[2]);
  assign mux_493_nl = MUX_s_1_2_2(or_469_cse, mux_tmp_130, fsm_output[4]);
  assign mux_3595_nl = MUX_s_1_2_2(mux_498_cse, mux_493_nl, fsm_output[2]);
  assign mux_3597_nl = MUX_s_1_2_2(mux_3596_nl, mux_3595_nl, fsm_output[0]);
  assign mux_454_nl = MUX_s_1_2_2(mux_tmp_165, or_tmp_88, fsm_output[4]);
  assign mux_3591_nl = MUX_s_1_2_2(mux_454_nl, nand_tmp_4, fsm_output[2]);
  assign mux_3588_nl = MUX_s_1_2_2(mux_171_cse, nand_tmp_4, fsm_output[2]);
  assign mux_3592_nl = MUX_s_1_2_2(mux_3591_nl, mux_3588_nl, fsm_output[0]);
  assign mux_3598_nl = MUX_s_1_2_2(mux_3597_nl, mux_3592_nl, fsm_output[1]);
  assign mux_3600_nl = MUX_s_1_2_2(mux_3599_nl, mux_3598_nl, fsm_output[7]);
  assign mux_3584_nl = MUX_s_1_2_2(or_2387_cse, mux_tmp_130, fsm_output[4]);
  assign mux_3585_nl = MUX_s_1_2_2(mux_3584_nl, nand_tmp_4, or_2368_cse);
  assign and_364_nl = or_3388_cse & (fsm_output[2]) & (fsm_output[4]);
  assign mux_3583_nl = MUX_s_1_2_2(mux_tmp_130, mux_tmp_141, and_364_nl);
  assign mux_3586_nl = MUX_s_1_2_2(mux_3585_nl, mux_3583_nl, fsm_output[7]);
  assign mux_3601_nl = MUX_s_1_2_2(mux_3600_nl, mux_3586_nl, fsm_output[5]);
  assign mux_3615_nl = MUX_s_1_2_2(mux_3614_nl, mux_3601_nl, fsm_output[6]);
  assign mux_3578_nl = MUX_s_1_2_2(mux_tmp_3577, mux_tmp_3576, fsm_output[0]);
  assign mux_3579_nl = MUX_s_1_2_2(mux_3578_nl, mux_tmp_3574, fsm_output[1]);
  assign mux_3580_nl = MUX_s_1_2_2(mux_tmp_130, mux_3579_nl, fsm_output[7]);
  assign mux_481_nl = MUX_s_1_2_2(or_3008_cse, (fsm_output[8]), fsm_output[4]);
  assign mux_3569_nl = MUX_s_1_2_2(mux_340_cse, mux_481_nl, fsm_output[2]);
  assign mux_3565_nl = MUX_s_1_2_2(mux_tmp_141, mux_tmp_139, fsm_output[4]);
  assign mux_3566_nl = MUX_s_1_2_2(mux_3565_nl, or_163_cse, fsm_output[2]);
  assign mux_3570_nl = MUX_s_1_2_2(mux_3569_nl, mux_3566_nl, fsm_output[0]);
  assign mux_3562_nl = MUX_s_1_2_2(or_3008_cse, mux_tmp_139, fsm_output[4]);
  assign mux_3563_nl = MUX_s_1_2_2(mux_3562_nl, or_163_cse, fsm_output[2]);
  assign mux_3571_nl = MUX_s_1_2_2(mux_3570_nl, mux_3563_nl, fsm_output[1]);
  assign mux_3572_nl = MUX_s_1_2_2(mux_3571_nl, mux_tmp_139, fsm_output[7]);
  assign mux_3581_nl = MUX_s_1_2_2(mux_3580_nl, mux_3572_nl, fsm_output[5]);
  assign and_365_nl = (~((fsm_output[2]) & (fsm_output[4]))) & (fsm_output[9]);
  assign mux_3557_nl = MUX_s_1_2_2(or_tmp_93, (fsm_output[8]), and_365_nl);
  assign mux_3556_nl = MUX_s_1_2_2(mux_3555_cse, or_2387_cse, and_366_cse);
  assign mux_3558_nl = MUX_s_1_2_2(mux_3557_nl, mux_3556_nl, and_526_cse);
  assign mux_3554_nl = MUX_s_1_2_2(nand_tmp_4, mux_tmp_131, and_536_cse);
  assign mux_3559_nl = MUX_s_1_2_2(mux_3558_nl, mux_3554_nl, fsm_output[7]);
  assign or_3177_nl = (~((fsm_output[2]) | (fsm_output[4]))) | (fsm_output[9]);
  assign mux_3546_nl = MUX_s_1_2_2((~ (fsm_output[8])), or_tmp_88, or_3177_nl);
  assign mux_3548_nl = MUX_s_1_2_2(mux_tmp_3547, mux_3546_nl, fsm_output[0]);
  assign mux_3552_nl = MUX_s_1_2_2(mux_tmp_3551, mux_3548_nl, fsm_output[1]);
  assign mux_3545_nl = MUX_s_1_2_2(mux_161_cse, or_tmp_96, or_2377_cse);
  assign mux_3553_nl = MUX_s_1_2_2(mux_3552_nl, mux_3545_nl, fsm_output[7]);
  assign mux_3560_nl = MUX_s_1_2_2(mux_3559_nl, mux_3553_nl, fsm_output[5]);
  assign mux_3582_nl = MUX_s_1_2_2(mux_3581_nl, mux_3560_nl, fsm_output[6]);
  assign mux_3616_nl = MUX_s_1_2_2(mux_3615_nl, mux_3582_nl, fsm_output[3]);
  assign mux_3627_nl = MUX_s_1_2_2(mux_tmp_3618, or_tmp_3135, fsm_output[3]);
  assign nor_565_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | mux_3627_nl);
  assign or_3213_nl = (fsm_output[2]) | (~ (fsm_output[1])) | (fsm_output[8]) | not_tmp_49;
  assign or_3211_nl = (fsm_output[2]) | (~ (fsm_output[1])) | (~ (fsm_output[8]))
      | (fsm_output[6]) | (fsm_output[10]);
  assign mux_3626_nl = MUX_s_1_2_2(or_3213_nl, or_3211_nl, fsm_output[3]);
  assign nor_566_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | mux_3626_nl);
  assign mux_3628_nl = MUX_s_1_2_2(nor_565_nl, nor_566_nl, fsm_output[9]);
  assign nor_567_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (~ (fsm_output[2])) | (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[6])
      | (~ (fsm_output[10])));
  assign nor_568_nl = ~((fsm_output[7]) | (~ (fsm_output[3])) | (~ (fsm_output[2]))
      | (fsm_output[1]) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign nor_569_nl = ~((~ (fsm_output[7])) | (~ (fsm_output[3])) | (fsm_output[2])
      | (fsm_output[1]) | (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[10]));
  assign mux_3624_nl = MUX_s_1_2_2(nor_568_nl, nor_569_nl, fsm_output[5]);
  assign mux_3625_nl = MUX_s_1_2_2(nor_567_nl, mux_3624_nl, fsm_output[9]);
  assign mux_3629_nl = MUX_s_1_2_2(mux_3628_nl, mux_3625_nl, fsm_output[4]);
  assign or_3203_nl = (~ (fsm_output[2])) | (fsm_output[1]) | (~ (fsm_output[8]))
      | (fsm_output[6]) | (~ (fsm_output[10]));
  assign mux_3621_nl = MUX_s_1_2_2(or_tmp_3135, or_3203_nl, fsm_output[3]);
  assign nor_570_nl = ~((~ (fsm_output[5])) | (fsm_output[7]) | mux_3621_nl);
  assign nor_571_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (fsm_output[2]) | (~ (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[6]))
      | (fsm_output[10]));
  assign mux_3622_nl = MUX_s_1_2_2(nor_570_nl, nor_571_nl, fsm_output[9]);
  assign nor_572_nl = ~((fsm_output[7]) | (~ (fsm_output[3])) | mux_tmp_3618);
  assign nor_573_nl = ~((~ (fsm_output[2])) | (fsm_output[1]) | (~ (fsm_output[8]))
      | (~ (fsm_output[6])) | (fsm_output[10]));
  assign nor_574_nl = ~((fsm_output[2]) | (~((fsm_output[1]) & (fsm_output[8]) &
      (fsm_output[6]) & (fsm_output[10]))));
  assign mux_3617_nl = MUX_s_1_2_2(nor_573_nl, nor_574_nl, fsm_output[3]);
  assign and_362_nl = (fsm_output[7]) & mux_3617_nl;
  assign mux_3619_nl = MUX_s_1_2_2(nor_572_nl, and_362_nl, fsm_output[5]);
  assign nor_575_nl = ~((fsm_output[5]) | (~ (fsm_output[7])) | (fsm_output[3]) |
      (fsm_output[2]) | (fsm_output[1]) | (~ (fsm_output[8])) | (fsm_output[6]) |
      (fsm_output[10]));
  assign mux_3620_nl = MUX_s_1_2_2(mux_3619_nl, nor_575_nl, fsm_output[9]);
  assign mux_3623_nl = MUX_s_1_2_2(mux_3622_nl, mux_3620_nl, fsm_output[4]);
  assign mux_3630_nl = MUX_s_1_2_2(mux_3629_nl, mux_3623_nl, fsm_output[0]);
  assign COMP_LOOP_mux1h_474_nl = MUX1HOT_s_1_3_2(COMP_LOOP_nor_12_itm, COMP_LOOP_nor_134_itm,
      COMP_LOOP_nor_12_nl, {(~ mux_3616_nl) , mux_3630_nl , COMP_LOOP_or_32_cse});
  assign or_3171_nl = (fsm_output[4]) | (~ (fsm_output[9])) | (~ (fsm_output[6]))
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_3540_nl = MUX_s_1_2_2(or_tmp_3095, or_3171_nl, fsm_output[3]);
  assign nor_578_nl = ~((fsm_output[7]) | (~ (fsm_output[5])) | mux_3540_nl);
  assign nor_579_nl = ~((fsm_output[5]) | (fsm_output[3]) | (fsm_output[4]) | (fsm_output[9])
      | (fsm_output[6]) | nand_138_cse);
  assign nor_580_nl = ~((fsm_output[5]) | (~ (fsm_output[3])) | (fsm_output[4]) |
      (fsm_output[9]) | (~ (fsm_output[6])) | (~ (fsm_output[8])) | (fsm_output[10]));
  assign mux_3539_nl = MUX_s_1_2_2(nor_579_nl, nor_580_nl, fsm_output[7]);
  assign mux_3541_nl = MUX_s_1_2_2(nor_578_nl, mux_3539_nl, fsm_output[2]);
  assign nand_411_nl = ~((fsm_output[1]) & mux_3541_nl);
  assign nand_139_nl = ~((fsm_output[4]) & (fsm_output[9]) & (fsm_output[6]) & (fsm_output[8])
      & (~ (fsm_output[10])));
  assign mux_3537_nl = MUX_s_1_2_2(nand_139_nl, or_tmp_3095, fsm_output[3]);
  assign or_3166_nl = (~ (fsm_output[7])) | (fsm_output[5]) | mux_3537_nl;
  assign nor_582_nl = ~((~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[6])
      | (fsm_output[8]) | (fsm_output[10]));
  assign nor_583_nl = ~((fsm_output[4]) | (fsm_output[9]) | nand_142_cse);
  assign mux_3536_nl = MUX_s_1_2_2(nor_582_nl, nor_583_nl, fsm_output[3]);
  assign nand_104_nl = ~((~((fsm_output[7]) | (~ (fsm_output[5])))) & mux_3536_nl);
  assign mux_3538_nl = MUX_s_1_2_2(or_3166_nl, nand_104_nl, fsm_output[2]);
  assign or_3499_nl = (fsm_output[1]) | mux_3538_nl;
  assign mux_3542_nl = MUX_s_1_2_2(nand_411_nl, or_3499_nl, fsm_output[0]);
  assign or_3228_nl = (fsm_output[9]) | (fsm_output[6]) | mux_tmp_3632;
  assign or_3226_nl = (~ (fsm_output[6])) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (~((fsm_output[8]) & (fsm_output[4]) & (fsm_output[10])));
  assign or_3224_nl = (fsm_output[6]) | (fsm_output[5]) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[8]) | (~ (fsm_output[4])) | (fsm_output[10]);
  assign mux_3634_nl = MUX_s_1_2_2(or_3226_nl, or_3224_nl, fsm_output[9]);
  assign mux_3635_nl = MUX_s_1_2_2(or_3228_nl, mux_3634_nl, fsm_output[2]);
  assign nor_562_nl = ~((fsm_output[1]) | mux_3635_nl);
  assign nor_563_nl = ~((~ (fsm_output[9])) | (fsm_output[6]) | mux_tmp_3632);
  assign or_3217_nl = (fsm_output[5]) | (~ (fsm_output[7])) | (~ (fsm_output[3]))
      | (fsm_output[8]) | not_tmp_39;
  assign or_3215_nl = (~ (fsm_output[5])) | (fsm_output[7]) | (fsm_output[3]) | (~
      (fsm_output[8])) | (fsm_output[4]) | (fsm_output[10]);
  assign mux_3631_nl = MUX_s_1_2_2(or_3217_nl, or_3215_nl, fsm_output[6]);
  assign nor_564_nl = ~((fsm_output[9]) | mux_3631_nl);
  assign mux_3633_nl = MUX_s_1_2_2(nor_563_nl, nor_564_nl, fsm_output[2]);
  assign and_361_nl = (fsm_output[1]) & mux_3633_nl;
  assign mux_3636_nl = MUX_s_1_2_2(nor_562_nl, and_361_nl, fsm_output[0]);
  assign COMP_LOOP_nor_14_nl = ~((z_out_2_12_1[3]) | (z_out_2_12_1[1]) | (z_out_2_12_1[0]));
  assign mux_3637_nl = MUX_s_1_2_2(mux_tmp_3457, mux_tmp_3474, fsm_output[6]);
  assign mux_3638_nl = MUX_s_1_2_2((~ mux_3485_itm), mux_3637_nl, fsm_output[4]);
  assign mux_3639_nl = MUX_s_1_2_2(mux_3638_nl, mux_tmp_3481, fsm_output[1]);
  assign mux_3640_nl = MUX_s_1_2_2(mux_tmp_3491, mux_3639_nl, fsm_output[0]);
  assign mux_3641_nl = MUX_s_1_2_2(mux_3640_nl, mux_tmp_3472, fsm_output[9]);
  assign mux_3642_nl = MUX_s_1_2_2(mux_3641_nl, mux_tmp_3453, fsm_output[10]);
  assign COMP_LOOP_mux1h_477_nl = MUX1HOT_s_1_4_2((COMP_LOOP_k_9_4_sva_4_0[4]), COMP_LOOP_nor_137_itm,
      COMP_LOOP_nor_134_itm, COMP_LOOP_nor_14_nl, {and_dcpl_257 , not_tmp_701 , (~
      mux_3642_nl) , COMP_LOOP_or_32_cse});
  assign or_3240_nl = (fsm_output[9]) | (fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[8]))
      | (fsm_output[10]);
  assign or_3239_nl = (fsm_output[9]) | (~ (fsm_output[3])) | (~ (fsm_output[4]))
      | (fsm_output[8]) | (~ (fsm_output[10]));
  assign mux_3647_nl = MUX_s_1_2_2(or_3240_nl, or_3239_nl, fsm_output[5]);
  assign or_3241_nl = (fsm_output[7:6]!=2'b00) | mux_3647_nl;
  assign or_3236_nl = (~ (fsm_output[6])) | (fsm_output[5]) | (fsm_output[9]) | (~
      (fsm_output[3])) | (~ (fsm_output[4])) | (fsm_output[8]) | (fsm_output[10]);
  assign or_3235_nl = (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[3])) | (~
      (fsm_output[4])) | (fsm_output[8]) | (fsm_output[10]);
  assign or_3234_nl = (fsm_output[5]) | (~ (fsm_output[9])) | (fsm_output[3]) | (~
      (fsm_output[4])) | (~ (fsm_output[8])) | (fsm_output[10]);
  assign mux_3645_nl = MUX_s_1_2_2(or_3235_nl, or_3234_nl, fsm_output[6]);
  assign mux_3646_nl = MUX_s_1_2_2(or_3236_nl, mux_3645_nl, fsm_output[7]);
  assign mux_3648_nl = MUX_s_1_2_2(or_3241_nl, mux_3646_nl, fsm_output[0]);
  assign or_3497_nl = (fsm_output[2]) | mux_3648_nl;
  assign or_3498_nl = (fsm_output[0]) | (fsm_output[7]) | (~ (fsm_output[6])) | (~
      (fsm_output[5])) | (~ (fsm_output[9])) | (~ (fsm_output[3])) | (fsm_output[4])
      | (~ (fsm_output[8])) | (fsm_output[10]);
  assign nor_560_nl = ~((~ (fsm_output[6])) | (~ (fsm_output[5])) | (fsm_output[9])
      | (fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[8])) | (fsm_output[10]));
  assign nor_561_nl = ~((fsm_output[6]) | (fsm_output[5]) | (fsm_output[9]) | (~
      (fsm_output[3])) | (~ (fsm_output[4])) | (fsm_output[8]) | (~ (fsm_output[10])));
  assign mux_3643_nl = MUX_s_1_2_2(nor_560_nl, nor_561_nl, fsm_output[7]);
  assign nand_410_nl = ~((fsm_output[0]) & mux_3643_nl);
  assign mux_3644_nl = MUX_s_1_2_2(or_3498_nl, nand_410_nl, fsm_output[2]);
  assign mux_3649_nl = MUX_s_1_2_2(or_3497_nl, mux_3644_nl, fsm_output[1]);
  assign nor_555_nl = ~((fsm_output[5]) | (~ (fsm_output[2])) | (~ (fsm_output[1]))
      | (fsm_output[3]) | (fsm_output[4]) | (~ (fsm_output[8])) | (fsm_output[9])
      | (fsm_output[6]) | (~ (fsm_output[10])));
  assign or_3253_nl = (~ (fsm_output[4])) | (~ (fsm_output[8])) | (fsm_output[9])
      | not_tmp_49;
  assign mux_3653_nl = MUX_s_1_2_2(or_3253_nl, or_tmp_3176, fsm_output[3]);
  assign or_3251_nl = (~ (fsm_output[3])) | (fsm_output[4]) | (~ (fsm_output[8]))
      | (fsm_output[9]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_3654_nl = MUX_s_1_2_2(mux_3653_nl, or_3251_nl, fsm_output[1]);
  assign nor_556_nl = ~((fsm_output[5]) | (~ (fsm_output[2])) | mux_3654_nl);
  assign mux_3655_nl = MUX_s_1_2_2(nor_555_nl, nor_556_nl, fsm_output[7]);
  assign or_3249_nl = (fsm_output[2]) | (~ (fsm_output[1])) | (fsm_output[3]) | (fsm_output[4])
      | (~ (fsm_output[8])) | (~ (fsm_output[9])) | (fsm_output[6]) | (fsm_output[10]);
  assign nand_383_nl = ~((fsm_output[1]) & (fsm_output[3]) & (fsm_output[4]) & (~
      (fsm_output[8])) & (fsm_output[9]) & (~ (fsm_output[6])) & (fsm_output[10]));
  assign or_3244_nl = (fsm_output[4]) | (~ (fsm_output[8])) | (fsm_output[9]) | not_tmp_49;
  assign mux_3650_nl = MUX_s_1_2_2(or_tmp_3176, or_3244_nl, fsm_output[3]);
  assign or_3246_nl = (fsm_output[1]) | mux_3650_nl;
  assign mux_3651_nl = MUX_s_1_2_2(nand_383_nl, or_3246_nl, fsm_output[2]);
  assign mux_3652_nl = MUX_s_1_2_2(or_3249_nl, mux_3651_nl, fsm_output[5]);
  assign nor_557_nl = ~((fsm_output[7]) | mux_3652_nl);
  assign mux_3656_nl = MUX_s_1_2_2(mux_3655_nl, nor_557_nl, fsm_output[0]);
  assign COMP_LOOP_nor_17_nl = ~((z_out_2_12_1[2:0]!=3'b000));
  assign COMP_LOOP_mux1h_479_nl = MUX1HOT_s_1_3_2(COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      COMP_LOOP_nor_137_itm, COMP_LOOP_nor_17_nl, {not_tmp_701 , (~ mux_3494_itm)
      , COMP_LOOP_or_32_cse});
  assign or_3266_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[6]) | (~
      (fsm_output[9]));
  assign mux_3660_nl = MUX_s_1_2_2(or_3417_cse, or_3266_nl, fsm_output[0]);
  assign nand_130_nl = ~((fsm_output[0]) & (fsm_output[1]) & (fsm_output[2]) & (fsm_output[6])
      & (~ (fsm_output[9])));
  assign mux_3661_nl = MUX_s_1_2_2(mux_3660_nl, nand_130_nl, fsm_output[5]);
  assign nor_552_nl = ~((fsm_output[7]) | mux_3661_nl);
  assign nor_553_nl = ~((~ (fsm_output[7])) | (fsm_output[5]) | (fsm_output[0]) |
      (~ (fsm_output[1])) | (~ (fsm_output[2])) | (~ (fsm_output[6])) | (fsm_output[9]));
  assign mux_3662_nl = MUX_s_1_2_2(nor_552_nl, nor_553_nl, fsm_output[3]);
  assign nand_389_nl = ~((fsm_output[8]) & mux_3662_nl);
  assign or_3261_nl = (~ (fsm_output[1])) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[9]);
  assign mux_3658_nl = MUX_s_1_2_2(or_3261_nl, or_tmp_3190, fsm_output[0]);
  assign or_3353_nl = (fsm_output[7]) | (~ (fsm_output[5])) | mux_3658_nl;
  assign mux_3657_nl = MUX_s_1_2_2(or_tmp_3190, or_3417_cse, fsm_output[0]);
  assign or_3260_nl = (~ (fsm_output[7])) | (fsm_output[5]) | mux_3657_nl;
  assign mux_3659_nl = MUX_s_1_2_2(or_3353_nl, or_3260_nl, fsm_output[3]);
  assign or_3443_nl = (fsm_output[8]) | mux_3659_nl;
  assign mux_3663_nl = MUX_s_1_2_2(nand_389_nl, or_3443_nl, fsm_output[4]);
  assign nor_547_nl = ~((fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) |
      (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[4]) | (fsm_output[9]) |
      not_tmp_253);
  assign or_3282_nl = (fsm_output[0]) | (~ (fsm_output[4])) | (fsm_output[9]) | (fsm_output[2])
      | (~ (fsm_output[10]));
  assign nand_382_nl = ~((fsm_output[0]) & (fsm_output[4]) & (fsm_output[9]) & (~
      (fsm_output[2])) & (fsm_output[10]));
  assign mux_3667_nl = MUX_s_1_2_2(or_3282_nl, nand_382_nl, fsm_output[1]);
  assign nor_548_nl = ~((fsm_output[6]) | mux_3667_nl);
  assign nor_549_nl = ~((~ (fsm_output[0])) | (fsm_output[4]) | (fsm_output[9]) |
      not_tmp_253);
  assign nor_550_nl = ~((fsm_output[0]) | (fsm_output[4]) | (~ (fsm_output[9])) |
      (fsm_output[2]) | (fsm_output[10]));
  assign mux_3666_nl = MUX_s_1_2_2(nor_549_nl, nor_550_nl, fsm_output[1]);
  assign and_358_nl = (fsm_output[6]) & mux_3666_nl;
  assign mux_3668_nl = MUX_s_1_2_2(nor_548_nl, and_358_nl, fsm_output[8]);
  assign and_357_nl = (fsm_output[3]) & mux_3668_nl;
  assign mux_3669_nl = MUX_s_1_2_2(nor_547_nl, and_357_nl, fsm_output[5]);
  assign or_3273_nl = (~ (fsm_output[4])) | (fsm_output[9]) | not_tmp_253;
  assign or_3271_nl = (~ (fsm_output[4])) | (~ (fsm_output[9])) | (fsm_output[2])
      | (fsm_output[10]);
  assign mux_3664_nl = MUX_s_1_2_2(or_3273_nl, or_3271_nl, fsm_output[0]);
  assign or_3274_nl = (~ (fsm_output[8])) | (~ (fsm_output[6])) | (fsm_output[1])
      | mux_3664_nl;
  assign or_3269_nl = (fsm_output[8]) | (fsm_output[6]) | (~ (fsm_output[1])) | (~
      (fsm_output[0])) | (~ (fsm_output[4])) | (fsm_output[9]) | not_tmp_253;
  assign mux_3665_nl = MUX_s_1_2_2(or_3274_nl, or_3269_nl, fsm_output[3]);
  assign nor_551_nl = ~((fsm_output[5]) | mux_3665_nl);
  assign mux_3670_nl = MUX_s_1_2_2(mux_3669_nl, nor_551_nl, fsm_output[7]);
  assign mux_3761_nl = MUX_s_1_2_2((~ mux_tmp_236), mux_tmp_228, fsm_output[7]);
  assign mux_3762_nl = MUX_s_1_2_2(mux_3761_nl, mux_tmp_3720, fsm_output[1]);
  assign mux_3763_nl = MUX_s_1_2_2(mux_tmp_3724, mux_3762_nl, and_366_cse);
  assign mux_3755_nl = MUX_s_1_2_2(or_361_cse, and_757_cse, fsm_output[5]);
  assign mux_3756_nl = MUX_s_1_2_2(mux_3755_nl, or_tmp_114, fsm_output[7]);
  assign mux_3757_nl = MUX_s_1_2_2(mux_3756_nl, mux_tmp_3753, fsm_output[0]);
  assign mux_3758_nl = MUX_s_1_2_2(mux_3757_nl, mux_tmp_3674, fsm_output[1]);
  assign mux_3754_nl = MUX_s_1_2_2(mux_tmp_3753, mux_tmp_3705, and_526_cse);
  assign mux_3759_nl = MUX_s_1_2_2(mux_3758_nl, mux_3754_nl, fsm_output[2]);
  assign or_3302_nl = (fsm_output[5]) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign mux_3750_nl = MUX_s_1_2_2(mux_tmp_231, or_3302_nl, fsm_output[7]);
  assign mux_3751_nl = MUX_s_1_2_2(mux_tmp_3698, mux_3750_nl, or_3388_cse);
  assign mux_3752_nl = MUX_s_1_2_2(mux_3751_nl, or_tmp_3224, fsm_output[2]);
  assign mux_3760_nl = MUX_s_1_2_2(mux_3759_nl, mux_3752_nl, fsm_output[4]);
  assign mux_3764_nl = MUX_s_1_2_2(mux_3763_nl, mux_3760_nl, fsm_output[8]);
  assign mux_3744_nl = MUX_s_1_2_2((~ nand_tmp_7), mux_tmp_3736, fsm_output[7]);
  assign nor_546_nl = ~((~ (fsm_output[5])) | (fsm_output[10]));
  assign mux_3743_nl = MUX_s_1_2_2(nor_546_nl, mux_tmp_3736, fsm_output[7]);
  assign mux_3745_nl = MUX_s_1_2_2(mux_3744_nl, mux_3743_nl, fsm_output[0]);
  assign mux_3742_nl = MUX_s_1_2_2(mux_tmp_3737, mux_tmp_3739, fsm_output[0]);
  assign mux_3746_nl = MUX_s_1_2_2(mux_3745_nl, mux_3742_nl, fsm_output[1]);
  assign mux_3740_nl = MUX_s_1_2_2(mux_tmp_3739, mux_tmp_3737, fsm_output[0]);
  assign mux_3741_nl = MUX_s_1_2_2(mux_3740_nl, mux_tmp_3691, fsm_output[1]);
  assign mux_3747_nl = MUX_s_1_2_2(mux_3746_nl, mux_3741_nl, fsm_output[2]);
  assign mux_3748_nl = MUX_s_1_2_2(mux_3747_nl, mux_tmp_3691, fsm_output[4]);
  assign or_3298_nl = (fsm_output[5]) | (fsm_output[9]) | (fsm_output[10]);
  assign mux_3733_nl = MUX_s_1_2_2(or_3298_nl, nand_tmp_7, fsm_output[7]);
  assign mux_3734_nl = MUX_s_1_2_2(mux_tmp_3681, mux_3733_nl, and_529_cse);
  assign and_349_nl = (fsm_output[1]) & (fsm_output[7]);
  assign mux_3731_nl = MUX_s_1_2_2(mux_tmp_215, nor_tmp_23, and_349_nl);
  assign mux_3729_nl = MUX_s_1_2_2(mux_tmp_215, nor_tmp_23, fsm_output[7]);
  assign mux_3728_nl = MUX_s_1_2_2(mux_tmp_215, mux_tmp_236, fsm_output[7]);
  assign mux_3730_nl = MUX_s_1_2_2(mux_3729_nl, mux_3728_nl, or_3388_cse);
  assign mux_3732_nl = MUX_s_1_2_2(mux_3731_nl, mux_3730_nl, fsm_output[2]);
  assign mux_3735_nl = MUX_s_1_2_2(mux_3734_nl, mux_3732_nl, fsm_output[4]);
  assign mux_3749_nl = MUX_s_1_2_2(mux_3748_nl, mux_3735_nl, fsm_output[8]);
  assign mux_3765_nl = MUX_s_1_2_2(mux_3764_nl, mux_3749_nl, fsm_output[6]);
  assign mux_3719_nl = MUX_s_1_2_2((~ or_tmp_114), mux_tmp_228, fsm_output[7]);
  assign mux_3721_nl = MUX_s_1_2_2(mux_tmp_3720, mux_3719_nl, fsm_output[0]);
  assign mux_3716_nl = MUX_s_1_2_2((~ and_757_cse), and_757_cse, fsm_output[5]);
  assign mux_3717_nl = MUX_s_1_2_2(mux_3716_nl, mux_259_cse, fsm_output[7]);
  assign mux_3722_nl = MUX_s_1_2_2(mux_3721_nl, mux_3717_nl, fsm_output[1]);
  assign mux_3713_nl = MUX_s_1_2_2((~ or_tmp_114), mux_259_cse, fsm_output[7]);
  assign mux_3711_nl = MUX_s_1_2_2((~ or_tmp_114), and_757_cse, fsm_output[7]);
  assign mux_3714_nl = MUX_s_1_2_2(mux_3713_nl, mux_3711_nl, fsm_output[0]);
  assign mux_3710_nl = MUX_s_1_2_2((~ or_tmp_114), nor_tmp_23, fsm_output[7]);
  assign mux_3715_nl = MUX_s_1_2_2(mux_3714_nl, mux_3710_nl, fsm_output[1]);
  assign mux_3723_nl = MUX_s_1_2_2(mux_3722_nl, mux_3715_nl, fsm_output[2]);
  assign mux_3725_nl = MUX_s_1_2_2(mux_tmp_3724, mux_3723_nl, fsm_output[4]);
  assign or_3295_nl = and_350_cse | and_757_cse;
  assign mux_3706_nl = MUX_s_1_2_2(mux_tmp_3705, or_3295_nl, fsm_output[0]);
  assign mux_3707_nl = MUX_s_1_2_2(mux_3706_nl, mux_tmp_3701, fsm_output[1]);
  assign mux_3699_nl = MUX_s_1_2_2(mux_tmp_231, or_tmp_114, fsm_output[7]);
  assign mux_3702_nl = MUX_s_1_2_2(mux_tmp_3701, mux_3699_nl, fsm_output[0]);
  assign mux_3703_nl = MUX_s_1_2_2(mux_3702_nl, mux_tmp_3698, fsm_output[1]);
  assign mux_3708_nl = MUX_s_1_2_2(mux_3707_nl, mux_3703_nl, fsm_output[2]);
  assign mux_3709_nl = MUX_s_1_2_2(mux_3708_nl, or_tmp_3224, fsm_output[4]);
  assign mux_3726_nl = MUX_s_1_2_2(mux_3725_nl, mux_3709_nl, fsm_output[8]);
  assign mux_3689_nl = MUX_s_1_2_2((~ or_2414_cse), or_tmp_104, fsm_output[5]);
  assign mux_3690_nl = MUX_s_1_2_2(mux_3689_nl, or_361_cse, fsm_output[7]);
  assign mux_3692_nl = MUX_s_1_2_2(mux_tmp_3691, mux_3690_nl, fsm_output[1]);
  assign nand_380_nl = ~((~((fsm_output[5]) & (fsm_output[9]))) & (fsm_output[10]));
  assign mux_3687_nl = MUX_s_1_2_2(nand_380_nl, or_361_cse, fsm_output[7]);
  assign mux_3685_nl = MUX_s_1_2_2((~ and_757_cse), or_tmp_104, fsm_output[5]);
  assign mux_3686_nl = MUX_s_1_2_2(mux_3685_nl, or_361_cse, fsm_output[7]);
  assign mux_3688_nl = MUX_s_1_2_2(mux_3687_nl, mux_3686_nl, and_526_cse);
  assign mux_3693_nl = MUX_s_1_2_2(mux_3692_nl, mux_3688_nl, fsm_output[2]);
  assign mux_3694_nl = MUX_s_1_2_2(mux_tmp_3691, mux_3693_nl, fsm_output[4]);
  assign mux_3682_nl = MUX_s_1_2_2(mux_tmp_3681, mux_tmp_3679, and_526_cse);
  assign nor_527_nl = ~((fsm_output[0]) | (~ (fsm_output[7])));
  assign mux_3678_nl = MUX_s_1_2_2(mux_tmp_215, nand_tmp_7, nor_527_nl);
  assign mux_3680_nl = MUX_s_1_2_2(mux_tmp_3679, mux_3678_nl, fsm_output[1]);
  assign mux_3683_nl = MUX_s_1_2_2(mux_3682_nl, mux_3680_nl, fsm_output[2]);
  assign mux_3676_nl = MUX_s_1_2_2(mux_tmp_3673, mux_tmp_3674, and_526_cse);
  assign mux_3675_nl = MUX_s_1_2_2(mux_tmp_3674, mux_tmp_3673, or_3388_cse);
  assign mux_3677_nl = MUX_s_1_2_2(mux_3676_nl, mux_3675_nl, fsm_output[2]);
  assign mux_3684_nl = MUX_s_1_2_2(mux_3683_nl, mux_3677_nl, fsm_output[4]);
  assign mux_3695_nl = MUX_s_1_2_2(mux_3694_nl, mux_3684_nl, fsm_output[8]);
  assign mux_3727_nl = MUX_s_1_2_2(mux_3726_nl, mux_3695_nl, fsm_output[6]);
  assign mux_3766_nl = MUX_s_1_2_2(mux_3765_nl, mux_3727_nl, fsm_output[3]);
  assign COMP_LOOP_or_28_nl = and_dcpl_140 | and_dcpl_197;
  assign COMP_LOOP_mux1h_480_nl = MUX1HOT_s_1_6_2(modExp_exp_1_4_1_sva, COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm,
      (COMP_LOOP_k_9_4_sva_4_0[0]), (z_out_6[7]), (z_out_7[6]), (z_out_7[5]), {not_tmp_701
      , (~ mux_3766_nl) , not_tmp_688 , COMP_LOOP_or_28_nl , and_dcpl_171 , and_dcpl_226});
  assign or_3396_nl = (fsm_output[5]) | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[10]);
  assign nand_175_nl = ~((fsm_output[0]) & (fsm_output[5]) & (fsm_output[7]) & (fsm_output[9])
      & (fsm_output[10]));
  assign mux_2449_nl = MUX_s_1_2_2(or_3396_nl, nand_175_nl, fsm_output[1]);
  assign mux_2450_nl = MUX_s_1_2_2(mux_2449_nl, nand_356_cse, or_491_cse);
  assign mux_2451_nl = MUX_s_1_2_2(mux_2450_nl, nand_357_cse, fsm_output[6]);
  assign mux_2452_nl = MUX_s_1_2_2(mux_2451_nl, nand_358_cse, fsm_output[8]);
  assign or_3549_nl = (fsm_output[2]) | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[9])
      | (fsm_output[10]);
  assign mux_3885_nl = MUX_s_1_2_2(or_3549_nl, mux_tmp_3864, fsm_output[3]);
  assign nor_1705_nl = ~((fsm_output[6]) | (~ mux_3885_nl));
  assign nor_1706_nl = ~((fsm_output[2:1]!=2'b00) | (~ and_757_cse));
  assign and_1165_nl = (fsm_output[2]) & (~ or_tmp_3347);
  assign mux_3883_nl = MUX_s_1_2_2(nor_1706_nl, and_1165_nl, fsm_output[3]);
  assign and_1166_nl = (fsm_output[3:2]==2'b11) & (~ or_tmp_3352);
  assign mux_3884_nl = MUX_s_1_2_2(mux_3883_nl, and_1166_nl, fsm_output[6]);
  assign mux_3886_nl = MUX_s_1_2_2(nor_1705_nl, mux_3884_nl, fsm_output[4]);
  assign or_3619_nl = (fsm_output[3:2]!=2'b00) | (~ nor_tmp_552);
  assign or_3543_nl = (fsm_output[1:0]!=2'b00) | (~ and_757_cse);
  assign mux_3880_nl = MUX_s_1_2_2((~ nor_tmp_554), or_3543_nl, fsm_output[2]);
  assign or_3620_nl = (fsm_output[3]) | mux_3880_nl;
  assign mux_3881_nl = MUX_s_1_2_2(or_3619_nl, or_3620_nl, fsm_output[6]);
  assign or_3541_nl = (~((fsm_output[1:0]!=2'b01))) | (fsm_output[10:9]!=2'b00);
  assign mux_3877_nl = MUX_s_1_2_2(or_3541_nl, or_tmp_3339, fsm_output[2]);
  assign mux_3878_nl = MUX_s_1_2_2(mux_3877_nl, (~ or_tmp_3357), fsm_output[3]);
  assign nor_1708_nl = ~((fsm_output[2:0]!=3'b000) | (~ and_757_cse));
  assign mux_3876_nl = MUX_s_1_2_2(mux_tmp_3856, nor_1708_nl, fsm_output[3]);
  assign mux_3879_nl = MUX_s_1_2_2(mux_3878_nl, mux_3876_nl, fsm_output[6]);
  assign mux_3882_nl = MUX_s_1_2_2(mux_3881_nl, mux_3879_nl, fsm_output[4]);
  assign mux_3887_nl = MUX_s_1_2_2(mux_3886_nl, mux_3882_nl, fsm_output[5]);
  assign or_3537_nl = (~ (fsm_output[1])) | (fsm_output[9]) | (fsm_output[10]);
  assign mux_3871_nl = MUX_s_1_2_2(or_3537_nl, or_tmp_3339, fsm_output[2]);
  assign mux_3872_nl = MUX_s_1_2_2((~ mux_3871_nl), or_tmp_3357, fsm_output[3]);
  assign mux_3868_nl = MUX_s_1_2_2(and_757_cse, mux_tmp_227, and_526_cse);
  assign mux_3869_nl = MUX_s_1_2_2(mux_3868_nl, mux_tmp_3830, fsm_output[2]);
  assign or_3534_nl = (fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[9])
      | (~ (fsm_output[10]));
  assign mux_3870_nl = MUX_s_1_2_2(mux_3869_nl, or_3534_nl, fsm_output[3]);
  assign mux_3873_nl = MUX_s_1_2_2(mux_3872_nl, mux_3870_nl, fsm_output[6]);
  assign nand_417_nl = ~((fsm_output[3]) & (~ mux_tmp_3864));
  assign mux_3867_nl = MUX_s_1_2_2(nand_417_nl, mux_tmp_3848, fsm_output[6]);
  assign mux_3874_nl = MUX_s_1_2_2(mux_3873_nl, mux_3867_nl, fsm_output[4]);
  assign and_1168_nl = (fsm_output[6]) & (fsm_output[3]);
  assign mux_3864_nl = MUX_s_1_2_2(and_757_cse, mux_tmp_3841, and_1168_nl);
  assign mux_3865_nl = MUX_s_1_2_2(mux_3864_nl, or_3532_cse, fsm_output[4]);
  assign mux_3875_nl = MUX_s_1_2_2(mux_3874_nl, mux_3865_nl, fsm_output[5]);
  assign mux_3888_nl = MUX_s_1_2_2(mux_3887_nl, mux_3875_nl, fsm_output[7]);
  assign mux_3859_nl = MUX_s_1_2_2(mux_tmp_3856, and_757_cse, fsm_output[3]);
  assign mux_3860_nl = MUX_s_1_2_2(mux_3859_nl, mux_tmp_3839, fsm_output[6]);
  assign or_3529_nl = (fsm_output[3]) | mux_tmp_3828;
  assign mux_3857_nl = MUX_s_1_2_2(and_757_cse, or_3529_nl, fsm_output[6]);
  assign mux_3861_nl = MUX_s_1_2_2(mux_3860_nl, mux_3857_nl, fsm_output[4]);
  assign mux_3852_nl = MUX_s_1_2_2(and_757_cse, mux_tmp_227, fsm_output[1]);
  assign mux_3851_nl = MUX_s_1_2_2(mux_tmp_227, or_tmp_104, or_3388_cse);
  assign mux_3853_nl = MUX_s_1_2_2(mux_3852_nl, mux_3851_nl, fsm_output[2]);
  assign mux_3854_nl = MUX_s_1_2_2(and_757_cse, mux_3853_nl, fsm_output[3]);
  assign mux_3855_nl = MUX_s_1_2_2(mux_3854_nl, mux_tmp_3848, fsm_output[6]);
  assign mux_3848_nl = MUX_s_1_2_2(or_tmp_3344, and_757_cse, fsm_output[6]);
  assign mux_3856_nl = MUX_s_1_2_2(mux_3855_nl, mux_3848_nl, fsm_output[4]);
  assign mux_3862_nl = MUX_s_1_2_2(mux_3861_nl, mux_3856_nl, fsm_output[5]);
  assign mux_3845_nl = MUX_s_1_2_2(and_757_cse, or_tmp_3344, fsm_output[6]);
  assign or_3522_nl = (fsm_output[3]) | mux_tmp_3841;
  assign mux_3844_nl = MUX_s_1_2_2(or_3522_nl, mux_tmp_3839, fsm_output[6]);
  assign mux_3846_nl = MUX_s_1_2_2(mux_3845_nl, mux_3844_nl, fsm_output[4]);
  assign nand_416_nl = ~((fsm_output[2]) & (~ or_tmp_3337));
  assign mux_3837_nl = MUX_s_1_2_2(nor_tmp_549, and_757_cse, fsm_output[2]);
  assign mux_3838_nl = MUX_s_1_2_2(nand_416_nl, mux_3837_nl, fsm_output[3]);
  assign mux_3839_nl = MUX_s_1_2_2(mux_3838_nl, and_757_cse, fsm_output[6]);
  assign mux_3834_nl = MUX_s_1_2_2(and_757_cse, mux_tmp_227, and_536_cse);
  assign or_3513_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[9]) | (~ (fsm_output[10]));
  assign mux_3833_nl = MUX_s_1_2_2(mux_tmp_3830, or_3513_nl, fsm_output[2]);
  assign mux_3835_nl = MUX_s_1_2_2(mux_3834_nl, mux_3833_nl, fsm_output[3]);
  assign mux_3831_nl = MUX_s_1_2_2(and_757_cse, mux_tmp_3828, fsm_output[3]);
  assign mux_3836_nl = MUX_s_1_2_2(mux_3835_nl, mux_3831_nl, fsm_output[6]);
  assign mux_3840_nl = MUX_s_1_2_2(mux_3839_nl, mux_3836_nl, fsm_output[4]);
  assign mux_3847_nl = MUX_s_1_2_2(mux_3846_nl, mux_3840_nl, fsm_output[5]);
  assign mux_3863_nl = MUX_s_1_2_2(mux_3862_nl, mux_3847_nl, fsm_output[7]);
  assign mux_3889_nl = MUX_s_1_2_2(mux_3888_nl, mux_3863_nl, fsm_output[8]);
  assign or_3612_nl = (~ (fsm_output[1])) | (fsm_output[10]) | (~ COMP_LOOP_nor_11_itm)
      | (~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign or_3611_nl = (fsm_output[1]) | (fsm_output[10]) | (fsm_output[6]) | (fsm_output[2])
      | (fsm_output[9]);
  assign mux_3938_nl = MUX_s_1_2_2(or_3612_nl, or_3611_nl, fsm_output[0]);
  assign mux_3936_nl = MUX_s_1_2_2(or_tmp_3409, or_2965_cse, fsm_output[1]);
  assign mux_3937_nl = MUX_s_1_2_2(mux_3936_nl, mux_3935_cse, fsm_output[0]);
  assign mux_3939_nl = MUX_s_1_2_2(mux_3938_nl, mux_3937_nl, fsm_output[3]);
  assign or_3608_nl = (fsm_output[3]) | (fsm_output[0]) | (~ (fsm_output[1])) | (~
      (fsm_output[10])) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[6])) | (fsm_output[2])
      | (~ (fsm_output[9]));
  assign mux_3940_nl = MUX_s_1_2_2(mux_3939_nl, or_3608_nl, fsm_output[5]);
  assign or_3606_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (~ (fsm_output[10]))
      | (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[9]));
  assign or_3604_nl = (fsm_output[1]) | (fsm_output[10]) | not_tmp_882;
  assign nand_423_nl = ~((fsm_output[1]) & (fsm_output[10]) & COMP_LOOP_nor_11_itm
      & (fsm_output[6]) & (fsm_output[2]) & (~ (fsm_output[9])));
  assign mux_3932_nl = MUX_s_1_2_2(or_3604_nl, nand_423_nl, fsm_output[0]);
  assign mux_3933_nl = MUX_s_1_2_2(or_3606_nl, mux_3932_nl, fsm_output[3]);
  assign or_3601_nl = (fsm_output[10]) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_3929_nl = MUX_s_1_2_2(or_3601_nl, mux_tmp_3906, fsm_output[1]);
  assign mux_3925_nl = MUX_s_1_2_2((fsm_output[9]), (~ (fsm_output[9])), fsm_output[2]);
  assign mux_3926_nl = MUX_s_1_2_2(mux_3925_nl, or_2855_cse, fsm_output[6]);
  assign mux_3927_nl = MUX_s_1_2_2(or_tmp_3402, mux_3926_nl, COMP_LOOP_nor_11_itm);
  assign or_3600_nl = (fsm_output[10]) | mux_3927_nl;
  assign mux_3928_nl = MUX_s_1_2_2(or_tmp_3409, or_3600_nl, fsm_output[1]);
  assign mux_3930_nl = MUX_s_1_2_2(mux_3929_nl, mux_3928_nl, fsm_output[0]);
  assign or_3599_nl = (~ (fsm_output[10])) | (fsm_output[6]) | (fsm_output[2]) |
      (fsm_output[9]);
  assign or_3598_nl = (~ (fsm_output[10])) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[6])
      | (fsm_output[2]) | (fsm_output[9]);
  assign mux_3923_nl = MUX_s_1_2_2(or_3599_nl, or_3598_nl, fsm_output[1]);
  assign nand_420_nl = ~((fsm_output[10]) & (~ mux_tmp_3903));
  assign or_3597_nl = (~ (fsm_output[10])) | (fsm_output[6]) | (fsm_output[2]) |
      (~ (fsm_output[9]));
  assign mux_3922_nl = MUX_s_1_2_2(nand_420_nl, or_3597_nl, fsm_output[1]);
  assign mux_3924_nl = MUX_s_1_2_2(mux_3923_nl, mux_3922_nl, fsm_output[0]);
  assign mux_3931_nl = MUX_s_1_2_2(mux_3930_nl, mux_3924_nl, fsm_output[3]);
  assign mux_3934_nl = MUX_s_1_2_2(mux_3933_nl, mux_3931_nl, fsm_output[5]);
  assign mux_3941_nl = MUX_s_1_2_2(mux_3940_nl, mux_3934_nl, fsm_output[4]);
  assign or_3594_nl = (fsm_output[10]) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[6]))
      | (fsm_output[2]) | (fsm_output[9]);
  assign mux_3918_nl = MUX_s_1_2_2(or_3594_nl, or_tmp_3382, fsm_output[1]);
  assign or_3593_nl = (~ (fsm_output[1])) | (fsm_output[10]) | (~ COMP_LOOP_nor_11_itm)
      | (~ (fsm_output[6])) | (fsm_output[2]) | (~ (fsm_output[9]));
  assign mux_3919_nl = MUX_s_1_2_2(mux_3918_nl, or_3593_nl, fsm_output[0]);
  assign or_3595_nl = (fsm_output[3]) | mux_3919_nl;
  assign or_3591_nl = (fsm_output[3]) | (~ (fsm_output[0])) | (fsm_output[1]) | (~
      (fsm_output[10])) | (~ COMP_LOOP_nor_11_itm) | (fsm_output[6]) | (fsm_output[2])
      | (fsm_output[9]);
  assign mux_3920_nl = MUX_s_1_2_2(or_3595_nl, or_3591_nl, fsm_output[5]);
  assign or_3589_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[10])
      | (~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign mux_3915_nl = MUX_s_1_2_2(or_tmp_3409, or_tmp_3403, fsm_output[1]);
  assign mux_3916_nl = MUX_s_1_2_2(mux_3915_nl, mux_tmp_3907, fsm_output[0]);
  assign mux_3917_nl = MUX_s_1_2_2(or_3589_nl, mux_3916_nl, fsm_output[3]);
  assign or_3590_nl = (fsm_output[5]) | mux_3917_nl;
  assign mux_3921_nl = MUX_s_1_2_2(mux_3920_nl, or_3590_nl, fsm_output[4]);
  assign mux_3942_nl = MUX_s_1_2_2(mux_3941_nl, mux_3921_nl, fsm_output[7]);
  assign or_3578_nl = (fsm_output[10]) | (fsm_output[6]) | (fsm_output[2]) | (~ (fsm_output[9]));
  assign mux_3906_nl = MUX_s_1_2_2(or_tmp_3403, or_3578_nl, fsm_output[1]);
  assign mux_3910_nl = MUX_s_1_2_2(mux_tmp_3907, mux_3906_nl, fsm_output[0]);
  assign or_3576_nl = (fsm_output[0]) | (fsm_output[1]) | (~ (fsm_output[10])) |
      (~ COMP_LOOP_nor_11_itm) | (fsm_output[6]) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_3911_nl = MUX_s_1_2_2(mux_3910_nl, or_3576_nl, fsm_output[3]);
  assign or_3575_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[10])
      | or_tmp_3384;
  assign or_3573_nl = (fsm_output[10]) | not_tmp_882;
  assign mux_3901_nl = MUX_s_1_2_2(or_3573_nl, or_tmp_3381, fsm_output[1]);
  assign mux_3902_nl = MUX_s_1_2_2(mux_3901_nl, mux_tmp_3892, fsm_output[0]);
  assign mux_3903_nl = MUX_s_1_2_2(or_3575_nl, mux_3902_nl, fsm_output[3]);
  assign mux_3912_nl = MUX_s_1_2_2(mux_3911_nl, mux_3903_nl, fsm_output[5]);
  assign or_3572_nl = (~ (fsm_output[5])) | (~ (fsm_output[3])) | (fsm_output[0])
      | (~ (fsm_output[1])) | (fsm_output[10]) | (fsm_output[6]) | (~ (fsm_output[2]))
      | (fsm_output[9]);
  assign mux_3913_nl = MUX_s_1_2_2(mux_3912_nl, or_3572_nl, fsm_output[4]);
  assign or_3571_nl = (~ (fsm_output[3])) | (fsm_output[0]) | (~ (fsm_output[1]))
      | (fsm_output[10]) | or_tmp_3384;
  assign or_3569_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[10]) |
      (fsm_output[6]) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign or_3568_nl = (fsm_output[1]) | (fsm_output[10]) | (fsm_output[6]) | (fsm_output[2])
      | (~ (fsm_output[9]));
  assign mux_3897_nl = MUX_s_1_2_2(or_3568_nl, or_2914_cse, fsm_output[0]);
  assign mux_3898_nl = MUX_s_1_2_2(or_3569_nl, mux_3897_nl, fsm_output[3]);
  assign mux_3899_nl = MUX_s_1_2_2(or_3571_nl, mux_3898_nl, fsm_output[5]);
  assign or_3556_nl = (fsm_output[10]) | (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[6]))
      | (fsm_output[2]) | (~ (fsm_output[9]));
  assign mux_3892_nl = MUX_s_1_2_2(or_tmp_3381, or_3556_nl, fsm_output[1]);
  assign mux_3895_nl = MUX_s_1_2_2(mux_tmp_3892, mux_3892_nl, fsm_output[0]);
  assign or_3565_nl = (fsm_output[3]) | mux_3895_nl;
  assign or_3554_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[10]) |
      (~ COMP_LOOP_nor_11_itm) | (~ (fsm_output[6])) | (~ (fsm_output[2])) | (fsm_output[9]);
  assign or_3553_nl = (fsm_output[1]) | (fsm_output[10]) | (~ COMP_LOOP_nor_11_itm)
      | (~ (fsm_output[6])) | (fsm_output[2]) | (~ (fsm_output[9]));
  assign or_3551_nl = (~ (fsm_output[1])) | (~ (fsm_output[10])) | (~ COMP_LOOP_nor_11_itm)
      | (~ (fsm_output[6])) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_3890_nl = MUX_s_1_2_2(or_3553_nl, or_3551_nl, fsm_output[0]);
  assign mux_3891_nl = MUX_s_1_2_2(or_3554_nl, mux_3890_nl, fsm_output[3]);
  assign mux_3896_nl = MUX_s_1_2_2(or_3565_nl, mux_3891_nl, fsm_output[5]);
  assign mux_3900_nl = MUX_s_1_2_2(mux_3899_nl, mux_3896_nl, fsm_output[4]);
  assign mux_3914_nl = MUX_s_1_2_2(mux_3913_nl, mux_3900_nl, fsm_output[7]);
  assign mux_3943_nl = MUX_s_1_2_2(mux_3942_nl, mux_3914_nl, fsm_output[8]);
  assign or_2641_nl = (fsm_output[1]) | (~ (fsm_output[4])) | (fsm_output[7]) | (~
      (fsm_output[5])) | (fsm_output[3]);
  assign or_2640_nl = (fsm_output[1]) | (fsm_output[4]) | (fsm_output[7]) | (fsm_output[5])
      | (~ (fsm_output[3]));
  assign mux_2638_nl = MUX_s_1_2_2(or_2641_nl, or_2640_nl, fsm_output[0]);
  assign or_2642_nl = (fsm_output[9]) | mux_2638_nl;
  assign or_2638_nl = (~ (fsm_output[9])) | (fsm_output[0]) | (~ (fsm_output[1]))
      | (fsm_output[4]) | (~ (fsm_output[7])) | (~ (fsm_output[5])) | (fsm_output[3]);
  assign mux_2639_nl = MUX_s_1_2_2(or_2642_nl, or_2638_nl, fsm_output[10]);
  assign or_3508_nl = mux_2639_nl | (fsm_output[2]) | (fsm_output[8]) | (fsm_output[6]);
  assign nor_1700_nl = ~((~ (fsm_output[3])) | (fsm_output[4]) | (~ (fsm_output[0]))
      | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[10]) | (fsm_output[9]) |
      (fsm_output[1]));
  assign or_3616_nl = (fsm_output[6]) | (~((fsm_output[7]) & (fsm_output[10]) & (fsm_output[9])
      & (fsm_output[1])));
  assign or_3615_nl = (~ (fsm_output[6])) | (fsm_output[7]) | (~((fsm_output[10])
      & (fsm_output[9]) & (fsm_output[1])));
  assign mux_3944_nl = MUX_s_1_2_2(or_3616_nl, or_3615_nl, fsm_output[0]);
  assign or_3613_nl = (fsm_output[0]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[10])
      | (fsm_output[9]) | (fsm_output[1]);
  assign mux_3945_nl = MUX_s_1_2_2(mux_3944_nl, or_3613_nl, fsm_output[4]);
  assign nor_1701_nl = ~((fsm_output[3]) | mux_3945_nl);
  assign mux_3946_nl = MUX_s_1_2_2(nor_1700_nl, nor_1701_nl, fsm_output[5]);
  assign nor_690_nl = ~((fsm_output[5]) | (fsm_output[7]) | (fsm_output[9]) | (fsm_output[10]));
  assign mux_2663_nl = MUX_s_1_2_2(nor_690_nl, mux_tmp_2659, and_526_cse);
  assign mux_2662_nl = MUX_s_1_2_2(mux_tmp_2659, and_465_cse, fsm_output[1]);
  assign mux_2664_nl = MUX_s_1_2_2(mux_2663_nl, mux_2662_nl, fsm_output[3]);
  assign mux_2661_nl = MUX_s_1_2_2(mux_tmp_2659, and_465_cse, fsm_output[3]);
  assign mux_2665_nl = MUX_s_1_2_2(mux_2664_nl, mux_2661_nl, fsm_output[2]);
  assign nand_170_nl = ~((fsm_output[3:0]==4'b1101));
  assign mux_2660_nl = MUX_s_1_2_2(mux_tmp_2659, and_465_cse, nand_170_nl);
  assign mux_2666_nl = MUX_s_1_2_2(mux_2665_nl, mux_2660_nl, fsm_output[4]);
  assign mux_2667_nl = MUX_s_1_2_2(mux_2666_nl, and_756_cse, fsm_output[6]);
  assign mux_2668_nl = MUX_s_1_2_2(mux_2667_nl, and_757_cse, fsm_output[8]);
  assign COMP_LOOP_or_8_nl = (COMP_LOOP_COMP_LOOP_nor_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_311_m1c);
  assign COMP_LOOP_or_9_nl = (COMP_LOOP_COMP_LOOP_and_305_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_311_m1c);
  assign COMP_LOOP_or_10_nl = (COMP_LOOP_COMP_LOOP_and_62_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_311_m1c);
  assign COMP_LOOP_or_11_nl = (COMP_LOOP_COMP_LOOP_and_2_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_311_m1c);
  assign COMP_LOOP_or_12_nl = (COMP_LOOP_COMP_LOOP_and_64_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_311_m1c);
  assign COMP_LOOP_or_13_nl = (COMP_LOOP_COMP_LOOP_and_4_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_311_m1c);
  assign COMP_LOOP_or_14_nl = (COMP_LOOP_COMP_LOOP_and_5_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_311_m1c);
  assign COMP_LOOP_or_15_nl = (COMP_LOOP_COMP_LOOP_and_6_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_311_m1c);
  assign COMP_LOOP_or_16_nl = (COMP_LOOP_COMP_LOOP_and_68_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_311_m1c);
  assign COMP_LOOP_or_17_nl = (COMP_LOOP_COMP_LOOP_and_8_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_311_m1c);
  assign COMP_LOOP_or_18_nl = (COMP_LOOP_COMP_LOOP_and_9_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_311_m1c);
  assign COMP_LOOP_or_19_nl = (COMP_LOOP_COMP_LOOP_and_10_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_311_m1c);
  assign COMP_LOOP_or_20_nl = (COMP_LOOP_COMP_LOOP_and_11_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_311_m1c);
  assign COMP_LOOP_or_21_nl = (COMP_LOOP_COMP_LOOP_and_12_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_311_m1c);
  assign COMP_LOOP_or_22_nl = (COMP_LOOP_COMP_LOOP_and_13_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_12_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_and_14_itm
      & and_311_m1c);
  assign COMP_LOOP_or_23_nl = (COMP_LOOP_COMP_LOOP_and_14_itm & and_dcpl_257) | (COMP_LOOP_COMP_LOOP_and_13_itm
      & and_279_m1c) | (COMP_LOOP_COMP_LOOP_and_12_itm & and_281_m1c) | (COMP_LOOP_COMP_LOOP_and_11_itm
      & and_284_m1c) | (COMP_LOOP_COMP_LOOP_and_10_itm & and_286_m1c) | (COMP_LOOP_COMP_LOOP_and_9_itm
      & and_288_m1c) | (COMP_LOOP_COMP_LOOP_and_8_itm & and_291_m1c) | (COMP_LOOP_COMP_LOOP_and_68_itm
      & and_292_m1c) | (COMP_LOOP_COMP_LOOP_and_6_itm & and_295_m1c) | (COMP_LOOP_COMP_LOOP_and_5_itm
      & and_297_m1c) | (COMP_LOOP_COMP_LOOP_and_4_itm & and_299_m1c) | (COMP_LOOP_COMP_LOOP_and_64_itm
      & and_302_m1c) | (COMP_LOOP_COMP_LOOP_and_2_itm & and_304_m1c) | (COMP_LOOP_COMP_LOOP_and_62_itm
      & and_307_m1c) | (COMP_LOOP_COMP_LOOP_and_305_itm & and_309_m1c) | (COMP_LOOP_COMP_LOOP_nor_itm
      & and_311_m1c);
  assign and_276_nl = (fsm_output[7]) & mux_tmp_2669;
  assign mux_2737_nl = MUX_s_1_2_2(mux_tmp_2736, and_276_nl, fsm_output[1]);
  assign nor_687_nl = ~((~ (fsm_output[9])) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_2734_nl = MUX_s_1_2_2(nor_687_nl, mux_tmp_2669, fsm_output[7]);
  assign mux_2735_nl = MUX_s_1_2_2(mux_2734_nl, mux_tmp_2709, and_526_cse);
  assign mux_2738_nl = MUX_s_1_2_2(mux_2737_nl, mux_2735_nl, fsm_output[2]);
  assign mux_2739_nl = MUX_s_1_2_2(mux_tmp_2736, mux_2738_nl, fsm_output[3]);
  assign mux_2730_nl = MUX_s_1_2_2(mux_tmp_2702, mux_tmp_2675, fsm_output[7]);
  assign mux_2729_nl = MUX_s_1_2_2(or_tmp_2604, mux_tmp_2675, fsm_output[7]);
  assign mux_2731_nl = MUX_s_1_2_2(mux_2730_nl, mux_2729_nl, or_3388_cse);
  assign or_2666_nl = (~(and_526_cse | (fsm_output[7]))) | (fsm_output[9]);
  assign mux_2728_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_167, or_2666_nl);
  assign mux_2732_nl = MUX_s_1_2_2(mux_2731_nl, mux_2728_nl, fsm_output[2]);
  assign and_454_nl = (fsm_output[2]) & (fsm_output[0]) & (fsm_output[1]) & (fsm_output[7]);
  assign mux_2727_nl = MUX_s_1_2_2(mux_tmp_2675, mux_tmp_2693, and_454_nl);
  assign mux_2733_nl = MUX_s_1_2_2(mux_2732_nl, mux_2727_nl, fsm_output[3]);
  assign mux_2740_nl = MUX_s_1_2_2(mux_2739_nl, mux_2733_nl, fsm_output[8]);
  assign mux_2725_nl = MUX_s_1_2_2((~ mux_2698_itm), mux_tmp_2675, fsm_output[7]);
  assign mux_2721_nl = MUX_s_1_2_2(mux_tmp_2675, mux_544_cse, fsm_output[7]);
  assign mux_2722_nl = MUX_s_1_2_2(mux_tmp_2690, mux_2721_nl, or_3388_cse);
  assign mux_2723_nl = MUX_s_1_2_2(mux_tmp_2690, mux_2722_nl, fsm_output[2]);
  assign mux_2717_nl = MUX_s_1_2_2((~ or_tmp_167), or_352_cse, fsm_output[9]);
  assign mux_2718_nl = MUX_s_1_2_2(mux_tmp_2693, mux_2717_nl, fsm_output[7]);
  assign mux_2719_nl = MUX_s_1_2_2(mux_2718_nl, mux_tmp_2715, and_526_cse);
  assign mux_2716_nl = MUX_s_1_2_2(mux_tmp_2715, mux_tmp_2672, fsm_output[1]);
  assign mux_2720_nl = MUX_s_1_2_2(mux_2719_nl, mux_2716_nl, fsm_output[2]);
  assign mux_2724_nl = MUX_s_1_2_2(mux_2723_nl, mux_2720_nl, fsm_output[3]);
  assign mux_2726_nl = MUX_s_1_2_2(mux_2725_nl, mux_2724_nl, fsm_output[8]);
  assign mux_2741_nl = MUX_s_1_2_2(mux_2740_nl, mux_2726_nl, fsm_output[5]);
  assign mux_2710_nl = MUX_s_1_2_2(mux_tmp_2709, mux_tmp_2706, fsm_output[1]);
  assign mux_2707_nl = MUX_s_1_2_2(mux_tmp_2706, mux_tmp_2703, and_526_cse);
  assign mux_2711_nl = MUX_s_1_2_2(mux_2710_nl, mux_2707_nl, fsm_output[2]);
  assign mux_2704_nl = MUX_s_1_2_2(mux_tmp_2703, mux_tmp_2700, fsm_output[1]);
  assign mux_2699_nl = MUX_s_1_2_2((~ mux_2698_itm), or_tmp_167, fsm_output[7]);
  assign mux_2701_nl = MUX_s_1_2_2(mux_tmp_2700, mux_2699_nl, or_3388_cse);
  assign mux_2705_nl = MUX_s_1_2_2(mux_2704_nl, mux_2701_nl, fsm_output[2]);
  assign mux_2712_nl = MUX_s_1_2_2(mux_2711_nl, mux_2705_nl, fsm_output[3]);
  assign mux_2694_nl = MUX_s_1_2_2(mux_tmp_2675, mux_tmp_2693, fsm_output[7]);
  assign mux_2695_nl = MUX_s_1_2_2(mux_2694_nl, mux_tmp_2691, fsm_output[1]);
  assign mux_2692_nl = MUX_s_1_2_2(mux_tmp_2691, mux_tmp_2690, or_3388_cse);
  assign mux_2696_nl = MUX_s_1_2_2(mux_2695_nl, mux_2692_nl, fsm_output[2]);
  assign mux_2697_nl = MUX_s_1_2_2(mux_2696_nl, mux_tmp_2690, fsm_output[3]);
  assign mux_2713_nl = MUX_s_1_2_2(mux_2712_nl, mux_2697_nl, fsm_output[8]);
  assign mux_2684_nl = MUX_s_1_2_2(nor_tmp_48, (fsm_output[6]), fsm_output[9]);
  assign mux_2685_nl = MUX_s_1_2_2((~ mux_2684_nl), mux_tmp_2675, fsm_output[7]);
  assign mux_2686_nl = MUX_s_1_2_2(mux_2685_nl, mux_tmp_2682, and_526_cse);
  assign mux_2680_nl = MUX_s_1_2_2(not_tmp_500, mux_tmp_2675, fsm_output[7]);
  assign mux_2683_nl = MUX_s_1_2_2(mux_tmp_2682, mux_2680_nl, fsm_output[1]);
  assign mux_2687_nl = MUX_s_1_2_2(mux_2686_nl, mux_2683_nl, fsm_output[2]);
  assign or_2658_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[7]);
  assign mux_2678_nl = MUX_s_1_2_2(not_tmp_500, mux_tmp_2675, or_2658_nl);
  assign mux_2674_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_167, and_458_cse);
  assign mux_2679_nl = MUX_s_1_2_2(mux_2678_nl, mux_2674_nl, fsm_output[2]);
  assign mux_2688_nl = MUX_s_1_2_2(mux_2687_nl, mux_2679_nl, fsm_output[3]);
  assign mux_2671_nl = MUX_s_1_2_2(mux_544_cse, mux_tmp_2669, fsm_output[7]);
  assign mux_2673_nl = MUX_s_1_2_2(mux_tmp_2672, mux_2671_nl, and_459_cse);
  assign mux_2689_nl = MUX_s_1_2_2(mux_2688_nl, mux_2673_nl, fsm_output[8]);
  assign mux_2714_nl = MUX_s_1_2_2(mux_2713_nl, mux_2689_nl, fsm_output[5]);
  assign and_312_nl = and_dcpl_236 & and_dcpl_127;
  assign COMP_LOOP_or_29_nl = ((~ (modulo_result_rem_cmp_z[63])) & and_317_m1c) |
      (~(mux_2840_itm | (modulo_result_rem_cmp_z[63])));
  assign COMP_LOOP_or_30_nl = ((modulo_result_rem_cmp_z[63]) & and_317_m1c) | ((~
      mux_2840_itm) & (modulo_result_rem_cmp_z[63]));
  assign COMP_LOOP_and_277_nl = COMP_LOOP_COMP_LOOP_nor_1_itm & mux_2771_m1c;
  assign COMP_LOOP_COMP_LOOP_and_932_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[0]) &
      COMP_LOOP_nor_11_itm & mux_2771_m1c;
  assign COMP_LOOP_COMP_LOOP_and_934_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[1]) &
      COMP_LOOP_nor_12_itm & mux_2771_m1c;
  assign COMP_LOOP_and_1_nl = COMP_LOOP_COMP_LOOP_and_137_itm & mux_2771_m1c;
  assign COMP_LOOP_COMP_LOOP_and_936_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[2]) &
      COMP_LOOP_nor_134_itm & mux_2771_m1c;
  assign COMP_LOOP_and_2_nl = COMP_LOOP_COMP_LOOP_and_139_itm & mux_2771_m1c;
  assign COMP_LOOP_and_3_nl = COMP_LOOP_COMP_LOOP_and_140_itm & mux_2771_m1c;
  assign COMP_LOOP_and_4_nl = COMP_LOOP_COMP_LOOP_and_141_itm & mux_2771_m1c;
  assign COMP_LOOP_COMP_LOOP_and_930_nl = (COMP_LOOP_acc_10_cse_12_1_1_sva[3]) &
      COMP_LOOP_nor_137_itm & mux_2771_m1c;
  assign COMP_LOOP_and_5_nl = COMP_LOOP_COMP_LOOP_and_143_itm & mux_2771_m1c;
  assign COMP_LOOP_and_6_nl = COMP_LOOP_COMP_LOOP_and_144_itm & mux_2771_m1c;
  assign COMP_LOOP_and_7_nl = COMP_LOOP_COMP_LOOP_and_145_itm & mux_2771_m1c;
  assign COMP_LOOP_and_8_nl = COMP_LOOP_COMP_LOOP_and_146_itm & mux_2771_m1c;
  assign COMP_LOOP_and_9_nl = COMP_LOOP_COMP_LOOP_and_147_itm & mux_2771_m1c;
  assign COMP_LOOP_and_10_nl = COMP_LOOP_COMP_LOOP_and_148_itm & mux_2771_m1c;
  assign COMP_LOOP_and_11_nl = COMP_LOOP_COMP_LOOP_and_149_itm & mux_2771_m1c;
  assign nand_2_nl = ~((fsm_output[5]) & mux_125_cse);
  assign mux_126_nl = MUX_s_1_2_2(nand_2_nl, or_tmp_68, fsm_output[2]);
  assign or_92_nl = (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[7])) |
      (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_127_nl = MUX_s_1_2_2(mux_126_nl, or_92_nl, fsm_output[9]);
  assign nand_3_nl = ~((fsm_output[4]) & (~ mux_127_nl));
  assign or_91_nl = (fsm_output[2]) | (~ (fsm_output[5])) | (fsm_output[7]) | mux_tmp_119;
  assign or_89_nl = (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[7])) |
      (fsm_output[3]) | (fsm_output[8]) | (~ (fsm_output[6])) | (fsm_output[10]);
  assign mux_123_nl = MUX_s_1_2_2(or_91_nl, or_89_nl, fsm_output[9]);
  assign or_88_nl = (fsm_output[9]) | (~((fsm_output[2]) & (fsm_output[5]) & (fsm_output[7])
      & (fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]) & (fsm_output[10])));
  assign mux_124_nl = MUX_s_1_2_2(mux_123_nl, or_88_nl, fsm_output[4]);
  assign mux_128_nl = MUX_s_1_2_2(nand_3_nl, mux_124_nl, fsm_output[1]);
  assign or_87_nl = (fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[7])) | (~
      (fsm_output[3])) | (fsm_output[8]) | not_tmp_49;
  assign or_85_nl = (~ (fsm_output[2])) | (~ (fsm_output[5])) | (fsm_output[7]) |
      mux_tmp_119;
  assign mux_120_nl = MUX_s_1_2_2(or_87_nl, or_85_nl, fsm_output[9]);
  assign or_81_nl = (fsm_output[9]) | (fsm_output[2]) | (fsm_output[5]) | (~ (fsm_output[7]))
      | (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) | (fsm_output[10]);
  assign mux_121_nl = MUX_s_1_2_2(mux_120_nl, or_81_nl, fsm_output[4]);
  assign or_79_nl = (~ (fsm_output[2])) | (fsm_output[5]) | (~ (fsm_output[7])) |
      (fsm_output[3]) | (~ (fsm_output[8])) | (fsm_output[6]) | (~ (fsm_output[10]));
  assign nand_373_nl = ~((fsm_output[5]) & (fsm_output[7]) & (fsm_output[3]) & (fsm_output[8])
      & (fsm_output[6]) & (~ (fsm_output[10])));
  assign mux_116_nl = MUX_s_1_2_2(nand_373_nl, or_tmp_68, fsm_output[2]);
  assign mux_117_nl = MUX_s_1_2_2(or_79_nl, mux_116_nl, fsm_output[9]);
  assign mux_118_nl = MUX_s_1_2_2(or_80_cse, mux_117_nl, fsm_output[4]);
  assign mux_122_nl = MUX_s_1_2_2(mux_121_nl, mux_118_nl, fsm_output[1]);
  assign mux_129_nl = MUX_s_1_2_2(mux_128_nl, mux_122_nl, fsm_output[0]);
  assign mux_2975_nl = MUX_s_1_2_2(mux_2203_cse, mux_tmp_2159, fsm_output[6]);
  assign mux_2976_nl = MUX_s_1_2_2(mux_2975_nl, mux_tmp_2920, fsm_output[0]);
  assign mux_2973_nl = MUX_s_1_2_2(or_tmp_2280, or_tmp_2729, fsm_output[6]);
  assign mux_2972_nl = MUX_s_1_2_2(or_tmp_2731, or_tmp_2729, fsm_output[6]);
  assign mux_2974_nl = MUX_s_1_2_2(mux_2973_nl, mux_2972_nl, fsm_output[0]);
  assign mux_2977_nl = MUX_s_1_2_2(mux_2976_nl, mux_2974_nl, fsm_output[8]);
  assign mux_2971_nl = MUX_s_1_2_2(mux_tmp_2879, or_tmp_2734, fsm_output[8]);
  assign mux_2978_nl = MUX_s_1_2_2(mux_2977_nl, mux_2971_nl, fsm_output[3]);
  assign mux_2967_nl = MUX_s_1_2_2(or_tmp_2749, mux_tmp_2912, fsm_output[6]);
  assign mux_2968_nl = MUX_s_1_2_2(mux_2967_nl, nand_tmp_71, fsm_output[0]);
  assign mux_2969_nl = MUX_s_1_2_2(mux_2968_nl, or_3532_cse, fsm_output[8]);
  assign mux_2963_nl = MUX_s_1_2_2((~ (fsm_output[10])), or_tmp_2276, fsm_output[9]);
  assign mux_2964_nl = MUX_s_1_2_2(mux_2963_nl, or_tmp_2731, fsm_output[6]);
  assign mux_2965_nl = MUX_s_1_2_2(mux_2964_nl, mux_tmp_2906, fsm_output[0]);
  assign mux_2966_nl = MUX_s_1_2_2(or_tmp_2740, mux_2965_nl, fsm_output[8]);
  assign mux_2970_nl = MUX_s_1_2_2(mux_2969_nl, mux_2966_nl, fsm_output[3]);
  assign mux_2979_nl = MUX_s_1_2_2(mux_2978_nl, mux_2970_nl, fsm_output[5]);
  assign or_2810_nl = (fsm_output[6]) | mux_tmp_2848;
  assign mux_2960_nl = MUX_s_1_2_2(nand_tmp_69, or_2810_nl, fsm_output[8]);
  assign nand_72_nl = ~((fsm_output[6]) & (~ mux_tmp_2895));
  assign mux_2959_nl = MUX_s_1_2_2(nand_72_nl, or_tmp_2743, fsm_output[8]);
  assign mux_2961_nl = MUX_s_1_2_2(mux_2960_nl, mux_2959_nl, fsm_output[3]);
  assign mux_2956_nl = MUX_s_1_2_2(mux_tmp_2867, mux_tmp_2890, fsm_output[0]);
  assign mux_2955_nl = MUX_s_1_2_2(mux_tmp_2862, mux_tmp_2888, fsm_output[0]);
  assign mux_2957_nl = MUX_s_1_2_2(mux_2956_nl, mux_2955_nl, fsm_output[8]);
  assign mux_2953_nl = MUX_s_1_2_2(mux_tmp_2850, mux_tmp_2886, fsm_output[0]);
  assign mux_2954_nl = MUX_s_1_2_2(mux_tmp_2878, mux_2953_nl, fsm_output[8]);
  assign mux_2958_nl = MUX_s_1_2_2(mux_2957_nl, mux_2954_nl, fsm_output[3]);
  assign mux_2962_nl = MUX_s_1_2_2(mux_2961_nl, mux_2958_nl, fsm_output[5]);
  assign mux_2980_nl = MUX_s_1_2_2(mux_2979_nl, mux_2962_nl, fsm_output[4]);
  assign or_2809_nl = (fsm_output[6]) | mux_tmp_2851;
  assign mux_2948_nl = MUX_s_1_2_2(or_2809_nl, or_tmp_2734, fsm_output[0]);
  assign mux_2949_nl = MUX_s_1_2_2(mux_tmp_2880, mux_2948_nl, fsm_output[8]);
  assign mux_2946_nl = MUX_s_1_2_2(mux_tmp_2916, mux_tmp_2876, fsm_output[0]);
  assign mux_2947_nl = MUX_s_1_2_2(mux_2946_nl, or_tmp_2734, fsm_output[8]);
  assign mux_2950_nl = MUX_s_1_2_2(mux_2949_nl, mux_2947_nl, fsm_output[3]);
  assign mux_2944_nl = MUX_s_1_2_2(nand_tmp_70, mux_tmp_2910, fsm_output[8]);
  assign mux_2942_nl = MUX_s_1_2_2(or_tmp_258, mux_tmp_2159, fsm_output[6]);
  assign mux_2943_nl = MUX_s_1_2_2(or_tmp_2740, mux_2942_nl, fsm_output[8]);
  assign mux_2945_nl = MUX_s_1_2_2(mux_2944_nl, mux_2943_nl, fsm_output[3]);
  assign mux_2951_nl = MUX_s_1_2_2(mux_2950_nl, mux_2945_nl, fsm_output[5]);
  assign mux_2938_nl = MUX_s_1_2_2(nand_tmp_69, nand_tmp_67, fsm_output[0]);
  assign mux_2936_nl = MUX_s_1_2_2(or_tmp_2731, or_tmp_2749, fsm_output[6]);
  assign mux_2937_nl = MUX_s_1_2_2(or_tmp_2745, mux_2936_nl, fsm_output[0]);
  assign mux_2939_nl = MUX_s_1_2_2(mux_2938_nl, mux_2937_nl, fsm_output[8]);
  assign mux_2933_nl = MUX_s_1_2_2(or_tmp_2746, mux_tmp_2856, fsm_output[6]);
  assign mux_2934_nl = MUX_s_1_2_2(nand_tmp_68, mux_2933_nl, fsm_output[0]);
  assign mux_2935_nl = MUX_s_1_2_2(mux_2934_nl, or_3532_cse, fsm_output[8]);
  assign mux_2940_nl = MUX_s_1_2_2(mux_2939_nl, mux_2935_nl, fsm_output[3]);
  assign mux_2930_nl = MUX_s_1_2_2(mux_tmp_2159, or_tmp_2736, fsm_output[6]);
  assign mux_2931_nl = MUX_s_1_2_2(mux_2930_nl, mux_tmp_2888, fsm_output[8]);
  assign mux_2927_nl = MUX_s_1_2_2((~ (fsm_output[7])), mux_2926_cse, fsm_output[9]);
  assign or_2807_nl = (fsm_output[6]) | mux_2927_nl;
  assign mux_2928_nl = MUX_s_1_2_2(or_2807_nl, or_tmp_2734, fsm_output[0]);
  assign mux_2929_nl = MUX_s_1_2_2(mux_2928_nl, mux_tmp_2844, fsm_output[8]);
  assign mux_2932_nl = MUX_s_1_2_2(mux_2931_nl, mux_2929_nl, fsm_output[3]);
  assign mux_2941_nl = MUX_s_1_2_2(mux_2940_nl, mux_2932_nl, fsm_output[5]);
  assign mux_2952_nl = MUX_s_1_2_2(mux_2951_nl, mux_2941_nl, fsm_output[4]);
  assign mux_2981_nl = MUX_s_1_2_2(mux_2980_nl, mux_2952_nl, fsm_output[2]);
  assign mux_2921_nl = MUX_s_1_2_2(mux_tmp_2920, or_tmp_2734, fsm_output[8]);
  assign mux_2917_nl = MUX_s_1_2_2(mux_tmp_2856, mux_tmp_2851, fsm_output[6]);
  assign mux_2918_nl = MUX_s_1_2_2(mux_2917_nl, mux_tmp_2916, fsm_output[0]);
  assign mux_2919_nl = MUX_s_1_2_2(mux_2918_nl, or_tmp_2734, fsm_output[8]);
  assign mux_2922_nl = MUX_s_1_2_2(mux_2921_nl, mux_2919_nl, fsm_output[3]);
  assign mux_2913_nl = MUX_s_1_2_2(nand_tmp_71, nand_tmp_70, fsm_output[0]);
  assign mux_2911_nl = MUX_s_1_2_2(or_3532_cse, mux_tmp_2910, fsm_output[0]);
  assign mux_2914_nl = MUX_s_1_2_2(mux_2913_nl, mux_2911_nl, fsm_output[8]);
  assign mux_2905_nl = MUX_s_1_2_2(or_tmp_258, mux_tmp_2851, fsm_output[6]);
  assign mux_2907_nl = MUX_s_1_2_2(mux_tmp_2906, mux_2905_nl, fsm_output[0]);
  assign mux_2908_nl = MUX_s_1_2_2(or_tmp_2740, mux_2907_nl, fsm_output[8]);
  assign mux_2915_nl = MUX_s_1_2_2(mux_2914_nl, mux_2908_nl, fsm_output[3]);
  assign mux_2923_nl = MUX_s_1_2_2(mux_2922_nl, mux_2915_nl, fsm_output[5]);
  assign mux_2899_nl = MUX_s_1_2_2(or_tmp_2742, or_tmp_2746, fsm_output[6]);
  assign mux_2900_nl = MUX_s_1_2_2(mux_2899_nl, or_tmp_2745, fsm_output[0]);
  assign mux_2902_nl = MUX_s_1_2_2(nand_tmp_69, mux_2900_nl, fsm_output[8]);
  assign mux_2896_nl = MUX_s_1_2_2(or_tmp_2739, mux_tmp_2895, fsm_output[6]);
  assign mux_2897_nl = MUX_s_1_2_2(mux_2896_nl, nand_tmp_68, fsm_output[0]);
  assign mux_2894_nl = MUX_s_1_2_2(or_tmp_2743, or_3532_cse, fsm_output[0]);
  assign mux_2898_nl = MUX_s_1_2_2(mux_2897_nl, mux_2894_nl, fsm_output[8]);
  assign mux_2903_nl = MUX_s_1_2_2(mux_2902_nl, mux_2898_nl, fsm_output[3]);
  assign mux_2889_nl = MUX_s_1_2_2(or_tmp_2731, or_tmp_2281, fsm_output[6]);
  assign mux_2891_nl = MUX_s_1_2_2(mux_tmp_2890, mux_2889_nl, fsm_output[0]);
  assign mux_2892_nl = MUX_s_1_2_2(mux_2891_nl, mux_tmp_2888, fsm_output[8]);
  assign mux_2887_nl = MUX_s_1_2_2(or_tmp_2734, mux_tmp_2886, fsm_output[8]);
  assign mux_2893_nl = MUX_s_1_2_2(mux_2892_nl, mux_2887_nl, fsm_output[3]);
  assign mux_2904_nl = MUX_s_1_2_2(mux_2903_nl, mux_2893_nl, fsm_output[5]);
  assign mux_2924_nl = MUX_s_1_2_2(mux_2923_nl, mux_2904_nl, fsm_output[4]);
  assign mux_2881_nl = MUX_s_1_2_2(mux_tmp_2880, mux_tmp_2879, fsm_output[0]);
  assign mux_2882_nl = MUX_s_1_2_2(mux_2881_nl, mux_tmp_2878, fsm_output[8]);
  assign mux_2873_nl = MUX_s_1_2_2(mux_tmp_2848, or_tmp_2739, fsm_output[6]);
  assign mux_2874_nl = MUX_s_1_2_2(or_tmp_2734, mux_2873_nl, fsm_output[0]);
  assign mux_2877_nl = MUX_s_1_2_2(mux_tmp_2876, mux_2874_nl, fsm_output[8]);
  assign mux_2883_nl = MUX_s_1_2_2(mux_2882_nl, mux_2877_nl, fsm_output[3]);
  assign mux_2869_nl = MUX_s_1_2_2((~ or_tmp_2280), or_tmp_2276, fsm_output[9]);
  assign mux_2870_nl = MUX_s_1_2_2(mux_2869_nl, or_tmp_2280, fsm_output[6]);
  assign mux_2871_nl = MUX_s_1_2_2(or_tmp_2740, mux_2870_nl, fsm_output[8]);
  assign mux_2864_nl = MUX_s_1_2_2(or_tmp_2276, mux_tmp_2863, fsm_output[6]);
  assign mux_2865_nl = MUX_s_1_2_2(mux_2864_nl, mux_tmp_2862, fsm_output[0]);
  assign mux_2868_nl = MUX_s_1_2_2(mux_tmp_2867, mux_2865_nl, fsm_output[8]);
  assign mux_2872_nl = MUX_s_1_2_2(mux_2871_nl, mux_2868_nl, fsm_output[3]);
  assign mux_2884_nl = MUX_s_1_2_2(mux_2883_nl, mux_2872_nl, fsm_output[5]);
  assign or_2797_nl = (fsm_output[6]) | or_tmp_2731;
  assign mux_2859_nl = MUX_s_1_2_2(nand_tmp_67, or_2797_nl, fsm_output[8]);
  assign nand_66_nl = ~((fsm_output[6]) & (~ mux_tmp_2856));
  assign mux_2857_nl = MUX_s_1_2_2(nand_66_nl, or_3532_cse, fsm_output[8]);
  assign mux_2860_nl = MUX_s_1_2_2(mux_2859_nl, mux_2857_nl, fsm_output[3]);
  assign mux_2852_nl = MUX_s_1_2_2(mux_tmp_2851, or_tmp_2736, fsm_output[6]);
  assign mux_2853_nl = MUX_s_1_2_2(mux_2852_nl, or_tmp_2734, fsm_output[0]);
  assign mux_2854_nl = MUX_s_1_2_2(mux_2853_nl, mux_tmp_2850, fsm_output[8]);
  assign mux_2842_nl = MUX_s_1_2_2(or_tmp_2729, mux_tmp_2841, fsm_output[6]);
  assign mux_2845_nl = MUX_s_1_2_2(mux_tmp_2844, mux_2842_nl, fsm_output[0]);
  assign mux_2847_nl = MUX_s_1_2_2(or_tmp_2734, mux_2845_nl, fsm_output[8]);
  assign mux_2855_nl = MUX_s_1_2_2(mux_2854_nl, mux_2847_nl, fsm_output[3]);
  assign mux_2861_nl = MUX_s_1_2_2(mux_2860_nl, mux_2855_nl, fsm_output[5]);
  assign mux_2885_nl = MUX_s_1_2_2(mux_2884_nl, mux_2861_nl, fsm_output[4]);
  assign mux_2925_nl = MUX_s_1_2_2(mux_2924_nl, mux_2885_nl, fsm_output[2]);
  assign COMP_LOOP_COMP_LOOP_and_17_nl = (z_out_2_12_1[3:0]==4'b0011);
  assign nl_COMP_LOOP_1_acc_8_nl = tmp_10_lpi_4_dfm - COMP_LOOP_10_mul_mut;
  assign COMP_LOOP_1_acc_8_nl = nl_COMP_LOOP_1_acc_8_nl[63:0];
  assign nor_631_nl = ~((~ (fsm_output[3])) | (~ (fsm_output[0])) | (~ (fsm_output[1]))
      | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[10]));
  assign mux_3284_nl = MUX_s_1_2_2(or_2921_cse, mux_3935_cse, fsm_output[0]);
  assign nor_632_nl = ~((fsm_output[3]) | mux_3284_nl);
  assign mux_3285_nl = MUX_s_1_2_2(nor_631_nl, nor_632_nl, fsm_output[8]);
  assign and_417_nl = (fsm_output[8]) & (fsm_output[3]) & (~ mux_3245_cse);
  assign mux_3286_nl = MUX_s_1_2_2(mux_3285_nl, and_417_nl, fsm_output[5]);
  assign or_2958_nl = (fsm_output[9]) | (~ (fsm_output[2])) | (fsm_output[6]) | (fsm_output[10]);
  assign or_2957_nl = (~ (fsm_output[9])) | (~ (fsm_output[2])) | (fsm_output[6])
      | (fsm_output[10]);
  assign mux_3279_nl = MUX_s_1_2_2(or_2958_nl, or_2957_nl, fsm_output[1]);
  assign or_2959_nl = (fsm_output[0]) | mux_3279_nl;
  assign or_2954_nl = (fsm_output[1]) | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[6])
      | (~ (fsm_output[10]));
  assign mux_3278_nl = MUX_s_1_2_2(or_2912_cse, or_2954_nl, fsm_output[0]);
  assign mux_3280_nl = MUX_s_1_2_2(or_2959_nl, mux_3278_nl, fsm_output[3]);
  assign nor_633_nl = ~((~ (fsm_output[5])) | (fsm_output[8]) | mux_3280_nl);
  assign mux_3287_nl = MUX_s_1_2_2(mux_3286_nl, nor_633_nl, fsm_output[4]);
  assign and_418_nl = (fsm_output[8]) & (fsm_output[3]) & (fsm_output[0]) & (fsm_output[1])
      & (~ (fsm_output[9])) & (fsm_output[2]) & (fsm_output[6]) & (~ (fsm_output[10]));
  assign nor_634_nl = ~((fsm_output[8]) | (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1])
      | (fsm_output[9]) | (fsm_output[2]) | (fsm_output[6]) | (~ (fsm_output[10])));
  assign mux_3276_nl = MUX_s_1_2_2(and_418_nl, nor_634_nl, fsm_output[5]);
  assign nand_92_nl = ~((fsm_output[3]) & (~ mux_3254_cse));
  assign or_2943_nl = (fsm_output[1]) | (fsm_output[9]) | nand_367_cse;
  assign mux_3273_nl = MUX_s_1_2_2(or_2905_cse, or_2943_nl, fsm_output[0]);
  assign or_2945_nl = (fsm_output[3]) | mux_3273_nl;
  assign mux_3275_nl = MUX_s_1_2_2(nand_92_nl, or_2945_nl, fsm_output[8]);
  assign nor_635_nl = ~((fsm_output[5]) | mux_3275_nl);
  assign mux_3277_nl = MUX_s_1_2_2(mux_3276_nl, nor_635_nl, fsm_output[4]);
  assign mux_3288_nl = MUX_s_1_2_2(mux_3287_nl, mux_3277_nl, fsm_output[7]);
  assign COMP_LOOP_COMP_LOOP_and_10_nl = (VEC_LOOP_j_sva_11_0[3:0]==4'b1011);
  assign nl_COMP_LOOP_1_acc_nl = ({(z_out_1[5:0]) , 4'b0000}) + ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:1]))})
      + 10'b0000000001;
  assign COMP_LOOP_1_acc_nl = nl_COMP_LOOP_1_acc_nl[9:0];
  assign or_2647_nl = (fsm_output[7:6]!=2'b00);
  assign mux_2642_nl = MUX_s_1_2_2(nor_609_cse, and_757_cse, or_2647_nl);
  assign mux_3330_nl = MUX_s_1_2_2(mux_tmp_3329, mux_2642_nl, or_3388_cse);
  assign mux_3331_nl = MUX_s_1_2_2(mux_3330_nl, mux_2643_cse, fsm_output[3]);
  assign or_3032_nl = (fsm_output[1]) | (fsm_output[6]);
  assign mux_3326_nl = MUX_s_1_2_2(mux_tmp_2640, and_756_cse, or_3032_nl);
  assign and_410_nl = ((~((~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[6])))
      | (fsm_output[7])) & (fsm_output[10:9]==2'b11);
  assign mux_3327_nl = MUX_s_1_2_2(mux_3326_nl, and_410_nl, fsm_output[3]);
  assign mux_3332_nl = MUX_s_1_2_2(mux_3331_nl, mux_3327_nl, fsm_output[4]);
  assign and_411_nl = ((~((~ (fsm_output[3])) | (fsm_output[6]))) | (fsm_output[7]))
      & (fsm_output[10:9]==2'b11);
  assign mux_3325_nl = MUX_s_1_2_2(mux_2643_cse, and_411_nl, fsm_output[4]);
  assign mux_3333_nl = MUX_s_1_2_2(mux_3332_nl, mux_3325_nl, fsm_output[2]);
  assign mux_3334_nl = MUX_s_1_2_2(mux_tmp_3329, mux_3333_nl, fsm_output[5]);
  assign or_3037_nl = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[2]) | (fsm_output[9]);
  assign mux_3337_nl = MUX_s_1_2_2((fsm_output[9]), or_3037_nl, and_407_cse);
  assign and_408_nl = (fsm_output[0]) & (fsm_output[1]) & (fsm_output[2]) & (fsm_output[9]);
  assign or_3036_nl = (fsm_output[5:3]!=3'b000);
  assign mux_3336_nl = MUX_s_1_2_2(and_408_nl, (fsm_output[9]), or_3036_nl);
  assign mux_3338_nl = MUX_s_1_2_2((~ mux_3337_nl), mux_3336_nl, fsm_output[7]);
  assign mux_3339_nl = MUX_s_1_2_2(mux_3338_nl, and_458_cse, fsm_output[6]);
  assign mux_3340_nl = MUX_s_1_2_2(mux_3339_nl, (fsm_output[9]), fsm_output[8]);
  assign mux_3346_nl = MUX_s_1_2_2(mux_tmp_3341, nor_tmp_457, fsm_output[3]);
  assign mux_3347_nl = MUX_s_1_2_2(not_tmp_90, mux_3346_nl, fsm_output[4]);
  assign mux_3344_nl = MUX_s_1_2_2(not_tmp_90, nor_tmp_457, fsm_output[4]);
  assign mux_3345_nl = MUX_s_1_2_2(mux_3344_nl, mux_tmp_3343, fsm_output[0]);
  assign mux_3348_nl = MUX_s_1_2_2(mux_3347_nl, mux_3345_nl, fsm_output[1]);
  assign mux_3349_nl = MUX_s_1_2_2(mux_3348_nl, mux_tmp_3343, fsm_output[2]);
  assign mux_3350_nl = MUX_s_1_2_2(not_tmp_90, mux_3349_nl, fsm_output[5]);
  assign nl_COMP_LOOP_acc_11_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b001});
  assign nor_623_nl = ~((fsm_output[5]) | (fsm_output[8]));
  assign mux_3351_nl = MUX_s_1_2_2(nor_623_nl, (fsm_output[8]), fsm_output[6]);
  assign mux_3353_nl = MUX_s_1_2_2(mux_648_cse, mux_3351_nl, or_3039_cse);
  assign mux_3354_nl = MUX_s_1_2_2(mux_648_cse, mux_3353_nl, fsm_output[4]);
  assign mux_3355_nl = MUX_s_1_2_2(mux_3354_nl, (fsm_output[8]), fsm_output[7]);
  assign and_401_nl = (fsm_output[0]) & (fsm_output[7]) & (fsm_output[8]);
  assign mux_3356_nl = MUX_s_1_2_2(not_tmp_133, and_401_nl, fsm_output[3]);
  assign and_402_nl = (fsm_output[3]) & (fsm_output[7]) & (fsm_output[8]);
  assign mux_3357_nl = MUX_s_1_2_2(mux_3356_nl, and_402_nl, or_2368_cse);
  assign mux_3358_nl = MUX_s_1_2_2(not_tmp_133, mux_3357_nl, and_407_cse);
  assign mux_3359_nl = MUX_s_1_2_2(mux_3358_nl, and_404_cse, fsm_output[6]);
  assign or_3045_nl = (fsm_output[8:6]!=3'b000) | mux_tmp_3361;
  assign mux_3362_nl = MUX_s_1_2_2(or_3079_cse, or_3045_nl, fsm_output[4]);
  assign mux_3360_nl = MUX_s_1_2_2(or_3079_cse, or_3074_cse, fsm_output[4]);
  assign mux_3363_nl = MUX_s_1_2_2(mux_3362_nl, mux_3360_nl, fsm_output[1]);
  assign mux_3364_nl = MUX_s_1_2_2(mux_3363_nl, (~ or_3074_cse), fsm_output[9]);
  assign nl_COMP_LOOP_acc_14_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b011});
  assign or_3048_nl = (or_3039_cse & (fsm_output[4])) | (fsm_output[9]);
  assign mux_3365_nl = MUX_s_1_2_2((fsm_output[9]), or_3048_nl, fsm_output[5]);
  assign nor_621_nl = ~((fsm_output[7]) | mux_3365_nl);
  assign and_334_nl = (fsm_output[7]) & (fsm_output[5]) & (and_459_cse | (fsm_output[4]))
      & (fsm_output[9]);
  assign mux_3366_nl = MUX_s_1_2_2(nor_621_nl, and_334_nl, fsm_output[6]);
  assign mux_3367_nl = MUX_s_1_2_2(mux_3366_nl, (fsm_output[9]), fsm_output[8]);
  assign nl_COMP_LOOP_acc_1_cse_8_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b0111});
  assign nor_619_nl = ~((fsm_output[9:8]!=2'b00));
  assign nor_620_nl = ~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[8])
      | (fsm_output[9]));
  assign mux_3370_nl = MUX_s_1_2_2(nor_619_nl, nor_620_nl, and_407_cse);
  assign and_30_nl = (fsm_output[8]) & (fsm_output[2]) & or_3388_cse & (fsm_output[9]);
  assign mux_3368_nl = MUX_s_1_2_2(and_30_nl, nor_tmp_82, fsm_output[3]);
  assign and_337_nl = (fsm_output[4]) & mux_3368_nl;
  assign mux_3369_nl = MUX_s_1_2_2(and_337_nl, nor_tmp_82, fsm_output[5]);
  assign mux_3371_nl = MUX_s_1_2_2(mux_3370_nl, mux_3369_nl, fsm_output[6]);
  assign mux_3372_nl = MUX_s_1_2_2(mux_3371_nl, nor_tmp_82, fsm_output[7]);
  assign nor_1596_nl = ~((fsm_output[9:7]!=3'b000));
  assign nor_1597_nl = ~((fsm_output[3]) | (fsm_output[1]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[9]));
  assign and_749_nl = (fsm_output[3]) & (fsm_output[7]) & (fsm_output[8]) & (fsm_output[9]);
  assign mux_3373_nl = MUX_s_1_2_2(nor_1597_nl, and_749_nl, fsm_output[2]);
  assign mux_3374_nl = MUX_s_1_2_2(nor_1596_nl, mux_3373_nl, and_407_cse);
  assign and_750_nl = (fsm_output[9:7]==3'b111);
  assign mux_3375_nl = MUX_s_1_2_2(mux_3374_nl, and_750_nl, fsm_output[6]);
  assign nl_COMP_LOOP_acc_1_cse_10_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1001});
  assign or_3060_nl = (~((fsm_output[9:6]!=4'b0000))) | (fsm_output[10]);
  assign mux_3379_nl = MUX_s_1_2_2(mux_tmp_3378, or_3060_nl, fsm_output[4]);
  assign or_3058_nl = (fsm_output[4]) | (fsm_output[6]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[9]);
  assign mux_3376_nl = MUX_s_1_2_2((~ (fsm_output[10])), (fsm_output[10]), or_3058_nl);
  assign mux_3377_nl = MUX_s_1_2_2(mux_3376_nl, or_tmp_2988, fsm_output[0]);
  assign mux_3380_nl = MUX_s_1_2_2(mux_3379_nl, mux_3377_nl, fsm_output[1]);
  assign mux_3381_nl = MUX_s_1_2_2(mux_3380_nl, or_tmp_2988, or_2644_cse);
  assign nl_COMP_LOOP_acc_17_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b101});
  assign or_3065_nl = (fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[10]);
  assign mux_3384_nl = MUX_s_1_2_2((fsm_output[10]), or_3065_nl, and_407_cse);
  assign and_394_nl = or_2368_cse & (fsm_output[3]) & (fsm_output[10]);
  assign mux_3383_nl = MUX_s_1_2_2(and_394_nl, (fsm_output[10]), or_3063_cse);
  assign mux_3385_nl = MUX_s_1_2_2((~ mux_3384_nl), mux_3383_nl, fsm_output[7]);
  assign mux_3386_nl = MUX_s_1_2_2(mux_3385_nl, and_395_cse, fsm_output[6]);
  assign nl_COMP_LOOP_acc_1_cse_12_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1011});
  assign nor_615_nl = ~((fsm_output[7]) | (fsm_output[10]));
  assign mux_3388_nl = MUX_s_1_2_2(nor_615_nl, and_395_cse, fsm_output[6]);
  assign mux_3389_nl = MUX_s_1_2_2(not_tmp_647, mux_3388_nl, fsm_output[0]);
  assign and_391_nl = (fsm_output[6]) & (fsm_output[7]) & (fsm_output[10]);
  assign mux_3390_nl = MUX_s_1_2_2(mux_3389_nl, and_391_nl, or_3039_cse);
  assign mux_3391_nl = MUX_s_1_2_2(not_tmp_647, mux_3390_nl, and_407_cse);
  assign nor_613_nl = ~((fsm_output[8]) | (fsm_output[10]));
  assign nor_614_nl = ~((fsm_output[1]) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[8])
      | (fsm_output[10]));
  assign mux_3394_nl = MUX_s_1_2_2(nor_613_nl, nor_614_nl, and_407_cse);
  assign and_388_nl = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[8]) & (fsm_output[10]);
  assign mux_3393_nl = MUX_s_1_2_2(and_388_nl, nor_tmp_405, fsm_output[5]);
  assign mux_3395_nl = MUX_s_1_2_2(mux_3394_nl, mux_3393_nl, fsm_output[6]);
  assign mux_3396_nl = MUX_s_1_2_2(mux_3395_nl, nor_tmp_405, fsm_output[7]);
  assign nl_COMP_LOOP_acc_1_cse_14_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1101});
  assign nor_611_nl = ~((fsm_output[7]) | (fsm_output[8]) | (fsm_output[10]));
  assign nor_612_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[7]) | (fsm_output[8])
      | (fsm_output[10]));
  assign and_384_nl = (fsm_output[2]) & (fsm_output[3]) & (fsm_output[0]) & (fsm_output[7])
      & (fsm_output[8]) & (fsm_output[10]);
  assign mux_3398_nl = MUX_s_1_2_2(nor_612_nl, and_384_nl, fsm_output[1]);
  assign mux_3399_nl = MUX_s_1_2_2(nor_611_nl, mux_3398_nl, and_407_cse);
  assign and_386_nl = (fsm_output[7]) & (fsm_output[8]) & (fsm_output[10]);
  assign mux_3400_nl = MUX_s_1_2_2(mux_3399_nl, and_386_nl, fsm_output[6]);
  assign nl_COMP_LOOP_acc_20_psp_sva  = (VEC_LOOP_j_sva_11_0[11:1]) + conv_u2u_8_11({COMP_LOOP_k_9_4_sva_4_0
      , 3'b111});
  assign or_3078_nl = (or_3039_cse & (fsm_output[5])) | (fsm_output[8:6]!=3'b000);
  assign mux_3403_nl = MUX_s_1_2_2(or_3079_cse, or_3078_nl, fsm_output[4]);
  assign nor_1680_nl = ~((fsm_output[10]) | mux_3403_nl);
  assign or_3076_nl = ((and_529_cse | (fsm_output[3])) & (fsm_output[5])) | (fsm_output[8:6]!=3'b000);
  assign mux_3402_nl = MUX_s_1_2_2(or_3076_nl, or_3074_cse, fsm_output[4]);
  assign and_1162_nl = (fsm_output[10]) & mux_3402_nl;
  assign nl_COMP_LOOP_acc_1_cse_sva  = VEC_LOOP_j_sva_11_0 + conv_u2u_9_12({COMP_LOOP_k_9_4_sva_4_0
      , 4'b1111});
  assign nor_610_nl = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[9])
      | (fsm_output[10]));
  assign mux_3406_nl = MUX_s_1_2_2(nor_609_cse, nor_610_nl, and_407_cse);
  assign and_341_nl = (fsm_output[3:2]==2'b11) & or_3388_cse & (fsm_output[10:9]==2'b11);
  assign mux_3405_nl = MUX_s_1_2_2(and_341_nl, and_757_cse, or_3063_cse);
  assign mux_3407_nl = MUX_s_1_2_2(mux_3406_nl, mux_3405_nl, fsm_output[7]);
  assign mux_3408_nl = MUX_s_1_2_2(mux_3407_nl, and_756_cse, fsm_output[6]);
  assign operator_64_false_1_mux_2_nl = MUX_v_12_2_2(({7'b0000001 , (~ COMP_LOOP_k_9_4_sva_4_0)}),
      VEC_LOOP_j_sva_11_0, and_dcpl_332);
  assign operator_64_false_1_mux_3_nl = MUX_v_10_2_2(10'b0000000001, STAGE_LOOP_lshift_psp_sva,
      and_dcpl_332);
  assign nl_z_out = conv_u2u_12_13(operator_64_false_1_mux_2_nl) + conv_u2u_10_13(operator_64_false_1_mux_3_nl);
  assign z_out = nl_z_out[12:0];
  assign COMP_LOOP_COMP_LOOP_or_72_nl = (~(and_dcpl_342 | and_dcpl_356)) | and_dcpl_350
      | and_dcpl_359;
  assign COMP_LOOP_COMP_LOOP_or_73_nl = (~((operator_66_true_div_cmp_z[63]) | and_dcpl_342
      | and_dcpl_356)) | and_dcpl_350;
  assign COMP_LOOP_mux1h_575_nl = MUX1HOT_v_63_4_2(({54'b000000000000000000000000000000000000000000000000000000
      , (VEC_LOOP_j_sva_11_0[11:3])}), (~ (operator_64_false_acc_mut_63_0[62:0])),
      ({58'b0000000000000000000000000000000000000000000000000000000000 , COMP_LOOP_k_9_4_sva_4_0}),
      (~ (operator_66_true_div_cmp_z[62:0])), {and_dcpl_342 , and_dcpl_350 , and_dcpl_356
      , and_dcpl_359});
  assign COMP_LOOP_nor_695_nl = ~(and_dcpl_350 | and_dcpl_356 | and_dcpl_359);
  assign COMP_LOOP_COMP_LOOP_and_938_nl = MUX_v_5_2_2(5'b00000, COMP_LOOP_k_9_4_sva_4_0,
      COMP_LOOP_nor_695_nl);
  assign nl_z_out_1 = ({COMP_LOOP_COMP_LOOP_or_72_nl , COMP_LOOP_COMP_LOOP_or_73_nl
      , COMP_LOOP_mux1h_575_nl}) + conv_u2u_6_65({COMP_LOOP_COMP_LOOP_and_938_nl
      , 1'b1});
  assign z_out_1 = nl_z_out_1[64:0];
  assign COMP_LOOP_mux1h_576_nl = MUX1HOT_v_7_4_2(({(z_out_7[5:0]) , (STAGE_LOOP_lshift_psp_sva[3])}),
      (z_out_5[9:3]), (z_out_4[9:3]), z_out_7, {and_824_ssc , COMP_LOOP_or_54_ssc
      , COMP_LOOP_or_55_ssc , and_872_ssc});
  assign COMP_LOOP_or_69_nl = and_824_ssc | and_872_ssc;
  assign COMP_LOOP_mux1h_577_nl = MUX1HOT_v_3_3_2((STAGE_LOOP_lshift_psp_sva[2:0]),
      (z_out_5[2:0]), (z_out_4[2:0]), {COMP_LOOP_or_69_nl , COMP_LOOP_or_54_ssc ,
      COMP_LOOP_or_55_ssc});
  assign nl_COMP_LOOP_acc_105_nl = conv_u2u_12_13(VEC_LOOP_j_sva_11_0) + conv_u2u_10_13({COMP_LOOP_mux1h_576_nl
      , COMP_LOOP_mux1h_577_nl});
  assign COMP_LOOP_acc_105_nl = nl_COMP_LOOP_acc_105_nl[12:0];
  assign z_out_2_12_1 = readslicef_13_12_1(COMP_LOOP_acc_105_nl);
  assign COMP_LOOP_COMP_LOOP_or_74_nl = (VEC_LOOP_j_sva_11_0[11]) | and_dcpl_460
      | and_dcpl_468 | and_dcpl_475 | and_dcpl_481 | and_dcpl_486 | and_dcpl_495
      | and_dcpl_500 | and_dcpl_503 | and_dcpl_507 | and_dcpl_510 | and_dcpl_513;
  assign COMP_LOOP_COMP_LOOP_mux_18_nl = MUX_v_9_2_2((VEC_LOOP_j_sva_11_0[10:2]),
      (~ (STAGE_LOOP_lshift_psp_sva[9:1])), COMP_LOOP_or_61_itm);
  assign COMP_LOOP_or_70_nl = (~ and_dcpl_453) | and_dcpl_460 | and_dcpl_468 | and_dcpl_475
      | and_dcpl_481 | and_dcpl_486 | and_dcpl_495 | and_dcpl_500 | and_dcpl_503
      | and_dcpl_507 | and_dcpl_510 | and_dcpl_513;
  assign COMP_LOOP_COMP_LOOP_mux_19_nl = MUX_v_5_2_2(({2'b00 , (COMP_LOOP_k_9_4_sva_4_0[4:2])}),
      COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_61_itm);
  assign COMP_LOOP_COMP_LOOP_or_75_nl = ((COMP_LOOP_k_9_4_sva_4_0[1]) & (~(and_dcpl_460
      | and_dcpl_468 | and_dcpl_475 | and_dcpl_481 | and_dcpl_486))) | and_dcpl_495
      | and_dcpl_500 | and_dcpl_503 | and_dcpl_507 | and_dcpl_510 | and_dcpl_513;
  assign COMP_LOOP_COMP_LOOP_or_76_nl = ((COMP_LOOP_k_9_4_sva_4_0[0]) & (~(and_dcpl_460
      | and_dcpl_468 | and_dcpl_495 | and_dcpl_500 | and_dcpl_503))) | and_dcpl_475
      | and_dcpl_481 | and_dcpl_486 | and_dcpl_507 | and_dcpl_510 | and_dcpl_513;
  assign COMP_LOOP_COMP_LOOP_or_77_nl = (~(and_dcpl_453 | and_dcpl_460 | and_dcpl_475
      | and_dcpl_481 | and_dcpl_495 | and_dcpl_500 | and_dcpl_507 | and_dcpl_510))
      | and_dcpl_468 | and_dcpl_486 | and_dcpl_503 | and_dcpl_513;
  assign COMP_LOOP_COMP_LOOP_or_78_nl = (~(and_dcpl_468 | and_dcpl_475 | and_dcpl_486
      | and_dcpl_495 | and_dcpl_503 | and_dcpl_507 | and_dcpl_513)) | and_dcpl_453
      | and_dcpl_460 | and_dcpl_481 | and_dcpl_500 | and_dcpl_510;
  assign nl_acc_3_nl = ({COMP_LOOP_COMP_LOOP_or_74_nl , COMP_LOOP_COMP_LOOP_mux_18_nl
      , COMP_LOOP_or_70_nl}) + conv_u2u_10_11({COMP_LOOP_COMP_LOOP_mux_19_nl , COMP_LOOP_COMP_LOOP_or_75_nl
      , COMP_LOOP_COMP_LOOP_or_76_nl , COMP_LOOP_COMP_LOOP_or_77_nl , COMP_LOOP_COMP_LOOP_or_78_nl
      , 1'b1});
  assign acc_3_nl = nl_acc_3_nl[10:0];
  assign z_out_3 = readslicef_11_10_1(acc_3_nl);
  assign COMP_LOOP_mux_82_nl = MUX_v_10_2_2((VEC_LOOP_j_sva_11_0[11:2]), STAGE_LOOP_lshift_psp_sva,
      COMP_LOOP_or_24_itm);
  assign COMP_LOOP_COMP_LOOP_mux_20_nl = MUX_v_5_2_2(({2'b00 , (COMP_LOOP_k_9_4_sva_4_0[4:2])}),
      COMP_LOOP_k_9_4_sva_4_0, COMP_LOOP_or_24_itm);
  assign COMP_LOOP_COMP_LOOP_or_79_nl = ((COMP_LOOP_k_9_4_sva_4_0[1]) & (~(and_dcpl_531
      | and_dcpl_540))) | and_dcpl_544 | and_dcpl_553 | and_dcpl_557 | and_dcpl_561;
  assign COMP_LOOP_COMP_LOOP_or_80_nl = ((COMP_LOOP_k_9_4_sva_4_0[0]) & (~(and_dcpl_544
      | and_dcpl_553))) | and_dcpl_531 | and_dcpl_540 | and_dcpl_557 | and_dcpl_561;
  assign COMP_LOOP_COMP_LOOP_or_81_nl = (~(and_dcpl_531 | and_dcpl_544 | and_dcpl_557
      | and_dcpl_561)) | and_978_ssc | and_dcpl_540 | and_dcpl_553;
  assign COMP_LOOP_COMP_LOOP_or_82_nl = (~(and_dcpl_531 | and_dcpl_557)) | and_978_ssc
      | and_dcpl_540 | and_dcpl_544 | and_dcpl_553 | and_dcpl_561;
  assign nl_z_out_4 = COMP_LOOP_mux_82_nl + conv_u2u_9_10({COMP_LOOP_COMP_LOOP_mux_20_nl
      , COMP_LOOP_COMP_LOOP_or_79_nl , COMP_LOOP_COMP_LOOP_or_80_nl , COMP_LOOP_COMP_LOOP_or_81_nl
      , COMP_LOOP_COMP_LOOP_or_82_nl});
  assign z_out_4 = nl_z_out_4[9:0];
  assign and_1178_nl = and_dcpl_569 & and_dcpl_567 & and_827_cse & and_825_cse;
  assign and_1179_nl = and_dcpl_569 & and_dcpl_383 & and_835_cse & (~ (fsm_output[6]))
      & (~ (fsm_output[0]));
  assign and_1180_nl = and_dcpl_472 & (~ (fsm_output[10])) & and_dcpl_114 & (fsm_output[8])
      & and_dcpl_371 & (fsm_output[1]) & (~ (fsm_output[6])) & (fsm_output[0]);
  assign and_1181_nl = and_dcpl_594 & and_dcpl_114 & (~ (fsm_output[8])) & (fsm_output[4])
      & (~ (fsm_output[7])) & (~ (fsm_output[1])) & and_825_cse;
  assign and_1182_nl = and_dcpl_594 & and_dcpl_567 & and_827_cse & and_815_cse;
  assign and_1183_nl = and_dcpl_568 & (fsm_output[10]) & and_dcpl_338 & and_835_cse
      & and_815_cse;
  assign and_1184_nl = and_dcpl_472 & (fsm_output[10]) & and_dcpl_383 & (fsm_output[4])
      & (fsm_output[7]) & (~ (fsm_output[1])) & and_815_cse;
  assign COMP_LOOP_mux1h_578_nl = MUX1HOT_v_4_7_2(4'b0001, 4'b0010, 4'b0011, 4'b0101,
      4'b0110, 4'b1010, 4'b1110, {and_1178_nl , and_1179_nl , and_1180_nl , and_1181_nl
      , and_1182_nl , and_1183_nl , and_1184_nl});
  assign and_1185_nl = (~ (fsm_output[2])) & (fsm_output[9]) & (fsm_output[10]) &
      and_dcpl_338 & and_dcpl_344 & (fsm_output[1]) & and_825_cse;
  assign COMP_LOOP_or_71_nl = MUX_v_4_2_2(COMP_LOOP_mux1h_578_nl, 4'b1111, and_1185_nl);
  assign nl_z_out_5 = STAGE_LOOP_lshift_psp_sva + conv_u2u_9_10({COMP_LOOP_k_9_4_sva_4_0
      , COMP_LOOP_or_71_nl});
  assign z_out_5 = nl_z_out_5[9:0];
  assign COMP_LOOP_COMP_LOOP_or_83_nl = ((p_sva[63]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_84_nl = ((p_sva[62]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_85_nl = ((p_sva[61]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_86_nl = ((p_sva[60]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_87_nl = ((p_sva[59]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_88_nl = ((p_sva[58]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_89_nl = ((p_sva[57]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_90_nl = ((p_sva[56]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_91_nl = ((p_sva[55]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_92_nl = ((p_sva[54]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_93_nl = ((p_sva[53]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_94_nl = ((p_sva[52]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_95_nl = ((p_sva[51]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_96_nl = ((p_sva[50]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_97_nl = ((p_sva[49]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_98_nl = ((p_sva[48]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_99_nl = ((p_sva[47]) & COMP_LOOP_nor_633_itm) | not_tmp_838
      | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_100_nl = ((p_sva[46]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_101_nl = ((p_sva[45]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_102_nl = ((p_sva[44]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_103_nl = ((p_sva[43]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_104_nl = ((p_sva[42]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_105_nl = ((p_sva[41]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_106_nl = ((p_sva[40]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_107_nl = ((p_sva[39]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_108_nl = ((p_sva[38]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_109_nl = ((p_sva[37]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_110_nl = ((p_sva[36]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_111_nl = ((p_sva[35]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_112_nl = ((p_sva[34]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_113_nl = ((p_sva[33]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_114_nl = ((p_sva[32]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_115_nl = ((p_sva[31]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_116_nl = ((p_sva[30]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_117_nl = ((p_sva[29]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_118_nl = ((p_sva[28]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_119_nl = ((p_sva[27]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_120_nl = ((p_sva[26]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_121_nl = ((p_sva[25]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_122_nl = ((p_sva[24]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_123_nl = ((p_sva[23]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_124_nl = ((p_sva[22]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_125_nl = ((p_sva[21]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_126_nl = ((p_sva[20]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_127_nl = ((p_sva[19]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_128_nl = ((p_sva[18]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_129_nl = ((p_sva[17]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_130_nl = ((p_sva[16]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_131_nl = ((p_sva[15]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_132_nl = ((p_sva[14]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_133_nl = ((p_sva[13]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_134_nl = ((p_sva[12]) & COMP_LOOP_nor_633_itm) |
      not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_mux_83_nl = MUX_v_4_2_2((VEC_LOOP_j_sva_11_0[11:8]), (p_sva[11:8]),
      and_dcpl_647);
  assign COMP_LOOP_and_398_nl = MUX_v_4_2_2(4'b0000, COMP_LOOP_mux_83_nl, COMP_LOOP_nor_685_itm);
  assign COMP_LOOP_or_72_nl = not_tmp_838 | and_dcpl_650;
  assign COMP_LOOP_COMP_LOOP_or_135_nl = MUX_v_4_2_2(COMP_LOOP_and_398_nl, 4'b1111,
      COMP_LOOP_or_72_nl);
  assign COMP_LOOP_mux1h_579_nl = MUX1HOT_s_1_4_2((VEC_LOOP_j_sva_11_0[7]), (~ modExp_exp_1_7_1_sva),
      (p_sva[7]), (~ COMP_LOOP_nor_134_itm), {and_dcpl_628 , not_tmp_838 , and_dcpl_647
      , and_dcpl_650});
  assign COMP_LOOP_or_73_nl = COMP_LOOP_mux1h_579_nl | and_dcpl_636 | and_dcpl_642;
  assign COMP_LOOP_mux1h_580_nl = MUX1HOT_v_7_5_2((VEC_LOOP_j_sva_11_0[6:0]), (~
      (STAGE_LOOP_lshift_psp_sva[9:3])), ({(~ modExp_exp_1_6_1_sva) , (~ modExp_exp_1_5_1_sva)
      , (~ modExp_exp_1_4_1_sva) , (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) , (~
      COMP_LOOP_nor_137_itm) , (~ COMP_LOOP_nor_134_itm) , (~ COMP_LOOP_nor_12_itm)}),
      (p_sva[6:0]), ({(~ modExp_exp_1_7_1_sva) , (~ modExp_exp_1_6_1_sva) , (~ modExp_exp_1_5_1_sva)
      , (~ modExp_exp_1_4_1_sva) , (~ COMP_LOOP_slc_COMP_LOOP_acc_12_7_itm) , (~
      COMP_LOOP_nor_137_itm) , (~ COMP_LOOP_nor_12_itm)}), {and_dcpl_628 , COMP_LOOP_or_65_itm
      , not_tmp_838 , and_dcpl_647 , and_dcpl_650});
  assign COMP_LOOP_or_74_nl = (~(and_dcpl_628 | not_tmp_838 | and_dcpl_647 | and_dcpl_650))
      | and_dcpl_636 | and_dcpl_642;
  assign COMP_LOOP_COMP_LOOP_or_136_nl = (~(and_dcpl_628 | and_dcpl_636 | and_dcpl_642
      | not_tmp_838 | and_dcpl_650)) | and_dcpl_647;
  assign COMP_LOOP_COMP_LOOP_or_137_nl = ((COMP_LOOP_k_9_4_sva_4_0[4]) & COMP_LOOP_nor_687_itm)
      | and_dcpl_647;
  assign COMP_LOOP_COMP_LOOP_or_138_nl = ((COMP_LOOP_k_9_4_sva_4_0[3]) & COMP_LOOP_nor_687_itm)
      | and_dcpl_647;
  assign COMP_LOOP_COMP_LOOP_mux_21_nl = MUX_v_3_2_2((COMP_LOOP_k_9_4_sva_4_0[2:0]),
      (COMP_LOOP_k_9_4_sva_4_0[4:2]), COMP_LOOP_or_65_itm);
  assign COMP_LOOP_nor_706_nl = ~(not_tmp_838 | and_dcpl_650);
  assign COMP_LOOP_and_401_nl = MUX_v_3_2_2(3'b000, COMP_LOOP_COMP_LOOP_mux_21_nl,
      COMP_LOOP_nor_706_nl);
  assign COMP_LOOP_or_75_nl = MUX_v_3_2_2(COMP_LOOP_and_401_nl, 3'b111, and_dcpl_647);
  assign COMP_LOOP_nor_707_nl = ~(and_dcpl_628 | not_tmp_838 | and_dcpl_650);
  assign COMP_LOOP_and_402_nl = MUX_v_2_2_2(2'b00, (COMP_LOOP_k_9_4_sva_4_0[1:0]),
      COMP_LOOP_nor_707_nl);
  assign COMP_LOOP_COMP_LOOP_or_139_nl = MUX_v_2_2_2(COMP_LOOP_and_402_nl, 2'b11,
      and_dcpl_647);
  assign COMP_LOOP_COMP_LOOP_or_140_nl = (~(and_dcpl_636 | not_tmp_838 | and_dcpl_650))
      | and_dcpl_628 | and_dcpl_642 | and_dcpl_647;
  assign COMP_LOOP_COMP_LOOP_or_141_nl = COMP_LOOP_nor_685_itm | and_dcpl_628 | not_tmp_838
      | and_dcpl_647 | and_dcpl_650;
  assign nl_acc_6_nl = conv_u2u_65_66({COMP_LOOP_COMP_LOOP_or_83_nl , COMP_LOOP_COMP_LOOP_or_84_nl
      , COMP_LOOP_COMP_LOOP_or_85_nl , COMP_LOOP_COMP_LOOP_or_86_nl , COMP_LOOP_COMP_LOOP_or_87_nl
      , COMP_LOOP_COMP_LOOP_or_88_nl , COMP_LOOP_COMP_LOOP_or_89_nl , COMP_LOOP_COMP_LOOP_or_90_nl
      , COMP_LOOP_COMP_LOOP_or_91_nl , COMP_LOOP_COMP_LOOP_or_92_nl , COMP_LOOP_COMP_LOOP_or_93_nl
      , COMP_LOOP_COMP_LOOP_or_94_nl , COMP_LOOP_COMP_LOOP_or_95_nl , COMP_LOOP_COMP_LOOP_or_96_nl
      , COMP_LOOP_COMP_LOOP_or_97_nl , COMP_LOOP_COMP_LOOP_or_98_nl , COMP_LOOP_COMP_LOOP_or_99_nl
      , COMP_LOOP_COMP_LOOP_or_100_nl , COMP_LOOP_COMP_LOOP_or_101_nl , COMP_LOOP_COMP_LOOP_or_102_nl
      , COMP_LOOP_COMP_LOOP_or_103_nl , COMP_LOOP_COMP_LOOP_or_104_nl , COMP_LOOP_COMP_LOOP_or_105_nl
      , COMP_LOOP_COMP_LOOP_or_106_nl , COMP_LOOP_COMP_LOOP_or_107_nl , COMP_LOOP_COMP_LOOP_or_108_nl
      , COMP_LOOP_COMP_LOOP_or_109_nl , COMP_LOOP_COMP_LOOP_or_110_nl , COMP_LOOP_COMP_LOOP_or_111_nl
      , COMP_LOOP_COMP_LOOP_or_112_nl , COMP_LOOP_COMP_LOOP_or_113_nl , COMP_LOOP_COMP_LOOP_or_114_nl
      , COMP_LOOP_COMP_LOOP_or_115_nl , COMP_LOOP_COMP_LOOP_or_116_nl , COMP_LOOP_COMP_LOOP_or_117_nl
      , COMP_LOOP_COMP_LOOP_or_118_nl , COMP_LOOP_COMP_LOOP_or_119_nl , COMP_LOOP_COMP_LOOP_or_120_nl
      , COMP_LOOP_COMP_LOOP_or_121_nl , COMP_LOOP_COMP_LOOP_or_122_nl , COMP_LOOP_COMP_LOOP_or_123_nl
      , COMP_LOOP_COMP_LOOP_or_124_nl , COMP_LOOP_COMP_LOOP_or_125_nl , COMP_LOOP_COMP_LOOP_or_126_nl
      , COMP_LOOP_COMP_LOOP_or_127_nl , COMP_LOOP_COMP_LOOP_or_128_nl , COMP_LOOP_COMP_LOOP_or_129_nl
      , COMP_LOOP_COMP_LOOP_or_130_nl , COMP_LOOP_COMP_LOOP_or_131_nl , COMP_LOOP_COMP_LOOP_or_132_nl
      , COMP_LOOP_COMP_LOOP_or_133_nl , COMP_LOOP_COMP_LOOP_or_134_nl , COMP_LOOP_COMP_LOOP_or_135_nl
      , COMP_LOOP_or_73_nl , COMP_LOOP_mux1h_580_nl , COMP_LOOP_or_74_nl}) + conv_s2u_11_66({COMP_LOOP_COMP_LOOP_or_136_nl
      , COMP_LOOP_COMP_LOOP_or_137_nl , COMP_LOOP_COMP_LOOP_or_138_nl , COMP_LOOP_or_75_nl
      , COMP_LOOP_COMP_LOOP_or_139_nl , COMP_LOOP_COMP_LOOP_or_140_nl , COMP_LOOP_COMP_LOOP_or_141_nl
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[65:0];
  assign z_out_6 = readslicef_66_65_1(acc_6_nl);
  assign COMP_LOOP_COMP_LOOP_or_142_nl = ((STAGE_LOOP_lshift_psp_sva[9]) & (~(and_dcpl_669
      | and_dcpl_678))) | and_dcpl_660;
  assign COMP_LOOP_mux1h_581_nl = MUX1HOT_v_6_4_2((~ (STAGE_LOOP_lshift_psp_sva[9:4])),
      ({1'b1 , (~ (STAGE_LOOP_lshift_psp_sva[9:5]))}), (STAGE_LOOP_lshift_psp_sva[9:4]),
      (STAGE_LOOP_lshift_psp_sva[8:3]), {and_dcpl_660 , and_dcpl_669 , and_dcpl_678
      , and_dcpl_686});
  assign COMP_LOOP_or_76_nl = (~(and_dcpl_678 | and_dcpl_686)) | and_dcpl_660 | and_dcpl_669;
  assign COMP_LOOP_or_77_nl = and_dcpl_669 | and_dcpl_678;
  assign COMP_LOOP_COMP_LOOP_mux_22_nl = MUX_v_5_2_2(COMP_LOOP_k_9_4_sva_4_0, ({1'b0
      , (COMP_LOOP_k_9_4_sva_4_0[4:1])}), COMP_LOOP_or_77_nl);
  assign COMP_LOOP_COMP_LOOP_or_143_nl = ((COMP_LOOP_k_9_4_sva_4_0[0]) & (~ and_dcpl_660))
      | and_dcpl_686;
  assign nl_acc_7_nl = ({COMP_LOOP_COMP_LOOP_or_142_nl , COMP_LOOP_mux1h_581_nl ,
      COMP_LOOP_or_76_nl}) + conv_u2u_7_8({COMP_LOOP_COMP_LOOP_mux_22_nl , COMP_LOOP_COMP_LOOP_or_143_nl
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[7:0];
  assign z_out_7 = readslicef_8_7_1(acc_7_nl);
  assign mux_3950_nl = MUX_s_1_2_2(or_tmp_3307, or_tmp_3326, fsm_output[0]);
  assign or_3639_nl = (~ (fsm_output[8])) | (fsm_output[6]) | mux_3950_nl;
  assign or_3640_nl = (fsm_output[8]) | (fsm_output[6]) | (~ (fsm_output[0])) | (fsm_output[9])
      | (fsm_output[10]) | (~ (fsm_output[1])) | (fsm_output[2]);
  assign mux_3949_nl = MUX_s_1_2_2(or_3639_nl, or_3640_nl, fsm_output[3]);
  assign nor_1711_nl = ~((fsm_output[4]) | mux_3949_nl);
  assign mux_3952_nl = MUX_s_1_2_2(or_tmp_3326, or_tmp_3312, fsm_output[0]);
  assign and_1186_nl = (fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]) & (~ mux_3952_nl);
  assign or_3641_nl = (fsm_output[10]) | (fsm_output[1]) | (~ (fsm_output[2]));
  assign or_3642_nl = (fsm_output[10]) | (~ and_529_cse);
  assign mux_3954_nl = MUX_s_1_2_2(or_3641_nl, or_3642_nl, fsm_output[9]);
  assign nor_1712_nl = ~((fsm_output[8]) | (fsm_output[6]) | (fsm_output[0]) | mux_3954_nl);
  assign nand_428_nl = ~((fsm_output[9]) & (fsm_output[10]) & (~ (fsm_output[1]))
      & (fsm_output[2]));
  assign or_3643_nl = (fsm_output[9]) | (~ (fsm_output[10])) | (fsm_output[1]) |
      (fsm_output[2]);
  assign mux_3955_nl = MUX_s_1_2_2(nand_428_nl, or_3643_nl, fsm_output[0]);
  assign nor_1713_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_3955_nl);
  assign mux_3953_nl = MUX_s_1_2_2(nor_1712_nl, nor_1713_nl, fsm_output[3]);
  assign mux_3951_nl = MUX_s_1_2_2(and_1186_nl, mux_3953_nl, fsm_output[4]);
  assign mux_3948_nl = MUX_s_1_2_2(nor_1711_nl, mux_3951_nl, fsm_output[5]);
  assign and_1187_nl = (fsm_output[3]) & (fsm_output[8]) & (fsm_output[6]) & (fsm_output[0])
      & (~ (fsm_output[9])) & (~ (fsm_output[10])) & and_529_cse;
  assign or_3644_nl = (fsm_output[9]) | (~ (fsm_output[10])) | (fsm_output[1]) |
      (~ (fsm_output[2]));
  assign mux_3959_nl = MUX_s_1_2_2(or_tmp_3312, or_3644_nl, fsm_output[0]);
  assign and_1188_nl = (fsm_output[8]) & (fsm_output[6]) & (~ mux_3959_nl);
  assign or_3645_nl = (fsm_output[9]) | (fsm_output[10]) | (~ (fsm_output[1])) |
      (fsm_output[2]);
  assign mux_3960_nl = MUX_s_1_2_2(or_3645_nl, or_tmp_3307, fsm_output[0]);
  assign nor_1714_nl = ~((fsm_output[8]) | (fsm_output[6]) | mux_3960_nl);
  assign mux_3958_nl = MUX_s_1_2_2(and_1188_nl, nor_1714_nl, fsm_output[3]);
  assign mux_3957_nl = MUX_s_1_2_2(and_1187_nl, mux_3958_nl, fsm_output[4]);
  assign mux_3956_nl = MUX_s_1_2_2(mux_3957_nl, nor_1657_cse, fsm_output[5]);
  assign mux_3947_nl = MUX_s_1_2_2(mux_3948_nl, mux_3956_nl, fsm_output[7]);
  assign modExp_while_if_mux_1_nl = MUX_v_64_2_2(modExp_result_sva, COMP_LOOP_10_mul_mut,
      mux_3947_nl);
  assign nl_z_out_8 = $signed(conv_u2s_64_65(modExp_while_if_mux_1_nl)) * $signed(COMP_LOOP_10_mul_mut);
  assign z_out_8 = nl_z_out_8[63:0];

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_6_2;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [5:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    result = result | ( input_3 & {4{sel[3]}});
    result = result | ( input_4 & {4{sel[4]}});
    result = result | ( input_5 & {4{sel[5]}});
    result = result | ( input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [62:0] MUX1HOT_v_63_4_2;
    input [62:0] input_3;
    input [62:0] input_2;
    input [62:0] input_1;
    input [62:0] input_0;
    input [3:0] sel;
    reg [62:0] result;
  begin
    result = input_0 & {63{sel[0]}};
    result = result | ( input_1 & {63{sel[1]}});
    result = result | ( input_2 & {63{sel[2]}});
    result = result | ( input_3 & {63{sel[3]}});
    MUX1HOT_v_63_4_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_17_2;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [16:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    MUX1HOT_v_64_17_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_21_2;
    input [63:0] input_20;
    input [63:0] input_19;
    input [63:0] input_18;
    input [63:0] input_17;
    input [63:0] input_16;
    input [63:0] input_15;
    input [63:0] input_14;
    input [63:0] input_13;
    input [63:0] input_12;
    input [63:0] input_11;
    input [63:0] input_10;
    input [63:0] input_9;
    input [63:0] input_8;
    input [63:0] input_7;
    input [63:0] input_6;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [20:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    result = result | ( input_6 & {64{sel[6]}});
    result = result | ( input_7 & {64{sel[7]}});
    result = result | ( input_8 & {64{sel[8]}});
    result = result | ( input_9 & {64{sel[9]}});
    result = result | ( input_10 & {64{sel[10]}});
    result = result | ( input_11 & {64{sel[11]}});
    result = result | ( input_12 & {64{sel[12]}});
    result = result | ( input_13 & {64{sel[13]}});
    result = result | ( input_14 & {64{sel[14]}});
    result = result | ( input_15 & {64{sel[15]}});
    result = result | ( input_16 & {64{sel[16]}});
    result = result | ( input_17 & {64{sel[17]}});
    result = result | ( input_18 & {64{sel[18]}});
    result = result | ( input_19 & {64{sel[19]}});
    result = result | ( input_20 & {64{sel[20]}});
    MUX1HOT_v_64_21_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_3_2;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [2:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    MUX1HOT_v_64_3_2 = result;
  end
  endfunction


  function automatic [63:0] MUX1HOT_v_64_6_2;
    input [63:0] input_5;
    input [63:0] input_4;
    input [63:0] input_3;
    input [63:0] input_2;
    input [63:0] input_1;
    input [63:0] input_0;
    input [5:0] sel;
    reg [63:0] result;
  begin
    result = input_0 & {64{sel[0]}};
    result = result | ( input_1 & {64{sel[1]}});
    result = result | ( input_2 & {64{sel[2]}});
    result = result | ( input_3 & {64{sel[3]}});
    result = result | ( input_4 & {64{sel[4]}});
    result = result | ( input_5 & {64{sel[5]}});
    MUX1HOT_v_64_6_2 = result;
  end
  endfunction


  function automatic [64:0] MUX1HOT_v_65_3_2;
    input [64:0] input_2;
    input [64:0] input_1;
    input [64:0] input_0;
    input [2:0] sel;
    reg [64:0] result;
  begin
    result = input_0 & {65{sel[0]}};
    result = result | ( input_1 & {65{sel[1]}});
    result = result | ( input_2 & {65{sel[2]}});
    MUX1HOT_v_65_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_5_2;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [4:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    result = result | ( input_4 & {7{sel[4]}});
    MUX1HOT_v_7_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_19_2;
    input [7:0] input_18;
    input [7:0] input_17;
    input [7:0] input_16;
    input [7:0] input_15;
    input [7:0] input_14;
    input [7:0] input_13;
    input [7:0] input_12;
    input [7:0] input_11;
    input [7:0] input_10;
    input [7:0] input_9;
    input [7:0] input_8;
    input [7:0] input_7;
    input [7:0] input_6;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [18:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | ( input_1 & {8{sel[1]}});
    result = result | ( input_2 & {8{sel[2]}});
    result = result | ( input_3 & {8{sel[3]}});
    result = result | ( input_4 & {8{sel[4]}});
    result = result | ( input_5 & {8{sel[5]}});
    result = result | ( input_6 & {8{sel[6]}});
    result = result | ( input_7 & {8{sel[7]}});
    result = result | ( input_8 & {8{sel[8]}});
    result = result | ( input_9 & {8{sel[9]}});
    result = result | ( input_10 & {8{sel[10]}});
    result = result | ( input_11 & {8{sel[11]}});
    result = result | ( input_12 & {8{sel[12]}});
    result = result | ( input_13 & {8{sel[13]}});
    result = result | ( input_14 & {8{sel[14]}});
    result = result | ( input_15 & {8{sel[15]}});
    result = result | ( input_16 & {8{sel[16]}});
    result = result | ( input_17 & {8{sel[17]}});
    result = result | ( input_18 & {8{sel[18]}});
    MUX1HOT_v_8_19_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [0:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input [0:0] sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [62:0] MUX_v_63_2_2;
    input [62:0] input_0;
    input [62:0] input_1;
    input [0:0] sel;
    reg [62:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_63_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [64:0] MUX_v_65_2_2;
    input [64:0] input_0;
    input [64:0] input_1;
    input [0:0] sel;
    reg [64:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_65_2_2 = result;
  end
  endfunction


  function automatic [8:0] MUX_v_9_2_2;
    input [8:0] input_0;
    input [8:0] input_1;
    input [0:0] sel;
    reg [8:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_9_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_10_1_9;
    input [9:0] vector;
    reg [9:0] tmp;
  begin
    tmp = vector >> 9;
    readslicef_10_1_9 = tmp[0:0];
  end
  endfunction


  function automatic [9:0] readslicef_11_10_1;
    input [10:0] vector;
    reg [10:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_11_10_1 = tmp[9:0];
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [64:0] readslicef_66_65_1;
    input [65:0] vector;
    reg [65:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_66_65_1 = tmp[64:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [65:0] conv_s2u_11_66 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_66 = {{55{vector[10]}}, vector};
  end
  endfunction


  function automatic [64:0] conv_u2s_64_65 ;
    input [63:0]  vector ;
  begin
    conv_u2s_64_65 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_5_8 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_8 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [64:0] conv_u2u_6_65 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_65 = {{59{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_8_11 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_11 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_9_10 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_10 = {1'b0, vector};
  end
  endfunction


  function automatic [11:0] conv_u2u_9_12 ;
    input [8:0]  vector ;
  begin
    conv_u2u_9_12 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [10:0] conv_u2u_10_11 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_11 = {1'b0, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_10_13 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_13 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [12:0] conv_u2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_u2u_12_13 = {1'b0, vector};
  end
  endfunction


  function automatic [65:0] conv_u2u_65_66 ;
    input [64:0]  vector ;
  begin
    conv_u2u_65_66 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    inPlaceNTT_DIT
// ------------------------------------------------------------------


module inPlaceNTT_DIT (
  clk, rst, vec_rsc_0_0_adra, vec_rsc_0_0_da, vec_rsc_0_0_wea, vec_rsc_0_0_qa, vec_rsc_triosy_0_0_lz,
      vec_rsc_0_1_adra, vec_rsc_0_1_da, vec_rsc_0_1_wea, vec_rsc_0_1_qa, vec_rsc_triosy_0_1_lz,
      vec_rsc_0_2_adra, vec_rsc_0_2_da, vec_rsc_0_2_wea, vec_rsc_0_2_qa, vec_rsc_triosy_0_2_lz,
      vec_rsc_0_3_adra, vec_rsc_0_3_da, vec_rsc_0_3_wea, vec_rsc_0_3_qa, vec_rsc_triosy_0_3_lz,
      vec_rsc_0_4_adra, vec_rsc_0_4_da, vec_rsc_0_4_wea, vec_rsc_0_4_qa, vec_rsc_triosy_0_4_lz,
      vec_rsc_0_5_adra, vec_rsc_0_5_da, vec_rsc_0_5_wea, vec_rsc_0_5_qa, vec_rsc_triosy_0_5_lz,
      vec_rsc_0_6_adra, vec_rsc_0_6_da, vec_rsc_0_6_wea, vec_rsc_0_6_qa, vec_rsc_triosy_0_6_lz,
      vec_rsc_0_7_adra, vec_rsc_0_7_da, vec_rsc_0_7_wea, vec_rsc_0_7_qa, vec_rsc_triosy_0_7_lz,
      vec_rsc_0_8_adra, vec_rsc_0_8_da, vec_rsc_0_8_wea, vec_rsc_0_8_qa, vec_rsc_triosy_0_8_lz,
      vec_rsc_0_9_adra, vec_rsc_0_9_da, vec_rsc_0_9_wea, vec_rsc_0_9_qa, vec_rsc_triosy_0_9_lz,
      vec_rsc_0_10_adra, vec_rsc_0_10_da, vec_rsc_0_10_wea, vec_rsc_0_10_qa, vec_rsc_triosy_0_10_lz,
      vec_rsc_0_11_adra, vec_rsc_0_11_da, vec_rsc_0_11_wea, vec_rsc_0_11_qa, vec_rsc_triosy_0_11_lz,
      vec_rsc_0_12_adra, vec_rsc_0_12_da, vec_rsc_0_12_wea, vec_rsc_0_12_qa, vec_rsc_triosy_0_12_lz,
      vec_rsc_0_13_adra, vec_rsc_0_13_da, vec_rsc_0_13_wea, vec_rsc_0_13_qa, vec_rsc_triosy_0_13_lz,
      vec_rsc_0_14_adra, vec_rsc_0_14_da, vec_rsc_0_14_wea, vec_rsc_0_14_qa, vec_rsc_triosy_0_14_lz,
      vec_rsc_0_15_adra, vec_rsc_0_15_da, vec_rsc_0_15_wea, vec_rsc_0_15_qa, vec_rsc_triosy_0_15_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_dat, r_rsc_triosy_lz
);
  input clk;
  input rst;
  output [7:0] vec_rsc_0_0_adra;
  output [63:0] vec_rsc_0_0_da;
  output vec_rsc_0_0_wea;
  input [63:0] vec_rsc_0_0_qa;
  output vec_rsc_triosy_0_0_lz;
  output [7:0] vec_rsc_0_1_adra;
  output [63:0] vec_rsc_0_1_da;
  output vec_rsc_0_1_wea;
  input [63:0] vec_rsc_0_1_qa;
  output vec_rsc_triosy_0_1_lz;
  output [7:0] vec_rsc_0_2_adra;
  output [63:0] vec_rsc_0_2_da;
  output vec_rsc_0_2_wea;
  input [63:0] vec_rsc_0_2_qa;
  output vec_rsc_triosy_0_2_lz;
  output [7:0] vec_rsc_0_3_adra;
  output [63:0] vec_rsc_0_3_da;
  output vec_rsc_0_3_wea;
  input [63:0] vec_rsc_0_3_qa;
  output vec_rsc_triosy_0_3_lz;
  output [7:0] vec_rsc_0_4_adra;
  output [63:0] vec_rsc_0_4_da;
  output vec_rsc_0_4_wea;
  input [63:0] vec_rsc_0_4_qa;
  output vec_rsc_triosy_0_4_lz;
  output [7:0] vec_rsc_0_5_adra;
  output [63:0] vec_rsc_0_5_da;
  output vec_rsc_0_5_wea;
  input [63:0] vec_rsc_0_5_qa;
  output vec_rsc_triosy_0_5_lz;
  output [7:0] vec_rsc_0_6_adra;
  output [63:0] vec_rsc_0_6_da;
  output vec_rsc_0_6_wea;
  input [63:0] vec_rsc_0_6_qa;
  output vec_rsc_triosy_0_6_lz;
  output [7:0] vec_rsc_0_7_adra;
  output [63:0] vec_rsc_0_7_da;
  output vec_rsc_0_7_wea;
  input [63:0] vec_rsc_0_7_qa;
  output vec_rsc_triosy_0_7_lz;
  output [7:0] vec_rsc_0_8_adra;
  output [63:0] vec_rsc_0_8_da;
  output vec_rsc_0_8_wea;
  input [63:0] vec_rsc_0_8_qa;
  output vec_rsc_triosy_0_8_lz;
  output [7:0] vec_rsc_0_9_adra;
  output [63:0] vec_rsc_0_9_da;
  output vec_rsc_0_9_wea;
  input [63:0] vec_rsc_0_9_qa;
  output vec_rsc_triosy_0_9_lz;
  output [7:0] vec_rsc_0_10_adra;
  output [63:0] vec_rsc_0_10_da;
  output vec_rsc_0_10_wea;
  input [63:0] vec_rsc_0_10_qa;
  output vec_rsc_triosy_0_10_lz;
  output [7:0] vec_rsc_0_11_adra;
  output [63:0] vec_rsc_0_11_da;
  output vec_rsc_0_11_wea;
  input [63:0] vec_rsc_0_11_qa;
  output vec_rsc_triosy_0_11_lz;
  output [7:0] vec_rsc_0_12_adra;
  output [63:0] vec_rsc_0_12_da;
  output vec_rsc_0_12_wea;
  input [63:0] vec_rsc_0_12_qa;
  output vec_rsc_triosy_0_12_lz;
  output [7:0] vec_rsc_0_13_adra;
  output [63:0] vec_rsc_0_13_da;
  output vec_rsc_0_13_wea;
  input [63:0] vec_rsc_0_13_qa;
  output vec_rsc_triosy_0_13_lz;
  output [7:0] vec_rsc_0_14_adra;
  output [63:0] vec_rsc_0_14_da;
  output vec_rsc_0_14_wea;
  input [63:0] vec_rsc_0_14_qa;
  output vec_rsc_triosy_0_14_lz;
  output [7:0] vec_rsc_0_15_adra;
  output [63:0] vec_rsc_0_15_da;
  output vec_rsc_0_15_wea;
  input [63:0] vec_rsc_0_15_qa;
  output vec_rsc_triosy_0_15_lz;
  input [63:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [63:0] r_rsc_dat;
  output r_rsc_triosy_lz;


  // Interconnect Declarations
  wire [63:0] vec_rsc_0_0_i_qa_d;
  wire vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_1_i_qa_d;
  wire vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_2_i_qa_d;
  wire vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_3_i_qa_d;
  wire vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_4_i_qa_d;
  wire vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_5_i_qa_d;
  wire vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_6_i_qa_d;
  wire vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_7_i_qa_d;
  wire vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_8_i_qa_d;
  wire vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_9_i_qa_d;
  wire vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_10_i_qa_d;
  wire vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_11_i_qa_d;
  wire vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_12_i_qa_d;
  wire vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_13_i_qa_d;
  wire vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_14_i_qa_d;
  wire vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [63:0] vec_rsc_0_15_i_qa_d;
  wire vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] vec_rsc_0_0_i_adra_d_iff;
  wire [63:0] vec_rsc_0_0_i_da_d_iff;
  wire vec_rsc_0_0_i_wea_d_iff;
  wire vec_rsc_0_1_i_wea_d_iff;
  wire vec_rsc_0_2_i_wea_d_iff;
  wire vec_rsc_0_3_i_wea_d_iff;
  wire vec_rsc_0_4_i_wea_d_iff;
  wire vec_rsc_0_5_i_wea_d_iff;
  wire vec_rsc_0_6_i_wea_d_iff;
  wire vec_rsc_0_7_i_wea_d_iff;
  wire vec_rsc_0_8_i_wea_d_iff;
  wire vec_rsc_0_9_i_wea_d_iff;
  wire vec_rsc_0_10_i_wea_d_iff;
  wire vec_rsc_0_11_i_wea_d_iff;
  wire vec_rsc_0_12_i_wea_d_iff;
  wire vec_rsc_0_13_i_wea_d_iff;
  wire vec_rsc_0_14_i_wea_d_iff;
  wire vec_rsc_0_15_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_4_8_64_256_256_64_1_gen vec_rsc_0_0_i
      (
      .qa(vec_rsc_0_0_qa),
      .wea(vec_rsc_0_0_wea),
      .da(vec_rsc_0_0_da),
      .adra(vec_rsc_0_0_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_0_i_qa_d),
      .wea_d(vec_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_0_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_5_8_64_256_256_64_1_gen vec_rsc_0_1_i
      (
      .qa(vec_rsc_0_1_qa),
      .wea(vec_rsc_0_1_wea),
      .da(vec_rsc_0_1_da),
      .adra(vec_rsc_0_1_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_1_i_qa_d),
      .wea_d(vec_rsc_0_1_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_1_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_6_8_64_256_256_64_1_gen vec_rsc_0_2_i
      (
      .qa(vec_rsc_0_2_qa),
      .wea(vec_rsc_0_2_wea),
      .da(vec_rsc_0_2_da),
      .adra(vec_rsc_0_2_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_2_i_qa_d),
      .wea_d(vec_rsc_0_2_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_2_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_7_8_64_256_256_64_1_gen vec_rsc_0_3_i
      (
      .qa(vec_rsc_0_3_qa),
      .wea(vec_rsc_0_3_wea),
      .da(vec_rsc_0_3_da),
      .adra(vec_rsc_0_3_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_3_i_qa_d),
      .wea_d(vec_rsc_0_3_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_3_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_8_8_64_256_256_64_1_gen vec_rsc_0_4_i
      (
      .qa(vec_rsc_0_4_qa),
      .wea(vec_rsc_0_4_wea),
      .da(vec_rsc_0_4_da),
      .adra(vec_rsc_0_4_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_4_i_qa_d),
      .wea_d(vec_rsc_0_4_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_4_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_9_8_64_256_256_64_1_gen vec_rsc_0_5_i
      (
      .qa(vec_rsc_0_5_qa),
      .wea(vec_rsc_0_5_wea),
      .da(vec_rsc_0_5_da),
      .adra(vec_rsc_0_5_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_5_i_qa_d),
      .wea_d(vec_rsc_0_5_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_5_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_10_8_64_256_256_64_1_gen
      vec_rsc_0_6_i (
      .qa(vec_rsc_0_6_qa),
      .wea(vec_rsc_0_6_wea),
      .da(vec_rsc_0_6_da),
      .adra(vec_rsc_0_6_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_6_i_qa_d),
      .wea_d(vec_rsc_0_6_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_6_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_11_8_64_256_256_64_1_gen
      vec_rsc_0_7_i (
      .qa(vec_rsc_0_7_qa),
      .wea(vec_rsc_0_7_wea),
      .da(vec_rsc_0_7_da),
      .adra(vec_rsc_0_7_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_7_i_qa_d),
      .wea_d(vec_rsc_0_7_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_7_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_12_8_64_256_256_64_1_gen
      vec_rsc_0_8_i (
      .qa(vec_rsc_0_8_qa),
      .wea(vec_rsc_0_8_wea),
      .da(vec_rsc_0_8_da),
      .adra(vec_rsc_0_8_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_8_i_qa_d),
      .wea_d(vec_rsc_0_8_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_8_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_13_8_64_256_256_64_1_gen
      vec_rsc_0_9_i (
      .qa(vec_rsc_0_9_qa),
      .wea(vec_rsc_0_9_wea),
      .da(vec_rsc_0_9_da),
      .adra(vec_rsc_0_9_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_9_i_qa_d),
      .wea_d(vec_rsc_0_9_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_9_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_14_8_64_256_256_64_1_gen
      vec_rsc_0_10_i (
      .qa(vec_rsc_0_10_qa),
      .wea(vec_rsc_0_10_wea),
      .da(vec_rsc_0_10_da),
      .adra(vec_rsc_0_10_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_10_i_qa_d),
      .wea_d(vec_rsc_0_10_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_10_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_15_8_64_256_256_64_1_gen
      vec_rsc_0_11_i (
      .qa(vec_rsc_0_11_qa),
      .wea(vec_rsc_0_11_wea),
      .da(vec_rsc_0_11_da),
      .adra(vec_rsc_0_11_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_11_i_qa_d),
      .wea_d(vec_rsc_0_11_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_11_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_16_8_64_256_256_64_1_gen
      vec_rsc_0_12_i (
      .qa(vec_rsc_0_12_qa),
      .wea(vec_rsc_0_12_wea),
      .da(vec_rsc_0_12_da),
      .adra(vec_rsc_0_12_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_12_i_qa_d),
      .wea_d(vec_rsc_0_12_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_12_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_17_8_64_256_256_64_1_gen
      vec_rsc_0_13_i (
      .qa(vec_rsc_0_13_qa),
      .wea(vec_rsc_0_13_wea),
      .da(vec_rsc_0_13_da),
      .adra(vec_rsc_0_13_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_13_i_qa_d),
      .wea_d(vec_rsc_0_13_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_13_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_18_8_64_256_256_64_1_gen
      vec_rsc_0_14_i (
      .qa(vec_rsc_0_14_qa),
      .wea(vec_rsc_0_14_wea),
      .da(vec_rsc_0_14_da),
      .adra(vec_rsc_0_14_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_14_i_qa_d),
      .wea_d(vec_rsc_0_14_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_14_i_wea_d_iff)
    );
  inPlaceNTT_DIT_Xilinx_RAMS_BLOCK_2R1W_RBW_DUAL_rwport_19_8_64_256_256_64_1_gen
      vec_rsc_0_15_i (
      .qa(vec_rsc_0_15_qa),
      .wea(vec_rsc_0_15_wea),
      .da(vec_rsc_0_15_da),
      .adra(vec_rsc_0_15_adra),
      .adra_d(vec_rsc_0_0_i_adra_d_iff),
      .da_d(vec_rsc_0_0_i_da_d_iff),
      .qa_d(vec_rsc_0_15_i_qa_d),
      .wea_d(vec_rsc_0_15_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(vec_rsc_0_15_i_wea_d_iff)
    );
  inPlaceNTT_DIT_core inPlaceNTT_DIT_core_inst (
      .clk(clk),
      .rst(rst),
      .vec_rsc_triosy_0_0_lz(vec_rsc_triosy_0_0_lz),
      .vec_rsc_triosy_0_1_lz(vec_rsc_triosy_0_1_lz),
      .vec_rsc_triosy_0_2_lz(vec_rsc_triosy_0_2_lz),
      .vec_rsc_triosy_0_3_lz(vec_rsc_triosy_0_3_lz),
      .vec_rsc_triosy_0_4_lz(vec_rsc_triosy_0_4_lz),
      .vec_rsc_triosy_0_5_lz(vec_rsc_triosy_0_5_lz),
      .vec_rsc_triosy_0_6_lz(vec_rsc_triosy_0_6_lz),
      .vec_rsc_triosy_0_7_lz(vec_rsc_triosy_0_7_lz),
      .vec_rsc_triosy_0_8_lz(vec_rsc_triosy_0_8_lz),
      .vec_rsc_triosy_0_9_lz(vec_rsc_triosy_0_9_lz),
      .vec_rsc_triosy_0_10_lz(vec_rsc_triosy_0_10_lz),
      .vec_rsc_triosy_0_11_lz(vec_rsc_triosy_0_11_lz),
      .vec_rsc_triosy_0_12_lz(vec_rsc_triosy_0_12_lz),
      .vec_rsc_triosy_0_13_lz(vec_rsc_triosy_0_13_lz),
      .vec_rsc_triosy_0_14_lz(vec_rsc_triosy_0_14_lz),
      .vec_rsc_triosy_0_15_lz(vec_rsc_triosy_0_15_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_dat(r_rsc_dat),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .vec_rsc_0_0_i_qa_d(vec_rsc_0_0_i_qa_d),
      .vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_1_i_qa_d(vec_rsc_0_1_i_qa_d),
      .vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_2_i_qa_d(vec_rsc_0_2_i_qa_d),
      .vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_3_i_qa_d(vec_rsc_0_3_i_qa_d),
      .vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_4_i_qa_d(vec_rsc_0_4_i_qa_d),
      .vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_5_i_qa_d(vec_rsc_0_5_i_qa_d),
      .vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_6_i_qa_d(vec_rsc_0_6_i_qa_d),
      .vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_7_i_qa_d(vec_rsc_0_7_i_qa_d),
      .vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_8_i_qa_d(vec_rsc_0_8_i_qa_d),
      .vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_9_i_qa_d(vec_rsc_0_9_i_qa_d),
      .vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_10_i_qa_d(vec_rsc_0_10_i_qa_d),
      .vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_11_i_qa_d(vec_rsc_0_11_i_qa_d),
      .vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_12_i_qa_d(vec_rsc_0_12_i_qa_d),
      .vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_13_i_qa_d(vec_rsc_0_13_i_qa_d),
      .vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_14_i_qa_d(vec_rsc_0_14_i_qa_d),
      .vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_15_i_qa_d(vec_rsc_0_15_i_qa_d),
      .vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(vec_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .vec_rsc_0_0_i_adra_d_pff(vec_rsc_0_0_i_adra_d_iff),
      .vec_rsc_0_0_i_da_d_pff(vec_rsc_0_0_i_da_d_iff),
      .vec_rsc_0_0_i_wea_d_pff(vec_rsc_0_0_i_wea_d_iff),
      .vec_rsc_0_1_i_wea_d_pff(vec_rsc_0_1_i_wea_d_iff),
      .vec_rsc_0_2_i_wea_d_pff(vec_rsc_0_2_i_wea_d_iff),
      .vec_rsc_0_3_i_wea_d_pff(vec_rsc_0_3_i_wea_d_iff),
      .vec_rsc_0_4_i_wea_d_pff(vec_rsc_0_4_i_wea_d_iff),
      .vec_rsc_0_5_i_wea_d_pff(vec_rsc_0_5_i_wea_d_iff),
      .vec_rsc_0_6_i_wea_d_pff(vec_rsc_0_6_i_wea_d_iff),
      .vec_rsc_0_7_i_wea_d_pff(vec_rsc_0_7_i_wea_d_iff),
      .vec_rsc_0_8_i_wea_d_pff(vec_rsc_0_8_i_wea_d_iff),
      .vec_rsc_0_9_i_wea_d_pff(vec_rsc_0_9_i_wea_d_iff),
      .vec_rsc_0_10_i_wea_d_pff(vec_rsc_0_10_i_wea_d_iff),
      .vec_rsc_0_11_i_wea_d_pff(vec_rsc_0_11_i_wea_d_iff),
      .vec_rsc_0_12_i_wea_d_pff(vec_rsc_0_12_i_wea_d_iff),
      .vec_rsc_0_13_i_wea_d_pff(vec_rsc_0_13_i_wea_d_iff),
      .vec_rsc_0_14_i_wea_d_pff(vec_rsc_0_14_i_wea_d_iff),
      .vec_rsc_0_15_i_wea_d_pff(vec_rsc_0_15_i_wea_d_iff)
    );
endmodule



