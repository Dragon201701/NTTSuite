
//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v 
//
// File:      $Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.v
//
// BASELINE:  Catapult-C version 2006b.63
// MODIFIED:  2007-04-03, tnagler
//
// Note: this file uses Verilog2001 features; 
//       please enable Verilog2001 in the flow!

module mgc_mul_pipe (a, b, clk, en, a_rst, s_rst, z);

    // Parameters:
    parameter integer width_a = 32'd4;  // input a bit width
    parameter         signd_a =  1'b1;  // input a type (1=signed, 0=unsigned)
    parameter integer width_b = 32'd4;  // input b bit width
    parameter         signd_b =  1'b1;  // input b type (1=signed, 0=unsigned)
    parameter integer width_z = 32'd8;  // result bit width (= width_a + width_b)
    parameter      clock_edge =  1'b0;  // clock polarity (1=posedge, 0=negedge)
    parameter   enable_active =  1'b0;  // enable polarity (1=posedge, 0=negedge)
    parameter    a_rst_active =  1'b1;  // unused
    parameter    s_rst_active =  1'b1;  // unused
    parameter integer  stages = 32'd2;  // number of output registers + 1 (careful!)
    parameter integer n_inreg = 32'd0;  // number of input registers
   
    localparam integer width_ab = width_a + width_b;  // multiplier result width
    localparam integer n_inreg_min = (n_inreg > 1) ? (n_inreg-1) : 0; // for Synopsys DC
   
    // I/O ports:
    input  [width_a-1:0] a;      // input A
    input  [width_b-1:0] b;      // input B
    input                clk;    // clock
    input                en;     // enable
    input                a_rst;  // async reset (unused)
    input                s_rst;  // sync reset (unused)
    output [width_z-1:0] z;      // output


    // Input registers:

    wire [width_a-1:0] a_f;
    wire [width_b-1:0] b_f;

    integer i;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a, 
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(negedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    else
    begin: POS_EDGE1
        case (n_inreg)
        32'd0: begin: B1
            assign a_f = a, 
                   b_f = b;
        end
        default: begin: B2
            reg [width_a-1:0] a_reg [n_inreg_min:0];
            reg [width_b-1:0] b_reg [n_inreg_min:0];
            always @(posedge clk)
            if (en == enable_active)
            begin: B21
                a_reg[0] <= a;
                b_reg[0] <= b;
                for (i = 0; i < n_inreg_min; i = i + 1)
                begin: B3
                    a_reg[i+1] <= a_reg[i];
                    b_reg[i+1] <= b_reg[i];
                end
            end
            assign a_f = a_reg[n_inreg_min],
                   b_f = b_reg[n_inreg_min];
        end
        endcase
    end
    endgenerate


    // Output:
    wire [width_z-1:0]  xz;

    function signed [width_z-1:0] conv_signed;
      input signed [width_ab-1:0] res;
      conv_signed = res[width_z-1:0];
    endfunction

    generate
      wire signed [width_ab-1:0] res;
      if ( (signd_a == 1'b1) && (signd_b == 1'b1) )
      begin: SIGNED_AB
              assign res = $signed(a_f) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b1) && (signd_b == 1'b0) )
      begin: SIGNED_A
              assign res = $signed(a_f) * $signed({1'b0, b_f});
              assign xz = conv_signed(res);
      end
      else if ( (signd_a == 1'b0) && (signd_b == 1'b1) )
      begin: SIGNED_B
              assign res = $signed({1'b0,a_f}) * $signed(b_f);
              assign xz = conv_signed(res);
      end
      else
      begin: UNSIGNED_AB
              assign res = a_f * b_f;
	      assign xz = res[width_z-1:0];
      end
    endgenerate


    // Output registers:

    reg  [width_z-1:0] reg_array[stages-2:0];
    wire [width_z-1:0] z;

    generate
    if (clock_edge == 1'b0)
    begin: NEG_EDGE2
        always @(negedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    else
    begin: POS_EDGE2
        always @(posedge clk)
        if (en == enable_active)
            for (i = stages-2; i >= 0; i = i-1)
                if (i == 0)
                    reg_array[i] <= xz;
                else
                    reg_array[i] <= reg_array[i-1];
    end
    endgenerate

    assign z = reg_array[stages-2];
endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v5.v 
module mgc_shift_bl_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate if ( signd_a )
   begin: SGNED
     assign z = fshl_s(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
     assign z = fshl_s(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift left - signed shift argument
   function [width_z-1:0] fshl_s;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      reg [width_a:0] sbit_arg1;
      begin
        // Ignoring the possibility that arg2[width_s-1] could be X
        // because of customer complaints regarding X'es in simulation results
        if ( arg2[width_s-1] == 1'b0 )
        begin
          sbit_arg1[width_a:0] = {(width_a+1){1'b0}};
          fshl_s = fshl_u(arg1, arg2, sbit);
        end
        else
        begin
          sbit_arg1[width_a] = sbit;
          sbit_arg1[width_a-1:0] = arg1;
          fshl_s = fshr_u(sbit_arg1[width_a:1], ~arg2, sbit);
        end
      end
   endfunction

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_DPRAM_RBW_DUAL.v 
// Memory Type:            BLOCK
// Operating Mode:         True Dual Port (2-Port)
// Clock Mode:             Dual Clock
// 
// RTL Code RW Resolution: RBW
// Catapult RW Resolution: RBW
// 
// HDL Work Library:       Xilinx_RAMS_lib
// Component Name:         BLOCK_DPRAM_RBW_DUAL
// Latency = 1:            RAM with no registers on inputs or outputs
//         = 2:            adds embedded register on RAM output
//         = 3:            adds fabric registers to non-clock input RAM pins
//         = 4:            adds fabric register to output (driven by embedded register from latency=2)

module BLOCK_DPRAM_RBW_DUAL #(
  parameter addr_width = 8 ,
  parameter data_width = 7 ,
  parameter depth = 256 ,
  parameter latency = 1 
  
)( adra,adrb,clka,clka_en,clkb,clkb_en,da,db,qa,qb,wea,web);

  input [addr_width-1:0] adra;
  input [addr_width-1:0] adrb;
  input  clka;
  input  clka_en;
  input  clkb;
  input  clkb_en;
  input [data_width-1:0] da;
  input [data_width-1:0] db;
  output [data_width-1:0] qa;
  output [data_width-1:0] qb;
  input  wea;
  input  web;
  
  (* ram_style = "block" *)
  reg [data_width-1:0] mem [depth-1:0];// synthesis syn_ramstyle="block"
  
  reg [data_width-1:0] ramqa;
  reg [data_width-1:0] ramqb;
  
  // Port Map
  // rwA :: ADDRESS adra CLOCK clka ENABLE clka_en DATA_IN da DATA_OUT qa WRITE_ENABLE wea
  // rwB :: ADDRESS adrb CLOCK clkb ENABLE clkb_en DATA_IN db DATA_OUT qb WRITE_ENABLE web

  generate
    // Register all non-clock inputs (latency < 3)
    if (latency > 2 ) begin
      reg [addr_width-1:0] adra_reg;
      reg [data_width-1:0] da_reg;
      reg wea_reg;
      reg [addr_width-1:0] adrb_reg;
      reg [data_width-1:0] db_reg;
      reg web_reg;
      
      always @(posedge clka) begin
        if (clka_en) begin
          adra_reg <= adra;
          da_reg <= da;
          wea_reg <= wea;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          adrb_reg <= adrb;
          db_reg <= db;
          web_reg <= web;
        end
      end
      
    // Access memory with registered inputs
      always @(posedge clka) begin
        if (clka_en) begin
            ramqa <= mem[adra_reg];
            if (wea_reg) begin
              mem[adra_reg] <= da_reg;
            end
        end
      end
      always @(posedge clka) begin
        if (clka_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
            ramqb <= mem[adrb_reg];
            if (web_reg) begin
              mem[adrb_reg] <= db_reg;
            end
        end
      end
      
    end // END register inputs

    else begin
    // latency = 1||2: Access memory with non-registered inputs
      always @(posedge clka) begin
        if (clka_en) begin
            ramqa <= mem[adra];
            if (wea) begin
              mem[adra] <= da;
            end
        end
      end
      always @(posedge clka) begin
        if (clka_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
            ramqb <= mem[adrb];
            if (web) begin
              mem[adrb] <= db;
            end
        end
      end
      
    end
  endgenerate //END input port generate 

  generate
    // latency=1: sequential RAM outputs drive module outputs
    if (latency == 1) begin
      assign qa = ramqa;
      assign qb = ramqb;
      
    end

    else if (latency == 2 || latency == 3) begin
    // latency=2: sequential (RAM output => tmp register => module output)
      reg [data_width-1:0] tmpqa;
      reg [data_width-1:0] tmpqb;
      
      always @(posedge clka) begin
        if (clka_en) begin
          tmpqa <= ramqa;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          tmpqb <= ramqb;
        end
      end
      
      assign qa = tmpqa;
      assign qb = tmpqb;
      
    end
    else if (latency == 4) begin
    // latency=4: (RAM => tmp1 register => tmp2 fabric register => module output)
      reg [data_width-1:0] tmp1qa;
      reg [data_width-1:0] tmp1qb;
      
      reg [data_width-1:0] tmp2qa;
      reg [data_width-1:0] tmp2qb;
      
      always @(posedge clka) begin
        if (clka_en) begin
          tmp1qa <= ramqa;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          tmp1qb <= ramqb;
        end
      end
      
      always @(posedge clka) begin
        if (clka_en) begin
          tmp2qa <= tmp1qa;
        end
      end
      always @(posedge clkb) begin
        if (clkb_en) begin
          tmp2qb <= tmp1qb;
        end
      end
      
      assign qa = tmp2qa;
      assign qb = tmp2qb;
      
    end
    else begin
      //Add error check if latency > 4 or add N-pipeline regs
    end
  endgenerate //END output port generate

endmodule

//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.5c/896140 Production Release
//  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
// 
//  Generated by:   yl7897@newnano.poly.edu
//  Generated date: Tue Sep 14 21:33:32 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen
    (
  qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en, da_d, qa_d, wea_d,
      rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
// ------------------------------------------------------------------


module peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen
    (
  clkb_en, clka_en, qb, web, db, adrb, qa, wea, da, adra, adra_d, clka, clka_en_d,
      clkb_en_d, da_d, qa_d, wea_d, rwA_rw_ram_ir_internal_RMASK_B_d, rwA_rw_ram_ir_internal_WMASK_B_d
);
  output clkb_en;
  output clka_en;
  input [31:0] qb;
  output web;
  output [31:0] db;
  output [7:0] adrb;
  input [31:0] qa;
  output wea;
  output [31:0] da;
  output [7:0] adra;
  input [15:0] adra_d;
  input clka;
  input clka_en_d;
  input clkb_en_d;
  input [63:0] da_d;
  output [63:0] qa_d;
  input [1:0] wea_d;
  input [1:0] rwA_rw_ram_ir_internal_RMASK_B_d;
  input [1:0] rwA_rw_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clkb_en = clkb_en_d;
  assign clka_en = clka_en_d;
  assign qa_d[63:32] = qb;
  assign web = (rwA_rw_ram_ir_internal_WMASK_B_d[1]);
  assign db = (da_d[63:32]);
  assign adrb = (adra_d[15:8]);
  assign qa_d[31:0] = qa;
  assign wea = (rwA_rw_ram_ir_internal_WMASK_B_d[0]);
  assign da = (da_d[31:0]);
  assign adra = (adra_d[7:0]);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module peaseNTT_core_core_fsm (
  clk, rst, fsm_output, INNER_LOOP1_C_0_tr0, INNER_LOOP2_C_0_tr0, STAGE_LOOP_C_2_tr0,
      INNER_LOOP3_C_0_tr0, INNER_LOOP4_C_0_tr0, INNER_LOOP4_C_0_tr1
);
  input clk;
  input rst;
  output [10:0] fsm_output;
  reg [10:0] fsm_output;
  input INNER_LOOP1_C_0_tr0;
  input INNER_LOOP2_C_0_tr0;
  input STAGE_LOOP_C_2_tr0;
  input INNER_LOOP3_C_0_tr0;
  input INNER_LOOP4_C_0_tr0;
  input INNER_LOOP4_C_0_tr1;


  // FSM State Type Declaration for peaseNTT_core_core_fsm_1
  parameter
    main_C_0 = 4'd0,
    STAGE_LOOP_C_0 = 4'd1,
    INNER_LOOP1_C_0 = 4'd2,
    STAGE_LOOP_C_1 = 4'd3,
    INNER_LOOP2_C_0 = 4'd4,
    STAGE_LOOP_C_2 = 4'd5,
    STAGE_LOOP1_C_0 = 4'd6,
    INNER_LOOP3_C_0 = 4'd7,
    STAGE_LOOP1_C_1 = 4'd8,
    INNER_LOOP4_C_0 = 4'd9,
    main_C_1 = 4'd10;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : peaseNTT_core_core_fsm_1
    case (state_var)
      STAGE_LOOP_C_0 : begin
        fsm_output = 11'b00000000010;
        state_var_NS = INNER_LOOP1_C_0;
      end
      INNER_LOOP1_C_0 : begin
        fsm_output = 11'b00000000100;
        if ( INNER_LOOP1_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_1;
        end
        else begin
          state_var_NS = INNER_LOOP1_C_0;
        end
      end
      STAGE_LOOP_C_1 : begin
        fsm_output = 11'b00000001000;
        state_var_NS = INNER_LOOP2_C_0;
      end
      INNER_LOOP2_C_0 : begin
        fsm_output = 11'b00000010000;
        if ( INNER_LOOP2_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP_C_2;
        end
        else begin
          state_var_NS = INNER_LOOP2_C_0;
        end
      end
      STAGE_LOOP_C_2 : begin
        fsm_output = 11'b00000100000;
        if ( STAGE_LOOP_C_2_tr0 ) begin
          state_var_NS = STAGE_LOOP1_C_0;
        end
        else begin
          state_var_NS = STAGE_LOOP_C_0;
        end
      end
      STAGE_LOOP1_C_0 : begin
        fsm_output = 11'b00001000000;
        state_var_NS = INNER_LOOP3_C_0;
      end
      INNER_LOOP3_C_0 : begin
        fsm_output = 11'b00010000000;
        if ( INNER_LOOP3_C_0_tr0 ) begin
          state_var_NS = STAGE_LOOP1_C_1;
        end
        else begin
          state_var_NS = INNER_LOOP3_C_0;
        end
      end
      STAGE_LOOP1_C_1 : begin
        fsm_output = 11'b00100000000;
        state_var_NS = INNER_LOOP4_C_0;
      end
      INNER_LOOP4_C_0 : begin
        fsm_output = 11'b01000000000;
        if ( INNER_LOOP4_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else if ( INNER_LOOP4_C_0_tr1 ) begin
          state_var_NS = INNER_LOOP4_C_0;
        end
        else begin
          state_var_NS = STAGE_LOOP1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 11'b10000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 11'b00000000001;
        state_var_NS = STAGE_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_core_wait_dp
// ------------------------------------------------------------------


module peaseNTT_core_wait_dp (
  yt_rsc_0_0_cgo_iro, yt_rsc_0_0_i_clka_en_d, yt_rsc_0_16_cgo_iro, yt_rsc_0_16_i_clka_en_d,
      ensig_cgo_iro, ensig_cgo_iro_17, yt_rsc_0_0_cgo, yt_rsc_0_16_cgo, ensig_cgo,
      mult_t_mul_cmp_en, ensig_cgo_17, mult_z_mul_cmp_1_en
);
  input yt_rsc_0_0_cgo_iro;
  output yt_rsc_0_0_i_clka_en_d;
  input yt_rsc_0_16_cgo_iro;
  output yt_rsc_0_16_i_clka_en_d;
  input ensig_cgo_iro;
  input ensig_cgo_iro_17;
  input yt_rsc_0_0_cgo;
  input yt_rsc_0_16_cgo;
  input ensig_cgo;
  output mult_t_mul_cmp_en;
  input ensig_cgo_17;
  output mult_z_mul_cmp_1_en;



  // Interconnect Declarations for Component Instantiations 
  assign yt_rsc_0_0_i_clka_en_d = yt_rsc_0_0_cgo | yt_rsc_0_0_cgo_iro;
  assign yt_rsc_0_16_i_clka_en_d = yt_rsc_0_16_cgo | yt_rsc_0_16_cgo_iro;
  assign mult_t_mul_cmp_en = ensig_cgo | ensig_cgo_iro;
  assign mult_z_mul_cmp_1_en = ensig_cgo_17 | ensig_cgo_iro_17;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT_core
// ------------------------------------------------------------------


module peaseNTT_core (
  clk, rst, xt_rsc_triosy_0_0_lz, xt_rsc_triosy_0_1_lz, xt_rsc_triosy_0_2_lz, xt_rsc_triosy_0_3_lz,
      xt_rsc_triosy_0_4_lz, xt_rsc_triosy_0_5_lz, xt_rsc_triosy_0_6_lz, xt_rsc_triosy_0_7_lz,
      xt_rsc_triosy_0_8_lz, xt_rsc_triosy_0_9_lz, xt_rsc_triosy_0_10_lz, xt_rsc_triosy_0_11_lz,
      xt_rsc_triosy_0_12_lz, xt_rsc_triosy_0_13_lz, xt_rsc_triosy_0_14_lz, xt_rsc_triosy_0_15_lz,
      xt_rsc_triosy_0_16_lz, xt_rsc_triosy_0_17_lz, xt_rsc_triosy_0_18_lz, xt_rsc_triosy_0_19_lz,
      xt_rsc_triosy_0_20_lz, xt_rsc_triosy_0_21_lz, xt_rsc_triosy_0_22_lz, xt_rsc_triosy_0_23_lz,
      xt_rsc_triosy_0_24_lz, xt_rsc_triosy_0_25_lz, xt_rsc_triosy_0_26_lz, xt_rsc_triosy_0_27_lz,
      xt_rsc_triosy_0_28_lz, xt_rsc_triosy_0_29_lz, xt_rsc_triosy_0_30_lz, xt_rsc_triosy_0_31_lz,
      p_rsc_dat, p_rsc_triosy_lz, r_rsc_triosy_lz, twiddle_rsc_triosy_0_0_lz, twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_triosy_0_2_lz, twiddle_rsc_triosy_0_3_lz, twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_triosy_0_5_lz, twiddle_rsc_triosy_0_6_lz, twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_triosy_0_8_lz, twiddle_rsc_triosy_0_9_lz, twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_triosy_0_11_lz, twiddle_rsc_triosy_0_12_lz, twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_triosy_0_14_lz, twiddle_rsc_triosy_0_15_lz, twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_triosy_0_1_lz, twiddle_h_rsc_triosy_0_2_lz, twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_triosy_0_4_lz, twiddle_h_rsc_triosy_0_5_lz, twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_triosy_0_7_lz, twiddle_h_rsc_triosy_0_8_lz, twiddle_h_rsc_triosy_0_9_lz,
      twiddle_h_rsc_triosy_0_10_lz, twiddle_h_rsc_triosy_0_11_lz, twiddle_h_rsc_triosy_0_12_lz,
      twiddle_h_rsc_triosy_0_13_lz, twiddle_h_rsc_triosy_0_14_lz, twiddle_h_rsc_triosy_0_15_lz,
      yt_rsc_0_0_i_adra_d, yt_rsc_0_0_i_clka_en_d, yt_rsc_0_0_i_da_d, yt_rsc_0_0_i_qa_d,
      yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d, yt_rsc_0_1_i_adra_d, yt_rsc_0_1_i_da_d,
      yt_rsc_0_1_i_qa_d, yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d, yt_rsc_0_2_i_adra_d,
      yt_rsc_0_2_i_da_d, yt_rsc_0_2_i_qa_d, yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_3_i_adra_d, yt_rsc_0_3_i_da_d, yt_rsc_0_3_i_qa_d, yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_4_i_adra_d, yt_rsc_0_4_i_da_d, yt_rsc_0_4_i_qa_d, yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_5_i_adra_d, yt_rsc_0_5_i_da_d, yt_rsc_0_5_i_qa_d, yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_6_i_adra_d, yt_rsc_0_6_i_da_d, yt_rsc_0_6_i_qa_d, yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_7_i_adra_d, yt_rsc_0_7_i_da_d, yt_rsc_0_7_i_qa_d, yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_8_i_adra_d, yt_rsc_0_8_i_da_d, yt_rsc_0_8_i_qa_d, yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_9_i_adra_d, yt_rsc_0_9_i_da_d, yt_rsc_0_9_i_qa_d, yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_10_i_adra_d, yt_rsc_0_10_i_da_d, yt_rsc_0_10_i_qa_d, yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_11_i_adra_d, yt_rsc_0_11_i_da_d, yt_rsc_0_11_i_qa_d, yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_12_i_adra_d, yt_rsc_0_12_i_da_d, yt_rsc_0_12_i_qa_d, yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_13_i_adra_d, yt_rsc_0_13_i_da_d, yt_rsc_0_13_i_qa_d, yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_14_i_adra_d, yt_rsc_0_14_i_da_d, yt_rsc_0_14_i_qa_d, yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_15_i_adra_d, yt_rsc_0_15_i_da_d, yt_rsc_0_15_i_qa_d, yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_16_i_adra_d, yt_rsc_0_16_i_clka_en_d, yt_rsc_0_16_i_da_d, yt_rsc_0_16_i_qa_d,
      yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d, yt_rsc_0_17_i_adra_d, yt_rsc_0_17_i_da_d,
      yt_rsc_0_17_i_qa_d, yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d, yt_rsc_0_18_i_adra_d,
      yt_rsc_0_18_i_da_d, yt_rsc_0_18_i_qa_d, yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_19_i_adra_d, yt_rsc_0_19_i_da_d, yt_rsc_0_19_i_qa_d, yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_20_i_adra_d, yt_rsc_0_20_i_da_d, yt_rsc_0_20_i_qa_d, yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_21_i_adra_d, yt_rsc_0_21_i_da_d, yt_rsc_0_21_i_qa_d, yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_22_i_adra_d, yt_rsc_0_22_i_da_d, yt_rsc_0_22_i_qa_d, yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_23_i_adra_d, yt_rsc_0_23_i_da_d, yt_rsc_0_23_i_qa_d, yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_24_i_adra_d, yt_rsc_0_24_i_da_d, yt_rsc_0_24_i_qa_d, yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_25_i_adra_d, yt_rsc_0_25_i_da_d, yt_rsc_0_25_i_qa_d, yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_26_i_adra_d, yt_rsc_0_26_i_da_d, yt_rsc_0_26_i_qa_d, yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_27_i_adra_d, yt_rsc_0_27_i_da_d, yt_rsc_0_27_i_qa_d, yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_28_i_adra_d, yt_rsc_0_28_i_da_d, yt_rsc_0_28_i_qa_d, yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_29_i_adra_d, yt_rsc_0_29_i_da_d, yt_rsc_0_29_i_qa_d, yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_30_i_adra_d, yt_rsc_0_30_i_da_d, yt_rsc_0_30_i_qa_d, yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_31_i_adra_d, yt_rsc_0_31_i_da_d, yt_rsc_0_31_i_qa_d, yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_0_i_adra_d, xt_rsc_0_0_i_da_d, xt_rsc_0_0_i_qa_d, xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_1_i_adra_d, xt_rsc_0_1_i_da_d, xt_rsc_0_1_i_qa_d, xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_2_i_adra_d, xt_rsc_0_2_i_da_d, xt_rsc_0_2_i_qa_d, xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_3_i_adra_d, xt_rsc_0_3_i_da_d, xt_rsc_0_3_i_qa_d, xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_4_i_adra_d, xt_rsc_0_4_i_da_d, xt_rsc_0_4_i_qa_d, xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_5_i_adra_d, xt_rsc_0_5_i_da_d, xt_rsc_0_5_i_qa_d, xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_6_i_adra_d, xt_rsc_0_6_i_da_d, xt_rsc_0_6_i_qa_d, xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_7_i_adra_d, xt_rsc_0_7_i_da_d, xt_rsc_0_7_i_qa_d, xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_8_i_adra_d, xt_rsc_0_8_i_da_d, xt_rsc_0_8_i_qa_d, xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_9_i_adra_d, xt_rsc_0_9_i_da_d, xt_rsc_0_9_i_qa_d, xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_10_i_adra_d, xt_rsc_0_10_i_da_d, xt_rsc_0_10_i_qa_d, xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_11_i_adra_d, xt_rsc_0_11_i_da_d, xt_rsc_0_11_i_qa_d, xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_12_i_adra_d, xt_rsc_0_12_i_da_d, xt_rsc_0_12_i_qa_d, xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_13_i_adra_d, xt_rsc_0_13_i_da_d, xt_rsc_0_13_i_qa_d, xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_14_i_adra_d, xt_rsc_0_14_i_da_d, xt_rsc_0_14_i_qa_d, xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_15_i_adra_d, xt_rsc_0_15_i_da_d, xt_rsc_0_15_i_qa_d, xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_16_i_adra_d, xt_rsc_0_16_i_da_d, xt_rsc_0_16_i_qa_d, xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_17_i_adra_d, xt_rsc_0_17_i_da_d, xt_rsc_0_17_i_qa_d, xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_18_i_adra_d, xt_rsc_0_18_i_da_d, xt_rsc_0_18_i_qa_d, xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_19_i_adra_d, xt_rsc_0_19_i_da_d, xt_rsc_0_19_i_qa_d, xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_20_i_adra_d, xt_rsc_0_20_i_da_d, xt_rsc_0_20_i_qa_d, xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_21_i_adra_d, xt_rsc_0_21_i_da_d, xt_rsc_0_21_i_qa_d, xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_22_i_adra_d, xt_rsc_0_22_i_da_d, xt_rsc_0_22_i_qa_d, xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_23_i_adra_d, xt_rsc_0_23_i_da_d, xt_rsc_0_23_i_qa_d, xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_24_i_adra_d, xt_rsc_0_24_i_da_d, xt_rsc_0_24_i_qa_d, xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_25_i_adra_d, xt_rsc_0_25_i_da_d, xt_rsc_0_25_i_qa_d, xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_26_i_adra_d, xt_rsc_0_26_i_da_d, xt_rsc_0_26_i_qa_d, xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_27_i_adra_d, xt_rsc_0_27_i_da_d, xt_rsc_0_27_i_qa_d, xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_28_i_adra_d, xt_rsc_0_28_i_da_d, xt_rsc_0_28_i_qa_d, xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_29_i_adra_d, xt_rsc_0_29_i_da_d, xt_rsc_0_29_i_qa_d, xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_30_i_adra_d, xt_rsc_0_30_i_da_d, xt_rsc_0_30_i_qa_d, xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_31_i_adra_d, xt_rsc_0_31_i_da_d, xt_rsc_0_31_i_qa_d, xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_0_i_adra_d, twiddle_rsc_0_0_i_qa_d, twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_1_i_adra_d, twiddle_rsc_0_1_i_qa_d, twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_2_i_adra_d, twiddle_rsc_0_2_i_qa_d, twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_3_i_adra_d, twiddle_rsc_0_3_i_qa_d, twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_4_i_adra_d, twiddle_rsc_0_4_i_qa_d, twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_5_i_adra_d, twiddle_rsc_0_5_i_qa_d, twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_6_i_adra_d, twiddle_rsc_0_6_i_qa_d, twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_7_i_adra_d, twiddle_rsc_0_7_i_qa_d, twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_8_i_adra_d, twiddle_rsc_0_8_i_qa_d, twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_9_i_adra_d, twiddle_rsc_0_9_i_qa_d, twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_10_i_adra_d, twiddle_rsc_0_10_i_qa_d, twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_11_i_adra_d, twiddle_rsc_0_11_i_qa_d, twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_12_i_adra_d, twiddle_rsc_0_12_i_qa_d, twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_13_i_adra_d, twiddle_rsc_0_13_i_qa_d, twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_14_i_adra_d, twiddle_rsc_0_14_i_qa_d, twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_rsc_0_15_i_adra_d, twiddle_rsc_0_15_i_qa_d, twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_0_i_adra_d, twiddle_h_rsc_0_0_i_qa_d, twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_1_i_adra_d, twiddle_h_rsc_0_1_i_qa_d, twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_2_i_adra_d, twiddle_h_rsc_0_2_i_qa_d, twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_3_i_adra_d, twiddle_h_rsc_0_3_i_qa_d, twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_4_i_adra_d, twiddle_h_rsc_0_4_i_qa_d, twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_5_i_adra_d, twiddle_h_rsc_0_5_i_qa_d, twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_6_i_adra_d, twiddle_h_rsc_0_6_i_qa_d, twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_7_i_adra_d, twiddle_h_rsc_0_7_i_qa_d, twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_8_i_adra_d, twiddle_h_rsc_0_8_i_qa_d, twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_9_i_adra_d, twiddle_h_rsc_0_9_i_qa_d, twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_10_i_adra_d, twiddle_h_rsc_0_10_i_qa_d, twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_11_i_adra_d, twiddle_h_rsc_0_11_i_qa_d, twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_12_i_adra_d, twiddle_h_rsc_0_12_i_qa_d, twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_13_i_adra_d, twiddle_h_rsc_0_13_i_qa_d, twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_14_i_adra_d, twiddle_h_rsc_0_14_i_qa_d, twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      twiddle_h_rsc_0_15_i_adra_d, twiddle_h_rsc_0_15_i_qa_d, twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_0_i_wea_d_pff, yt_rsc_0_16_i_wea_d_pff, xt_rsc_0_0_i_wea_d_pff, xt_rsc_0_16_i_wea_d_pff
);
  input clk;
  input rst;
  output xt_rsc_triosy_0_0_lz;
  output xt_rsc_triosy_0_1_lz;
  output xt_rsc_triosy_0_2_lz;
  output xt_rsc_triosy_0_3_lz;
  output xt_rsc_triosy_0_4_lz;
  output xt_rsc_triosy_0_5_lz;
  output xt_rsc_triosy_0_6_lz;
  output xt_rsc_triosy_0_7_lz;
  output xt_rsc_triosy_0_8_lz;
  output xt_rsc_triosy_0_9_lz;
  output xt_rsc_triosy_0_10_lz;
  output xt_rsc_triosy_0_11_lz;
  output xt_rsc_triosy_0_12_lz;
  output xt_rsc_triosy_0_13_lz;
  output xt_rsc_triosy_0_14_lz;
  output xt_rsc_triosy_0_15_lz;
  output xt_rsc_triosy_0_16_lz;
  output xt_rsc_triosy_0_17_lz;
  output xt_rsc_triosy_0_18_lz;
  output xt_rsc_triosy_0_19_lz;
  output xt_rsc_triosy_0_20_lz;
  output xt_rsc_triosy_0_21_lz;
  output xt_rsc_triosy_0_22_lz;
  output xt_rsc_triosy_0_23_lz;
  output xt_rsc_triosy_0_24_lz;
  output xt_rsc_triosy_0_25_lz;
  output xt_rsc_triosy_0_26_lz;
  output xt_rsc_triosy_0_27_lz;
  output xt_rsc_triosy_0_28_lz;
  output xt_rsc_triosy_0_29_lz;
  output xt_rsc_triosy_0_30_lz;
  output xt_rsc_triosy_0_31_lz;
  input [31:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  output r_rsc_triosy_lz;
  output twiddle_rsc_triosy_0_0_lz;
  output twiddle_rsc_triosy_0_1_lz;
  output twiddle_rsc_triosy_0_2_lz;
  output twiddle_rsc_triosy_0_3_lz;
  output twiddle_rsc_triosy_0_4_lz;
  output twiddle_rsc_triosy_0_5_lz;
  output twiddle_rsc_triosy_0_6_lz;
  output twiddle_rsc_triosy_0_7_lz;
  output twiddle_rsc_triosy_0_8_lz;
  output twiddle_rsc_triosy_0_9_lz;
  output twiddle_rsc_triosy_0_10_lz;
  output twiddle_rsc_triosy_0_11_lz;
  output twiddle_rsc_triosy_0_12_lz;
  output twiddle_rsc_triosy_0_13_lz;
  output twiddle_rsc_triosy_0_14_lz;
  output twiddle_rsc_triosy_0_15_lz;
  output twiddle_h_rsc_triosy_0_0_lz;
  output twiddle_h_rsc_triosy_0_1_lz;
  output twiddle_h_rsc_triosy_0_2_lz;
  output twiddle_h_rsc_triosy_0_3_lz;
  output twiddle_h_rsc_triosy_0_4_lz;
  output twiddle_h_rsc_triosy_0_5_lz;
  output twiddle_h_rsc_triosy_0_6_lz;
  output twiddle_h_rsc_triosy_0_7_lz;
  output twiddle_h_rsc_triosy_0_8_lz;
  output twiddle_h_rsc_triosy_0_9_lz;
  output twiddle_h_rsc_triosy_0_10_lz;
  output twiddle_h_rsc_triosy_0_11_lz;
  output twiddle_h_rsc_triosy_0_12_lz;
  output twiddle_h_rsc_triosy_0_13_lz;
  output twiddle_h_rsc_triosy_0_14_lz;
  output twiddle_h_rsc_triosy_0_15_lz;
  output [15:0] yt_rsc_0_0_i_adra_d;
  output yt_rsc_0_0_i_clka_en_d;
  output [63:0] yt_rsc_0_0_i_da_d;
  input [63:0] yt_rsc_0_0_i_qa_d;
  output [1:0] yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_1_i_adra_d;
  output [63:0] yt_rsc_0_1_i_da_d;
  input [63:0] yt_rsc_0_1_i_qa_d;
  output [1:0] yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_2_i_adra_d;
  output [63:0] yt_rsc_0_2_i_da_d;
  input [63:0] yt_rsc_0_2_i_qa_d;
  output [1:0] yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_3_i_adra_d;
  output [63:0] yt_rsc_0_3_i_da_d;
  input [63:0] yt_rsc_0_3_i_qa_d;
  output [1:0] yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_4_i_adra_d;
  output [63:0] yt_rsc_0_4_i_da_d;
  input [63:0] yt_rsc_0_4_i_qa_d;
  output [1:0] yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_5_i_adra_d;
  output [63:0] yt_rsc_0_5_i_da_d;
  input [63:0] yt_rsc_0_5_i_qa_d;
  output [1:0] yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_6_i_adra_d;
  output [63:0] yt_rsc_0_6_i_da_d;
  input [63:0] yt_rsc_0_6_i_qa_d;
  output [1:0] yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_7_i_adra_d;
  output [63:0] yt_rsc_0_7_i_da_d;
  input [63:0] yt_rsc_0_7_i_qa_d;
  output [1:0] yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_8_i_adra_d;
  output [63:0] yt_rsc_0_8_i_da_d;
  input [63:0] yt_rsc_0_8_i_qa_d;
  output [1:0] yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_9_i_adra_d;
  output [63:0] yt_rsc_0_9_i_da_d;
  input [63:0] yt_rsc_0_9_i_qa_d;
  output [1:0] yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_10_i_adra_d;
  output [63:0] yt_rsc_0_10_i_da_d;
  input [63:0] yt_rsc_0_10_i_qa_d;
  output [1:0] yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_11_i_adra_d;
  output [63:0] yt_rsc_0_11_i_da_d;
  input [63:0] yt_rsc_0_11_i_qa_d;
  output [1:0] yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_12_i_adra_d;
  output [63:0] yt_rsc_0_12_i_da_d;
  input [63:0] yt_rsc_0_12_i_qa_d;
  output [1:0] yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_13_i_adra_d;
  output [63:0] yt_rsc_0_13_i_da_d;
  input [63:0] yt_rsc_0_13_i_qa_d;
  output [1:0] yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_14_i_adra_d;
  output [63:0] yt_rsc_0_14_i_da_d;
  input [63:0] yt_rsc_0_14_i_qa_d;
  output [1:0] yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_15_i_adra_d;
  output [63:0] yt_rsc_0_15_i_da_d;
  input [63:0] yt_rsc_0_15_i_qa_d;
  output [1:0] yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_16_i_adra_d;
  output yt_rsc_0_16_i_clka_en_d;
  output [63:0] yt_rsc_0_16_i_da_d;
  input [63:0] yt_rsc_0_16_i_qa_d;
  output [1:0] yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_17_i_adra_d;
  output [63:0] yt_rsc_0_17_i_da_d;
  input [63:0] yt_rsc_0_17_i_qa_d;
  output [1:0] yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_18_i_adra_d;
  output [63:0] yt_rsc_0_18_i_da_d;
  input [63:0] yt_rsc_0_18_i_qa_d;
  output [1:0] yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_19_i_adra_d;
  output [63:0] yt_rsc_0_19_i_da_d;
  input [63:0] yt_rsc_0_19_i_qa_d;
  output [1:0] yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_20_i_adra_d;
  output [63:0] yt_rsc_0_20_i_da_d;
  input [63:0] yt_rsc_0_20_i_qa_d;
  output [1:0] yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_21_i_adra_d;
  output [63:0] yt_rsc_0_21_i_da_d;
  input [63:0] yt_rsc_0_21_i_qa_d;
  output [1:0] yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_22_i_adra_d;
  output [63:0] yt_rsc_0_22_i_da_d;
  input [63:0] yt_rsc_0_22_i_qa_d;
  output [1:0] yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_23_i_adra_d;
  output [63:0] yt_rsc_0_23_i_da_d;
  input [63:0] yt_rsc_0_23_i_qa_d;
  output [1:0] yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_24_i_adra_d;
  output [63:0] yt_rsc_0_24_i_da_d;
  input [63:0] yt_rsc_0_24_i_qa_d;
  output [1:0] yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_25_i_adra_d;
  output [63:0] yt_rsc_0_25_i_da_d;
  input [63:0] yt_rsc_0_25_i_qa_d;
  output [1:0] yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_26_i_adra_d;
  output [63:0] yt_rsc_0_26_i_da_d;
  input [63:0] yt_rsc_0_26_i_qa_d;
  output [1:0] yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_27_i_adra_d;
  output [63:0] yt_rsc_0_27_i_da_d;
  input [63:0] yt_rsc_0_27_i_qa_d;
  output [1:0] yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_28_i_adra_d;
  output [63:0] yt_rsc_0_28_i_da_d;
  input [63:0] yt_rsc_0_28_i_qa_d;
  output [1:0] yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_29_i_adra_d;
  output [63:0] yt_rsc_0_29_i_da_d;
  input [63:0] yt_rsc_0_29_i_qa_d;
  output [1:0] yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_30_i_adra_d;
  output [63:0] yt_rsc_0_30_i_da_d;
  input [63:0] yt_rsc_0_30_i_qa_d;
  output [1:0] yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] yt_rsc_0_31_i_adra_d;
  output [63:0] yt_rsc_0_31_i_da_d;
  input [63:0] yt_rsc_0_31_i_qa_d;
  output [1:0] yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_0_i_adra_d;
  output [63:0] xt_rsc_0_0_i_da_d;
  input [63:0] xt_rsc_0_0_i_qa_d;
  output [1:0] xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_1_i_adra_d;
  output [63:0] xt_rsc_0_1_i_da_d;
  input [63:0] xt_rsc_0_1_i_qa_d;
  output [1:0] xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_2_i_adra_d;
  output [63:0] xt_rsc_0_2_i_da_d;
  input [63:0] xt_rsc_0_2_i_qa_d;
  output [1:0] xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_3_i_adra_d;
  output [63:0] xt_rsc_0_3_i_da_d;
  input [63:0] xt_rsc_0_3_i_qa_d;
  output [1:0] xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_4_i_adra_d;
  output [63:0] xt_rsc_0_4_i_da_d;
  input [63:0] xt_rsc_0_4_i_qa_d;
  output [1:0] xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_5_i_adra_d;
  output [63:0] xt_rsc_0_5_i_da_d;
  input [63:0] xt_rsc_0_5_i_qa_d;
  output [1:0] xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_6_i_adra_d;
  output [63:0] xt_rsc_0_6_i_da_d;
  input [63:0] xt_rsc_0_6_i_qa_d;
  output [1:0] xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_7_i_adra_d;
  output [63:0] xt_rsc_0_7_i_da_d;
  input [63:0] xt_rsc_0_7_i_qa_d;
  output [1:0] xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_8_i_adra_d;
  output [63:0] xt_rsc_0_8_i_da_d;
  input [63:0] xt_rsc_0_8_i_qa_d;
  output [1:0] xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_9_i_adra_d;
  output [63:0] xt_rsc_0_9_i_da_d;
  input [63:0] xt_rsc_0_9_i_qa_d;
  output [1:0] xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_10_i_adra_d;
  output [63:0] xt_rsc_0_10_i_da_d;
  input [63:0] xt_rsc_0_10_i_qa_d;
  output [1:0] xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_11_i_adra_d;
  output [63:0] xt_rsc_0_11_i_da_d;
  input [63:0] xt_rsc_0_11_i_qa_d;
  output [1:0] xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_12_i_adra_d;
  output [63:0] xt_rsc_0_12_i_da_d;
  input [63:0] xt_rsc_0_12_i_qa_d;
  output [1:0] xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_13_i_adra_d;
  output [63:0] xt_rsc_0_13_i_da_d;
  input [63:0] xt_rsc_0_13_i_qa_d;
  output [1:0] xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_14_i_adra_d;
  output [63:0] xt_rsc_0_14_i_da_d;
  input [63:0] xt_rsc_0_14_i_qa_d;
  output [1:0] xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_15_i_adra_d;
  output [63:0] xt_rsc_0_15_i_da_d;
  input [63:0] xt_rsc_0_15_i_qa_d;
  output [1:0] xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_16_i_adra_d;
  output [63:0] xt_rsc_0_16_i_da_d;
  input [63:0] xt_rsc_0_16_i_qa_d;
  output [1:0] xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_17_i_adra_d;
  output [63:0] xt_rsc_0_17_i_da_d;
  input [63:0] xt_rsc_0_17_i_qa_d;
  output [1:0] xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_18_i_adra_d;
  output [63:0] xt_rsc_0_18_i_da_d;
  input [63:0] xt_rsc_0_18_i_qa_d;
  output [1:0] xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_19_i_adra_d;
  output [63:0] xt_rsc_0_19_i_da_d;
  input [63:0] xt_rsc_0_19_i_qa_d;
  output [1:0] xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_20_i_adra_d;
  output [63:0] xt_rsc_0_20_i_da_d;
  input [63:0] xt_rsc_0_20_i_qa_d;
  output [1:0] xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_21_i_adra_d;
  output [63:0] xt_rsc_0_21_i_da_d;
  input [63:0] xt_rsc_0_21_i_qa_d;
  output [1:0] xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_22_i_adra_d;
  output [63:0] xt_rsc_0_22_i_da_d;
  input [63:0] xt_rsc_0_22_i_qa_d;
  output [1:0] xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_23_i_adra_d;
  output [63:0] xt_rsc_0_23_i_da_d;
  input [63:0] xt_rsc_0_23_i_qa_d;
  output [1:0] xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_24_i_adra_d;
  output [63:0] xt_rsc_0_24_i_da_d;
  input [63:0] xt_rsc_0_24_i_qa_d;
  output [1:0] xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_25_i_adra_d;
  output [63:0] xt_rsc_0_25_i_da_d;
  input [63:0] xt_rsc_0_25_i_qa_d;
  output [1:0] xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_26_i_adra_d;
  output [63:0] xt_rsc_0_26_i_da_d;
  input [63:0] xt_rsc_0_26_i_qa_d;
  output [1:0] xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_27_i_adra_d;
  output [63:0] xt_rsc_0_27_i_da_d;
  input [63:0] xt_rsc_0_27_i_qa_d;
  output [1:0] xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_28_i_adra_d;
  output [63:0] xt_rsc_0_28_i_da_d;
  input [63:0] xt_rsc_0_28_i_qa_d;
  output [1:0] xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_29_i_adra_d;
  output [63:0] xt_rsc_0_29_i_da_d;
  input [63:0] xt_rsc_0_29_i_qa_d;
  output [1:0] xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_30_i_adra_d;
  output [63:0] xt_rsc_0_30_i_da_d;
  input [63:0] xt_rsc_0_30_i_qa_d;
  output [1:0] xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [15:0] xt_rsc_0_31_i_adra_d;
  output [63:0] xt_rsc_0_31_i_da_d;
  input [63:0] xt_rsc_0_31_i_qa_d;
  output [1:0] xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_0_i_adra_d;
  input [63:0] twiddle_rsc_0_0_i_qa_d;
  output [1:0] twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_1_i_adra_d;
  input [63:0] twiddle_rsc_0_1_i_qa_d;
  output [1:0] twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_2_i_adra_d;
  input [63:0] twiddle_rsc_0_2_i_qa_d;
  output [1:0] twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_3_i_adra_d;
  input [63:0] twiddle_rsc_0_3_i_qa_d;
  output [1:0] twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_4_i_adra_d;
  input [63:0] twiddle_rsc_0_4_i_qa_d;
  output [1:0] twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_5_i_adra_d;
  input [63:0] twiddle_rsc_0_5_i_qa_d;
  output [1:0] twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_6_i_adra_d;
  input [63:0] twiddle_rsc_0_6_i_qa_d;
  output [1:0] twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_7_i_adra_d;
  input [63:0] twiddle_rsc_0_7_i_qa_d;
  output [1:0] twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_8_i_adra_d;
  input [63:0] twiddle_rsc_0_8_i_qa_d;
  output [1:0] twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_9_i_adra_d;
  input [63:0] twiddle_rsc_0_9_i_qa_d;
  output [1:0] twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_10_i_adra_d;
  input [63:0] twiddle_rsc_0_10_i_qa_d;
  output [1:0] twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_11_i_adra_d;
  input [63:0] twiddle_rsc_0_11_i_qa_d;
  output [1:0] twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_12_i_adra_d;
  input [63:0] twiddle_rsc_0_12_i_qa_d;
  output [1:0] twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_13_i_adra_d;
  input [63:0] twiddle_rsc_0_13_i_qa_d;
  output [1:0] twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_14_i_adra_d;
  input [63:0] twiddle_rsc_0_14_i_qa_d;
  output [1:0] twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_rsc_0_15_i_adra_d;
  input [63:0] twiddle_rsc_0_15_i_qa_d;
  output [1:0] twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_0_i_adra_d;
  input [63:0] twiddle_h_rsc_0_0_i_qa_d;
  output [1:0] twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_1_i_adra_d;
  input [63:0] twiddle_h_rsc_0_1_i_qa_d;
  output [1:0] twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_2_i_adra_d;
  input [63:0] twiddle_h_rsc_0_2_i_qa_d;
  output [1:0] twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_3_i_adra_d;
  input [63:0] twiddle_h_rsc_0_3_i_qa_d;
  output [1:0] twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_4_i_adra_d;
  input [63:0] twiddle_h_rsc_0_4_i_qa_d;
  output [1:0] twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_5_i_adra_d;
  input [63:0] twiddle_h_rsc_0_5_i_qa_d;
  output [1:0] twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_6_i_adra_d;
  input [63:0] twiddle_h_rsc_0_6_i_qa_d;
  output [1:0] twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_7_i_adra_d;
  input [63:0] twiddle_h_rsc_0_7_i_qa_d;
  output [1:0] twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_8_i_adra_d;
  input [63:0] twiddle_h_rsc_0_8_i_qa_d;
  output [1:0] twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_9_i_adra_d;
  input [63:0] twiddle_h_rsc_0_9_i_qa_d;
  output [1:0] twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_10_i_adra_d;
  input [63:0] twiddle_h_rsc_0_10_i_qa_d;
  output [1:0] twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_11_i_adra_d;
  input [63:0] twiddle_h_rsc_0_11_i_qa_d;
  output [1:0] twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_12_i_adra_d;
  input [63:0] twiddle_h_rsc_0_12_i_qa_d;
  output [1:0] twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_13_i_adra_d;
  input [63:0] twiddle_h_rsc_0_13_i_qa_d;
  output [1:0] twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_14_i_adra_d;
  input [63:0] twiddle_h_rsc_0_14_i_qa_d;
  output [1:0] twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [7:0] twiddle_h_rsc_0_15_i_adra_d;
  input [63:0] twiddle_h_rsc_0_15_i_qa_d;
  output [1:0] twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  output [1:0] yt_rsc_0_0_i_wea_d_pff;
  output [1:0] yt_rsc_0_16_i_wea_d_pff;
  output [1:0] xt_rsc_0_0_i_wea_d_pff;
  output [1:0] xt_rsc_0_16_i_wea_d_pff;


  // Interconnect Declarations
  wire [31:0] p_rsci_idat;
  wire mult_t_mul_cmp_en;
  wire [63:0] mult_t_mul_cmp_z;
  wire [63:0] mult_t_mul_cmp_1_z;
  wire [63:0] mult_t_mul_cmp_2_z;
  wire [63:0] mult_t_mul_cmp_3_z;
  wire [63:0] mult_t_mul_cmp_4_z;
  wire [63:0] mult_t_mul_cmp_5_z;
  wire [63:0] mult_t_mul_cmp_6_z;
  wire [63:0] mult_t_mul_cmp_7_z;
  wire [63:0] mult_t_mul_cmp_8_z;
  wire [63:0] mult_t_mul_cmp_9_z;
  wire [63:0] mult_t_mul_cmp_10_z;
  wire [63:0] mult_t_mul_cmp_11_z;
  wire [63:0] mult_t_mul_cmp_12_z;
  wire [63:0] mult_t_mul_cmp_13_z;
  wire [63:0] mult_t_mul_cmp_14_z;
  wire [63:0] mult_t_mul_cmp_15_z;
  wire [31:0] mult_z_mul_cmp_z;
  wire mult_z_mul_cmp_1_en;
  wire [31:0] mult_z_mul_cmp_1_z;
  wire [31:0] mult_z_mul_cmp_2_z;
  wire [31:0] mult_z_mul_cmp_3_z;
  wire [31:0] mult_z_mul_cmp_4_z;
  wire [31:0] mult_z_mul_cmp_5_z;
  wire [31:0] mult_z_mul_cmp_6_z;
  wire [31:0] mult_z_mul_cmp_7_z;
  wire [31:0] mult_z_mul_cmp_8_z;
  wire [31:0] mult_z_mul_cmp_9_z;
  wire [31:0] mult_z_mul_cmp_10_z;
  wire [31:0] mult_z_mul_cmp_11_z;
  wire [31:0] mult_z_mul_cmp_12_z;
  wire [31:0] mult_z_mul_cmp_13_z;
  wire [31:0] mult_z_mul_cmp_14_z;
  wire [31:0] mult_z_mul_cmp_15_z;
  wire [31:0] mult_z_mul_cmp_16_z;
  wire [31:0] mult_z_mul_cmp_17_z;
  wire [31:0] mult_z_mul_cmp_18_z;
  wire [31:0] mult_z_mul_cmp_19_z;
  wire [31:0] mult_z_mul_cmp_20_z;
  wire [31:0] mult_z_mul_cmp_21_z;
  wire [31:0] mult_z_mul_cmp_22_z;
  wire [31:0] mult_z_mul_cmp_23_z;
  wire [31:0] mult_z_mul_cmp_24_z;
  wire [31:0] mult_z_mul_cmp_25_z;
  wire [31:0] mult_z_mul_cmp_26_z;
  wire [31:0] mult_z_mul_cmp_27_z;
  wire [31:0] mult_z_mul_cmp_28_z;
  wire [31:0] mult_z_mul_cmp_29_z;
  wire [31:0] mult_z_mul_cmp_30_z;
  wire [31:0] mult_z_mul_cmp_31_z;
  wire [10:0] fsm_output;
  wire INNER_LOOP4_nor_tmp;
  wire or_dcpl_13;
  wire or_dcpl_22;
  wire or_dcpl_45;
  wire or_dcpl_65;
  wire or_dcpl_101;
  wire or_dcpl_121;
  wire and_dcpl_51;
  wire and_dcpl_56;
  wire and_dcpl_57;
  wire or_dcpl_194;
  wire and_dcpl_58;
  wire and_dcpl_59;
  wire or_dcpl_197;
  wire or_dcpl_198;
  wire or_dcpl_199;
  wire or_dcpl_200;
  wire and_dcpl_67;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_70;
  wire or_dcpl_205;
  wire or_dcpl_206;
  wire or_dcpl_207;
  wire or_dcpl_208;
  wire or_dcpl_210;
  wire or_dcpl_212;
  wire or_dcpl_214;
  wire and_dcpl_79;
  wire and_dcpl_81;
  wire and_dcpl_82;
  wire or_dcpl_217;
  wire or_dcpl_218;
  wire and_dcpl_90;
  wire or_dcpl_233;
  wire or_tmp_21;
  wire or_tmp_22;
  wire or_tmp_25;
  wire or_tmp_26;
  wire or_tmp_203;
  wire or_tmp_204;
  wire or_tmp_207;
  wire or_tmp_208;
  wire or_tmp_771;
  wire or_tmp_779;
  wire or_tmp_782;
  wire or_tmp_790;
  wire or_tmp_792;
  wire or_tmp_809;
  wire or_tmp_819;
  wire or_tmp_885;
  wire or_tmp_894;
  wire or_tmp_1134;
  wire or_tmp_1138;
  wire or_tmp_1189;
  wire and_167_cse;
  wire and_192_cse;
  wire and_1445_cse;
  wire and_1454_cse;
  wire and_1463_cse;
  wire and_1700_cse;
  wire and_1719_cse;
  wire and_1725_cse;
  wire and_1763_cse;
  wire and_1783_cse;
  reg [6:0] INNER_LOOP4_r_11_4_sva_6_0;
  reg [6:0] INNER_LOOP3_r_11_4_sva_6_0;
  reg [6:0] INNER_LOOP2_r_11_4_sva_6_0;
  reg [6:0] INNER_LOOP1_r_11_4_sva_6_0;
  reg [1:0] butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm;
  reg c_1_sva;
  reg INNER_LOOP1_stage_0_10;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10;
  reg INNER_LOOP1_stage_0;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8;
  reg INNER_LOOP1_stage_0_9;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm;
  reg INNER_LOOP1_stage_0_11;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7;
  reg [2:0] operator_20_false_acc_cse_sva;
  reg [1:0] operator_33_true_3_lshift_psp_1_0_sva;
  reg INNER_LOOP1_stage_0_4;
  reg INNER_LOOP1_stage_0_2;
  reg INNER_LOOP1_stage_0_3;
  reg INNER_LOOP1_stage_0_6;
  reg INNER_LOOP1_stage_0_7;
  reg INNER_LOOP1_stage_0_5;
  reg [31:0] p_sva;
  reg reg_yt_rsc_0_0_cgo_cse;
  reg reg_yt_rsc_0_16_cgo_cse;
  reg reg_xt_rsc_triosy_0_31_obj_ld_cse;
  reg reg_ensig_cgo_cse;
  wire mult_15_t_and_49_cse;
  wire mult_15_t_and_51_cse;
  wire mult_15_t_and_53_cse;
  wire mult_15_t_and_55_cse;
  wire mult_15_t_and_44_cse;
  wire mult_15_t_and_45_cse;
  wire mult_15_t_and_46_cse;
  wire mult_15_t_and_47_cse;
  wire mult_15_t_and_48_cse;
  wire mult_15_t_and_50_cse;
  wire mult_15_t_and_52_cse;
  wire mult_15_t_and_54_cse;
  reg reg_ensig_cgo_17_cse;
  wire butterFly1_or_5_cse;
  wire butterFly1_or_1_cse;
  wire butterFly1_mux_17_cse;
  wire butterFly1_or_4_cse;
  wire butterFly1_or_cse;
  wire [31:0] mult_15_res_sva_1;
  wire [32:0] nl_mult_15_res_sva_1;
  wire [31:0] mult_14_res_sva_1;
  wire [32:0] nl_mult_14_res_sva_1;
  wire [31:0] mult_13_res_sva_1;
  wire [32:0] nl_mult_13_res_sva_1;
  wire [31:0] mult_12_res_sva_1;
  wire [32:0] nl_mult_12_res_sva_1;
  wire [31:0] mult_11_res_sva_1;
  wire [32:0] nl_mult_11_res_sva_1;
  wire [31:0] mult_10_res_sva_1;
  wire [32:0] nl_mult_10_res_sva_1;
  wire [31:0] mult_9_res_sva_1;
  wire [32:0] nl_mult_9_res_sva_1;
  wire [31:0] mult_8_res_sva_1;
  wire [32:0] nl_mult_8_res_sva_1;
  wire [31:0] mult_7_res_sva_1;
  wire [32:0] nl_mult_7_res_sva_1;
  wire [31:0] mult_6_res_sva_1;
  wire [32:0] nl_mult_6_res_sva_1;
  wire [31:0] mult_5_res_sva_1;
  wire [32:0] nl_mult_5_res_sva_1;
  wire [31:0] mult_4_res_sva_1;
  wire [32:0] nl_mult_4_res_sva_1;
  wire [31:0] mult_3_res_sva_1;
  wire [32:0] nl_mult_3_res_sva_1;
  wire [31:0] mult_2_res_sva_1;
  wire [32:0] nl_mult_2_res_sva_1;
  wire [31:0] mult_1_res_sva_1;
  wire [32:0] nl_mult_1_res_sva_1;
  wire [31:0] mult_res_sva_1;
  wire [32:0] nl_mult_res_sva_1;
  wire butterFly2_7_tw_nor_cse;
  wire butterFly2_7_tw_nor_1_cse;
  wire butterFly2_7_tw_nor_2_cse;
  wire mult_15_t_or_9_cse;
  wire mult_15_t_or_10_cse;
  wire mult_15_t_or_11_cse;
  wire mult_15_t_or_12_cse;
  wire mult_15_t_and_41_cse;
  wire mult_15_t_and_42_cse;
  wire mult_15_t_and_43_cse;
  wire mult_15_t_and_37_cse;
  wire mult_15_t_and_38_cse;
  wire mult_15_t_and_39_cse;
  wire mult_15_t_and_30_cse;
  wire mult_15_t_and_31_cse;
  wire mult_15_t_and_32_cse;
  wire mult_15_t_or_3_cse;
  wire mult_15_t_and_40_cse;
  wire mult_15_t_and_36_cse;
  wire mult_15_t_and_29_cse;
  wire nor_7_cse;
  wire mult_15_t_or_1_cse;
  wire mult_15_t_or_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse;
  reg [5:0] reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse;
  wire or_261_rmff;
  wire butterFly1_nor_7_rmff;
  wire butterFly1_butterFly1_or_1_rmff;
  wire [5:0] butterFly1_butterFly1_mux_3_rmff;
  wire butterFly1_butterFly1_and_17_rmff;
  wire [5:0] butterFly1_mux1h_15_rmff;
  wire and_202_rmff;
  wire [5:0] butterFly1_1_butterFly1_1_mux_3_rmff;
  wire [5:0] butterFly1_1_mux1h_11_rmff;
  wire [5:0] butterFly1_2_butterFly1_2_mux_3_rmff;
  wire [5:0] butterFly1_2_mux1h_11_rmff;
  wire [5:0] butterFly1_3_butterFly1_3_mux_3_rmff;
  wire [5:0] butterFly1_3_mux1h_11_rmff;
  wire [5:0] butterFly1_4_butterFly1_4_mux_3_rmff;
  wire [5:0] butterFly1_4_mux1h_11_rmff;
  wire [5:0] butterFly1_7_butterFly1_7_mux_3_rmff;
  wire [5:0] butterFly1_8_butterFly1_8_mux_3_rmff;
  wire [5:0] butterFly1_8_mux1h_11_rmff;
  wire or_443_rmff;
  wire butterFly1_nor_4_rmff;
  wire butterFly1_butterFly1_or_rmff;
  wire [5:0] butterFly1_butterFly1_mux_4_rmff;
  wire butterFly1_butterFly1_and_15_rmff;
  wire [5:0] butterFly1_mux1h_13_rmff;
  wire [5:0] butterFly1_1_butterFly1_1_mux_4_rmff;
  wire [5:0] butterFly1_1_mux1h_9_rmff;
  wire [5:0] butterFly1_2_butterFly1_2_mux_4_rmff;
  wire [5:0] butterFly1_2_mux1h_9_rmff;
  wire [5:0] butterFly1_3_butterFly1_3_mux_4_rmff;
  wire [5:0] butterFly1_3_mux1h_9_rmff;
  wire [5:0] butterFly1_4_butterFly1_4_mux_4_rmff;
  wire [5:0] butterFly1_4_mux1h_9_rmff;
  wire [5:0] butterFly1_7_butterFly1_7_mux_4_rmff;
  wire [5:0] butterFly1_8_butterFly1_8_mux_4_rmff;
  wire [5:0] butterFly1_8_mux1h_9_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_65_rmff;
  wire [31:0] butterFly1_f1_butterFly1_f1_mux_2_rmff;
  wire [31:0] butterFly1_f1_butterFly1_f1_mux_3_rmff;
  wire butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff;
  wire and_921_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_64_rmff;
  wire [31:0] butterFly1_f2_butterFly1_f2_mux_2_rmff;
  wire [31:0] butterFly1_f2_butterFly1_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_63_rmff;
  wire [31:0] butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff;
  wire [31:0] butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_62_rmff;
  wire [31:0] butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff;
  wire [31:0] butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_61_rmff;
  wire [31:0] butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff;
  wire [31:0] butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_60_rmff;
  wire [31:0] butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff;
  wire [31:0] butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_59_rmff;
  wire [31:0] butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff;
  wire [31:0] butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_58_rmff;
  wire [31:0] butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff;
  wire [31:0] butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_57_rmff;
  wire [31:0] butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff;
  wire [31:0] butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_56_rmff;
  wire [31:0] butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff;
  wire [31:0] butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_55_rmff;
  wire [31:0] butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff;
  wire [31:0] butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_54_rmff;
  wire [31:0] butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff;
  wire [31:0] butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_53_rmff;
  wire [31:0] butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff;
  wire [31:0] butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_52_rmff;
  wire [31:0] butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff;
  wire [31:0] butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_51_rmff;
  wire [31:0] butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff;
  wire [31:0] butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff;
  wire [6:0] butterFly1_15_f2_mux1h_50_rmff;
  wire [31:0] butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff;
  wire [31:0] butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff;
  wire butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff;
  wire [6:0] INNER_LOOP1_tw_h_mux1h_4_rmff;
  wire and_1435_rmff;
  wire [6:0] butterFly2_1_tw_butterFly2_1_tw_mux_rmff;
  wire or_896_rmff;
  wire or_900_rmff;
  wire or_904_rmff;
  wire or_908_rmff;
  wire or_912_rmff;
  wire or_916_rmff;
  wire or_920_rmff;
  wire and_1506_rmff;
  wire or_997_rmff;
  wire or_1156_rmff;
  wire [31:0] mult_4_t_mux1h_1_rmff;
  wire [31:0] yt_rsc_0_15_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_15_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_15_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_31_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_14_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_14_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_14_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_30_qr_lpi_3_dfm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1;
  wire [31:0] yt_rsc_0_13_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_13_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_13_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_29_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_12_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_12_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_12_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_28_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_11_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_11_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_11_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_27_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_10_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_10_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_10_qr_lpi_3_dfm_1;
  reg [31:0] modulo_add_26_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_9_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_9_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_25_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_8_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_8_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_24_qr_lpi_3_dfm_1;
  wire [31:0] yt_rsc_0_7_i_da_d_mx0w0_63_32;
  reg [31:0] modulo_add_23_qr_lpi_3_dfm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9;
  wire [31:0] yt_rsc_0_6_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_6_i_da_d_mx0w2_63_32;
  reg [31:0] modulo_add_1_qr_lpi_3_dfm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1;
  wire [31:0] yt_rsc_0_5_i_da_d_mx0w2_63_32;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1;
  wire [31:0] yt_rsc_0_4_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_4_i_da_d_mx0w2_63_32;
  wire [31:0] yt_rsc_0_3_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_3_i_da_d_mx0w2_63_32;
  wire [31:0] yt_rsc_0_2_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_2_i_da_d_mx0w2_63_32;
  wire [31:0] yt_rsc_0_1_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_1_i_da_d_mx0w2_63_32;
  wire [31:0] yt_rsc_0_0_i_da_d_mx0w0_63_32;
  wire [31:0] yt_rsc_0_0_i_da_d_mx0w2_63_32;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8;
  wire yt_rsc_0_0_i_wea_d_mx0c2;
  wire yt_rsc_0_0_i_wea_d_mx0c0;
  wire yt_rsc_0_16_i_wea_d_mx0c2;
  wire yt_rsc_0_16_i_wea_d_mx0c0;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2;
  wire [10:0] z_out;
  wire [2:0] z_out_1;
  wire [3:0] nl_z_out_1;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  wire [31:0] z_out_4;
  wire [32:0] nl_z_out_4;
  wire [31:0] z_out_5;
  wire [32:0] nl_z_out_5;
  wire [31:0] z_out_8;
  wire [32:0] nl_z_out_8;
  wire [31:0] z_out_9;
  wire [32:0] nl_z_out_9;
  wire [31:0] z_out_10;
  wire [32:0] nl_z_out_10;
  wire [31:0] z_out_12;
  wire [32:0] nl_z_out_12;
  wire [31:0] z_out_13;
  wire [32:0] nl_z_out_13;
  wire [31:0] z_out_14;
  wire [32:0] nl_z_out_14;
  wire [31:0] z_out_16;
  wire [32:0] nl_z_out_16;
  wire [31:0] z_out_17;
  wire [32:0] nl_z_out_17;
  wire [31:0] z_out_18;
  wire [32:0] nl_z_out_18;
  wire [31:0] z_out_20;
  wire [32:0] nl_z_out_20;
  wire [31:0] z_out_21;
  wire [32:0] nl_z_out_21;
  wire [31:0] z_out_22;
  wire [32:0] nl_z_out_22;
  wire [31:0] z_out_24;
  wire [32:0] nl_z_out_24;
  wire [31:0] z_out_25;
  wire [32:0] nl_z_out_25;
  wire [31:0] z_out_26;
  wire [32:0] nl_z_out_26;
  wire [31:0] z_out_28;
  wire [32:0] nl_z_out_28;
  wire [31:0] z_out_29;
  wire [32:0] nl_z_out_29;
  wire [31:0] z_out_31;
  wire [32:0] nl_z_out_31;
  wire [31:0] z_out_32;
  wire [32:0] nl_z_out_32;
  wire [31:0] z_out_34;
  wire [32:0] nl_z_out_34;
  wire [31:0] z_out_36;
  wire [32:0] nl_z_out_36;
  wire [31:0] z_out_37;
  wire [32:0] nl_z_out_37;
  wire [31:0] z_out_39;
  wire [32:0] nl_z_out_39;
  wire [31:0] z_out_41;
  wire [32:0] nl_z_out_41;
  wire [31:0] z_out_42;
  wire [32:0] nl_z_out_42;
  wire [31:0] z_out_44;
  wire [32:0] nl_z_out_44;
  wire [31:0] z_out_46;
  wire [32:0] nl_z_out_46;
  wire [31:0] z_out_47;
  wire [32:0] nl_z_out_47;
  wire [31:0] z_out_49;
  wire [32:0] nl_z_out_49;
  wire [31:0] z_out_51;
  wire [31:0] z_out_52;
  wire [31:0] z_out_53;
  wire [31:0] z_out_54;
  wire [31:0] z_out_55;
  wire [31:0] z_out_56;
  wire [31:0] z_out_57;
  wire [31:0] z_out_58;
  wire [31:0] z_out_59;
  wire [31:0] z_out_60;
  wire [31:0] z_out_61;
  wire [31:0] z_out_62;
  wire [31:0] z_out_63;
  wire [31:0] z_out_64;
  wire [31:0] z_out_65;
  wire [31:0] z_out_66;
  wire [31:0] z_out_67;
  wire [32:0] nl_z_out_67;
  wire [31:0] z_out_68;
  wire [32:0] nl_z_out_68;
  wire [31:0] z_out_69;
  wire [32:0] nl_z_out_69;
  wire [31:0] z_out_70;
  wire [32:0] nl_z_out_70;
  wire [31:0] z_out_71;
  wire [32:0] nl_z_out_71;
  wire [31:0] z_out_72;
  wire [32:0] nl_z_out_72;
  wire [31:0] z_out_73;
  wire [32:0] nl_z_out_73;
  wire [31:0] z_out_74;
  wire [32:0] nl_z_out_74;
  wire [31:0] z_out_75;
  wire [32:0] nl_z_out_75;
  wire [31:0] z_out_76;
  wire [32:0] nl_z_out_76;
  wire [31:0] z_out_77;
  wire [32:0] nl_z_out_77;
  wire [31:0] z_out_78;
  wire [32:0] nl_z_out_78;
  wire [31:0] z_out_79;
  wire [32:0] nl_z_out_79;
  wire [31:0] z_out_80;
  wire [32:0] nl_z_out_80;
  wire [31:0] z_out_81;
  wire [32:0] nl_z_out_81;
  wire [31:0] z_out_82;
  wire [32:0] nl_z_out_82;
  reg [5:0] operator_33_true_1_lshift_psp_9_4_sva;
  reg INNER_LOOP1_stage_0_8;
  reg [31:0] mult_res_lpi_3_dfm_1;
  reg [31:0] mult_1_res_lpi_3_dfm_1;
  reg [31:0] mult_2_res_lpi_3_dfm_1;
  reg [31:0] mult_3_res_lpi_3_dfm_1;
  reg [31:0] mult_4_res_lpi_3_dfm_1;
  reg [31:0] mult_5_res_lpi_3_dfm_1;
  reg [31:0] mult_6_res_lpi_3_dfm_1;
  reg [31:0] mult_7_res_lpi_3_dfm_1;
  reg [31:0] mult_8_res_lpi_3_dfm_1;
  reg [31:0] mult_9_res_lpi_3_dfm_1;
  reg [31:0] mult_10_res_lpi_3_dfm_1;
  reg [31:0] mult_11_res_lpi_3_dfm_1;
  reg [31:0] mult_12_res_lpi_3_dfm_1;
  reg [31:0] mult_13_res_lpi_3_dfm_1;
  reg [31:0] mult_14_res_lpi_3_dfm_1;
  reg [31:0] mult_15_res_lpi_3_dfm_1;
  reg [31:0] mult_1_z_asn_itm_1;
  reg [31:0] mult_1_z_asn_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_7;
  reg [31:0] mult_10_z_asn_itm_1;
  reg [31:0] mult_10_z_asn_itm_2;
  reg [31:0] mult_10_z_asn_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_7;
  reg [31:0] mult_11_z_asn_itm_1;
  reg [31:0] mult_11_z_asn_itm_2;
  reg [31:0] mult_11_z_asn_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_7;
  reg [31:0] mult_12_z_asn_itm_1;
  reg [31:0] mult_12_z_asn_itm_2;
  reg [31:0] mult_12_z_asn_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_7;
  reg [31:0] mult_13_z_asn_itm_1;
  reg [31:0] mult_13_z_asn_itm_2;
  reg [31:0] mult_13_z_asn_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_7;
  reg [31:0] mult_14_z_asn_itm_1;
  reg [31:0] mult_14_z_asn_itm_2;
  reg [31:0] mult_14_z_asn_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_1;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_7;
  reg [31:0] mult_15_z_asn_itm_1;
  reg [31:0] mult_15_z_asn_itm_2;
  reg [31:0] mult_15_z_asn_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_7;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_8;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_2;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_3;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_4;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_5;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_6;
  reg [5:0] INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_7;
  reg INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2;
  reg [31:0] tmp_10_sva_1;
  reg [31:0] tmp_10_sva_2;
  reg [31:0] tmp_10_sva_3;
  reg [31:0] tmp_10_sva_4;
  reg [31:0] tmp_10_sva_5;
  reg [31:0] tmp_10_sva_6;
  reg [31:0] tmp_10_sva_7;
  reg [31:0] mult_16_z_asn_itm_3;
  reg [31:0] mult_17_z_asn_itm_3;
  reg [31:0] mult_18_z_asn_itm_3;
  reg [31:0] mult_19_z_asn_itm_3;
  reg [31:0] mult_20_z_asn_itm_3;
  reg [31:0] mult_21_z_asn_itm_3;
  reg [31:0] mult_22_z_asn_itm_3;
  reg [31:0] mult_23_z_asn_itm_1;
  reg [31:0] mult_23_z_asn_itm_2;
  reg [31:0] mult_23_z_asn_itm_3;
  reg [31:0] mult_24_z_asn_itm_1;
  reg [31:0] mult_24_z_asn_itm_2;
  reg [31:0] mult_24_z_asn_itm_3;
  reg [31:0] mult_25_z_asn_itm_1;
  reg [31:0] mult_25_z_asn_itm_2;
  reg [31:0] mult_25_z_asn_itm_3;
  reg [31:0] mult_26_z_asn_itm_1;
  reg [31:0] mult_26_z_asn_itm_2;
  reg [31:0] mult_27_z_asn_itm_1;
  reg [31:0] mult_27_z_asn_itm_2;
  reg [31:0] mult_28_z_asn_itm_1;
  reg [31:0] mult_28_z_asn_itm_2;
  reg [31:0] mult_29_z_asn_itm_1;
  reg [31:0] mult_29_z_asn_itm_2;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_3;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_4;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_5;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_6;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_7;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_8;
  reg [31:0] mult_30_z_asn_itm_1;
  reg [31:0] mult_30_z_asn_itm_2;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_1;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_2;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_3;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_4;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_5;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_6;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_7;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_8;
  reg [5:0] INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9;
  reg [31:0] mult_31_z_asn_itm_1;
  reg [31:0] mult_31_z_asn_itm_2;
  reg [31:0] tmp_102_sva_1;
  reg [31:0] tmp_102_sva_2;
  reg [31:0] tmp_102_sva_3;
  reg [31:0] tmp_102_sva_4;
  reg [31:0] tmp_102_sva_5;
  reg [31:0] tmp_102_sva_6;
  reg [31:0] tmp_102_sva_7;
  reg [31:0] tmp_104_sva_1;
  reg [31:0] tmp_104_sva_2;
  reg [31:0] tmp_104_sva_3;
  reg [31:0] tmp_104_sva_4;
  reg [31:0] tmp_104_sva_5;
  reg [31:0] tmp_104_sva_6;
  reg [31:0] tmp_104_sva_7;
  reg [31:0] tmp_106_sva_1;
  reg [31:0] tmp_106_sva_2;
  reg [31:0] tmp_106_sva_3;
  reg [31:0] tmp_106_sva_4;
  reg [31:0] tmp_106_sva_5;
  reg [31:0] tmp_106_sva_6;
  reg [31:0] tmp_106_sva_7;
  reg [31:0] tmp_108_sva_1;
  reg [31:0] tmp_108_sva_2;
  reg [31:0] tmp_108_sva_3;
  reg [31:0] tmp_108_sva_4;
  reg [31:0] tmp_108_sva_5;
  reg [31:0] tmp_108_sva_6;
  reg [31:0] tmp_108_sva_7;
  reg [31:0] tmp_110_sva_1;
  reg [31:0] tmp_110_sva_2;
  reg [31:0] tmp_110_sva_3;
  reg [31:0] tmp_110_sva_4;
  reg [31:0] tmp_110_sva_5;
  reg [31:0] tmp_110_sva_6;
  reg [31:0] tmp_110_sva_7;
  reg [31:0] tmp_112_sva_1;
  reg [31:0] tmp_112_sva_2;
  reg [31:0] tmp_112_sva_3;
  reg [31:0] tmp_112_sva_4;
  reg [31:0] tmp_112_sva_5;
  reg [31:0] tmp_112_sva_6;
  reg [31:0] tmp_112_sva_7;
  reg [31:0] tmp_114_sva_1;
  reg [31:0] tmp_114_sva_2;
  reg [31:0] tmp_114_sva_3;
  reg [31:0] tmp_114_sva_4;
  reg [31:0] tmp_114_sva_5;
  reg [31:0] tmp_114_sva_6;
  reg [31:0] tmp_114_sva_7;
  reg [31:0] tmp_116_sva_1;
  reg [31:0] tmp_116_sva_2;
  reg [31:0] tmp_116_sva_3;
  reg [31:0] tmp_116_sva_4;
  reg [31:0] tmp_116_sva_5;
  reg [31:0] tmp_116_sva_6;
  reg [31:0] tmp_116_sva_7;
  reg [31:0] tmp_118_sva_1;
  reg [31:0] tmp_118_sva_2;
  reg [31:0] tmp_118_sva_3;
  reg [31:0] tmp_118_sva_4;
  reg [31:0] tmp_118_sva_5;
  reg [31:0] tmp_118_sva_6;
  reg [31:0] tmp_118_sva_7;
  reg [31:0] tmp_120_sva_1;
  reg [31:0] tmp_120_sva_2;
  reg [31:0] tmp_120_sva_3;
  reg [31:0] tmp_120_sva_4;
  reg [31:0] tmp_120_sva_5;
  reg [31:0] tmp_120_sva_6;
  reg [31:0] tmp_120_sva_7;
  reg [31:0] tmp_122_sva_1;
  reg [31:0] tmp_122_sva_2;
  reg [31:0] tmp_122_sva_3;
  reg [31:0] tmp_122_sva_4;
  reg [31:0] tmp_122_sva_5;
  reg [31:0] tmp_122_sva_6;
  reg [31:0] tmp_122_sva_7;
  reg [31:0] tmp_124_sva_1;
  reg [31:0] tmp_124_sva_2;
  reg [31:0] tmp_124_sva_3;
  reg [31:0] tmp_124_sva_4;
  reg [31:0] tmp_124_sva_5;
  reg [31:0] tmp_124_sva_6;
  reg [31:0] tmp_124_sva_7;
  reg [31:0] tmp_126_sva_1;
  reg [31:0] tmp_126_sva_2;
  reg [31:0] tmp_126_sva_3;
  reg [31:0] tmp_126_sva_4;
  reg [31:0] tmp_126_sva_5;
  reg [31:0] tmp_126_sva_6;
  reg [31:0] tmp_126_sva_7;
  reg butterFly2_15_tw_equal_tmp_1;
  reg butterFly2_15_tw_equal_tmp_3_1;
  reg butterFly2_15_tw_equal_tmp_5_1;
  reg butterFly2_15_tw_equal_tmp_6_1;
  reg butterFly2_15_tw_equal_tmp_7_1;
  reg [31:0] tmp_60_sva_1;
  reg [31:0] tmp_60_sva_2;
  reg [31:0] tmp_60_sva_3;
  reg [31:0] tmp_60_sva_4;
  reg [31:0] tmp_60_sva_5;
  reg [31:0] tmp_60_sva_6;
  reg [31:0] tmp_60_sva_7;
  reg [31:0] tmp_62_sva_1;
  reg [31:0] tmp_62_sva_2;
  reg [31:0] tmp_62_sva_3;
  reg [31:0] tmp_62_sva_4;
  reg [31:0] tmp_62_sva_5;
  reg [31:0] tmp_62_sva_6;
  reg [31:0] tmp_62_sva_7;
  wire [1:0] operator_33_true_3_lshift_psp_1_0_sva_mx0w3;
  wire [31:0] mult_15_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_14_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_13_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_12_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_11_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_10_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_9_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_8_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_7_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_6_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_5_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_4_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_3_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_2_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_1_res_lpi_3_dfm_1_mx0;
  wire [31:0] mult_res_lpi_3_dfm_1_mx0;
  wire modulo_sub_31_qelse_and_ssc;
  wire modulo_sub_31_qelse_and_ssc_1;
  reg reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_30_qelse_and_ssc;
  wire modulo_sub_30_qelse_and_ssc_1;
  reg reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_29_qelse_and_ssc;
  wire modulo_sub_29_qelse_and_ssc_1;
  reg reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_28_qelse_and_ssc;
  wire modulo_sub_28_qelse_and_ssc_1;
  reg reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_27_qelse_and_ssc;
  wire modulo_sub_27_qelse_and_ssc_1;
  reg reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_26_qelse_and_ssc;
  wire modulo_sub_26_qelse_and_ssc_1;
  reg reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_25_qelse_and_ssc;
  wire modulo_sub_25_qelse_and_ssc_1;
  reg reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_24_qelse_and_ssc;
  wire modulo_sub_24_qelse_and_ssc_1;
  reg reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_23_qelse_and_ssc;
  wire modulo_sub_23_qelse_and_ssc_1;
  reg reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_22_qelse_and_ssc;
  wire modulo_sub_22_qelse_and_ssc_1;
  reg reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_21_qelse_and_ssc;
  wire modulo_sub_21_qelse_and_ssc_1;
  reg reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_20_qelse_and_ssc;
  wire modulo_sub_20_qelse_and_ssc_1;
  reg reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_19_qelse_and_ssc;
  wire modulo_sub_19_qelse_and_ssc_1;
  reg reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_18_qelse_and_ssc;
  wire modulo_sub_18_qelse_and_ssc_1;
  reg reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_17_qelse_and_ssc;
  wire modulo_sub_17_qelse_and_ssc_1;
  reg reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_sub_16_qelse_and_ssc;
  wire modulo_sub_16_qelse_and_ssc_1;
  reg reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd;
  reg [30:0] reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1;
  wire modulo_add_1_qelse_or_m1c;
  reg [31:0] reg_mult_17_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_25_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_28_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_20_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_22_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_30_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_26_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_18_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_19_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_23_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_27_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_31_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_29_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_24_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_21_res_lpi_3_dfm_1_cse;
  reg [31:0] reg_mult_16_res_lpi_3_dfm_1_cse;
  wire or_12_cse;
  wire or_44_cse;
  wire or_64_cse;
  wire or_84_cse;
  wire or_103_cse;
  wire or_123_cse;
  wire or_143_cse;
  wire or_142_cse;
  wire [31:0] modulo_sub_5_qelse_mux_cse;
  wire z_out_83_32;
  wire z_out_84_32;
  wire z_out_85_32;
  wire z_out_86_32;
  wire z_out_87_32;
  wire z_out_88_32;
  wire z_out_89_32;
  wire z_out_90_32;
  wire z_out_91_32;
  wire z_out_92_32;
  wire z_out_93_32;
  wire z_out_94_32;
  wire z_out_95_32;
  wire z_out_96_32;
  wire z_out_97_32;
  wire z_out_98_32;

  wire[0:0] c_mux_nl;
  wire[0:0] butterFly2_21_tw_butterFly2_21_tw_or_nl;
  wire[1:0] STAGE_LOOP_mux1h_nl;
  wire[0:0] STAGE_LOOP_and_nl;
  wire[0:0] nor_4_nl;
  wire[0:0] INNER_LOOP1_r_mux_44_nl;
  wire[32:0] acc_2_nl;
  wire[33:0] nl_acc_2_nl;
  wire[31:0] modulo_add_1_qif_mux1h_2_nl;
  wire[0:0] modulo_add_1_qelse_and_nl;
  wire[0:0] modulo_add_1_qelse_or_1_nl;
  wire[0:0] modulo_add_1_qelse_and_4_nl;
  wire[0:0] modulo_add_1_qelse_and_5_nl;
  wire[32:0] acc_6_nl;
  wire[33:0] nl_acc_6_nl;
  wire[31:0] modulo_add_10_qif_mux1h_2_nl;
  wire[0:0] modulo_add_10_qelse_and_nl;
  wire[0:0] modulo_add_10_qelse_or_nl;
  wire[0:0] modulo_add_10_qelse_and_5_nl;
  wire[0:0] modulo_add_10_qelse_and_6_nl;
  wire[0:0] modulo_add_10_qelse_and_7_nl;
  wire[32:0] acc_10_nl;
  wire[33:0] nl_acc_10_nl;
  wire[31:0] modulo_add_11_qif_mux1h_2_nl;
  wire[0:0] modulo_add_11_qelse_and_nl;
  wire[0:0] modulo_add_11_qelse_or_nl;
  wire[0:0] modulo_add_11_qelse_and_5_nl;
  wire[0:0] modulo_add_11_qelse_and_6_nl;
  wire[0:0] modulo_add_11_qelse_and_7_nl;
  wire[32:0] acc_14_nl;
  wire[33:0] nl_acc_14_nl;
  wire[31:0] modulo_add_12_qif_mux1h_2_nl;
  wire[0:0] modulo_add_12_qelse_and_nl;
  wire[0:0] modulo_add_12_qelse_or_1_nl;
  wire[0:0] modulo_add_12_qelse_and_4_nl;
  wire[0:0] modulo_add_12_qelse_and_5_nl;
  wire[32:0] acc_18_nl;
  wire[33:0] nl_acc_18_nl;
  wire[31:0] modulo_add_13_qif_mux1h_2_nl;
  wire[0:0] modulo_add_13_qelse_and_nl;
  wire[0:0] modulo_add_13_qelse_or_1_nl;
  wire[0:0] modulo_add_13_qelse_and_4_nl;
  wire[0:0] modulo_add_13_qelse_and_5_nl;
  wire[32:0] acc_22_nl;
  wire[33:0] nl_acc_22_nl;
  wire[31:0] modulo_add_14_qif_mux1h_2_nl;
  wire[0:0] modulo_add_14_qelse_and_nl;
  wire[0:0] modulo_add_14_qelse_or_1_nl;
  wire[0:0] modulo_add_14_qelse_and_4_nl;
  wire[0:0] modulo_add_14_qelse_and_5_nl;
  wire[32:0] acc_26_nl;
  wire[33:0] nl_acc_26_nl;
  wire[31:0] modulo_add_15_qif_mux1h_2_nl;
  wire[0:0] modulo_add_15_qelse_and_nl;
  wire[0:0] modulo_add_15_qelse_or_nl;
  wire[0:0] modulo_add_15_qelse_and_5_nl;
  wire[0:0] modulo_add_15_qelse_and_6_nl;
  wire[0:0] modulo_add_15_qelse_and_7_nl;
  wire[0:0] INNER_LOOP1_r_mux_45_nl;
  wire[0:0] INNER_LOOP1_mux_nl;
  wire[0:0] INNER_LOOP1_r_mux1h_46_nl;
  wire[0:0] INNER_LOOP1_r_INNER_LOOP1_r_and_1_nl;
  wire[0:0] INNER_LOOP1_r_INNER_LOOP1_r_and_3_nl;
  wire[0:0] or_1465_nl;
  wire[0:0] INNER_LOOP1_mux_11_nl;
  wire[0:0] INNER_LOOP1_r_INNER_LOOP1_r_and_2_nl;
  wire[0:0] INNER_LOOP1_r_INNER_LOOP1_r_and_nl;
  wire[6:0] STAGE_LOOP_base_STAGE_LOOP_base_mux_nl;
  wire[0:0] INNER_LOOP2_r_or_nl;
  wire[32:0] acc_29_nl;
  wire[33:0] nl_acc_29_nl;
  wire[31:0] modulo_add_2_qif_mux1h_2_nl;
  wire[0:0] modulo_add_23_qelse_and_nl;
  wire[0:0] modulo_add_23_qelse_or_1_nl;
  wire[0:0] modulo_add_23_qelse_and_4_nl;
  wire[0:0] modulo_add_23_qelse_and_5_nl;
  wire[32:0] acc_32_nl;
  wire[33:0] nl_acc_32_nl;
  wire[31:0] modulo_add_3_qif_mux1h_2_nl;
  wire[0:0] modulo_add_24_qelse_and_nl;
  wire[0:0] modulo_add_24_qelse_or_1_nl;
  wire[0:0] modulo_add_24_qelse_and_4_nl;
  wire[0:0] modulo_add_24_qelse_and_5_nl;
  wire[32:0] acc_34_nl;
  wire[33:0] nl_acc_34_nl;
  wire[31:0] modulo_add_4_qif_mux1h_2_nl;
  wire[0:0] modulo_add_25_qelse_and_nl;
  wire[0:0] modulo_add_25_qelse_or_1_nl;
  wire[0:0] modulo_add_25_qelse_and_4_nl;
  wire[0:0] modulo_add_25_qelse_and_5_nl;
  wire[32:0] acc_37_nl;
  wire[33:0] nl_acc_37_nl;
  wire[31:0] modulo_add_5_qif_mux1h_2_nl;
  wire[0:0] modulo_add_26_qelse_and_nl;
  wire[0:0] modulo_add_26_qelse_or_nl;
  wire[0:0] modulo_add_26_qelse_and_5_nl;
  wire[0:0] modulo_add_26_qelse_and_6_nl;
  wire[0:0] modulo_add_26_qelse_and_7_nl;
  wire[32:0] acc_39_nl;
  wire[33:0] nl_acc_39_nl;
  wire[31:0] modulo_add_6_qif_mux1h_2_nl;
  wire[0:0] modulo_add_27_qelse_and_nl;
  wire[0:0] modulo_add_27_qelse_or_nl;
  wire[0:0] modulo_add_27_qelse_and_5_nl;
  wire[0:0] modulo_add_27_qelse_and_6_nl;
  wire[0:0] modulo_add_27_qelse_and_7_nl;
  wire[32:0] acc_42_nl;
  wire[33:0] nl_acc_42_nl;
  wire[31:0] modulo_add_7_qif_mux1h_2_nl;
  wire[0:0] modulo_add_28_qelse_and_nl;
  wire[0:0] modulo_add_28_qelse_or_nl;
  wire[0:0] modulo_add_28_qelse_and_5_nl;
  wire[0:0] modulo_add_28_qelse_and_6_nl;
  wire[0:0] modulo_add_28_qelse_and_7_nl;
  wire[32:0] acc_44_nl;
  wire[33:0] nl_acc_44_nl;
  wire[31:0] modulo_add_8_qif_mux1h_2_nl;
  wire[0:0] modulo_add_29_qelse_and_nl;
  wire[0:0] modulo_add_29_qelse_or_nl;
  wire[0:0] modulo_add_29_qelse_and_5_nl;
  wire[0:0] modulo_add_29_qelse_and_6_nl;
  wire[0:0] modulo_add_29_qelse_and_7_nl;
  wire[32:0] acc_47_nl;
  wire[33:0] nl_acc_47_nl;
  wire[31:0] modulo_add_9_qif_mux1h_2_nl;
  wire[0:0] modulo_add_30_qelse_and_nl;
  wire[0:0] modulo_add_30_qelse_or_nl;
  wire[0:0] modulo_add_30_qelse_and_5_nl;
  wire[0:0] modulo_add_30_qelse_and_6_nl;
  wire[0:0] modulo_add_30_qelse_and_7_nl;
  wire[32:0] acc_49_nl;
  wire[33:0] nl_acc_49_nl;
  wire[31:0] modulo_add_qif_mux1h_2_nl;
  wire[0:0] modulo_add_31_qelse_and_nl;
  wire[0:0] modulo_add_31_qelse_or_nl;
  wire[0:0] modulo_add_31_qelse_and_5_nl;
  wire[0:0] modulo_add_31_qelse_and_6_nl;
  wire[0:0] modulo_add_31_qelse_and_7_nl;
  wire[0:0] modulo_sub_16_qelse_or_nl;
  wire[0:0] modulo_sub_17_qelse_or_nl;
  wire[0:0] modulo_sub_18_qelse_or_nl;
  wire[0:0] modulo_sub_19_qelse_or_nl;
  wire[0:0] modulo_sub_20_qelse_or_nl;
  wire[0:0] modulo_sub_21_qelse_or_nl;
  wire[0:0] modulo_sub_22_qelse_or_nl;
  wire[0:0] modulo_sub_23_qelse_or_nl;
  wire[0:0] modulo_sub_24_qelse_or_nl;
  wire[0:0] modulo_sub_25_qelse_or_nl;
  wire[0:0] modulo_sub_26_qelse_or_nl;
  wire[0:0] modulo_sub_27_qelse_or_nl;
  wire[0:0] modulo_sub_28_qelse_or_nl;
  wire[0:0] modulo_sub_29_qelse_or_nl;
  wire[0:0] modulo_sub_30_qelse_or_nl;
  wire[0:0] modulo_sub_31_qelse_or_nl;
  wire[31:0] modulo_sub_5_qif_acc_nl;
  wire[32:0] nl_modulo_sub_5_qif_acc_nl;
  wire[31:0] mult_15_if_acc_nl;
  wire[32:0] nl_mult_15_if_acc_nl;
  wire[32:0] mult_31_acc_1_nl;
  wire[33:0] nl_mult_31_acc_1_nl;
  wire[31:0] mult_14_if_acc_nl;
  wire[32:0] nl_mult_14_if_acc_nl;
  wire[32:0] mult_30_acc_1_nl;
  wire[33:0] nl_mult_30_acc_1_nl;
  wire[31:0] mult_13_if_acc_nl;
  wire[32:0] nl_mult_13_if_acc_nl;
  wire[32:0] mult_29_acc_1_nl;
  wire[33:0] nl_mult_29_acc_1_nl;
  wire[31:0] mult_12_if_acc_nl;
  wire[32:0] nl_mult_12_if_acc_nl;
  wire[32:0] mult_28_acc_1_nl;
  wire[33:0] nl_mult_28_acc_1_nl;
  wire[31:0] mult_11_if_acc_nl;
  wire[32:0] nl_mult_11_if_acc_nl;
  wire[32:0] mult_27_acc_1_nl;
  wire[33:0] nl_mult_27_acc_1_nl;
  wire[31:0] mult_10_if_acc_nl;
  wire[32:0] nl_mult_10_if_acc_nl;
  wire[32:0] mult_26_acc_1_nl;
  wire[33:0] nl_mult_26_acc_1_nl;
  wire[31:0] mult_9_if_acc_nl;
  wire[32:0] nl_mult_9_if_acc_nl;
  wire[32:0] mult_25_acc_1_nl;
  wire[33:0] nl_mult_25_acc_1_nl;
  wire[31:0] mult_8_if_acc_nl;
  wire[32:0] nl_mult_8_if_acc_nl;
  wire[32:0] mult_24_acc_1_nl;
  wire[33:0] nl_mult_24_acc_1_nl;
  wire[31:0] mult_7_if_acc_nl;
  wire[32:0] nl_mult_7_if_acc_nl;
  wire[32:0] mult_23_acc_1_nl;
  wire[33:0] nl_mult_23_acc_1_nl;
  wire[31:0] mult_6_if_acc_nl;
  wire[32:0] nl_mult_6_if_acc_nl;
  wire[32:0] mult_22_acc_1_nl;
  wire[33:0] nl_mult_22_acc_1_nl;
  wire[31:0] mult_5_if_acc_nl;
  wire[32:0] nl_mult_5_if_acc_nl;
  wire[32:0] mult_21_acc_1_nl;
  wire[33:0] nl_mult_21_acc_1_nl;
  wire[31:0] mult_4_if_acc_nl;
  wire[32:0] nl_mult_4_if_acc_nl;
  wire[32:0] mult_20_acc_1_nl;
  wire[33:0] nl_mult_20_acc_1_nl;
  wire[31:0] mult_3_if_acc_nl;
  wire[32:0] nl_mult_3_if_acc_nl;
  wire[32:0] mult_19_acc_1_nl;
  wire[33:0] nl_mult_19_acc_1_nl;
  wire[31:0] mult_2_if_acc_nl;
  wire[32:0] nl_mult_2_if_acc_nl;
  wire[32:0] mult_18_acc_1_nl;
  wire[33:0] nl_mult_18_acc_1_nl;
  wire[31:0] mult_1_if_acc_nl;
  wire[32:0] nl_mult_1_if_acc_nl;
  wire[32:0] mult_17_acc_1_nl;
  wire[33:0] nl_mult_17_acc_1_nl;
  wire[31:0] mult_if_acc_nl;
  wire[32:0] nl_mult_if_acc_nl;
  wire[32:0] mult_16_acc_1_nl;
  wire[33:0] nl_mult_16_acc_1_nl;
  wire[6:0] INNER_LOOP1_tw_and_nl;
  wire[5:0] INNER_LOOP2_tw_and_nl;
  wire[31:0] butterFly1_butterFly1_mux_2_nl;
  wire[31:0] butterFly1_butterFly1_mux_6_nl;
  wire[0:0] butterFly1_butterFly1_nor_2_nl;
  wire[0:0] butterFly1_butterFly1_nor_3_nl;
  wire[0:0] butterFly1_mux_15_nl;
  wire[31:0] butterFly1_1_butterFly1_1_mux_2_nl;
  wire[31:0] butterFly1_1_butterFly1_1_mux_6_nl;
  wire[31:0] butterFly1_2_butterFly1_2_mux_2_nl;
  wire[31:0] butterFly1_2_butterFly1_2_mux_6_nl;
  wire[31:0] butterFly1_3_butterFly1_3_mux_2_nl;
  wire[31:0] butterFly1_3_butterFly1_3_mux_6_nl;
  wire[31:0] butterFly1_4_butterFly1_4_mux_2_nl;
  wire[31:0] butterFly1_4_butterFly1_4_mux_6_nl;
  wire[5:0] butterFly1_5_butterFly1_5_mux_3_nl;
  wire[5:0] butterFly1_5_mux1h_11_nl;
  wire[31:0] butterFly1_5_butterFly1_5_mux_2_nl;
  wire[31:0] butterFly1_5_butterFly1_5_mux_6_nl;
  wire[5:0] butterFly1_6_butterFly1_6_mux_3_nl;
  wire[5:0] butterFly1_6_mux1h_11_nl;
  wire[31:0] butterFly1_6_butterFly1_6_mux_2_nl;
  wire[31:0] butterFly1_6_butterFly1_6_mux_6_nl;
  wire[5:0] butterFly1_7_mux1h_11_nl;
  wire[31:0] butterFly1_7_butterFly1_7_mux_2_nl;
  wire[31:0] butterFly1_7_butterFly1_7_mux_6_nl;
  wire[31:0] butterFly1_8_butterFly1_8_mux_2_nl;
  wire[31:0] butterFly1_8_butterFly1_8_mux_6_nl;
  wire[31:0] butterFly1_9_butterFly1_9_mux_2_nl;
  wire[31:0] butterFly1_9_butterFly1_9_mux_6_nl;
  wire[31:0] butterFly1_10_butterFly1_10_mux_2_nl;
  wire[31:0] butterFly1_10_butterFly1_10_mux_6_nl;
  wire[31:0] butterFly1_11_butterFly1_11_mux_2_nl;
  wire[31:0] butterFly1_11_butterFly1_11_mux_6_nl;
  wire[31:0] butterFly1_12_butterFly1_12_mux_2_nl;
  wire[31:0] butterFly1_12_butterFly1_12_mux_6_nl;
  wire[31:0] butterFly1_13_butterFly1_13_mux_2_nl;
  wire[31:0] butterFly1_13_butterFly1_13_mux_6_nl;
  wire[5:0] butterFly1_14_mux1h_11_nl;
  wire[31:0] butterFly1_14_butterFly1_14_mux_2_nl;
  wire[31:0] butterFly1_14_butterFly1_14_mux_6_nl;
  wire[31:0] butterFly1_15_butterFly1_15_mux_2_nl;
  wire[31:0] butterFly1_15_butterFly1_15_mux_6_nl;
  wire[31:0] butterFly1_butterFly1_mux_nl;
  wire[31:0] butterFly1_butterFly1_mux_5_nl;
  wire[0:0] butterFly1_butterFly1_nor_nl;
  wire[0:0] butterFly1_butterFly1_nor_1_nl;
  wire[0:0] butterFly1_mux_nl;
  wire[31:0] butterFly1_1_butterFly1_1_mux_nl;
  wire[31:0] butterFly1_1_butterFly1_1_mux_5_nl;
  wire[31:0] butterFly1_2_butterFly1_2_mux_nl;
  wire[31:0] butterFly1_2_butterFly1_2_mux_5_nl;
  wire[31:0] butterFly1_3_butterFly1_3_mux_nl;
  wire[31:0] butterFly1_3_butterFly1_3_mux_5_nl;
  wire[31:0] butterFly1_4_butterFly1_4_mux_nl;
  wire[31:0] butterFly1_4_butterFly1_4_mux_5_nl;
  wire[5:0] butterFly1_5_butterFly1_5_mux_4_nl;
  wire[5:0] butterFly1_5_mux1h_9_nl;
  wire[31:0] butterFly1_5_butterFly1_5_mux_nl;
  wire[31:0] butterFly1_5_butterFly1_5_mux_5_nl;
  wire[5:0] butterFly1_6_butterFly1_6_mux_4_nl;
  wire[5:0] butterFly1_6_mux1h_9_nl;
  wire[31:0] butterFly1_6_butterFly1_6_mux_nl;
  wire[31:0] butterFly1_6_butterFly1_6_mux_5_nl;
  wire[5:0] butterFly1_7_mux1h_9_nl;
  wire[31:0] butterFly1_7_butterFly1_7_mux_nl;
  wire[31:0] butterFly1_7_butterFly1_7_mux_5_nl;
  wire[31:0] butterFly1_8_butterFly1_8_mux_nl;
  wire[31:0] butterFly1_8_butterFly1_8_mux_5_nl;
  wire[31:0] butterFly1_9_butterFly1_9_mux_nl;
  wire[31:0] butterFly1_9_butterFly1_9_mux_5_nl;
  wire[31:0] butterFly1_10_butterFly1_10_mux_nl;
  wire[31:0] butterFly1_10_butterFly1_10_mux_5_nl;
  wire[31:0] butterFly1_11_butterFly1_11_mux_nl;
  wire[31:0] butterFly1_11_butterFly1_11_mux_5_nl;
  wire[31:0] butterFly1_12_butterFly1_12_mux_nl;
  wire[31:0] butterFly1_12_butterFly1_12_mux_5_nl;
  wire[31:0] butterFly1_13_butterFly1_13_mux_nl;
  wire[31:0] butterFly1_13_butterFly1_13_mux_5_nl;
  wire[5:0] butterFly1_14_mux1h_9_nl;
  wire[31:0] butterFly1_14_butterFly1_14_mux_nl;
  wire[31:0] butterFly1_14_butterFly1_14_mux_5_nl;
  wire[31:0] butterFly1_15_butterFly1_15_mux_nl;
  wire[31:0] butterFly1_15_butterFly1_15_mux_5_nl;
  wire[2:0] operator_20_false_mux_2_nl;
  wire[6:0] operator_20_false_mux1h_2_nl;
  wire[30:0] modulo_sub_6_qif_mux_2_nl;
  wire[30:0] modulo_sub_37_qif_mux_2_nl;
  wire[30:0] modulo_sub_36_qif_mux_2_nl;
  wire[30:0] modulo_sub_4_qif_mux_2_nl;
  wire[30:0] modulo_sub_35_qif_mux_2_nl;
  wire[30:0] modulo_sub_3_qif_mux_2_nl;
  wire[30:0] modulo_sub_34_qif_mux_2_nl;
  wire[30:0] modulo_sub_2_qif_mux_2_nl;
  wire[30:0] modulo_sub_33_qif_mux_2_nl;
  wire[30:0] modulo_sub_1_qif_mux_2_nl;
  wire[30:0] modulo_sub_32_qif_mux_2_nl;
  wire[30:0] modulo_sub_qif_mux_2_nl;
  wire[30:0] modulo_sub_31_qif_mux_2_nl;
  wire[30:0] modulo_sub_13_qif_mux_2_nl;
  wire[30:0] modulo_sub_30_qif_mux_2_nl;
  wire[30:0] modulo_sub_45_qif_mux_2_nl;
  wire[30:0] modulo_sub_29_qif_mux_2_nl;
  wire[30:0] modulo_sub_15_qif_mux_2_nl;
  wire[30:0] modulo_sub_28_qif_mux_2_nl;
  wire[30:0] modulo_sub_27_qif_mux_2_nl;
  wire[30:0] modulo_sub_26_qif_mux_2_nl;
  wire[30:0] modulo_sub_25_qif_mux_2_nl;
  wire[30:0] modulo_sub_24_qif_mux_2_nl;
  wire[30:0] modulo_sub_23_qif_mux_2_nl;
  wire[30:0] modulo_sub_22_qif_mux_2_nl;
  wire[30:0] modulo_sub_21_qif_mux_2_nl;
  wire[30:0] modulo_sub_20_qif_mux_2_nl;
  wire[30:0] modulo_sub_19_qif_mux_2_nl;
  wire[30:0] modulo_sub_18_qif_mux_2_nl;
  wire[30:0] modulo_sub_17_qif_mux_2_nl;
  wire[30:0] modulo_sub_16_qif_mux_2_nl;
  wire[32:0] acc_50_nl;
  wire[33:0] nl_acc_50_nl;
  wire[31:0] butterFly1_mux1h_17_nl;
  wire[32:0] acc_51_nl;
  wire[33:0] nl_acc_51_nl;
  wire[31:0] butterFly1_1_mux1h_13_nl;
  wire[32:0] acc_52_nl;
  wire[33:0] nl_acc_52_nl;
  wire[31:0] butterFly1_2_mux1h_13_nl;
  wire[32:0] acc_53_nl;
  wire[33:0] nl_acc_53_nl;
  wire[31:0] butterFly1_3_mux1h_13_nl;
  wire[32:0] acc_54_nl;
  wire[33:0] nl_acc_54_nl;
  wire[31:0] butterFly1_4_mux1h_13_nl;
  wire[32:0] acc_55_nl;
  wire[33:0] nl_acc_55_nl;
  wire[31:0] butterFly1_5_mux1h_13_nl;
  wire[32:0] acc_56_nl;
  wire[33:0] nl_acc_56_nl;
  wire[31:0] butterFly1_6_mux1h_13_nl;
  wire[32:0] acc_57_nl;
  wire[33:0] nl_acc_57_nl;
  wire[31:0] butterFly1_7_mux1h_13_nl;
  wire[32:0] acc_58_nl;
  wire[33:0] nl_acc_58_nl;
  wire[31:0] butterFly1_8_mux1h_13_nl;
  wire[32:0] acc_59_nl;
  wire[33:0] nl_acc_59_nl;
  wire[31:0] butterFly1_9_mux1h_13_nl;
  wire[32:0] acc_60_nl;
  wire[33:0] nl_acc_60_nl;
  wire[31:0] butterFly1_10_mux1h_13_nl;
  wire[32:0] acc_61_nl;
  wire[33:0] nl_acc_61_nl;
  wire[31:0] butterFly1_11_mux1h_13_nl;
  wire[32:0] acc_62_nl;
  wire[33:0] nl_acc_62_nl;
  wire[31:0] butterFly1_12_mux1h_13_nl;
  wire[32:0] acc_63_nl;
  wire[33:0] nl_acc_63_nl;
  wire[31:0] butterFly1_13_mux1h_13_nl;
  wire[32:0] acc_64_nl;
  wire[33:0] nl_acc_64_nl;
  wire[31:0] butterFly1_14_mux1h_13_nl;
  wire[32:0] acc_65_nl;
  wire[33:0] nl_acc_65_nl;
  wire[31:0] butterFly1_15_mux1h_13_nl;
  wire[31:0] butterFly1_15_mux1h_14_nl;
  wire[31:0] butterFly1_14_mux1h_14_nl;
  wire[31:0] butterFly1_13_mux1h_14_nl;
  wire[31:0] butterFly1_12_mux1h_14_nl;
  wire[31:0] butterFly1_11_mux1h_14_nl;
  wire[31:0] butterFly1_10_mux1h_14_nl;
  wire[31:0] butterFly1_9_mux1h_14_nl;
  wire[31:0] butterFly1_8_mux1h_14_nl;
  wire[31:0] butterFly1_7_mux1h_14_nl;
  wire[31:0] butterFly1_6_mux1h_14_nl;
  wire[31:0] butterFly1_5_mux1h_14_nl;
  wire[31:0] butterFly1_4_mux1h_14_nl;
  wire[31:0] butterFly1_3_mux1h_14_nl;
  wire[31:0] butterFly1_2_mux1h_14_nl;
  wire[31:0] butterFly1_1_mux1h_14_nl;
  wire[31:0] butterFly1_mux1h_18_nl;
  wire[33:0] acc_82_nl;
  wire[34:0] nl_acc_82_nl;
  wire[31:0] modulo_add_1_mux1h_3_nl;
  wire[33:0] acc_83_nl;
  wire[34:0] nl_acc_83_nl;
  wire[31:0] modulo_add_10_mux1h_3_nl;
  wire[33:0] acc_84_nl;
  wire[34:0] nl_acc_84_nl;
  wire[31:0] modulo_add_54_mux1h_3_nl;
  wire[33:0] acc_85_nl;
  wire[34:0] nl_acc_85_nl;
  wire[31:0] modulo_add_48_mux1h_3_nl;
  wire[33:0] acc_86_nl;
  wire[34:0] nl_acc_86_nl;
  wire[31:0] modulo_add_33_mux1h_3_nl;
  wire[33:0] acc_87_nl;
  wire[34:0] nl_acc_87_nl;
  wire[31:0] modulo_add_34_mux1h_3_nl;
  wire[33:0] acc_88_nl;
  wire[34:0] nl_acc_88_nl;
  wire[31:0] modulo_add_6_mux1h_3_nl;
  wire[33:0] acc_89_nl;
  wire[34:0] nl_acc_89_nl;
  wire[31:0] modulo_add_50_mux1h_3_nl;
  wire[33:0] acc_90_nl;
  wire[34:0] nl_acc_90_nl;
  wire[31:0] modulo_add_51_mux1h_3_nl;
  wire[33:0] acc_91_nl;
  wire[34:0] nl_acc_91_nl;
  wire[31:0] modulo_add_14_mux1h_3_nl;
  wire[33:0] acc_92_nl;
  wire[34:0] nl_acc_92_nl;
  wire[31:0] modulo_add_36_mux1h_3_nl;
  wire[33:0] acc_93_nl;
  wire[34:0] nl_acc_93_nl;
  wire[31:0] modulo_add_52_mux1h_3_nl;
  wire[33:0] acc_94_nl;
  wire[34:0] nl_acc_94_nl;
  wire[31:0] modulo_add_41_mux1h_3_nl;
  wire[33:0] acc_95_nl;
  wire[34:0] nl_acc_95_nl;
  wire[31:0] modulo_add_2_mux1h_3_nl;
  wire[33:0] acc_96_nl;
  wire[34:0] nl_acc_96_nl;
  wire[31:0] modulo_add_53_mux1h_3_nl;
  wire[33:0] acc_97_nl;
  wire[34:0] nl_acc_97_nl;
  wire[31:0] modulo_add_55_mux1h_3_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_mult_t_mul_cmp_a;
  assign nl_mult_t_mul_cmp_a = MUX1HOT_v_32_4_2((xt_rsc_0_1_i_qa_d[31:0]), (yt_rsc_0_1_i_qa_d[31:0]),
      (xt_rsc_0_31_i_qa_d[31:0]), (yt_rsc_0_31_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_b;
  assign nl_mult_t_mul_cmp_b = MUX1HOT_v_32_9_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]),
      (twiddle_h_rsc_0_11_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]), (twiddle_h_rsc_0_13_i_qa_d[31:0]),
      (twiddle_h_rsc_0_14_i_qa_d[31:0]), (twiddle_h_rsc_0_15_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_44_cse , mult_15_t_and_45_cse , mult_15_t_and_46_cse , mult_15_t_and_47_cse
      , mult_15_t_or_9_cse , mult_15_t_or_10_cse , mult_15_t_or_11_cse , mult_15_t_or_12_cse});
  wire [31:0] nl_mult_t_mul_cmp_1_a;
  assign nl_mult_t_mul_cmp_1_a = MUX1HOT_v_32_4_2((xt_rsc_0_31_i_qa_d[31:0]), (yt_rsc_0_31_i_qa_d[31:0]),
      (xt_rsc_0_29_i_qa_d[31:0]), (yt_rsc_0_1_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_1_b;
  assign nl_mult_t_mul_cmp_1_b = MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]),
      (twiddle_h_rsc_0_14_i_qa_d[31:0]), {or_tmp_771 , mult_15_t_and_40_cse , mult_15_t_and_41_cse
      , mult_15_t_and_42_cse , mult_15_t_and_43_cse});
  wire [31:0] nl_mult_t_mul_cmp_2_a;
  assign nl_mult_t_mul_cmp_2_a = MUX1HOT_v_32_4_2((xt_rsc_0_29_i_qa_d[31:0]), (yt_rsc_0_29_i_qa_d[31:0]),
      (xt_rsc_0_27_i_qa_d[31:0]), (yt_rsc_0_3_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_2_b;
  assign nl_mult_t_mul_cmp_2_b = MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]),
      (twiddle_h_rsc_0_13_i_qa_d[31:0]), (twiddle_h_rsc_0_1_i_qa_d[31:0]), {or_tmp_779
      , mult_15_t_and_36_cse , mult_15_t_and_37_cse , mult_15_t_and_38_cse , mult_15_t_and_39_cse
      , or_tmp_782});
  wire [31:0] nl_mult_t_mul_cmp_3_a;
  assign nl_mult_t_mul_cmp_3_a = MUX1HOT_v_32_4_2((xt_rsc_0_27_i_qa_d[31:0]), (yt_rsc_0_27_i_qa_d[31:0]),
      (xt_rsc_0_25_i_qa_d[31:0]), (yt_rsc_0_5_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_1029_nl;
  wire [31:0] nl_mult_t_mul_cmp_3_b;
  assign or_1029_nl = and_1719_cse | modulo_add_1_qelse_or_m1c;
  assign nl_mult_t_mul_cmp_3_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_12_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]),
      {or_1029_nl , or_tmp_790 , and_1725_cse , or_tmp_792});
  wire [31:0] nl_mult_t_mul_cmp_4_a;
  assign nl_mult_t_mul_cmp_4_a = MUX1HOT_v_32_4_2((xt_rsc_0_25_i_qa_d[31:0]), (yt_rsc_0_25_i_qa_d[31:0]),
      (xt_rsc_0_23_i_qa_d[31:0]), (yt_rsc_0_7_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_t_or_8_nl;
  wire [31:0] nl_mult_t_mul_cmp_4_b;
  assign mult_15_t_or_8_nl = modulo_add_1_qelse_or_m1c | mult_15_t_and_49_cse;
  assign nl_mult_t_mul_cmp_4_b = MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]),
      (twiddle_h_rsc_0_11_i_qa_d[31:0]), (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]),
      (twiddle_h_rsc_0_3_i_qa_d[31:0]), {mult_15_t_or_8_nl , mult_15_t_and_29_cse
      , mult_15_t_and_30_cse , mult_15_t_and_31_cse , mult_15_t_and_32_cse , mult_15_t_and_51_cse
      , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_t_mul_cmp_5_a;
  assign nl_mult_t_mul_cmp_5_a = MUX1HOT_v_32_4_2((xt_rsc_0_23_i_qa_d[31:0]), (yt_rsc_0_23_i_qa_d[31:0]),
      (xt_rsc_0_21_i_qa_d[31:0]), (yt_rsc_0_9_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_5_b;
  assign nl_mult_t_mul_cmp_5_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_10_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]),
      {modulo_add_1_qelse_or_m1c , or_tmp_809 , and_1763_cse , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_6_a;
  assign nl_mult_t_mul_cmp_6_a = MUX1HOT_v_32_4_2((xt_rsc_0_21_i_qa_d[31:0]), (yt_rsc_0_21_i_qa_d[31:0]),
      (xt_rsc_0_19_i_qa_d[31:0]), (yt_rsc_0_11_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_6_b;
  assign nl_mult_t_mul_cmp_6_b = MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_5_i_qa_d[31:0]),
      (twiddle_h_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c , or_tmp_819 ,
      and_1783_cse , or_tmp_782 , and_1700_cse});
  wire [31:0] nl_mult_t_mul_cmp_7_a;
  assign nl_mult_t_mul_cmp_7_a = MUX1HOT_v_32_4_2((xt_rsc_0_19_i_qa_d[31:0]), (yt_rsc_0_19_i_qa_d[31:0]),
      (xt_rsc_0_17_i_qa_d[31:0]), (yt_rsc_0_13_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_7_b;
  assign nl_mult_t_mul_cmp_7_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_6_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]),
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , or_tmp_792 , and_1719_cse});
  wire [31:0] nl_mult_t_mul_cmp_8_a;
  assign nl_mult_t_mul_cmp_8_a = MUX1HOT_v_32_4_2((xt_rsc_0_17_i_qa_d[31:0]), (yt_rsc_0_17_i_qa_d[31:0]),
      (xt_rsc_0_15_i_qa_d[31:0]), (yt_rsc_0_15_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_8_b;
  assign nl_mult_t_mul_cmp_8_b = MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_3_i_qa_d[31:0]),
      (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_5_i_qa_d[31:0]), (twiddle_h_rsc_0_6_i_qa_d[31:0]),
      (twiddle_h_rsc_0_7_i_qa_d[31:0]), {mult_15_t_or_3_cse , mult_15_t_and_45_cse
      , mult_15_t_and_46_cse , mult_15_t_and_47_cse , mult_15_t_or_9_cse , mult_15_t_or_10_cse
      , mult_15_t_or_11_cse , mult_15_t_or_12_cse});
  wire [31:0] nl_mult_t_mul_cmp_9_a;
  assign nl_mult_t_mul_cmp_9_a = MUX1HOT_v_32_4_2((xt_rsc_0_15_i_qa_d[31:0]), (yt_rsc_0_15_i_qa_d[31:0]),
      (xt_rsc_0_13_i_qa_d[31:0]), (yt_rsc_0_17_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_t_or_2_nl;
  wire [31:0] nl_mult_t_mul_cmp_9_b;
  assign mult_15_t_or_2_nl = modulo_add_1_qelse_or_m1c | mult_15_t_and_40_cse;
  assign nl_mult_t_mul_cmp_9_b = MUX1HOT_v_32_5_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_6_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), {mult_15_t_or_2_nl , mult_15_t_and_41_cse
      , mult_15_t_and_42_cse , mult_15_t_and_43_cse , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_10_a;
  assign nl_mult_t_mul_cmp_10_a = MUX1HOT_v_32_4_2((xt_rsc_0_13_i_qa_d[31:0]), (yt_rsc_0_13_i_qa_d[31:0]),
      (xt_rsc_0_11_i_qa_d[31:0]), (yt_rsc_0_19_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_10_b;
  assign nl_mult_t_mul_cmp_10_b = MUX1HOT_v_32_6_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_5_i_qa_d[31:0]),
      (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]), {mult_15_t_or_1_cse
      , mult_15_t_and_37_cse , mult_15_t_and_38_cse , mult_15_t_and_39_cse , or_tmp_782
      , and_1700_cse});
  wire [31:0] nl_mult_t_mul_cmp_11_a;
  assign nl_mult_t_mul_cmp_11_a = MUX1HOT_v_32_4_2((xt_rsc_0_11_i_qa_d[31:0]), (yt_rsc_0_11_i_qa_d[31:0]),
      (xt_rsc_0_9_i_qa_d[31:0]), (yt_rsc_0_21_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_1107_nl;
  wire [31:0] nl_mult_t_mul_cmp_11_b;
  assign or_1107_nl = and_1725_cse | modulo_add_1_qelse_or_m1c;
  assign nl_mult_t_mul_cmp_11_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_4_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]), (twiddle_h_rsc_0_8_i_qa_d[31:0]),
      {or_1107_nl , or_tmp_790 , or_tmp_792 , and_1719_cse});
  wire [31:0] nl_mult_t_mul_cmp_12_b;
  assign nl_mult_t_mul_cmp_12_b = MUX1HOT_v_32_8_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_3_i_qa_d[31:0]),
      (twiddle_h_rsc_0_8_i_qa_d[31:0]), (twiddle_h_rsc_0_9_i_qa_d[31:0]), (twiddle_h_rsc_0_10_i_qa_d[31:0]),
      (twiddle_h_rsc_0_11_i_qa_d[31:0]), {mult_15_t_or_cse , mult_15_t_and_30_cse
      , mult_15_t_and_31_cse , mult_15_t_and_32_cse , mult_15_t_and_49_cse , mult_15_t_and_51_cse
      , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_t_mul_cmp_13_a;
  assign nl_mult_t_mul_cmp_13_a = MUX1HOT_v_32_4_2((xt_rsc_0_7_i_qa_d[31:0]), (yt_rsc_0_7_i_qa_d[31:0]),
      (xt_rsc_0_5_i_qa_d[31:0]), (yt_rsc_0_25_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_13_b;
  assign nl_mult_t_mul_cmp_13_b = MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_2_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]), {or_tmp_885
      , or_tmp_809 , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_14_a;
  assign nl_mult_t_mul_cmp_14_a = MUX1HOT_v_32_4_2((xt_rsc_0_5_i_qa_d[31:0]), (yt_rsc_0_5_i_qa_d[31:0]),
      (xt_rsc_0_3_i_qa_d[31:0]), (yt_rsc_0_27_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_t_mul_cmp_14_b;
  assign nl_mult_t_mul_cmp_14_b = MUX1HOT_v_32_4_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_1_i_qa_d[31:0]), (twiddle_h_rsc_0_13_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]),
      {or_tmp_894 , or_tmp_819 , or_tmp_782 , and_1700_cse});
  wire [31:0] nl_mult_t_mul_cmp_15_a;
  assign nl_mult_t_mul_cmp_15_a = MUX1HOT_v_32_4_2((xt_rsc_0_3_i_qa_d[31:0]), (yt_rsc_0_3_i_qa_d[31:0]),
      (xt_rsc_0_1_i_qa_d[31:0]), (yt_rsc_0_29_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_1145_nl;
  wire [31:0] nl_mult_t_mul_cmp_15_b;
  assign or_1145_nl = modulo_add_1_qelse_or_m1c | (fsm_output[7]);
  assign nl_mult_t_mul_cmp_15_b = MUX1HOT_v_32_3_2((twiddle_h_rsc_0_0_i_qa_d[31:0]),
      (twiddle_h_rsc_0_14_i_qa_d[31:0]), (twiddle_h_rsc_0_12_i_qa_d[31:0]), {or_1145_nl
      , or_tmp_792 , and_1719_cse});
  wire [31:0] nl_mult_z_mul_cmp_a;
  assign nl_mult_z_mul_cmp_a = MUX1HOT_v_32_3_2((xt_rsc_0_1_i_qa_d[31:0]), (yt_rsc_0_1_i_qa_d[31:0]),
      (xt_rsc_0_31_i_qa_d[31:0]), {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
  wire [31:0] nl_mult_z_mul_cmp_b;
  assign nl_mult_z_mul_cmp_b = MUX1HOT_v_32_9_2((twiddle_rsc_0_0_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]),
      (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]), (twiddle_rsc_0_11_i_qa_d[31:0]),
      (twiddle_rsc_0_12_i_qa_d[31:0]), (twiddle_rsc_0_13_i_qa_d[31:0]), (twiddle_rsc_0_14_i_qa_d[31:0]),
      (twiddle_rsc_0_15_i_qa_d[31:0]), {or_tmp_771 , mult_15_t_and_44_cse , mult_15_t_and_45_cse
      , mult_15_t_and_46_cse , mult_15_t_and_47_cse , mult_15_t_and_48_cse , mult_15_t_and_50_cse
      , mult_15_t_and_52_cse , mult_15_t_and_54_cse});
  wire [31:0] nl_mult_z_mul_cmp_1_a;
  assign nl_mult_z_mul_cmp_1_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_1_z[63:32]), (mult_t_mul_cmp_11_z[63:32]),
      (mult_t_mul_cmp_12_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_1_b;
  assign nl_mult_z_mul_cmp_1_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_2_a;
  assign nl_mult_z_mul_cmp_2_a = MUX1HOT_v_32_4_2((xt_rsc_0_31_i_qa_d[31:0]), (yt_rsc_0_31_i_qa_d[31:0]),
      (xt_rsc_0_1_i_qa_d[31:0]), (yt_rsc_0_17_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_2_b;
  assign nl_mult_z_mul_cmp_2_b = MUX_v_32_2_2((twiddle_rsc_0_0_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]),
      fsm_output[9]);
  wire [31:0] nl_mult_z_mul_cmp_3_a;
  assign nl_mult_z_mul_cmp_3_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_2_z[63:32]), (mult_t_mul_cmp_5_z[63:32]),
      (mult_t_mul_cmp_6_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_3_b;
  assign nl_mult_z_mul_cmp_3_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_4_a;
  assign nl_mult_z_mul_cmp_4_a = MUX1HOT_v_32_3_2((xt_rsc_0_29_i_qa_d[31:0]), (yt_rsc_0_29_i_qa_d[31:0]),
      (yt_rsc_0_9_i_qa_d[31:0]), {or_dcpl_210 , (fsm_output[4]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_4_b;
  assign nl_mult_z_mul_cmp_4_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]),
      (twiddle_rsc_0_14_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_40_cse , mult_15_t_and_41_cse , mult_15_t_and_42_cse , mult_15_t_and_43_cse
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_5_a;
  assign nl_mult_z_mul_cmp_5_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_3_z[63:32]), (mult_t_mul_cmp_12_z[63:32]),
      (mult_t_mul_cmp_13_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_5_b;
  assign nl_mult_z_mul_cmp_5_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_6_a;
  assign nl_mult_z_mul_cmp_6_a = MUX1HOT_v_32_4_2((xt_rsc_0_27_i_qa_d[31:0]), (yt_rsc_0_27_i_qa_d[31:0]),
      (xt_rsc_0_15_i_qa_d[31:0]), (yt_rsc_0_31_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_6_b;
  assign nl_mult_z_mul_cmp_6_b = MUX1HOT_v_32_12_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_3_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]), (twiddle_rsc_0_6_i_qa_d[31:0]),
      (twiddle_rsc_0_7_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]), (twiddle_rsc_0_13_i_qa_d[31:0]),
      (twiddle_rsc_0_14_i_qa_d[31:0]), (twiddle_rsc_0_15_i_qa_d[31:0]), {mult_15_t_or_3_cse
      , mult_15_t_and_45_cse , mult_15_t_and_46_cse , mult_15_t_and_47_cse , mult_15_t_and_48_cse
      , mult_15_t_and_50_cse , mult_15_t_and_52_cse , mult_15_t_and_54_cse , mult_15_t_and_49_cse
      , mult_15_t_and_51_cse , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_7_a;
  assign nl_mult_z_mul_cmp_7_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_4_z[63:32]), (mult_t_mul_cmp_2_z[63:32]),
      (mult_t_mul_cmp_3_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_7_b;
  assign nl_mult_z_mul_cmp_7_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_8_a;
  assign nl_mult_z_mul_cmp_8_a = MUX1HOT_v_32_4_2((xt_rsc_0_25_i_qa_d[31:0]), (yt_rsc_0_25_i_qa_d[31:0]),
      (xt_rsc_0_3_i_qa_d[31:0]), (yt_rsc_0_19_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_8_b;
  assign nl_mult_z_mul_cmp_8_b = MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]),
      {or_tmp_894 , or_tmp_819 , or_tmp_782 , and_1700_cse});
  wire [31:0] nl_mult_z_mul_cmp_9_a;
  assign nl_mult_z_mul_cmp_9_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_5_z[63:32]), (mult_t_mul_cmp_10_z[63:32]),
      (mult_t_mul_cmp_11_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_9_b;
  assign nl_mult_z_mul_cmp_9_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_10_a;
  assign nl_mult_z_mul_cmp_10_a = MUX1HOT_v_32_4_2((xt_rsc_0_23_i_qa_d[31:0]), (yt_rsc_0_23_i_qa_d[31:0]),
      (xt_rsc_0_17_i_qa_d[31:0]), (yt_rsc_0_15_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_10_b;
  assign nl_mult_z_mul_cmp_10_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]),
      (twiddle_rsc_0_6_i_qa_d[31:0]), (twiddle_rsc_0_7_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , mult_15_t_and_49_cse , mult_15_t_and_51_cse , mult_15_t_and_53_cse
      , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_11_a;
  assign nl_mult_z_mul_cmp_11_a = MUX_v_32_2_2((mult_t_mul_cmp_6_z[63:32]), (mult_t_mul_cmp_7_z[63:32]),
      fsm_output[9]);
  wire [31:0] nl_mult_z_mul_cmp_11_b;
  assign nl_mult_z_mul_cmp_11_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_12_a;
  assign nl_mult_z_mul_cmp_12_a = MUX1HOT_v_32_4_2((xt_rsc_0_21_i_qa_d[31:0]), (yt_rsc_0_21_i_qa_d[31:0]),
      (xt_rsc_0_5_i_qa_d[31:0]), (yt_rsc_0_7_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_z_or_3_nl;
  wire[0:0] mult_15_z_or_6_nl;
  wire [31:0] nl_mult_z_mul_cmp_12_b;
  assign mult_15_z_or_3_nl = or_tmp_885 | mult_15_t_and_49_cse;
  assign mult_15_z_or_6_nl = or_tmp_809 | mult_15_t_and_53_cse;
  assign nl_mult_z_mul_cmp_12_b = MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_3_i_qa_d[31:0]),
      {mult_15_z_or_3_nl , mult_15_z_or_6_nl , mult_15_t_and_51_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_13_a;
  assign nl_mult_z_mul_cmp_13_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_7_z[63:32]), (mult_t_mul_cmp_1_z[63:32]),
      (mult_t_mul_cmp_2_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) ,
      (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_13_b;
  assign nl_mult_z_mul_cmp_13_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_14_a;
  assign nl_mult_z_mul_cmp_14_a = MUX1HOT_v_32_4_2((xt_rsc_0_19_i_qa_d[31:0]), (yt_rsc_0_19_i_qa_d[31:0]),
      (xt_rsc_0_27_i_qa_d[31:0]), (yt_rsc_0_29_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_z_or_5_nl;
  wire [31:0] nl_mult_z_mul_cmp_14_b;
  assign mult_15_z_or_5_nl = mult_15_t_and_38_cse | and_1719_cse;
  assign nl_mult_z_mul_cmp_14_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]),
      (twiddle_rsc_0_13_i_qa_d[31:0]), (twiddle_rsc_0_14_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_36_cse , mult_15_t_and_37_cse , mult_15_z_or_5_nl , mult_15_t_and_39_cse
      , or_tmp_792});
  wire [31:0] nl_mult_z_mul_cmp_15_a;
  assign nl_mult_z_mul_cmp_15_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_8_z[63:32]), (mult_t_mul_cmp_13_z[63:32]),
      (mult_t_mul_cmp_14_z[63:32]), {modulo_add_1_qelse_or_m1c , (fsm_output[7])
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_15_b;
  assign nl_mult_z_mul_cmp_15_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_16_a;
  assign nl_mult_z_mul_cmp_16_a = MUX1HOT_v_32_4_2((xt_rsc_0_17_i_qa_d[31:0]), (yt_rsc_0_17_i_qa_d[31:0]),
      (xt_rsc_0_13_i_qa_d[31:0]), (yt_rsc_0_3_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] mult_15_z_or_2_nl;
  wire [31:0] nl_mult_z_mul_cmp_16_b;
  assign mult_15_z_or_2_nl = or_tmp_779 | mult_15_t_and_40_cse;
  assign nl_mult_z_mul_cmp_16_b = MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_6_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), {mult_15_z_or_2_nl , mult_15_t_and_41_cse ,
      mult_15_t_and_42_cse , mult_15_t_and_43_cse , or_tmp_782});
  wire [31:0] nl_mult_z_mul_cmp_17_a;
  assign nl_mult_z_mul_cmp_17_a = MUX_v_32_2_2((mult_t_mul_cmp_9_z[63:32]), (mult_t_mul_cmp_10_z[63:32]),
      fsm_output[9]);
  wire [31:0] nl_mult_z_mul_cmp_17_b;
  assign nl_mult_z_mul_cmp_17_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_18_a;
  assign nl_mult_z_mul_cmp_18_a = MUX1HOT_v_32_4_2((xt_rsc_0_15_i_qa_d[31:0]), (yt_rsc_0_15_i_qa_d[31:0]),
      (xt_rsc_0_19_i_qa_d[31:0]), (yt_rsc_0_21_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire[0:0] or_1280_nl;
  wire [31:0] nl_mult_z_mul_cmp_18_b;
  assign or_1280_nl = and_1783_cse | and_1719_cse;
  assign nl_mult_z_mul_cmp_18_b = MUX1HOT_v_32_4_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]),
      {modulo_add_1_qelse_or_m1c , or_tmp_819 , or_1280_nl , or_tmp_792});
  wire [31:0] nl_mult_z_mul_cmp_19_a;
  assign nl_mult_z_mul_cmp_19_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_10_z[63:32]),
      (mult_t_mul_cmp_4_z[63:32]), (mult_t_mul_cmp_5_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_19_b;
  assign nl_mult_z_mul_cmp_19_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_20_a;
  assign nl_mult_z_mul_cmp_20_a = MUX1HOT_v_32_4_2((xt_rsc_0_13_i_qa_d[31:0]), (yt_rsc_0_13_i_qa_d[31:0]),
      (xt_rsc_0_25_i_qa_d[31:0]), (yt_rsc_0_11_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_20_b;
  assign nl_mult_z_mul_cmp_20_b = MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_12_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c , or_tmp_790 , and_1725_cse
      , or_tmp_782 , and_1700_cse});
  wire [31:0] nl_mult_z_mul_cmp_21_a;
  assign nl_mult_z_mul_cmp_21_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_11_z[63:32]),
      (mult_t_mul_cmp_14_z[63:32]), (mult_t_mul_cmp_15_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_21_b;
  assign nl_mult_z_mul_cmp_21_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_22_a;
  assign nl_mult_z_mul_cmp_22_a = MUX1HOT_v_32_3_2((xt_rsc_0_11_i_qa_d[31:0]), (yt_rsc_0_11_i_qa_d[31:0]),
      (yt_rsc_0_27_i_qa_d[31:0]), {or_dcpl_210 , (fsm_output[4]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_22_b;
  assign nl_mult_z_mul_cmp_22_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_5_i_qa_d[31:0]),
      (twiddle_rsc_0_13_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]), {mult_15_t_or_1_cse
      , mult_15_t_and_37_cse , mult_15_t_and_38_cse , mult_15_t_and_39_cse , or_tmp_782
      , and_1700_cse});
  wire [31:0] nl_mult_z_mul_cmp_23_a;
  assign nl_mult_z_mul_cmp_23_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_12_z[63:32]),
      (mult_t_mul_cmp_3_z[63:32]), (mult_t_mul_cmp_4_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_23_b;
  assign nl_mult_z_mul_cmp_23_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_24_b;
  assign nl_mult_z_mul_cmp_24_b = MUX1HOT_v_32_8_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_1_i_qa_d[31:0]), (twiddle_rsc_0_2_i_qa_d[31:0]), (twiddle_rsc_0_3_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]),
      (twiddle_rsc_0_11_i_qa_d[31:0]), {mult_15_t_or_cse , mult_15_t_and_30_cse ,
      mult_15_t_and_31_cse , mult_15_t_and_32_cse , mult_15_t_and_49_cse , mult_15_t_and_51_cse
      , mult_15_t_and_53_cse , mult_15_t_and_55_cse});
  wire [31:0] nl_mult_z_mul_cmp_25_a;
  assign nl_mult_z_mul_cmp_25_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_13_z[63:32]),
      (mult_t_mul_cmp_8_z[63:32]), (mult_t_mul_cmp_9_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_25_b;
  assign nl_mult_z_mul_cmp_25_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_26_a;
  assign nl_mult_z_mul_cmp_26_a = MUX1HOT_v_32_4_2((xt_rsc_0_7_i_qa_d[31:0]), (yt_rsc_0_7_i_qa_d[31:0]),
      (xt_rsc_0_21_i_qa_d[31:0]), (yt_rsc_0_13_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_26_b;
  assign nl_mult_z_mul_cmp_26_b = MUX1HOT_v_32_5_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_10_i_qa_d[31:0]), (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_6_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c , or_tmp_809 , and_1763_cse
      , or_tmp_792 , and_1719_cse});
  wire [31:0] nl_mult_z_mul_cmp_27_a;
  assign nl_mult_z_mul_cmp_27_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_14_z[63:32]),
      (mult_t_mul_cmp_7_z[63:32]), (mult_t_mul_cmp_8_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_27_b;
  assign nl_mult_z_mul_cmp_27_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_28_a;
  assign nl_mult_z_mul_cmp_28_a = MUX1HOT_v_32_3_2((xt_rsc_0_5_i_qa_d[31:0]), (yt_rsc_0_5_i_qa_d[31:0]),
      (xt_rsc_0_9_i_qa_d[31:0]), {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
  wire[0:0] or_1351_nl;
  wire [31:0] nl_mult_z_mul_cmp_28_b;
  assign or_1351_nl = and_1725_cse | and_1719_cse | modulo_add_1_qelse_or_m1c;
  assign nl_mult_z_mul_cmp_28_b = MUX1HOT_v_32_3_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_4_i_qa_d[31:0]), (twiddle_rsc_0_2_i_qa_d[31:0]), {or_1351_nl
      , or_tmp_790 , or_tmp_792});
  wire [31:0] nl_mult_z_mul_cmp_29_a;
  assign nl_mult_z_mul_cmp_29_a = MUX1HOT_v_32_3_2((mult_t_mul_cmp_15_z[63:32]),
      (mult_t_mul_cmp_z[63:32]), (mult_t_mul_cmp_1_z[63:32]), {modulo_add_1_qelse_or_m1c
      , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_29_b;
  assign nl_mult_z_mul_cmp_29_b = p_sva;
  wire [31:0] nl_mult_z_mul_cmp_30_a;
  assign nl_mult_z_mul_cmp_30_a = MUX1HOT_v_32_4_2((xt_rsc_0_3_i_qa_d[31:0]), (yt_rsc_0_3_i_qa_d[31:0]),
      (xt_rsc_0_23_i_qa_d[31:0]), (yt_rsc_0_25_i_qa_d[31:0]), {(fsm_output[2]) ,
      (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_30_b;
  assign nl_mult_z_mul_cmp_30_b = MUX1HOT_v_32_6_2((twiddle_rsc_0_0_i_qa_d[31:0]),
      (twiddle_rsc_0_8_i_qa_d[31:0]), (twiddle_rsc_0_9_i_qa_d[31:0]), (twiddle_rsc_0_10_i_qa_d[31:0]),
      (twiddle_rsc_0_11_i_qa_d[31:0]), (twiddle_rsc_0_12_i_qa_d[31:0]), {modulo_add_1_qelse_or_m1c
      , mult_15_t_and_29_cse , mult_15_t_and_30_cse , mult_15_t_and_31_cse , mult_15_t_and_32_cse
      , (fsm_output[9])});
  wire [31:0] nl_mult_z_mul_cmp_31_a;
  assign nl_mult_z_mul_cmp_31_a = MUX_v_32_2_2((mult_t_mul_cmp_z[63:32]), (mult_t_mul_cmp_15_z[63:32]),
      fsm_output[7]);
  wire [31:0] nl_mult_z_mul_cmp_31_b;
  assign nl_mult_z_mul_cmp_31_b = p_sva;
  wire [2:0] nl_operator_33_true_3_lshift_rg_s;
  assign nl_operator_33_true_3_lshift_rg_s = {1'b0 , (~ c_1_sva) , 1'b0};
  wire[2:0] operator_33_true_mux1h_nl;
  wire[0:0] operator_33_true_operator_33_true_or_nl;
  wire [3:0] nl_operator_33_true_1_lshift_rg_s;
  assign operator_33_true_mux1h_nl = MUX1HOT_v_3_3_2(z_out_1, operator_20_false_acc_cse_sva,
      ({2'b00 , (~ c_1_sva)}), {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[6])});
  assign operator_33_true_operator_33_true_or_nl = (~ (fsm_output[3])) | (fsm_output[1])
      | (fsm_output[6]);
  assign nl_operator_33_true_1_lshift_rg_s = {operator_33_true_mux1h_nl , operator_33_true_operator_33_true_or_nl};
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0;
  assign nl_peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0 = ~(INNER_LOOP1_stage_0
      | INNER_LOOP1_stage_0_2 | INNER_LOOP1_stage_0_3 | INNER_LOOP1_stage_0_4 | INNER_LOOP1_stage_0_5
      | INNER_LOOP1_stage_0_6 | INNER_LOOP1_stage_0_7 | INNER_LOOP1_stage_0_8 | INNER_LOOP1_stage_0_9
      | INNER_LOOP1_stage_0_10);
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0;
  assign nl_peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0 = z_out_1[2];
  wire [0:0] nl_peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1;
  assign nl_peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 = ~ INNER_LOOP4_nor_tmp;
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd32)) p_rsci (
      .dat(p_rsc_dat),
      .idat(p_rsci_idat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_31_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_31_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_30_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_30_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_29_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_29_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_28_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_28_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_27_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_27_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_26_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_26_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_25_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_25_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_24_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_24_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_23_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_23_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_22_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_22_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_21_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_21_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_20_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_20_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_19_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_19_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_18_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_18_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_17_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_17_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_16_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_16_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_15_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_14_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_13_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_12_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_11_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_10_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_9_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_8_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_7_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_6_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_5_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_4_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_3_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_2_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_1_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) xt_rsc_triosy_0_0_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(xt_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) p_rsc_triosy_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(p_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) r_rsc_triosy_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(r_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_15_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_14_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_13_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_12_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_11_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_10_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_9_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_8_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_7_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_6_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_5_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_4_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_3_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_2_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_1_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_rsc_triosy_0_0_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_rsc_triosy_0_0_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_15_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_15_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_14_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_14_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_13_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_13_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_12_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_12_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_11_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_11_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_10_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_10_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_9_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_9_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_8_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_8_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_7_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_7_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_6_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_6_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_5_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_5_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_4_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_4_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_3_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_3_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_2_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_2_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_1_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_1_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) twiddle_h_rsc_triosy_0_0_obj (
      .ld(reg_xt_rsc_triosy_0_31_obj_ld_cse),
      .lz(twiddle_h_rsc_triosy_0_0_lz)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp (
      .a(nl_mult_t_mul_cmp_a[31:0]),
      .b(nl_mult_t_mul_cmp_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_1 (
      .a(nl_mult_t_mul_cmp_1_a[31:0]),
      .b(nl_mult_t_mul_cmp_1_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_1_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_2 (
      .a(nl_mult_t_mul_cmp_2_a[31:0]),
      .b(nl_mult_t_mul_cmp_2_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_2_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_3 (
      .a(nl_mult_t_mul_cmp_3_a[31:0]),
      .b(nl_mult_t_mul_cmp_3_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_3_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_4 (
      .a(nl_mult_t_mul_cmp_4_a[31:0]),
      .b(nl_mult_t_mul_cmp_4_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_4_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_5 (
      .a(nl_mult_t_mul_cmp_5_a[31:0]),
      .b(nl_mult_t_mul_cmp_5_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_5_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_6 (
      .a(nl_mult_t_mul_cmp_6_a[31:0]),
      .b(nl_mult_t_mul_cmp_6_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_6_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_7 (
      .a(nl_mult_t_mul_cmp_7_a[31:0]),
      .b(nl_mult_t_mul_cmp_7_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_7_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_8 (
      .a(nl_mult_t_mul_cmp_8_a[31:0]),
      .b(nl_mult_t_mul_cmp_8_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_8_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_9 (
      .a(nl_mult_t_mul_cmp_9_a[31:0]),
      .b(nl_mult_t_mul_cmp_9_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_9_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_10 (
      .a(nl_mult_t_mul_cmp_10_a[31:0]),
      .b(nl_mult_t_mul_cmp_10_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_10_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_11 (
      .a(nl_mult_t_mul_cmp_11_a[31:0]),
      .b(nl_mult_t_mul_cmp_11_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_11_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_12 (
      .a(mult_4_t_mux1h_1_rmff),
      .b(nl_mult_t_mul_cmp_12_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_12_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_13 (
      .a(nl_mult_t_mul_cmp_13_a[31:0]),
      .b(nl_mult_t_mul_cmp_13_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_13_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_14 (
      .a(nl_mult_t_mul_cmp_14_a[31:0]),
      .b(nl_mult_t_mul_cmp_14_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_14_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd64),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_t_mul_cmp_15 (
      .a(nl_mult_t_mul_cmp_15_a[31:0]),
      .b(nl_mult_t_mul_cmp_15_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_t_mul_cmp_15_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp (
      .a(nl_mult_z_mul_cmp_a[31:0]),
      .b(nl_mult_z_mul_cmp_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_1 (
      .a(nl_mult_z_mul_cmp_1_a[31:0]),
      .b(nl_mult_z_mul_cmp_1_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_1_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_2 (
      .a(nl_mult_z_mul_cmp_2_a[31:0]),
      .b(nl_mult_z_mul_cmp_2_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_2_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_3 (
      .a(nl_mult_z_mul_cmp_3_a[31:0]),
      .b(nl_mult_z_mul_cmp_3_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_3_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_4 (
      .a(nl_mult_z_mul_cmp_4_a[31:0]),
      .b(nl_mult_z_mul_cmp_4_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_4_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_5 (
      .a(nl_mult_z_mul_cmp_5_a[31:0]),
      .b(nl_mult_z_mul_cmp_5_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_5_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_6 (
      .a(nl_mult_z_mul_cmp_6_a[31:0]),
      .b(nl_mult_z_mul_cmp_6_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_6_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_7 (
      .a(nl_mult_z_mul_cmp_7_a[31:0]),
      .b(nl_mult_z_mul_cmp_7_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_7_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_8 (
      .a(nl_mult_z_mul_cmp_8_a[31:0]),
      .b(nl_mult_z_mul_cmp_8_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_8_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_9 (
      .a(nl_mult_z_mul_cmp_9_a[31:0]),
      .b(nl_mult_z_mul_cmp_9_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_9_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_10 (
      .a(nl_mult_z_mul_cmp_10_a[31:0]),
      .b(nl_mult_z_mul_cmp_10_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_10_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_11 (
      .a(nl_mult_z_mul_cmp_11_a[31:0]),
      .b(nl_mult_z_mul_cmp_11_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_11_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_12 (
      .a(nl_mult_z_mul_cmp_12_a[31:0]),
      .b(nl_mult_z_mul_cmp_12_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_12_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_13 (
      .a(nl_mult_z_mul_cmp_13_a[31:0]),
      .b(nl_mult_z_mul_cmp_13_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_13_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_14 (
      .a(nl_mult_z_mul_cmp_14_a[31:0]),
      .b(nl_mult_z_mul_cmp_14_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_14_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_15 (
      .a(nl_mult_z_mul_cmp_15_a[31:0]),
      .b(nl_mult_z_mul_cmp_15_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_15_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_16 (
      .a(nl_mult_z_mul_cmp_16_a[31:0]),
      .b(nl_mult_z_mul_cmp_16_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_16_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_17 (
      .a(nl_mult_z_mul_cmp_17_a[31:0]),
      .b(nl_mult_z_mul_cmp_17_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_17_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_18 (
      .a(nl_mult_z_mul_cmp_18_a[31:0]),
      .b(nl_mult_z_mul_cmp_18_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_18_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_19 (
      .a(nl_mult_z_mul_cmp_19_a[31:0]),
      .b(nl_mult_z_mul_cmp_19_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_19_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_20 (
      .a(nl_mult_z_mul_cmp_20_a[31:0]),
      .b(nl_mult_z_mul_cmp_20_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_20_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_21 (
      .a(nl_mult_z_mul_cmp_21_a[31:0]),
      .b(nl_mult_z_mul_cmp_21_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_21_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_22 (
      .a(nl_mult_z_mul_cmp_22_a[31:0]),
      .b(nl_mult_z_mul_cmp_22_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_22_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_23 (
      .a(nl_mult_z_mul_cmp_23_a[31:0]),
      .b(nl_mult_z_mul_cmp_23_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_23_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_24 (
      .a(mult_4_t_mux1h_1_rmff),
      .b(nl_mult_z_mul_cmp_24_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_24_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_25 (
      .a(nl_mult_z_mul_cmp_25_a[31:0]),
      .b(nl_mult_z_mul_cmp_25_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_25_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_26 (
      .a(nl_mult_z_mul_cmp_26_a[31:0]),
      .b(nl_mult_z_mul_cmp_26_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_26_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_27 (
      .a(nl_mult_z_mul_cmp_27_a[31:0]),
      .b(nl_mult_z_mul_cmp_27_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_27_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_28 (
      .a(nl_mult_z_mul_cmp_28_a[31:0]),
      .b(nl_mult_z_mul_cmp_28_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_28_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_29 (
      .a(nl_mult_z_mul_cmp_29_a[31:0]),
      .b(nl_mult_z_mul_cmp_29_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_29_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_30 (
      .a(nl_mult_z_mul_cmp_30_a[31:0]),
      .b(nl_mult_z_mul_cmp_30_b[31:0]),
      .clk(clk),
      .en(mult_t_mul_cmp_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_30_z)
    );
  mgc_mul_pipe #(.width_a(32'sd32),
  .signd_a(32'sd0),
  .width_b(32'sd32),
  .signd_b(32'sd0),
  .width_z(32'sd32),
  .clock_edge(32'sd1),
  .enable_active(32'sd1),
  .a_rst_active(32'sd0),
  .s_rst_active(32'sd1),
  .stages(32'sd3),
  .n_inreg(32'sd1)) mult_z_mul_cmp_31 (
      .a(nl_mult_z_mul_cmp_31_a[31:0]),
      .b(nl_mult_z_mul_cmp_31_b[31:0]),
      .clk(clk),
      .en(mult_z_mul_cmp_1_en),
      .a_rst(1'b1),
      .s_rst(rst),
      .z(mult_z_mul_cmp_31_z)
    );
  mgc_shift_bl_v5 #(.width_a(32'sd1),
  .signd_a(32'sd1),
  .width_s(32'sd3),
  .width_z(32'sd2)) operator_33_true_3_lshift_rg (
      .a(1'b1),
      .s(nl_operator_33_true_3_lshift_rg_s[2:0]),
      .z(operator_33_true_3_lshift_psp_1_0_sva_mx0w3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd11)) operator_33_true_1_lshift_rg (
      .a(1'b1),
      .s(nl_operator_33_true_1_lshift_rg_s[3:0]),
      .z(z_out)
    );
  peaseNTT_core_wait_dp peaseNTT_core_wait_dp_inst (
      .yt_rsc_0_0_cgo_iro(or_261_rmff),
      .yt_rsc_0_0_i_clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .yt_rsc_0_16_cgo_iro(or_443_rmff),
      .yt_rsc_0_16_i_clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .ensig_cgo_iro(or_997_rmff),
      .ensig_cgo_iro_17(or_1156_rmff),
      .yt_rsc_0_0_cgo(reg_yt_rsc_0_0_cgo_cse),
      .yt_rsc_0_16_cgo(reg_yt_rsc_0_16_cgo_cse),
      .ensig_cgo(reg_ensig_cgo_cse),
      .mult_t_mul_cmp_en(mult_t_mul_cmp_en),
      .ensig_cgo_17(reg_ensig_cgo_17_cse),
      .mult_z_mul_cmp_1_en(mult_z_mul_cmp_1_en)
    );
  peaseNTT_core_core_fsm peaseNTT_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .INNER_LOOP1_C_0_tr0(nl_peaseNTT_core_core_fsm_inst_INNER_LOOP1_C_0_tr0[0:0]),
      .INNER_LOOP2_C_0_tr0(INNER_LOOP4_nor_tmp),
      .STAGE_LOOP_C_2_tr0(nl_peaseNTT_core_core_fsm_inst_STAGE_LOOP_C_2_tr0[0:0]),
      .INNER_LOOP3_C_0_tr0(INNER_LOOP4_nor_tmp),
      .INNER_LOOP4_C_0_tr0(and_dcpl_51),
      .INNER_LOOP4_C_0_tr1(nl_peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1[0:0])
    );
  assign or_261_rmff = ((and_dcpl_57 | and_dcpl_56 | ((~ INNER_LOOP1_stage_0_10)
      & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8)) & (fsm_output[7])) |
      and_167_cse | (((INNER_LOOP1_stage_0_11 & (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10))
      | and_dcpl_59 | and_dcpl_58) & (fsm_output[2]));
  assign and_202_rmff = INNER_LOOP1_stage_0 & or_dcpl_194;
  assign or_443_rmff = ((and_dcpl_68 | and_dcpl_67 | (INNER_LOOP1_stage_0_10 & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8))
      & (fsm_output[7])) | and_167_cse | (((INNER_LOOP1_stage_0_11 & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10)
      | and_dcpl_70 | and_dcpl_69) & (fsm_output[2]));
  assign and_921_rmff = INNER_LOOP1_stage_0 & or_dcpl_210;
  assign and_1435_rmff = INNER_LOOP1_stage_0 & or_dcpl_214;
  assign butterFly2_1_tw_butterFly2_1_tw_mux_rmff = MUX_v_7_2_2(INNER_LOOP3_r_11_4_sva_6_0,
      INNER_LOOP4_r_11_4_sva_6_0, fsm_output[9]);
  assign or_896_rmff = (and_dcpl_79 & (fsm_output[7])) | and_1445_cse;
  assign or_900_rmff = (and_dcpl_81 & (fsm_output[7])) | and_1454_cse;
  assign or_904_rmff = (and_dcpl_79 & (operator_20_false_acc_cse_sva[1]) & (fsm_output[7]))
      | and_1463_cse;
  assign or_908_rmff = (INNER_LOOP1_stage_0 & (operator_20_false_acc_cse_sva[2])
      & (fsm_output[7])) | (INNER_LOOP1_stage_0 & (fsm_output[9]));
  assign or_912_rmff = (and_dcpl_79 & (operator_20_false_acc_cse_sva[2]) & (fsm_output[7]))
      | and_1445_cse;
  assign or_916_rmff = (and_dcpl_81 & (operator_20_false_acc_cse_sva[2]) & (fsm_output[7]))
      | and_1454_cse;
  assign or_920_rmff = (and_dcpl_79 & (operator_20_false_acc_cse_sva[2:1]==2'b11)
      & (fsm_output[7])) | and_1463_cse;
  assign and_1506_rmff = INNER_LOOP1_stage_0 & or_dcpl_212;
  assign or_997_rmff = ((INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2
      | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1) & or_dcpl_218) | ((INNER_LOOP1_stage_0_4
      | INNER_LOOP1_stage_0_2 | INNER_LOOP1_stage_0_3) & (fsm_output[2]));
  assign mult_15_t_and_49_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b00) &
      (fsm_output[9]);
  assign mult_15_t_and_51_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b01) &
      (fsm_output[9]);
  assign mult_15_t_and_53_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b10) &
      (fsm_output[9]);
  assign mult_15_t_and_55_cse = (operator_33_true_3_lshift_psp_1_0_sva==2'b11) &
      (fsm_output[9]);
  assign mult_15_t_and_44_cse = butterFly2_15_tw_equal_tmp_1 & (fsm_output[7]);
  assign butterFly2_7_tw_nor_cse = ~((operator_20_false_acc_cse_sva[2:1]!=2'b00));
  assign mult_15_t_and_45_cse = (operator_20_false_acc_cse_sva[0]) & butterFly2_7_tw_nor_cse
      & (fsm_output[7]);
  assign butterFly2_7_tw_nor_1_cse = ~((operator_20_false_acc_cse_sva[2]) | (operator_20_false_acc_cse_sva[0]));
  assign mult_15_t_and_46_cse = (operator_20_false_acc_cse_sva[1]) & butterFly2_7_tw_nor_1_cse
      & (fsm_output[7]);
  assign mult_15_t_and_47_cse = butterFly2_15_tw_equal_tmp_3_1 & (fsm_output[7]);
  assign butterFly2_7_tw_nor_2_cse = ~((operator_20_false_acc_cse_sva[1:0]!=2'b00));
  assign mult_15_t_and_48_cse = (operator_20_false_acc_cse_sva[2]) & butterFly2_7_tw_nor_2_cse
      & (fsm_output[7]);
  assign mult_15_t_and_50_cse = butterFly2_15_tw_equal_tmp_5_1 & (fsm_output[7]);
  assign mult_15_t_and_52_cse = butterFly2_15_tw_equal_tmp_6_1 & (fsm_output[7]);
  assign mult_15_t_and_54_cse = butterFly2_15_tw_equal_tmp_7_1 & (fsm_output[7]);
  assign mult_15_t_or_9_cse = mult_15_t_and_48_cse | mult_15_t_and_49_cse;
  assign mult_15_t_or_10_cse = mult_15_t_and_50_cse | mult_15_t_and_51_cse;
  assign mult_15_t_or_11_cse = mult_15_t_and_52_cse | mult_15_t_and_53_cse;
  assign mult_15_t_or_12_cse = mult_15_t_and_54_cse | mult_15_t_and_55_cse;
  assign mult_15_t_and_41_cse = (operator_20_false_acc_cse_sva[2:1]==2'b01) & (fsm_output[7]);
  assign mult_15_t_and_42_cse = (operator_20_false_acc_cse_sva[2:1]==2'b10) & (fsm_output[7]);
  assign mult_15_t_and_43_cse = (operator_20_false_acc_cse_sva[2:1]==2'b11) & (fsm_output[7]);
  assign mult_15_t_and_40_cse = butterFly2_7_tw_nor_cse & (fsm_output[7]);
  assign mult_15_t_and_37_cse = (operator_20_false_acc_cse_sva[0]) & (~ (operator_20_false_acc_cse_sva[2]))
      & (fsm_output[7]);
  assign mult_15_t_and_38_cse = (operator_20_false_acc_cse_sva[2]) & (~ (operator_20_false_acc_cse_sva[0]))
      & (fsm_output[7]);
  assign mult_15_t_and_39_cse = (operator_20_false_acc_cse_sva[2]) & (operator_20_false_acc_cse_sva[0])
      & (fsm_output[7]);
  assign mult_15_t_and_36_cse = butterFly2_7_tw_nor_1_cse & (fsm_output[7]);
  assign mult_15_t_and_30_cse = (operator_20_false_acc_cse_sva[1:0]==2'b01) & (fsm_output[7]);
  assign mult_15_t_and_31_cse = (operator_20_false_acc_cse_sva[1:0]==2'b10) & (fsm_output[7]);
  assign mult_15_t_and_32_cse = (operator_20_false_acc_cse_sva[1:0]==2'b11) & (fsm_output[7]);
  assign mult_15_t_and_29_cse = butterFly2_7_tw_nor_2_cse & (fsm_output[7]);
  assign mult_15_t_or_3_cse = modulo_add_1_qelse_or_m1c | mult_15_t_and_44_cse;
  assign mult_15_t_or_1_cse = modulo_add_1_qelse_or_m1c | mult_15_t_and_36_cse;
  assign mult_4_t_mux1h_1_rmff = MUX1HOT_v_32_4_2((xt_rsc_0_9_i_qa_d[31:0]), (yt_rsc_0_9_i_qa_d[31:0]),
      (xt_rsc_0_7_i_qa_d[31:0]), (yt_rsc_0_23_i_qa_d[31:0]), {(fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7]) , (fsm_output[9])});
  assign mult_15_t_or_cse = modulo_add_1_qelse_or_m1c | mult_15_t_and_29_cse;
  assign or_1156_rmff = ((INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4
      | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3) & or_dcpl_218) | ((INNER_LOOP1_stage_0_6
      | INNER_LOOP1_stage_0_7 | INNER_LOOP1_stage_0_5) & (fsm_output[2]));
  assign modulo_add_1_qelse_or_m1c = (fsm_output[2]) | (fsm_output[4]);
  assign or_12_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 | INNER_LOOP1_stage_0_9;
  assign or_44_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 | INNER_LOOP1_stage_0_8;
  assign or_64_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 | INNER_LOOP1_stage_0_7;
  assign or_84_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 | INNER_LOOP1_stage_0_6;
  assign or_103_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 | INNER_LOOP1_stage_0_5;
  assign or_123_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 | INNER_LOOP1_stage_0_4;
  assign or_142_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm | INNER_LOOP1_stage_0_3;
  assign or_143_cse = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm | INNER_LOOP1_stage_0_2;
  assign modulo_sub_16_qelse_and_ssc = ~((z_out_66[31]) | (fsm_output[9]));
  assign modulo_sub_16_qelse_and_ssc_1 = (~ (z_out_51[31])) & (fsm_output[9]);
  assign modulo_sub_17_qelse_and_ssc = ~((z_out_56[31]) | (fsm_output[9]));
  assign modulo_sub_17_qelse_and_ssc_1 = (~ (z_out_52[31])) & (fsm_output[9]);
  assign modulo_sub_18_qelse_and_ssc = ~((z_out_63[31]) | (fsm_output[9]));
  assign modulo_sub_18_qelse_and_ssc_1 = (~ (z_out_53[31])) & (fsm_output[9]);
  assign modulo_sub_19_qelse_and_ssc = ~((z_out_64[31]) | (fsm_output[9]));
  assign modulo_sub_19_qelse_and_ssc_1 = (~ (z_out_54[31])) & (fsm_output[9]);
  assign modulo_sub_20_qelse_and_ssc = ~((z_out_65[31]) | (fsm_output[9]));
  assign modulo_sub_20_qelse_and_ssc_1 = (~ (z_out_55[31])) & (fsm_output[9]);
  assign modulo_sub_21_qelse_and_ssc = ~((z_out_51[31]) | (fsm_output[9]));
  assign modulo_sub_21_qelse_and_ssc_1 = (~ (z_out_56[31])) & (fsm_output[9]);
  assign modulo_sub_22_qelse_and_ssc = ~((z_out_52[31]) | (fsm_output[9]));
  assign modulo_sub_22_qelse_and_ssc_1 = (~ (z_out_57[31])) & (fsm_output[9]);
  assign modulo_sub_23_qelse_and_ssc = ~((z_out_53[31]) | (fsm_output[9]));
  assign modulo_sub_23_qelse_and_ssc_1 = (~ (z_out_58[31])) & (fsm_output[9]);
  assign modulo_sub_24_qelse_and_ssc = ~((z_out_54[31]) | (fsm_output[9]));
  assign modulo_sub_24_qelse_and_ssc_1 = (~ (z_out_59[31])) & (fsm_output[9]);
  assign modulo_sub_25_qelse_and_ssc = ~((z_out_55[31]) | (fsm_output[9]));
  assign modulo_sub_25_qelse_and_ssc_1 = (~ (z_out_60[31])) & (fsm_output[9]);
  assign modulo_sub_26_qelse_and_ssc = ~((z_out_57[31]) | (fsm_output[9]));
  assign modulo_sub_26_qelse_and_ssc_1 = (~ (z_out_61[31])) & (fsm_output[9]);
  assign modulo_sub_27_qelse_and_ssc = ~((z_out_58[31]) | (fsm_output[9]));
  assign modulo_sub_27_qelse_and_ssc_1 = (~ (z_out_62[31])) & (fsm_output[9]);
  assign modulo_sub_28_qelse_and_ssc = ~((z_out_59[31]) | (fsm_output[9]));
  assign modulo_sub_28_qelse_and_ssc_1 = (~ (z_out_63[31])) & (fsm_output[9]);
  assign modulo_sub_29_qelse_and_ssc = ~((z_out_60[31]) | (fsm_output[9]));
  assign modulo_sub_29_qelse_and_ssc_1 = (~ (z_out_64[31])) & (fsm_output[9]);
  assign modulo_sub_30_qelse_and_ssc = ~((z_out_61[31]) | (fsm_output[9]));
  assign modulo_sub_30_qelse_and_ssc_1 = (~ (z_out_65[31])) & (fsm_output[9]);
  assign modulo_sub_31_qelse_and_ssc = ~((z_out_62[31]) | (fsm_output[9]));
  assign modulo_sub_31_qelse_and_ssc_1 = (~ (z_out_66[31])) & (fsm_output[9]);
  assign yt_rsc_0_0_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_51[30:0])}),
      z_out_20, z_out_51[31]);
  assign yt_rsc_0_0_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_65[30:0])}),
      z_out_18, z_out_65[31]);
  assign yt_rsc_0_1_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_52[30:0])}),
      z_out_17, z_out_52[31]);
  assign yt_rsc_0_1_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_66[30:0])}),
      z_out_16, z_out_66[31]);
  assign yt_rsc_0_2_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_53[30:0])}),
      z_out_14, z_out_53[31]);
  assign yt_rsc_0_2_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_51[30:0])}),
      z_out_13, z_out_51[31]);
  assign yt_rsc_0_3_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_54[30:0])}),
      z_out_12, z_out_54[31]);
  assign yt_rsc_0_3_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_52[30:0])}),
      z_out_10, z_out_52[31]);
  assign yt_rsc_0_4_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_55[30:0])}),
      z_out_9, z_out_55[31]);
  assign yt_rsc_0_4_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_53[30:0])}),
      z_out_8, z_out_53[31]);
  assign nl_modulo_sub_5_qif_acc_nl = ({1'b1 , (z_out_56[30:0])}) + p_sva;
  assign modulo_sub_5_qif_acc_nl = nl_modulo_sub_5_qif_acc_nl[31:0];
  assign modulo_sub_5_qelse_mux_cse = MUX_v_32_2_2(({1'b0 , (z_out_56[30:0])}), modulo_sub_5_qif_acc_nl,
      z_out_56[31]);
  assign yt_rsc_0_5_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_54[30:0])}),
      z_out_5, z_out_54[31]);
  assign yt_rsc_0_6_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_57[30:0])}),
      z_out_4, z_out_57[31]);
  assign yt_rsc_0_6_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_55[30:0])}),
      z_out_4, z_out_55[31]);
  assign yt_rsc_0_7_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_58[30:0])}),
      z_out_5, z_out_58[31]);
  assign yt_rsc_0_8_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_59[30:0])}),
      z_out_8, z_out_59[31]);
  assign yt_rsc_0_8_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_57[30:0])}),
      z_out_9, z_out_57[31]);
  assign yt_rsc_0_9_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_60[30:0])}),
      z_out_10, z_out_60[31]);
  assign yt_rsc_0_9_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_58[30:0])}),
      z_out_12, z_out_58[31]);
  assign yt_rsc_0_10_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_61[30:0])}),
      z_out_13, z_out_61[31]);
  assign yt_rsc_0_10_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_59[30:0])}),
      z_out_14, z_out_59[31]);
  assign yt_rsc_0_11_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_62[30:0])}),
      z_out_16, z_out_62[31]);
  assign yt_rsc_0_11_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_60[30:0])}),
      z_out_17, z_out_60[31]);
  assign yt_rsc_0_12_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_63[30:0])}),
      z_out_18, z_out_63[31]);
  assign yt_rsc_0_12_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_61[30:0])}),
      z_out_20, z_out_61[31]);
  assign yt_rsc_0_13_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_64[30:0])}),
      z_out_22, z_out_64[31]);
  assign yt_rsc_0_13_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_62[30:0])}),
      z_out_25, z_out_62[31]);
  assign yt_rsc_0_14_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_65[30:0])}),
      z_out_25, z_out_65[31]);
  assign yt_rsc_0_14_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_63[30:0])}),
      z_out_22, z_out_63[31]);
  assign yt_rsc_0_15_i_da_d_mx0w0_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_66[30:0])}),
      z_out_28, z_out_66[31]);
  assign yt_rsc_0_15_i_da_d_mx0w2_63_32 = MUX_v_32_2_2(({1'b0 , (z_out_64[30:0])}),
      z_out_28, z_out_64[31]);
  assign nl_mult_15_if_acc_nl = mult_15_res_sva_1 - p_sva;
  assign mult_15_if_acc_nl = nl_mult_15_if_acc_nl[31:0];
  assign nl_mult_31_acc_1_nl = ({1'b1 , mult_15_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_31_acc_1_nl = nl_mult_31_acc_1_nl[32:0];
  assign mult_15_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_15_if_acc_nl, mult_15_res_sva_1,
      readslicef_33_1_32(mult_31_acc_1_nl));
  assign nl_mult_14_if_acc_nl = mult_14_res_sva_1 - p_sva;
  assign mult_14_if_acc_nl = nl_mult_14_if_acc_nl[31:0];
  assign nl_mult_30_acc_1_nl = ({1'b1 , mult_14_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_30_acc_1_nl = nl_mult_30_acc_1_nl[32:0];
  assign mult_14_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_14_if_acc_nl, mult_14_res_sva_1,
      readslicef_33_1_32(mult_30_acc_1_nl));
  assign nl_mult_13_if_acc_nl = mult_13_res_sva_1 - p_sva;
  assign mult_13_if_acc_nl = nl_mult_13_if_acc_nl[31:0];
  assign nl_mult_29_acc_1_nl = ({1'b1 , mult_13_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_29_acc_1_nl = nl_mult_29_acc_1_nl[32:0];
  assign mult_13_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_13_if_acc_nl, mult_13_res_sva_1,
      readslicef_33_1_32(mult_29_acc_1_nl));
  assign nl_mult_12_if_acc_nl = mult_12_res_sva_1 - p_sva;
  assign mult_12_if_acc_nl = nl_mult_12_if_acc_nl[31:0];
  assign nl_mult_28_acc_1_nl = ({1'b1 , mult_12_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_28_acc_1_nl = nl_mult_28_acc_1_nl[32:0];
  assign mult_12_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_12_if_acc_nl, mult_12_res_sva_1,
      readslicef_33_1_32(mult_28_acc_1_nl));
  assign nl_mult_11_if_acc_nl = mult_11_res_sva_1 - p_sva;
  assign mult_11_if_acc_nl = nl_mult_11_if_acc_nl[31:0];
  assign nl_mult_27_acc_1_nl = ({1'b1 , mult_11_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_27_acc_1_nl = nl_mult_27_acc_1_nl[32:0];
  assign mult_11_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_11_if_acc_nl, mult_11_res_sva_1,
      readslicef_33_1_32(mult_27_acc_1_nl));
  assign nl_mult_10_if_acc_nl = mult_10_res_sva_1 - p_sva;
  assign mult_10_if_acc_nl = nl_mult_10_if_acc_nl[31:0];
  assign nl_mult_26_acc_1_nl = ({1'b1 , mult_10_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_26_acc_1_nl = nl_mult_26_acc_1_nl[32:0];
  assign mult_10_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_10_if_acc_nl, mult_10_res_sva_1,
      readslicef_33_1_32(mult_26_acc_1_nl));
  assign nl_mult_9_if_acc_nl = mult_9_res_sva_1 - p_sva;
  assign mult_9_if_acc_nl = nl_mult_9_if_acc_nl[31:0];
  assign nl_mult_25_acc_1_nl = ({1'b1 , mult_9_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_25_acc_1_nl = nl_mult_25_acc_1_nl[32:0];
  assign mult_9_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_9_if_acc_nl, mult_9_res_sva_1,
      readslicef_33_1_32(mult_25_acc_1_nl));
  assign nl_mult_8_if_acc_nl = mult_8_res_sva_1 - p_sva;
  assign mult_8_if_acc_nl = nl_mult_8_if_acc_nl[31:0];
  assign nl_mult_24_acc_1_nl = ({1'b1 , mult_8_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_24_acc_1_nl = nl_mult_24_acc_1_nl[32:0];
  assign mult_8_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_8_if_acc_nl, mult_8_res_sva_1,
      readslicef_33_1_32(mult_24_acc_1_nl));
  assign nl_mult_7_if_acc_nl = mult_7_res_sva_1 - p_sva;
  assign mult_7_if_acc_nl = nl_mult_7_if_acc_nl[31:0];
  assign nl_mult_23_acc_1_nl = ({1'b1 , mult_7_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_23_acc_1_nl = nl_mult_23_acc_1_nl[32:0];
  assign mult_7_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_7_if_acc_nl, mult_7_res_sva_1,
      readslicef_33_1_32(mult_23_acc_1_nl));
  assign nl_mult_6_if_acc_nl = mult_6_res_sva_1 - p_sva;
  assign mult_6_if_acc_nl = nl_mult_6_if_acc_nl[31:0];
  assign nl_mult_22_acc_1_nl = ({1'b1 , mult_6_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_22_acc_1_nl = nl_mult_22_acc_1_nl[32:0];
  assign mult_6_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_6_if_acc_nl, mult_6_res_sva_1,
      readslicef_33_1_32(mult_22_acc_1_nl));
  assign nl_mult_5_if_acc_nl = mult_5_res_sva_1 - p_sva;
  assign mult_5_if_acc_nl = nl_mult_5_if_acc_nl[31:0];
  assign nl_mult_21_acc_1_nl = ({1'b1 , mult_5_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_21_acc_1_nl = nl_mult_21_acc_1_nl[32:0];
  assign mult_5_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_5_if_acc_nl, mult_5_res_sva_1,
      readslicef_33_1_32(mult_21_acc_1_nl));
  assign nl_mult_4_if_acc_nl = mult_4_res_sva_1 - p_sva;
  assign mult_4_if_acc_nl = nl_mult_4_if_acc_nl[31:0];
  assign nl_mult_20_acc_1_nl = ({1'b1 , mult_4_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_20_acc_1_nl = nl_mult_20_acc_1_nl[32:0];
  assign mult_4_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_4_if_acc_nl, mult_4_res_sva_1,
      readslicef_33_1_32(mult_20_acc_1_nl));
  assign nl_mult_3_if_acc_nl = mult_3_res_sva_1 - p_sva;
  assign mult_3_if_acc_nl = nl_mult_3_if_acc_nl[31:0];
  assign nl_mult_19_acc_1_nl = ({1'b1 , mult_3_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_19_acc_1_nl = nl_mult_19_acc_1_nl[32:0];
  assign mult_3_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_3_if_acc_nl, mult_3_res_sva_1,
      readslicef_33_1_32(mult_19_acc_1_nl));
  assign nl_mult_2_if_acc_nl = mult_2_res_sva_1 - p_sva;
  assign mult_2_if_acc_nl = nl_mult_2_if_acc_nl[31:0];
  assign nl_mult_18_acc_1_nl = ({1'b1 , mult_2_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_18_acc_1_nl = nl_mult_18_acc_1_nl[32:0];
  assign mult_2_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_2_if_acc_nl, mult_2_res_sva_1,
      readslicef_33_1_32(mult_18_acc_1_nl));
  assign nl_mult_1_if_acc_nl = mult_1_res_sva_1 - p_sva;
  assign mult_1_if_acc_nl = nl_mult_1_if_acc_nl[31:0];
  assign nl_mult_17_acc_1_nl = ({1'b1 , mult_1_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_17_acc_1_nl = nl_mult_17_acc_1_nl[32:0];
  assign mult_1_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_1_if_acc_nl, mult_1_res_sva_1,
      readslicef_33_1_32(mult_17_acc_1_nl));
  assign nl_mult_if_acc_nl = mult_res_sva_1 - p_sva;
  assign mult_if_acc_nl = nl_mult_if_acc_nl[31:0];
  assign nl_mult_16_acc_1_nl = ({1'b1 , mult_res_sva_1}) + conv_u2u_32_33(~ p_sva)
      + 33'b000000000000000000000000000000001;
  assign mult_16_acc_1_nl = nl_mult_16_acc_1_nl[32:0];
  assign mult_res_lpi_3_dfm_1_mx0 = MUX_v_32_2_2(mult_if_acc_nl, mult_res_sva_1,
      readslicef_33_1_32(mult_16_acc_1_nl));
  assign nl_mult_15_res_sva_1 = mult_15_z_asn_itm_3 - mult_z_mul_cmp_1_z;
  assign mult_15_res_sva_1 = nl_mult_15_res_sva_1[31:0];
  assign nl_mult_14_res_sva_1 = mult_14_z_asn_itm_3 - mult_z_mul_cmp_3_z;
  assign mult_14_res_sva_1 = nl_mult_14_res_sva_1[31:0];
  assign nl_mult_13_res_sva_1 = mult_13_z_asn_itm_3 - mult_z_mul_cmp_5_z;
  assign mult_13_res_sva_1 = nl_mult_13_res_sva_1[31:0];
  assign nl_mult_12_res_sva_1 = mult_12_z_asn_itm_3 - mult_z_mul_cmp_7_z;
  assign mult_12_res_sva_1 = nl_mult_12_res_sva_1[31:0];
  assign nl_mult_11_res_sva_1 = mult_11_z_asn_itm_3 - mult_z_mul_cmp_9_z;
  assign mult_11_res_sva_1 = nl_mult_11_res_sva_1[31:0];
  assign nl_mult_10_res_sva_1 = mult_10_z_asn_itm_3 - mult_z_mul_cmp_11_z;
  assign mult_10_res_sva_1 = nl_mult_10_res_sva_1[31:0];
  assign nl_mult_9_res_sva_1 = mult_25_z_asn_itm_3 - mult_z_mul_cmp_13_z;
  assign mult_9_res_sva_1 = nl_mult_9_res_sva_1[31:0];
  assign nl_mult_8_res_sva_1 = mult_24_z_asn_itm_3 - mult_z_mul_cmp_15_z;
  assign mult_8_res_sva_1 = nl_mult_8_res_sva_1[31:0];
  assign nl_mult_7_res_sva_1 = mult_23_z_asn_itm_3 - mult_z_mul_cmp_17_z;
  assign mult_7_res_sva_1 = nl_mult_7_res_sva_1[31:0];
  assign nl_mult_6_res_sva_1 = mult_22_z_asn_itm_3 - mult_z_mul_cmp_19_z;
  assign mult_6_res_sva_1 = nl_mult_6_res_sva_1[31:0];
  assign nl_mult_5_res_sva_1 = mult_21_z_asn_itm_3 - mult_z_mul_cmp_21_z;
  assign mult_5_res_sva_1 = nl_mult_5_res_sva_1[31:0];
  assign nl_mult_4_res_sva_1 = mult_20_z_asn_itm_3 - mult_z_mul_cmp_23_z;
  assign mult_4_res_sva_1 = nl_mult_4_res_sva_1[31:0];
  assign nl_mult_3_res_sva_1 = mult_19_z_asn_itm_3 - mult_z_mul_cmp_25_z;
  assign mult_3_res_sva_1 = nl_mult_3_res_sva_1[31:0];
  assign nl_mult_2_res_sva_1 = mult_18_z_asn_itm_3 - mult_z_mul_cmp_27_z;
  assign mult_2_res_sva_1 = nl_mult_2_res_sva_1[31:0];
  assign nl_mult_1_res_sva_1 = mult_17_z_asn_itm_3 - mult_z_mul_cmp_29_z;
  assign mult_1_res_sva_1 = nl_mult_1_res_sva_1[31:0];
  assign nl_mult_res_sva_1 = mult_16_z_asn_itm_3 - mult_z_mul_cmp_31_z;
  assign mult_res_sva_1 = nl_mult_res_sva_1[31:0];
  assign INNER_LOOP4_nor_tmp = ~(INNER_LOOP1_stage_0 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm
      | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2
      | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4
      | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6
      | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10);
  assign or_dcpl_13 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 | INNER_LOOP1_stage_0_8;
  assign or_dcpl_22 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 | INNER_LOOP1_stage_0_7;
  assign or_dcpl_45 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 | INNER_LOOP1_stage_0_6;
  assign or_dcpl_65 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 | INNER_LOOP1_stage_0_5;
  assign or_dcpl_101 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 | INNER_LOOP1_stage_0_4;
  assign or_dcpl_121 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 | INNER_LOOP1_stage_0_3;
  assign and_dcpl_51 = INNER_LOOP4_nor_tmp & c_1_sva;
  assign and_dcpl_56 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 & (~ INNER_LOOP1_stage_0_9);
  assign and_dcpl_57 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 & (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9);
  assign or_dcpl_194 = (fsm_output[4]) | (fsm_output[9]);
  assign and_dcpl_58 = INNER_LOOP1_stage_0_9 & (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8);
  assign and_dcpl_59 = (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9) & INNER_LOOP1_stage_0_10;
  assign or_dcpl_197 = (~ INNER_LOOP1_stage_0_9) | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8;
  assign or_dcpl_198 = (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7) | INNER_LOOP1_stage_0_9;
  assign or_dcpl_199 = (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10) | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9;
  assign or_dcpl_200 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 | (~ INNER_LOOP1_stage_0_10);
  assign and_dcpl_67 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 & INNER_LOOP1_stage_0_9;
  assign and_dcpl_68 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9;
  assign and_dcpl_69 = INNER_LOOP1_stage_0_9 & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8;
  assign and_dcpl_70 = INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 & INNER_LOOP1_stage_0_10;
  assign or_dcpl_205 = ~(INNER_LOOP1_stage_0_9 & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8);
  assign or_dcpl_206 = ~(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 & INNER_LOOP1_stage_0_9);
  assign or_dcpl_207 = ~(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 & INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9);
  assign or_dcpl_208 = ~(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 & INNER_LOOP1_stage_0_10);
  assign or_dcpl_210 = (fsm_output[2]) | (fsm_output[7]);
  assign or_dcpl_212 = (fsm_output[7]) | (fsm_output[9]);
  assign or_dcpl_214 = modulo_add_1_qelse_or_m1c | or_dcpl_212;
  assign and_dcpl_79 = INNER_LOOP1_stage_0 & (operator_20_false_acc_cse_sva[0]);
  assign and_dcpl_81 = INNER_LOOP1_stage_0 & (operator_20_false_acc_cse_sva[1]);
  assign and_dcpl_82 = INNER_LOOP1_stage_0 & (operator_33_true_3_lshift_psp_1_0_sva[1]);
  assign or_dcpl_217 = (fsm_output[4]) | (fsm_output[7]);
  assign or_dcpl_218 = or_dcpl_217 | (fsm_output[9]);
  assign and_dcpl_90 = ~((fsm_output[7]) | (fsm_output[9]));
  assign or_dcpl_233 = (fsm_output[4:3]!=2'b00);
  assign and_167_cse = (INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm | INNER_LOOP1_stage_0)
      & or_dcpl_194;
  assign or_tmp_21 = and_dcpl_58 & (fsm_output[2]);
  assign or_tmp_22 = or_dcpl_197 & (fsm_output[2]);
  assign or_tmp_25 = and_dcpl_56 & (fsm_output[7]);
  assign or_tmp_26 = or_dcpl_198 & (fsm_output[7]);
  assign and_192_cse = ~((fsm_output[2]) | (fsm_output[7]));
  assign or_tmp_203 = and_dcpl_69 & (fsm_output[2]);
  assign or_tmp_204 = or_dcpl_205 & (fsm_output[2]);
  assign or_tmp_207 = and_dcpl_67 & (fsm_output[7]);
  assign or_tmp_208 = or_dcpl_206 & (fsm_output[7]);
  assign nor_7_cse = ~((fsm_output[4]) | (fsm_output[9]));
  assign and_1445_cse = INNER_LOOP1_stage_0 & (operator_33_true_3_lshift_psp_1_0_sva[0])
      & (fsm_output[9]);
  assign and_1454_cse = and_dcpl_82 & (fsm_output[9]);
  assign and_1463_cse = and_dcpl_82 & (operator_33_true_3_lshift_psp_1_0_sva[0])
      & (fsm_output[9]);
  assign or_tmp_771 = modulo_add_1_qelse_or_m1c | (fsm_output[9]);
  assign and_1700_cse = (~ (operator_33_true_3_lshift_psp_1_0_sva[0])) & (fsm_output[9]);
  assign or_tmp_779 = and_1700_cse | modulo_add_1_qelse_or_m1c;
  assign or_tmp_782 = (operator_33_true_3_lshift_psp_1_0_sva[0]) & (fsm_output[9]);
  assign and_1719_cse = (~ (operator_33_true_3_lshift_psp_1_0_sva[1])) & (fsm_output[9]);
  assign or_tmp_790 = (operator_20_false_acc_cse_sva[2]) & (fsm_output[7]);
  assign and_1725_cse = (~ (operator_20_false_acc_cse_sva[2])) & (fsm_output[7]);
  assign or_tmp_792 = (operator_33_true_3_lshift_psp_1_0_sva[1]) & (fsm_output[9]);
  assign or_tmp_809 = (operator_20_false_acc_cse_sva[1]) & (fsm_output[7]);
  assign and_1763_cse = (~ (operator_20_false_acc_cse_sva[1])) & (fsm_output[7]);
  assign or_tmp_819 = (operator_20_false_acc_cse_sva[0]) & (fsm_output[7]);
  assign and_1783_cse = (~ (operator_20_false_acc_cse_sva[0])) & (fsm_output[7]);
  assign or_tmp_885 = and_1763_cse | modulo_add_1_qelse_or_m1c;
  assign or_tmp_894 = and_1783_cse | modulo_add_1_qelse_or_m1c;
  assign or_tmp_1134 = (fsm_output[7:6]!=2'b00);
  assign or_tmp_1138 = (~ (fsm_output[4])) & (~ (fsm_output[2])) & and_dcpl_90;
  assign or_tmp_1189 = (fsm_output[2]) | (fsm_output[9]);
  assign yt_rsc_0_0_i_wea_d_mx0c0 = (or_dcpl_199 & or_dcpl_198 & (fsm_output[7]))
      | and_192_cse | (or_dcpl_200 & or_dcpl_197 & (fsm_output[2]));
  assign yt_rsc_0_0_i_wea_d_mx0c2 = (and_dcpl_57 & or_dcpl_198 & (fsm_output[7]))
      | (and_dcpl_59 & or_dcpl_197 & (fsm_output[2]));
  assign yt_rsc_0_16_i_wea_d_mx0c0 = (or_dcpl_207 & or_dcpl_206 & (fsm_output[7]))
      | and_192_cse | (or_dcpl_208 & or_dcpl_205 & (fsm_output[2]));
  assign yt_rsc_0_16_i_wea_d_mx0c2 = (and_dcpl_68 & or_dcpl_206 & (fsm_output[7]))
      | (and_dcpl_70 & or_dcpl_205 & (fsm_output[2]));
  assign butterFly1_nor_7_rmff = ~(or_tmp_21 | or_tmp_25);
  assign butterFly1_mux_17_cse = MUX_s_1_2_2((INNER_LOOP2_r_11_4_sva_6_0[6]), (INNER_LOOP4_r_11_4_sva_6_0[6]),
      fsm_output[9]);
  assign butterFly1_butterFly1_and_17_rmff = butterFly1_mux_17_cse & (~(or_tmp_21
      | or_tmp_22 | or_tmp_25 | or_tmp_26));
  assign butterFly1_or_5_cse = or_tmp_25 | or_tmp_26;
  assign butterFly1_or_1_cse = or_tmp_21 | or_tmp_22;
  assign butterFly1_mux1h_15_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign butterFly1_1_mux1h_11_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign butterFly1_2_mux1h_11_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign butterFly1_3_mux1h_11_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign butterFly1_4_mux1h_11_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign butterFly1_8_mux1h_11_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign butterFly1_nor_4_rmff = ~(or_tmp_203 | or_tmp_207);
  assign butterFly1_butterFly1_and_15_rmff = butterFly1_mux_17_cse & (~(or_tmp_203
      | or_tmp_204 | or_tmp_207 | or_tmp_208));
  assign butterFly1_or_4_cse = or_tmp_207 | or_tmp_208;
  assign butterFly1_or_cse = or_tmp_203 | or_tmp_204;
  assign butterFly1_mux1h_13_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign butterFly1_1_mux1h_9_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign butterFly1_2_mux1h_9_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign butterFly1_3_mux1h_9_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign butterFly1_4_mux1h_9_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign butterFly1_8_mux1h_9_rmff = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign butterFly1_15_f2_mux1h_65_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_f1_butterFly1_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1}), modulo_add_10_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_f1_butterFly1_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_64_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_f2_butterFly1_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1}), modulo_add_11_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_f2_butterFly1_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_63_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1}), modulo_add_12_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_62_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1}), modulo_add_13_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_61_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1}), modulo_add_14_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_60_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1}), modulo_add_15_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_59_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1}), modulo_add_1_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_58_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1}), modulo_add_23_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_57_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1}), modulo_add_24_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_56_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1}), modulo_add_25_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_55_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1}), modulo_add_26_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_54_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1}), modulo_add_27_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_53_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1}), modulo_add_28_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_52_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1}), modulo_add_29_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_51_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1}), modulo_add_30_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff = MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign butterFly1_15_f2_mux1h_50_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      ({1'b0 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1}), INNER_LOOP3_r_11_4_sva_6_0,
      ({1'b1 , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2}), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff = MUX_v_32_2_2(({reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd
      , reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1}), modulo_add_31_qr_lpi_3_dfm_1, fsm_output[9]);
  assign butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff = MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1,
      ({reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd , reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1}),
      fsm_output[9]);
  assign INNER_LOOP1_tw_and_nl = INNER_LOOP2_r_11_4_sva_6_0 & INNER_LOOP1_r_11_4_sva_6_0;
  assign INNER_LOOP2_tw_and_nl = operator_33_true_1_lshift_psp_9_4_sva & (INNER_LOOP2_r_11_4_sva_6_0[5:0]);
  assign INNER_LOOP1_tw_h_mux1h_4_rmff = MUX1HOT_v_7_4_2(INNER_LOOP1_tw_and_nl, ({(INNER_LOOP2_r_11_4_sva_6_0[6])
      , INNER_LOOP2_tw_and_nl}), INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign butterFly1_butterFly1_or_1_rmff = or_tmp_21 | or_tmp_25;
  assign butterFly1_butterFly1_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse, or_tmp_25);
  assign butterFly1_1_butterFly1_1_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse, or_tmp_25);
  assign butterFly1_2_butterFly1_2_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse, or_tmp_25);
  assign butterFly1_3_butterFly1_3_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse, or_tmp_25);
  assign butterFly1_4_butterFly1_4_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse, or_tmp_25);
  assign butterFly1_7_butterFly1_7_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse, or_tmp_25);
  assign butterFly1_8_butterFly1_8_mux_3_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse, or_tmp_25);
  assign butterFly1_butterFly1_or_rmff = or_tmp_203 | or_tmp_207;
  assign butterFly1_butterFly1_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse, or_tmp_207);
  assign butterFly1_1_butterFly1_1_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse, or_tmp_207);
  assign butterFly1_2_butterFly1_2_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse, or_tmp_207);
  assign butterFly1_3_butterFly1_3_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse, or_tmp_207);
  assign butterFly1_4_butterFly1_4_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse, or_tmp_207);
  assign butterFly1_7_butterFly1_7_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse, or_tmp_207);
  assign butterFly1_8_butterFly1_8_mux_4_rmff = MUX_v_6_2_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse,
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse, or_tmp_207);
  assign butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff = ~(nor_7_cse
      | (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10) | INNER_LOOP1_stage_0_9);
  assign butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff = ~(nor_7_cse
      | (~ INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10) | (~ INNER_LOOP1_stage_0_9));
  assign yt_rsc_0_0_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_butterFly1_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_mux1h_15_rmff};
  assign butterFly1_butterFly1_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_0_i_da_d_mx0w0_63_32,
      yt_rsc_0_0_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_butterFly1_mux_6_nl = MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1,
      modulo_add_10_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_0_i_da_d = {butterFly1_butterFly1_mux_2_nl , butterFly1_butterFly1_mux_6_nl};
  assign butterFly1_butterFly1_nor_2_nl = ~(yt_rsc_0_0_i_wea_d_mx0c2 | yt_rsc_0_0_i_wea_d_mx0c0);
  assign butterFly1_mux_15_nl = MUX_s_1_2_2((~ or_dcpl_200), (~ or_dcpl_199), or_tmp_25);
  assign butterFly1_butterFly1_nor_3_nl = ~((~(butterFly1_mux_15_nl | yt_rsc_0_0_i_wea_d_mx0c2))
      | yt_rsc_0_0_i_wea_d_mx0c0);
  assign yt_rsc_0_0_i_wea_d_pff = {butterFly1_butterFly1_nor_2_nl , butterFly1_butterFly1_nor_3_nl};
  assign yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_1_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_1_butterFly1_1_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_1_mux1h_11_rmff};
  assign butterFly1_1_butterFly1_1_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_1_i_da_d_mx0w0_63_32,
      yt_rsc_0_1_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_1_butterFly1_1_mux_6_nl = MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1,
      modulo_add_11_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_1_i_da_d = {butterFly1_1_butterFly1_1_mux_2_nl , butterFly1_1_butterFly1_1_mux_6_nl};
  assign yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_2_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_2_butterFly1_2_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_2_mux1h_11_rmff};
  assign butterFly1_2_butterFly1_2_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_2_i_da_d_mx0w0_63_32,
      yt_rsc_0_2_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_2_butterFly1_2_mux_6_nl = MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1,
      modulo_add_12_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_2_i_da_d = {butterFly1_2_butterFly1_2_mux_2_nl , butterFly1_2_butterFly1_2_mux_6_nl};
  assign yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_3_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_3_butterFly1_3_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_3_mux1h_11_rmff};
  assign butterFly1_3_butterFly1_3_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_3_i_da_d_mx0w0_63_32,
      yt_rsc_0_3_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_3_butterFly1_3_mux_6_nl = MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1,
      modulo_add_13_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_3_i_da_d = {butterFly1_3_butterFly1_3_mux_2_nl , butterFly1_3_butterFly1_3_mux_6_nl};
  assign yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_4_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_4_butterFly1_4_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_4_mux1h_11_rmff};
  assign butterFly1_4_butterFly1_4_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_4_i_da_d_mx0w0_63_32,
      yt_rsc_0_4_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_4_butterFly1_4_mux_6_nl = MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1,
      modulo_add_14_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_4_i_da_d = {butterFly1_4_butterFly1_4_mux_2_nl , butterFly1_4_butterFly1_4_mux_6_nl};
  assign yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_5_butterFly1_5_mux_3_nl = MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9, or_tmp_25);
  assign butterFly1_5_mux1h_11_nl = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign yt_rsc_0_5_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_5_butterFly1_5_mux_3_nl , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_5_mux1h_11_nl};
  assign butterFly1_5_butterFly1_5_mux_2_nl = MUX_v_32_2_2(modulo_sub_5_qelse_mux_cse,
      yt_rsc_0_5_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_5_butterFly1_5_mux_6_nl = MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1,
      modulo_add_15_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_5_i_da_d = {butterFly1_5_butterFly1_5_mux_2_nl , butterFly1_5_butterFly1_5_mux_6_nl};
  assign yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_6_butterFly1_6_mux_3_nl = MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9, or_tmp_25);
  assign butterFly1_6_mux1h_11_nl = MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign yt_rsc_0_6_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_6_butterFly1_6_mux_3_nl , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_6_mux1h_11_nl};
  assign butterFly1_6_butterFly1_6_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_6_i_da_d_mx0w0_63_32,
      yt_rsc_0_6_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_6_butterFly1_6_mux_6_nl = MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1,
      modulo_add_1_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_6_i_da_d = {butterFly1_6_butterFly1_6_mux_2_nl , butterFly1_6_butterFly1_6_mux_6_nl};
  assign yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_7_mux1h_11_nl = MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign yt_rsc_0_7_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_7_butterFly1_7_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_7_mux1h_11_nl};
  assign butterFly1_7_butterFly1_7_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_7_i_da_d_mx0w0_63_32,
      modulo_sub_5_qelse_mux_cse, or_tmp_25);
  assign butterFly1_7_butterFly1_7_mux_6_nl = MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1,
      modulo_add_23_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_7_i_da_d = {butterFly1_7_butterFly1_7_mux_2_nl , butterFly1_7_butterFly1_7_mux_6_nl};
  assign yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_8_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_8_butterFly1_8_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_8_mux1h_11_rmff};
  assign butterFly1_8_butterFly1_8_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_8_i_da_d_mx0w0_63_32,
      yt_rsc_0_8_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_8_butterFly1_8_mux_6_nl = MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1,
      modulo_add_24_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_8_i_da_d = {butterFly1_8_butterFly1_8_mux_2_nl , butterFly1_8_butterFly1_8_mux_6_nl};
  assign yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_9_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_butterFly1_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_mux1h_15_rmff};
  assign butterFly1_9_butterFly1_9_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_9_i_da_d_mx0w0_63_32,
      yt_rsc_0_9_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_9_butterFly1_9_mux_6_nl = MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1,
      modulo_add_25_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_9_i_da_d = {butterFly1_9_butterFly1_9_mux_2_nl , butterFly1_9_butterFly1_9_mux_6_nl};
  assign yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_10_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_1_butterFly1_1_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_1_mux1h_11_rmff};
  assign butterFly1_10_butterFly1_10_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_10_i_da_d_mx0w0_63_32,
      yt_rsc_0_10_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_10_butterFly1_10_mux_6_nl = MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1,
      modulo_add_26_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_10_i_da_d = {butterFly1_10_butterFly1_10_mux_2_nl , butterFly1_10_butterFly1_10_mux_6_nl};
  assign yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_11_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_2_butterFly1_2_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_2_mux1h_11_rmff};
  assign butterFly1_11_butterFly1_11_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_11_i_da_d_mx0w0_63_32,
      yt_rsc_0_11_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_11_butterFly1_11_mux_6_nl = MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1,
      modulo_add_27_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_11_i_da_d = {butterFly1_11_butterFly1_11_mux_2_nl , butterFly1_11_butterFly1_11_mux_6_nl};
  assign yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_12_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_3_butterFly1_3_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_3_mux1h_11_rmff};
  assign butterFly1_12_butterFly1_12_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_12_i_da_d_mx0w0_63_32,
      yt_rsc_0_12_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_12_butterFly1_12_mux_6_nl = MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1,
      modulo_add_28_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_12_i_da_d = {butterFly1_12_butterFly1_12_mux_2_nl , butterFly1_12_butterFly1_12_mux_6_nl};
  assign yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_13_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_4_butterFly1_4_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_4_mux1h_11_rmff};
  assign butterFly1_13_butterFly1_13_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_13_i_da_d_mx0w0_63_32,
      yt_rsc_0_13_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_13_butterFly1_13_mux_6_nl = MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1,
      modulo_add_29_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_13_i_da_d = {butterFly1_13_butterFly1_13_mux_2_nl , butterFly1_13_butterFly1_13_mux_6_nl};
  assign yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_14_mux1h_11_nl = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_1_cse , (fsm_output[4]) ,
      butterFly1_or_5_cse , (fsm_output[9])});
  assign yt_rsc_0_14_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_7_butterFly1_7_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_14_mux1h_11_nl};
  assign butterFly1_14_butterFly1_14_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_14_i_da_d_mx0w0_63_32,
      yt_rsc_0_14_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_14_butterFly1_14_mux_6_nl = MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1,
      modulo_add_30_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_14_i_da_d = {butterFly1_14_butterFly1_14_mux_2_nl , butterFly1_14_butterFly1_14_mux_6_nl};
  assign yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_15_i_adra_d = {butterFly1_nor_7_rmff , butterFly1_butterFly1_or_1_rmff
      , butterFly1_8_butterFly1_8_mux_3_rmff , 1'b0 , butterFly1_butterFly1_and_17_rmff
      , butterFly1_8_mux1h_11_rmff};
  assign butterFly1_15_butterFly1_15_mux_2_nl = MUX_v_32_2_2(yt_rsc_0_15_i_da_d_mx0w0_63_32,
      yt_rsc_0_15_i_da_d_mx0w2_63_32, or_tmp_25);
  assign butterFly1_15_butterFly1_15_mux_6_nl = MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1,
      modulo_add_31_qr_lpi_3_dfm_1, butterFly1_or_5_cse);
  assign yt_rsc_0_15_i_da_d = {butterFly1_15_butterFly1_15_mux_2_nl , butterFly1_15_butterFly1_15_mux_6_nl};
  assign yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_16_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_butterFly1_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_mux1h_13_rmff};
  assign butterFly1_butterFly1_mux_nl = MUX_v_32_2_2(yt_rsc_0_0_i_da_d_mx0w0_63_32,
      yt_rsc_0_0_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_butterFly1_mux_5_nl = MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1,
      modulo_add_10_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_16_i_da_d = {butterFly1_butterFly1_mux_nl , butterFly1_butterFly1_mux_5_nl};
  assign butterFly1_butterFly1_nor_nl = ~(yt_rsc_0_16_i_wea_d_mx0c2 | yt_rsc_0_16_i_wea_d_mx0c0);
  assign butterFly1_mux_nl = MUX_s_1_2_2((~ or_dcpl_208), (~ or_dcpl_207), or_tmp_207);
  assign butterFly1_butterFly1_nor_1_nl = ~((~(butterFly1_mux_nl | yt_rsc_0_16_i_wea_d_mx0c2))
      | yt_rsc_0_16_i_wea_d_mx0c0);
  assign yt_rsc_0_16_i_wea_d_pff = {butterFly1_butterFly1_nor_nl , butterFly1_butterFly1_nor_1_nl};
  assign yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_17_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_1_butterFly1_1_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_1_mux1h_9_rmff};
  assign butterFly1_1_butterFly1_1_mux_nl = MUX_v_32_2_2(yt_rsc_0_1_i_da_d_mx0w0_63_32,
      yt_rsc_0_1_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_1_butterFly1_1_mux_5_nl = MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1,
      modulo_add_11_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_17_i_da_d = {butterFly1_1_butterFly1_1_mux_nl , butterFly1_1_butterFly1_1_mux_5_nl};
  assign yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_18_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_2_butterFly1_2_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_2_mux1h_9_rmff};
  assign butterFly1_2_butterFly1_2_mux_nl = MUX_v_32_2_2(yt_rsc_0_2_i_da_d_mx0w0_63_32,
      yt_rsc_0_2_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_2_butterFly1_2_mux_5_nl = MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1,
      modulo_add_12_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_18_i_da_d = {butterFly1_2_butterFly1_2_mux_nl , butterFly1_2_butterFly1_2_mux_5_nl};
  assign yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_19_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_3_butterFly1_3_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_3_mux1h_9_rmff};
  assign butterFly1_3_butterFly1_3_mux_nl = MUX_v_32_2_2(yt_rsc_0_3_i_da_d_mx0w0_63_32,
      yt_rsc_0_3_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_3_butterFly1_3_mux_5_nl = MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1,
      modulo_add_13_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_19_i_da_d = {butterFly1_3_butterFly1_3_mux_nl , butterFly1_3_butterFly1_3_mux_5_nl};
  assign yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_20_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_4_butterFly1_4_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_4_mux1h_9_rmff};
  assign butterFly1_4_butterFly1_4_mux_nl = MUX_v_32_2_2(yt_rsc_0_4_i_da_d_mx0w0_63_32,
      yt_rsc_0_4_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_4_butterFly1_4_mux_5_nl = MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1,
      modulo_add_14_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_20_i_da_d = {butterFly1_4_butterFly1_4_mux_nl , butterFly1_4_butterFly1_4_mux_5_nl};
  assign yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_5_butterFly1_5_mux_4_nl = MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9, or_tmp_207);
  assign butterFly1_5_mux1h_9_nl = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign yt_rsc_0_21_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_5_butterFly1_5_mux_4_nl , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_5_mux1h_9_nl};
  assign butterFly1_5_butterFly1_5_mux_nl = MUX_v_32_2_2(modulo_sub_5_qelse_mux_cse,
      yt_rsc_0_5_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_5_butterFly1_5_mux_5_nl = MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1,
      modulo_add_15_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_21_i_da_d = {butterFly1_5_butterFly1_5_mux_nl , butterFly1_5_butterFly1_5_mux_5_nl};
  assign yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_6_butterFly1_6_mux_4_nl = MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9, or_tmp_207);
  assign butterFly1_6_mux1h_9_nl = MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign yt_rsc_0_22_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_6_butterFly1_6_mux_4_nl , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_6_mux1h_9_nl};
  assign butterFly1_6_butterFly1_6_mux_nl = MUX_v_32_2_2(yt_rsc_0_6_i_da_d_mx0w0_63_32,
      yt_rsc_0_6_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_6_butterFly1_6_mux_5_nl = MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1,
      modulo_add_1_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_22_i_da_d = {butterFly1_6_butterFly1_6_mux_nl , butterFly1_6_butterFly1_6_mux_5_nl};
  assign yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_7_mux1h_9_nl = MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign yt_rsc_0_23_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_7_butterFly1_7_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_7_mux1h_9_nl};
  assign butterFly1_7_butterFly1_7_mux_nl = MUX_v_32_2_2(yt_rsc_0_7_i_da_d_mx0w0_63_32,
      modulo_sub_5_qelse_mux_cse, or_tmp_207);
  assign butterFly1_7_butterFly1_7_mux_5_nl = MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1,
      modulo_add_23_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_23_i_da_d = {butterFly1_7_butterFly1_7_mux_nl , butterFly1_7_butterFly1_7_mux_5_nl};
  assign yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_24_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_8_butterFly1_8_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_8_mux1h_9_rmff};
  assign butterFly1_8_butterFly1_8_mux_nl = MUX_v_32_2_2(yt_rsc_0_8_i_da_d_mx0w0_63_32,
      yt_rsc_0_8_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_8_butterFly1_8_mux_5_nl = MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1,
      modulo_add_24_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_24_i_da_d = {butterFly1_8_butterFly1_8_mux_nl , butterFly1_8_butterFly1_8_mux_5_nl};
  assign yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_25_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_butterFly1_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_mux1h_13_rmff};
  assign butterFly1_9_butterFly1_9_mux_nl = MUX_v_32_2_2(yt_rsc_0_9_i_da_d_mx0w0_63_32,
      yt_rsc_0_9_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_9_butterFly1_9_mux_5_nl = MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1,
      modulo_add_25_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_25_i_da_d = {butterFly1_9_butterFly1_9_mux_nl , butterFly1_9_butterFly1_9_mux_5_nl};
  assign yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_26_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_1_butterFly1_1_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_1_mux1h_9_rmff};
  assign butterFly1_10_butterFly1_10_mux_nl = MUX_v_32_2_2(yt_rsc_0_10_i_da_d_mx0w0_63_32,
      yt_rsc_0_10_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_10_butterFly1_10_mux_5_nl = MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1,
      modulo_add_26_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_26_i_da_d = {butterFly1_10_butterFly1_10_mux_nl , butterFly1_10_butterFly1_10_mux_5_nl};
  assign yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_27_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_2_butterFly1_2_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_2_mux1h_9_rmff};
  assign butterFly1_11_butterFly1_11_mux_nl = MUX_v_32_2_2(yt_rsc_0_11_i_da_d_mx0w0_63_32,
      yt_rsc_0_11_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_11_butterFly1_11_mux_5_nl = MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1,
      modulo_add_27_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_27_i_da_d = {butterFly1_11_butterFly1_11_mux_nl , butterFly1_11_butterFly1_11_mux_5_nl};
  assign yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_28_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_3_butterFly1_3_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_3_mux1h_9_rmff};
  assign butterFly1_12_butterFly1_12_mux_nl = MUX_v_32_2_2(yt_rsc_0_12_i_da_d_mx0w0_63_32,
      yt_rsc_0_12_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_12_butterFly1_12_mux_5_nl = MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1,
      modulo_add_28_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_28_i_da_d = {butterFly1_12_butterFly1_12_mux_nl , butterFly1_12_butterFly1_12_mux_5_nl};
  assign yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_29_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_4_butterFly1_4_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_4_mux1h_9_rmff};
  assign butterFly1_13_butterFly1_13_mux_nl = MUX_v_32_2_2(yt_rsc_0_13_i_da_d_mx0w0_63_32,
      yt_rsc_0_13_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_13_butterFly1_13_mux_5_nl = MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1,
      modulo_add_29_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_29_i_da_d = {butterFly1_13_butterFly1_13_mux_nl , butterFly1_13_butterFly1_13_mux_5_nl};
  assign yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign butterFly1_14_mux1h_9_nl = MUX1HOT_v_6_4_2(reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse,
      (INNER_LOOP2_r_11_4_sva_6_0[5:0]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
      (INNER_LOOP4_r_11_4_sva_6_0[5:0]), {butterFly1_or_cse , (fsm_output[4]) , butterFly1_or_4_cse
      , (fsm_output[9])});
  assign yt_rsc_0_30_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_7_butterFly1_7_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_14_mux1h_9_nl};
  assign butterFly1_14_butterFly1_14_mux_nl = MUX_v_32_2_2(yt_rsc_0_14_i_da_d_mx0w0_63_32,
      yt_rsc_0_14_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_14_butterFly1_14_mux_5_nl = MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1,
      modulo_add_30_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_30_i_da_d = {butterFly1_14_butterFly1_14_mux_nl , butterFly1_14_butterFly1_14_mux_5_nl};
  assign yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign yt_rsc_0_31_i_adra_d = {butterFly1_nor_4_rmff , butterFly1_butterFly1_or_rmff
      , butterFly1_8_butterFly1_8_mux_4_rmff , 1'b0 , butterFly1_butterFly1_and_15_rmff
      , butterFly1_8_mux1h_9_rmff};
  assign butterFly1_15_butterFly1_15_mux_nl = MUX_v_32_2_2(yt_rsc_0_15_i_da_d_mx0w0_63_32,
      yt_rsc_0_15_i_da_d_mx0w2_63_32, or_tmp_207);
  assign butterFly1_15_butterFly1_15_mux_5_nl = MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1,
      modulo_add_31_qr_lpi_3_dfm_1, butterFly1_or_4_cse);
  assign yt_rsc_0_31_i_da_d = {butterFly1_15_butterFly1_15_mux_nl , butterFly1_15_butterFly1_15_mux_5_nl};
  assign yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_202_rmff};
  assign xt_rsc_0_0_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3
      , 1'b0 , butterFly1_15_f2_mux1h_65_rmff};
  assign xt_rsc_0_0_i_da_d = {butterFly1_f1_butterFly1_f1_mux_2_rmff , butterFly1_f1_butterFly1_f1_mux_3_rmff};
  assign xt_rsc_0_0_i_wea_d_pff = {butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff
      , butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_f1_nor_rmff};
  assign xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_1_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4
      , 1'b0 , butterFly1_15_f2_mux1h_64_rmff};
  assign xt_rsc_0_1_i_da_d = {butterFly1_f2_butterFly1_f2_mux_2_rmff , butterFly1_f2_butterFly1_f2_mux_3_rmff};
  assign xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_2_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5
      , 1'b0 , butterFly1_15_f2_mux1h_63_rmff};
  assign xt_rsc_0_2_i_da_d = {butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff , butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff};
  assign xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_3_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6
      , 1'b0 , butterFly1_15_f2_mux1h_62_rmff};
  assign xt_rsc_0_3_i_da_d = {butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff , butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff};
  assign xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_4_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7
      , 1'b0 , butterFly1_15_f2_mux1h_61_rmff};
  assign xt_rsc_0_4_i_da_d = {butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff , butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff};
  assign xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_5_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8
      , 1'b0 , butterFly1_15_f2_mux1h_60_rmff};
  assign xt_rsc_0_5_i_da_d = {butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff , butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff};
  assign xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_6_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9
      , 1'b0 , butterFly1_15_f2_mux1h_59_rmff};
  assign xt_rsc_0_6_i_da_d = {butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff , butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff};
  assign xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_7_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1
      , 1'b0 , butterFly1_15_f2_mux1h_58_rmff};
  assign xt_rsc_0_7_i_da_d = {butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff , butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff};
  assign xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_8_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2
      , 1'b0 , butterFly1_15_f2_mux1h_57_rmff};
  assign xt_rsc_0_8_i_da_d = {butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff , butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff};
  assign xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_9_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3
      , 1'b0 , butterFly1_15_f2_mux1h_56_rmff};
  assign xt_rsc_0_9_i_da_d = {butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff , butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff};
  assign xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_10_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4
      , 1'b0 , butterFly1_15_f2_mux1h_55_rmff};
  assign xt_rsc_0_10_i_da_d = {butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff , butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff};
  assign xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_11_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5
      , 1'b0 , butterFly1_15_f2_mux1h_54_rmff};
  assign xt_rsc_0_11_i_da_d = {butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff , butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff};
  assign xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_12_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6
      , 1'b0 , butterFly1_15_f2_mux1h_53_rmff};
  assign xt_rsc_0_12_i_da_d = {butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff , butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff};
  assign xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_13_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9
      , 1'b0 , butterFly1_15_f2_mux1h_52_rmff};
  assign xt_rsc_0_13_i_da_d = {butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff , butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff};
  assign xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_14_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1
      , 1'b0 , butterFly1_15_f2_mux1h_51_rmff};
  assign xt_rsc_0_14_i_da_d = {butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff , butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff};
  assign xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_15_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2
      , 1'b0 , butterFly1_15_f2_mux1h_50_rmff};
  assign xt_rsc_0_15_i_da_d = {butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff , butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff};
  assign xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_16_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3
      , 1'b0 , butterFly1_15_f2_mux1h_65_rmff};
  assign xt_rsc_0_16_i_da_d = {butterFly1_f1_butterFly1_f1_mux_2_rmff , butterFly1_f1_butterFly1_f1_mux_3_rmff};
  assign xt_rsc_0_16_i_wea_d_pff = {butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff
      , butterFly1_f1_butterFly1_f1_butterFly1_f1_butterFly1_8_f1_nor_rmff};
  assign xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_17_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4
      , 1'b0 , butterFly1_15_f2_mux1h_64_rmff};
  assign xt_rsc_0_17_i_da_d = {butterFly1_f2_butterFly1_f2_mux_2_rmff , butterFly1_f2_butterFly1_f2_mux_3_rmff};
  assign xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_18_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5
      , 1'b0 , butterFly1_15_f2_mux1h_63_rmff};
  assign xt_rsc_0_18_i_da_d = {butterFly1_1_f1_butterFly1_1_f1_mux_2_rmff , butterFly1_1_f1_butterFly1_1_f1_mux_3_rmff};
  assign xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_19_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6
      , 1'b0 , butterFly1_15_f2_mux1h_62_rmff};
  assign xt_rsc_0_19_i_da_d = {butterFly1_1_f2_butterFly1_1_f2_mux_2_rmff , butterFly1_1_f2_butterFly1_1_f2_mux_3_rmff};
  assign xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_20_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7
      , 1'b0 , butterFly1_15_f2_mux1h_61_rmff};
  assign xt_rsc_0_20_i_da_d = {butterFly1_2_f1_butterFly1_2_f1_mux_2_rmff , butterFly1_2_f1_butterFly1_2_f1_mux_3_rmff};
  assign xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_21_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8
      , 1'b0 , butterFly1_15_f2_mux1h_60_rmff};
  assign xt_rsc_0_21_i_da_d = {butterFly1_2_f2_butterFly1_2_f2_mux_2_rmff , butterFly1_2_f2_butterFly1_2_f2_mux_3_rmff};
  assign xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_22_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9
      , 1'b0 , butterFly1_15_f2_mux1h_59_rmff};
  assign xt_rsc_0_22_i_da_d = {butterFly1_3_f1_butterFly1_3_f1_mux_2_rmff , butterFly1_3_f1_butterFly1_3_f1_mux_3_rmff};
  assign xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_23_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1
      , 1'b0 , butterFly1_15_f2_mux1h_58_rmff};
  assign xt_rsc_0_23_i_da_d = {butterFly1_3_f2_butterFly1_3_f2_mux_2_rmff , butterFly1_3_f2_butterFly1_3_f2_mux_3_rmff};
  assign xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_24_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2
      , 1'b0 , butterFly1_15_f2_mux1h_57_rmff};
  assign xt_rsc_0_24_i_da_d = {butterFly1_4_f1_butterFly1_4_f1_mux_2_rmff , butterFly1_4_f1_butterFly1_4_f1_mux_3_rmff};
  assign xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_25_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3
      , 1'b0 , butterFly1_15_f2_mux1h_56_rmff};
  assign xt_rsc_0_25_i_da_d = {butterFly1_4_f2_butterFly1_4_f2_mux_2_rmff , butterFly1_4_f2_butterFly1_4_f2_mux_3_rmff};
  assign xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_26_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4
      , 1'b0 , butterFly1_15_f2_mux1h_55_rmff};
  assign xt_rsc_0_26_i_da_d = {butterFly1_5_f1_butterFly1_5_f1_mux_2_rmff , butterFly1_5_f1_butterFly1_5_f1_mux_3_rmff};
  assign xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_27_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5
      , 1'b0 , butterFly1_15_f2_mux1h_54_rmff};
  assign xt_rsc_0_27_i_da_d = {butterFly1_5_f2_butterFly1_5_f2_mux_2_rmff , butterFly1_5_f2_butterFly1_5_f2_mux_3_rmff};
  assign xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_28_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6
      , 1'b0 , butterFly1_15_f2_mux1h_53_rmff};
  assign xt_rsc_0_28_i_da_d = {butterFly1_6_f1_butterFly1_6_f1_mux_2_rmff , butterFly1_6_f1_butterFly1_6_f1_mux_3_rmff};
  assign xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_29_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9
      , 1'b0 , butterFly1_15_f2_mux1h_52_rmff};
  assign xt_rsc_0_29_i_da_d = {butterFly1_6_f2_butterFly1_6_f2_mux_2_rmff , butterFly1_6_f2_butterFly1_6_f2_mux_3_rmff};
  assign xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_30_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1
      , 1'b0 , butterFly1_15_f2_mux1h_51_rmff};
  assign xt_rsc_0_30_i_da_d = {butterFly1_7_f1_butterFly1_7_f1_mux_2_rmff , butterFly1_7_f1_butterFly1_7_f1_mux_3_rmff};
  assign xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign xt_rsc_0_31_i_adra_d = {nor_7_cse , (~ (fsm_output[9])) , INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2
      , 1'b0 , butterFly1_15_f2_mux1h_50_rmff};
  assign xt_rsc_0_31_i_da_d = {butterFly1_7_f2_butterFly1_7_f2_mux_2_rmff , butterFly1_7_f2_butterFly1_7_f2_mux_3_rmff};
  assign xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_921_rmff};
  assign twiddle_rsc_0_0_i_adra_d = {1'b0 , INNER_LOOP1_tw_h_mux1h_4_rmff};
  assign twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_1435_rmff};
  assign twiddle_rsc_0_1_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_896_rmff};
  assign twiddle_rsc_0_2_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_900_rmff};
  assign twiddle_rsc_0_3_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_904_rmff};
  assign twiddle_rsc_0_4_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_908_rmff};
  assign twiddle_rsc_0_5_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_912_rmff};
  assign twiddle_rsc_0_6_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_916_rmff};
  assign twiddle_rsc_0_7_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_920_rmff};
  assign twiddle_rsc_0_8_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_1506_rmff};
  assign twiddle_rsc_0_9_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_896_rmff};
  assign twiddle_rsc_0_10_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_900_rmff};
  assign twiddle_rsc_0_11_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_904_rmff};
  assign twiddle_rsc_0_12_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_908_rmff};
  assign twiddle_rsc_0_13_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_912_rmff};
  assign twiddle_rsc_0_14_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_916_rmff};
  assign twiddle_rsc_0_15_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_920_rmff};
  assign twiddle_h_rsc_0_0_i_adra_d = {1'b0 , INNER_LOOP1_tw_h_mux1h_4_rmff};
  assign twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_1435_rmff};
  assign twiddle_h_rsc_0_1_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_896_rmff};
  assign twiddle_h_rsc_0_2_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_900_rmff};
  assign twiddle_h_rsc_0_3_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_904_rmff};
  assign twiddle_h_rsc_0_4_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_908_rmff};
  assign twiddle_h_rsc_0_5_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_912_rmff};
  assign twiddle_h_rsc_0_6_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_916_rmff};
  assign twiddle_h_rsc_0_7_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_920_rmff};
  assign twiddle_h_rsc_0_8_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , and_1506_rmff};
  assign twiddle_h_rsc_0_9_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_896_rmff};
  assign twiddle_h_rsc_0_10_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_900_rmff};
  assign twiddle_h_rsc_0_11_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_904_rmff};
  assign twiddle_h_rsc_0_12_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_908_rmff};
  assign twiddle_h_rsc_0_13_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_912_rmff};
  assign twiddle_h_rsc_0_14_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_916_rmff};
  assign twiddle_h_rsc_0_15_i_adra_d = {1'b0 , butterFly2_1_tw_butterFly2_1_tw_mux_rmff};
  assign twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d = {1'b0 , or_920_rmff};
  always @(posedge clk) begin
    if ( (fsm_output[10]) | (fsm_output[0]) ) begin
      p_sva <= p_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      c_1_sva <= 1'b0;
    end
    else if ( (fsm_output[5]) | (fsm_output[0]) | (fsm_output[9]) ) begin
      c_1_sva <= c_mux_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_yt_rsc_0_0_cgo_cse <= 1'b0;
      reg_yt_rsc_0_16_cgo_cse <= 1'b0;
      reg_xt_rsc_triosy_0_31_obj_ld_cse <= 1'b0;
      reg_ensig_cgo_cse <= 1'b0;
      reg_ensig_cgo_17_cse <= 1'b0;
      butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm <= 2'b00;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8 <= 1'b0;
      INNER_LOOP1_stage_0 <= 1'b0;
      INNER_LOOP1_r_11_4_sva_6_0 <= 7'b0000000;
      INNER_LOOP1_stage_0_2 <= 1'b0;
      INNER_LOOP1_stage_0_3 <= 1'b0;
      INNER_LOOP1_stage_0_4 <= 1'b0;
      INNER_LOOP1_stage_0_5 <= 1'b0;
      INNER_LOOP1_stage_0_6 <= 1'b0;
      INNER_LOOP1_stage_0_7 <= 1'b0;
      INNER_LOOP1_stage_0_8 <= 1'b0;
      INNER_LOOP1_stage_0_9 <= 1'b0;
      INNER_LOOP1_stage_0_10 <= 1'b0;
      INNER_LOOP1_stage_0_11 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 <= 1'b0;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm <= 1'b0;
      INNER_LOOP3_r_11_4_sva_6_0 <= 7'b0000000;
      INNER_LOOP4_r_11_4_sva_6_0 <= 7'b0000000;
    end
    else begin
      reg_yt_rsc_0_0_cgo_cse <= or_261_rmff;
      reg_yt_rsc_0_16_cgo_cse <= or_443_rmff;
      reg_xt_rsc_triosy_0_31_obj_ld_cse <= and_dcpl_51 & (fsm_output[9]);
      reg_ensig_cgo_cse <= or_997_rmff;
      reg_ensig_cgo_17_cse <= or_1156_rmff;
      butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm <= MUX_v_2_2_2(STAGE_LOOP_mux1h_nl,
          2'b11, nor_4_nl);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10 <= INNER_LOOP1_r_mux_44_nl
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9 <= MUX_s_1_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8,
          INNER_LOOP1_stage_0_9, fsm_output[7]);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_8 <= INNER_LOOP1_r_mux_45_nl
          & (~ and_192_cse);
      INNER_LOOP1_stage_0 <= (INNER_LOOP1_stage_0 & (~ (z_out_2[7]))) | or_tmp_1138;
      INNER_LOOP1_r_11_4_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (z_out_2[6:0]), (fsm_output[2]));
      INNER_LOOP1_stage_0_2 <= INNER_LOOP1_mux_nl & (~ or_tmp_1138);
      INNER_LOOP1_stage_0_3 <= INNER_LOOP1_stage_0_2 & or_dcpl_214;
      INNER_LOOP1_stage_0_4 <= INNER_LOOP1_stage_0_3 & or_dcpl_214;
      INNER_LOOP1_stage_0_5 <= INNER_LOOP1_stage_0_4 & or_dcpl_214;
      INNER_LOOP1_stage_0_6 <= INNER_LOOP1_stage_0_5 & or_dcpl_214;
      INNER_LOOP1_stage_0_7 <= INNER_LOOP1_stage_0_6 & or_dcpl_214;
      INNER_LOOP1_stage_0_8 <= INNER_LOOP1_stage_0_7 & or_dcpl_214;
      INNER_LOOP1_stage_0_9 <= INNER_LOOP1_stage_0_8 & or_dcpl_214;
      INNER_LOOP1_stage_0_10 <= INNER_LOOP1_r_mux1h_46_nl & (~((fsm_output[10]) |
          (fsm_output[5]) | (fsm_output[6]) | (fsm_output[0]) | (fsm_output[1])));
      INNER_LOOP1_stage_0_11 <= INNER_LOOP1_mux_11_nl & ((fsm_output[6]) | (fsm_output[4])
          | (fsm_output[2]) | (~ and_dcpl_90));
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm
          & (~ or_tmp_1138);
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm <= MUX_s_1_2_2(INNER_LOOP1_r_INNER_LOOP1_r_and_nl,
          INNER_LOOP1_stage_0, or_dcpl_218);
      INNER_LOOP3_r_11_4_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (z_out_2[6:0]), (fsm_output[7]));
      INNER_LOOP4_r_11_4_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (z_out_2[6:0]), (fsm_output[9]));
    end
  end
  always @(posedge clk) begin
    modulo_add_1_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_81, (readslicef_33_32_1(acc_2_nl)),
        z_out_78, z_out_76, {modulo_add_1_qelse_and_nl , modulo_add_1_qelse_or_1_nl
        , modulo_add_1_qelse_and_4_nl , modulo_add_1_qelse_and_5_nl});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    modulo_add_10_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_72, (readslicef_33_32_1(acc_6_nl)),
        z_out_67, z_out_68, z_out_82, {modulo_add_10_qelse_and_nl , modulo_add_10_qelse_or_nl
        , modulo_add_10_qelse_and_5_nl , modulo_add_10_qelse_and_6_nl , modulo_add_10_qelse_and_7_nl});
    modulo_add_11_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_71, (readslicef_33_32_1(acc_10_nl)),
        z_out_77, z_out_67, z_out_81, {modulo_add_11_qelse_and_nl , modulo_add_11_qelse_or_nl
        , modulo_add_11_qelse_and_5_nl , modulo_add_11_qelse_and_6_nl , modulo_add_11_qelse_and_7_nl});
    modulo_add_12_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_70, (readslicef_33_32_1(acc_14_nl)),
        z_out_82, z_out_80, {modulo_add_12_qelse_and_nl , modulo_add_12_qelse_or_1_nl
        , modulo_add_12_qelse_and_4_nl , modulo_add_12_qelse_and_5_nl});
    modulo_add_13_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_69, (readslicef_33_32_1(acc_18_nl)),
        z_out_81, z_out_79, {modulo_add_13_qelse_and_nl , modulo_add_13_qelse_or_1_nl
        , modulo_add_13_qelse_and_4_nl , modulo_add_13_qelse_and_5_nl});
    modulo_add_14_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_68, (readslicef_33_32_1(acc_22_nl)),
        z_out_80, z_out_78, {modulo_add_14_qelse_and_nl , modulo_add_14_qelse_or_1_nl
        , modulo_add_14_qelse_and_4_nl , modulo_add_14_qelse_and_5_nl});
    modulo_add_15_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_67, (readslicef_33_32_1(acc_26_nl)),
        z_out_82, z_out_79, z_out_77, {modulo_add_15_qelse_and_nl , modulo_add_15_qelse_or_nl
        , modulo_add_15_qelse_and_5_nl , modulo_add_15_qelse_and_6_nl , modulo_add_15_qelse_and_7_nl});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    mult_15_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_15_z_asn_itm_2, mult_31_z_asn_itm_2,
        mult_14_z_asn_itm_2, mult_27_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_14_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_14_z_asn_itm_2, mult_30_z_asn_itm_2,
        mult_26_z_asn_itm_2, mult_15_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_13_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_13_z_asn_itm_2, mult_29_z_asn_itm_2,
        mult_28_z_asn_itm_2, {or_dcpl_210 , (fsm_output[4]) , (fsm_output[9])});
    mult_12_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_12_z_asn_itm_2, mult_28_z_asn_itm_2,
        mult_29_z_asn_itm_2, {or_tmp_1189 , (fsm_output[4]) , (fsm_output[7])});
    mult_11_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_11_z_asn_itm_2, mult_27_z_asn_itm_2,
        mult_15_z_asn_itm_2, mult_26_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_10_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_10_z_asn_itm_2, mult_26_z_asn_itm_2,
        mult_25_z_asn_itm_2, mult_1_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_8 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_7 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    mult_15_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_2_z, mult_z_mul_cmp_22_z,
        mult_z_mul_cmp_20_z, {(fsm_output[2]) , or_dcpl_217 , (fsm_output[9])});
    mult_14_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_4_z, mult_z_mul_cmp_24_z,
        mult_z_mul_cmp_28_z, {or_tmp_1189 , (fsm_output[4]) , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_7 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    mult_13_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_6_z, mult_z_mul_cmp_26_z,
        mult_z_mul_cmp_24_z, mult_z_mul_cmp_12_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_6 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    mult_12_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_8_z, mult_z_mul_cmp_28_z,
        mult_z_mul_cmp_12_z, {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    mult_11_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_10_z, mult_z_mul_cmp_30_z,
        mult_z_mul_cmp_8_z, mult_z_mul_cmp_16_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_10_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_12_z, mult_z_mul_cmp_z,
        mult_z_mul_cmp_2_z, {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    mult_1_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_30_z, mult_z_mul_cmp_20_z,
        mult_z_mul_cmp_16_z, mult_z_mul_cmp_26_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_6 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_5 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_5 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_4 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_4 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_3 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_2 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_3 <= MUX1HOT_v_6_3_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {or_dcpl_210
        , (fsm_output[4]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_2 <= MUX1HOT_v_6_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1,
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP3_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_1 <= MUX1HOT_v_6_4_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), (INNER_LOOP3_r_11_4_sva_6_0[6:1]), (INNER_LOOP4_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_9, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_2 <= MUX_v_6_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1,
        (INNER_LOOP3_r_11_4_sva_6_0[6:1]), fsm_output[7]);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_1 <= MUX1HOT_v_6_3_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse, (INNER_LOOP3_r_11_4_sva_6_0[6:1]),
        {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse, or_dcpl_218);
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_1 <= MUX1HOT_v_6_4_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        (INNER_LOOP2_r_11_4_sva_6_0[6:1]), INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8,
        (INNER_LOOP4_r_11_4_sva_6_0[6:1]), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
        , (fsm_output[9])});
    INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_1 <= MUX_v_6_2_2((INNER_LOOP1_r_11_4_sva_6_0[6:1]),
        INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_8, or_dcpl_218);
    mult_16_z_asn_itm_3 <= MUX_v_32_2_2(mult_31_z_asn_itm_2, mult_10_z_asn_itm_2,
        or_dcpl_217);
    mult_17_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_1_z_asn_itm_2, mult_11_z_asn_itm_2,
        mult_31_z_asn_itm_2, mult_10_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_18_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_23_z_asn_itm_2, mult_12_z_asn_itm_2,
        mult_24_z_asn_itm_2, {or_tmp_1189 , (fsm_output[4]) , (fsm_output[7])});
    mult_19_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_24_z_asn_itm_2, mult_13_z_asn_itm_2,
        mult_23_z_asn_itm_2, {or_tmp_1189 , (fsm_output[4]) , (fsm_output[7])});
    mult_20_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_25_z_asn_itm_2, mult_14_z_asn_itm_2,
        mult_28_z_asn_itm_2, mult_13_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_21_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_26_z_asn_itm_2, mult_15_z_asn_itm_2,
        mult_11_z_asn_itm_2, mult_30_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_22_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_27_z_asn_itm_2, mult_1_z_asn_itm_2,
        mult_14_z_asn_itm_2, {or_dcpl_210 , (fsm_output[4]) , (fsm_output[9])});
    mult_23_z_asn_itm_3 <= MUX1HOT_v_32_4_2(mult_28_z_asn_itm_2, mult_23_z_asn_itm_2,
        mult_1_z_asn_itm_2, mult_25_z_asn_itm_2, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_24_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_29_z_asn_itm_2, mult_24_z_asn_itm_2,
        mult_12_z_asn_itm_2, {or_tmp_1189 , (fsm_output[4]) , (fsm_output[7])});
    mult_25_z_asn_itm_3 <= MUX1HOT_v_32_3_2(mult_30_z_asn_itm_2, mult_25_z_asn_itm_2,
        mult_11_z_asn_itm_2, {or_dcpl_210 , (fsm_output[4]) , (fsm_output[9])});
    modulo_add_23_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_80, (readslicef_33_32_1(acc_29_nl)),
        z_out_77, z_out_75, {modulo_add_23_qelse_and_nl , modulo_add_23_qelse_or_1_nl
        , modulo_add_23_qelse_and_4_nl , modulo_add_23_qelse_and_5_nl});
    modulo_add_24_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_79, (readslicef_33_32_1(acc_32_nl)),
        z_out_76, z_out_74, {modulo_add_24_qelse_and_nl , modulo_add_24_qelse_or_1_nl
        , modulo_add_24_qelse_and_4_nl , modulo_add_24_qelse_and_5_nl});
    modulo_add_25_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_4_2(z_out_78, (readslicef_33_32_1(acc_34_nl)),
        z_out_75, z_out_73, {modulo_add_25_qelse_and_nl , modulo_add_25_qelse_or_1_nl
        , modulo_add_25_qelse_and_4_nl , modulo_add_25_qelse_and_5_nl});
    modulo_add_26_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_77, (readslicef_33_32_1(acc_37_nl)),
        z_out_76, z_out_74, z_out_72, {modulo_add_26_qelse_and_nl , modulo_add_26_qelse_or_nl
        , modulo_add_26_qelse_and_5_nl , modulo_add_26_qelse_and_6_nl , modulo_add_26_qelse_and_7_nl});
    modulo_add_27_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_76, (readslicef_33_32_1(acc_39_nl)),
        z_out_75, z_out_73, z_out_71, {modulo_add_27_qelse_and_nl , modulo_add_27_qelse_or_nl
        , modulo_add_27_qelse_and_5_nl , modulo_add_27_qelse_and_6_nl , modulo_add_27_qelse_and_7_nl});
    modulo_add_28_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_75, (readslicef_33_32_1(acc_42_nl)),
        z_out_74, z_out_72, z_out_70, {modulo_add_28_qelse_and_nl , modulo_add_28_qelse_or_nl
        , modulo_add_28_qelse_and_5_nl , modulo_add_28_qelse_and_6_nl , modulo_add_28_qelse_and_7_nl});
    modulo_add_29_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_74, (readslicef_33_32_1(acc_44_nl)),
        z_out_73, z_out_71, z_out_69, {modulo_add_29_qelse_and_nl , modulo_add_29_qelse_or_nl
        , modulo_add_29_qelse_and_5_nl , modulo_add_29_qelse_and_6_nl , modulo_add_29_qelse_and_7_nl});
    modulo_add_30_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_73, (readslicef_33_32_1(acc_47_nl)),
        z_out_72, z_out_70, z_out_68, {modulo_add_30_qelse_and_nl , modulo_add_30_qelse_or_nl
        , modulo_add_30_qelse_and_5_nl , modulo_add_30_qelse_and_6_nl , modulo_add_30_qelse_and_7_nl});
    modulo_add_31_qr_lpi_3_dfm_1 <= MUX1HOT_v_32_5_2(z_out_82, (readslicef_33_32_1(acc_49_nl)),
        z_out_71, z_out_69, z_out_67, {modulo_add_31_qelse_and_nl , modulo_add_31_qelse_or_nl
        , modulo_add_31_qelse_and_5_nl , modulo_add_31_qelse_and_6_nl , modulo_add_31_qelse_and_7_nl});
    mult_23_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_28_z, mult_z_mul_cmp_18_z,
        mult_z_mul_cmp_6_z, mult_z_mul_cmp_10_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_24_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_26_z, mult_z_mul_cmp_16_z,
        mult_z_mul_cmp_10_z, mult_z_mul_cmp_2_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_25_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_24_z, mult_z_mul_cmp_14_z,
        mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_26_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_22_z, mult_z_mul_cmp_12_z,
        mult_z_mul_cmp_26_z, mult_z_mul_cmp_18_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_27_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_20_z, mult_z_mul_cmp_10_z,
        mult_z_mul_cmp_30_z, mult_z_mul_cmp_24_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_28_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_18_z, mult_z_mul_cmp_8_z,
        mult_z_mul_cmp_20_z, mult_z_mul_cmp_30_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_29_z_asn_itm_1 <= MUX1HOT_v_32_4_2(mult_z_mul_cmp_16_z, mult_z_mul_cmp_6_z,
        mult_z_mul_cmp_14_z, mult_z_mul_cmp_22_z, {(fsm_output[2]) , (fsm_output[4])
        , (fsm_output[7]) , (fsm_output[9])});
    mult_30_z_asn_itm_1 <= MUX_v_32_2_2(mult_z_mul_cmp_14_z, mult_z_mul_cmp_4_z,
        or_dcpl_217);
    mult_31_z_asn_itm_1 <= MUX1HOT_v_32_3_2(mult_z_mul_cmp_z, mult_z_mul_cmp_2_z,
        mult_z_mul_cmp_6_z, {or_dcpl_210 , (fsm_output[4]) , (fsm_output[9])});
    tmp_10_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_0_i_qa_d[31:0]), (yt_rsc_0_10_i_qa_d[31:0]),
        (xt_rsc_0_4_i_qa_d[31:0]), (yt_rsc_0_0_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_102_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_2_i_qa_d[31:0]), (yt_rsc_0_12_i_qa_d[31:0]),
        (xt_rsc_0_6_i_qa_d[31:0]), (yt_rsc_0_2_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_104_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_4_i_qa_d[31:0]), (yt_rsc_0_14_i_qa_d[31:0]),
        (xt_rsc_0_8_i_qa_d[31:0]), (yt_rsc_0_4_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_106_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_6_i_qa_d[31:0]), (yt_rsc_0_16_i_qa_d[31:0]),
        (xt_rsc_0_10_i_qa_d[31:0]), (yt_rsc_0_6_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_108_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_8_i_qa_d[31:0]), (yt_rsc_0_18_i_qa_d[31:0]),
        (xt_rsc_0_12_i_qa_d[31:0]), (yt_rsc_0_8_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_110_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_10_i_qa_d[31:0]), (yt_rsc_0_2_i_qa_d[31:0]),
        (xt_rsc_0_14_i_qa_d[31:0]), (yt_rsc_0_10_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_112_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_12_i_qa_d[31:0]), (yt_rsc_0_20_i_qa_d[31:0]),
        (xt_rsc_0_16_i_qa_d[31:0]), (yt_rsc_0_12_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_114_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_14_i_qa_d[31:0]), (yt_rsc_0_22_i_qa_d[31:0]),
        (xt_rsc_0_18_i_qa_d[31:0]), (yt_rsc_0_14_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_116_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_16_i_qa_d[31:0]), (yt_rsc_0_24_i_qa_d[31:0]),
        (xt_rsc_0_20_i_qa_d[31:0]), (yt_rsc_0_16_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_118_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_18_i_qa_d[31:0]), (yt_rsc_0_26_i_qa_d[31:0]),
        (xt_rsc_0_22_i_qa_d[31:0]), (yt_rsc_0_18_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_120_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_20_i_qa_d[31:0]), (yt_rsc_0_28_i_qa_d[31:0]),
        (xt_rsc_0_24_i_qa_d[31:0]), (yt_rsc_0_20_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_122_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_22_i_qa_d[31:0]), (yt_rsc_0_30_i_qa_d[31:0]),
        (xt_rsc_0_26_i_qa_d[31:0]), (yt_rsc_0_22_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_124_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_24_i_qa_d[31:0]), (yt_rsc_0_4_i_qa_d[31:0]),
        (xt_rsc_0_28_i_qa_d[31:0]), (yt_rsc_0_24_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_126_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_26_i_qa_d[31:0]), (yt_rsc_0_6_i_qa_d[31:0]),
        (xt_rsc_0_30_i_qa_d[31:0]), (yt_rsc_0_26_i_qa_d[31:0]), {(fsm_output[2])
        , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_60_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_28_i_qa_d[31:0]), (yt_rsc_0_8_i_qa_d[31:0]),
        (xt_rsc_0_0_i_qa_d[31:0]), (yt_rsc_0_28_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    tmp_62_sva_1 <= MUX1HOT_v_32_4_2((xt_rsc_0_30_i_qa_d[31:0]), (yt_rsc_0_0_i_qa_d[31:0]),
        (xt_rsc_0_2_i_qa_d[31:0]), (yt_rsc_0_30_i_qa_d[31:0]), {(fsm_output[2]) ,
        (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
    reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd <= (z_out_49[31]) & (~(modulo_sub_16_qelse_and_ssc
        | modulo_sub_16_qelse_and_ssc_1));
    reg_modulo_sub_16_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_66[30:0]),
        (z_out_49[30:0]), (z_out_51[30:0]), {modulo_sub_16_qelse_and_ssc , modulo_sub_16_qelse_or_nl
        , modulo_sub_16_qelse_and_ssc_1});
    reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd <= (z_out_47[31]) & (~(modulo_sub_17_qelse_and_ssc
        | modulo_sub_17_qelse_and_ssc_1));
    reg_modulo_sub_17_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_56[30:0]),
        (z_out_47[30:0]), (z_out_52[30:0]), {modulo_sub_17_qelse_and_ssc , modulo_sub_17_qelse_or_nl
        , modulo_sub_17_qelse_and_ssc_1});
    reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd <= (z_out_46[31]) & (~(modulo_sub_18_qelse_and_ssc
        | modulo_sub_18_qelse_and_ssc_1));
    reg_modulo_sub_18_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_63[30:0]),
        (z_out_46[30:0]), (z_out_53[30:0]), {modulo_sub_18_qelse_and_ssc , modulo_sub_18_qelse_or_nl
        , modulo_sub_18_qelse_and_ssc_1});
    reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd <= (z_out_44[31]) & (~(modulo_sub_19_qelse_and_ssc
        | modulo_sub_19_qelse_and_ssc_1));
    reg_modulo_sub_19_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_64[30:0]),
        (z_out_44[30:0]), (z_out_54[30:0]), {modulo_sub_19_qelse_and_ssc , modulo_sub_19_qelse_or_nl
        , modulo_sub_19_qelse_and_ssc_1});
    reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd <= (z_out_42[31]) & (~(modulo_sub_20_qelse_and_ssc
        | modulo_sub_20_qelse_and_ssc_1));
    reg_modulo_sub_20_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_65[30:0]),
        (z_out_42[30:0]), (z_out_55[30:0]), {modulo_sub_20_qelse_and_ssc , modulo_sub_20_qelse_or_nl
        , modulo_sub_20_qelse_and_ssc_1});
    reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd <= (z_out_41[31]) & (~(modulo_sub_21_qelse_and_ssc
        | modulo_sub_21_qelse_and_ssc_1));
    reg_modulo_sub_21_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_51[30:0]),
        (z_out_41[30:0]), (z_out_56[30:0]), {modulo_sub_21_qelse_and_ssc , modulo_sub_21_qelse_or_nl
        , modulo_sub_21_qelse_and_ssc_1});
    reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd <= (z_out_39[31]) & (~(modulo_sub_22_qelse_and_ssc
        | modulo_sub_22_qelse_and_ssc_1));
    reg_modulo_sub_22_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_52[30:0]),
        (z_out_39[30:0]), (z_out_57[30:0]), {modulo_sub_22_qelse_and_ssc , modulo_sub_22_qelse_or_nl
        , modulo_sub_22_qelse_and_ssc_1});
    reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd <= (z_out_37[31]) & (~(modulo_sub_23_qelse_and_ssc
        | modulo_sub_23_qelse_and_ssc_1));
    reg_modulo_sub_23_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_53[30:0]),
        (z_out_37[30:0]), (z_out_58[30:0]), {modulo_sub_23_qelse_and_ssc , modulo_sub_23_qelse_or_nl
        , modulo_sub_23_qelse_and_ssc_1});
    reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd <= (z_out_36[31]) & (~(modulo_sub_24_qelse_and_ssc
        | modulo_sub_24_qelse_and_ssc_1));
    reg_modulo_sub_24_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_54[30:0]),
        (z_out_36[30:0]), (z_out_59[30:0]), {modulo_sub_24_qelse_and_ssc , modulo_sub_24_qelse_or_nl
        , modulo_sub_24_qelse_and_ssc_1});
    reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd <= (z_out_34[31]) & (~(modulo_sub_25_qelse_and_ssc
        | modulo_sub_25_qelse_and_ssc_1));
    reg_modulo_sub_25_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_55[30:0]),
        (z_out_34[30:0]), (z_out_60[30:0]), {modulo_sub_25_qelse_and_ssc , modulo_sub_25_qelse_or_nl
        , modulo_sub_25_qelse_and_ssc_1});
    reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd <= (z_out_32[31]) & (~(modulo_sub_26_qelse_and_ssc
        | modulo_sub_26_qelse_and_ssc_1));
    reg_modulo_sub_26_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_57[30:0]),
        (z_out_32[30:0]), (z_out_61[30:0]), {modulo_sub_26_qelse_and_ssc , modulo_sub_26_qelse_or_nl
        , modulo_sub_26_qelse_and_ssc_1});
    reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd <= (z_out_31[31]) & (~(modulo_sub_27_qelse_and_ssc
        | modulo_sub_27_qelse_and_ssc_1));
    reg_modulo_sub_27_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_58[30:0]),
        (z_out_31[30:0]), (z_out_62[30:0]), {modulo_sub_27_qelse_and_ssc , modulo_sub_27_qelse_or_nl
        , modulo_sub_27_qelse_and_ssc_1});
    reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd <= (z_out_29[31]) & (~(modulo_sub_28_qelse_and_ssc
        | modulo_sub_28_qelse_and_ssc_1));
    reg_modulo_sub_28_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_59[30:0]),
        (z_out_29[30:0]), (z_out_63[30:0]), {modulo_sub_28_qelse_and_ssc , modulo_sub_28_qelse_or_nl
        , modulo_sub_28_qelse_and_ssc_1});
    reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd <= (z_out_26[31]) & (~(modulo_sub_29_qelse_and_ssc
        | modulo_sub_29_qelse_and_ssc_1));
    reg_modulo_sub_29_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_60[30:0]),
        (z_out_26[30:0]), (z_out_64[30:0]), {modulo_sub_29_qelse_and_ssc , modulo_sub_29_qelse_or_nl
        , modulo_sub_29_qelse_and_ssc_1});
    reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd <= (z_out_24[31]) & (~(modulo_sub_30_qelse_and_ssc
        | modulo_sub_30_qelse_and_ssc_1));
    reg_modulo_sub_30_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_61[30:0]),
        (z_out_24[30:0]), (z_out_65[30:0]), {modulo_sub_30_qelse_and_ssc , modulo_sub_30_qelse_or_nl
        , modulo_sub_30_qelse_and_ssc_1});
    reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd <= (z_out_21[31]) & (~(modulo_sub_31_qelse_and_ssc
        | modulo_sub_31_qelse_and_ssc_1));
    reg_modulo_sub_31_qr_lpi_3_dfm_1_ftd_1 <= MUX1HOT_v_31_3_2((z_out_62[30:0]),
        (z_out_21[30:0]), (z_out_66[30:0]), {modulo_sub_31_qelse_and_ssc , modulo_sub_31_qelse_or_nl
        , modulo_sub_31_qelse_and_ssc_1});
    INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_3 <= reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse;
    INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_1 <= MUX_v_6_2_2((INNER_LOOP2_r_11_4_sva_6_0[6:1]),
        (INNER_LOOP4_r_11_4_sva_6_0[6:1]), fsm_output[9]);
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_114_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_161_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_224_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_287_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_350_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_413_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_9 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_12_cse ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_602_itm_9_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_129_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_192_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_255_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_318_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_381_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_570_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_7;
      tmp_10_sva_7 <= tmp_10_sva_6;
      tmp_102_sva_7 <= tmp_102_sva_6;
      tmp_104_sva_7 <= tmp_104_sva_6;
      tmp_106_sva_7 <= tmp_106_sva_6;
      tmp_108_sva_7 <= tmp_108_sva_6;
      tmp_110_sva_7 <= tmp_110_sva_6;
      tmp_112_sva_7 <= tmp_112_sva_6;
      tmp_114_sva_7 <= tmp_114_sva_6;
      tmp_116_sva_7 <= tmp_116_sva_6;
      tmp_118_sva_7 <= tmp_118_sva_6;
      tmp_120_sva_7 <= tmp_120_sva_6;
      tmp_122_sva_7 <= tmp_122_sva_6;
      tmp_124_sva_7 <= tmp_124_sva_6;
      tmp_126_sva_7 <= tmp_126_sva_6;
      tmp_60_sva_7 <= tmp_60_sva_6;
      tmp_62_sva_7 <= tmp_62_sva_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_13 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      reg_INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_633_itm_8_cse <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_stage_0_8 ) begin
      mult_15_res_lpi_3_dfm_1 <= mult_15_res_lpi_3_dfm_1_mx0;
      mult_14_res_lpi_3_dfm_1 <= mult_14_res_lpi_3_dfm_1_mx0;
      mult_13_res_lpi_3_dfm_1 <= mult_13_res_lpi_3_dfm_1_mx0;
      mult_12_res_lpi_3_dfm_1 <= mult_12_res_lpi_3_dfm_1_mx0;
      mult_11_res_lpi_3_dfm_1 <= mult_11_res_lpi_3_dfm_1_mx0;
      mult_10_res_lpi_3_dfm_1 <= mult_10_res_lpi_3_dfm_1_mx0;
      mult_9_res_lpi_3_dfm_1 <= mult_9_res_lpi_3_dfm_1_mx0;
      mult_8_res_lpi_3_dfm_1 <= mult_8_res_lpi_3_dfm_1_mx0;
      mult_7_res_lpi_3_dfm_1 <= mult_7_res_lpi_3_dfm_1_mx0;
      mult_6_res_lpi_3_dfm_1 <= mult_6_res_lpi_3_dfm_1_mx0;
      mult_5_res_lpi_3_dfm_1 <= mult_5_res_lpi_3_dfm_1_mx0;
      mult_4_res_lpi_3_dfm_1 <= mult_4_res_lpi_3_dfm_1_mx0;
      mult_3_res_lpi_3_dfm_1 <= mult_3_res_lpi_3_dfm_1_mx0;
      mult_2_res_lpi_3_dfm_1 <= mult_2_res_lpi_3_dfm_1_mx0;
      mult_1_res_lpi_3_dfm_1 <= mult_1_res_lpi_3_dfm_1_mx0;
      mult_res_lpi_3_dfm_1 <= mult_res_lpi_3_dfm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_20_false_acc_cse_sva <= 3'b000;
    end
    else if ( ~(or_dcpl_233 | or_dcpl_210) ) begin
      operator_20_false_acc_cse_sva <= MUX_v_3_2_2(z_out_1, (z_out[2:0]), fsm_output[6]);
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 ) begin
      mult_15_z_asn_itm_2 <= mult_15_z_asn_itm_1;
      mult_14_z_asn_itm_2 <= mult_14_z_asn_itm_1;
      mult_13_z_asn_itm_2 <= mult_13_z_asn_itm_1;
      mult_12_z_asn_itm_2 <= mult_12_z_asn_itm_1;
      mult_11_z_asn_itm_2 <= mult_11_z_asn_itm_1;
      mult_10_z_asn_itm_2 <= mult_10_z_asn_itm_1;
      mult_1_z_asn_itm_2 <= mult_1_z_asn_itm_1;
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_5;
      mult_23_z_asn_itm_2 <= mult_23_z_asn_itm_1;
      mult_24_z_asn_itm_2 <= mult_24_z_asn_itm_1;
      mult_25_z_asn_itm_2 <= mult_25_z_asn_itm_1;
      mult_26_z_asn_itm_2 <= mult_26_z_asn_itm_1;
      mult_27_z_asn_itm_2 <= mult_27_z_asn_itm_1;
      mult_28_z_asn_itm_2 <= mult_28_z_asn_itm_1;
      mult_29_z_asn_itm_2 <= mult_29_z_asn_itm_1;
      mult_30_z_asn_itm_2 <= mult_30_z_asn_itm_1;
      mult_31_z_asn_itm_2 <= mult_31_z_asn_itm_1;
      tmp_10_sva_5 <= tmp_10_sva_4;
      tmp_102_sva_5 <= tmp_102_sva_4;
      tmp_104_sva_5 <= tmp_104_sva_4;
      tmp_106_sva_5 <= tmp_106_sva_4;
      tmp_108_sva_5 <= tmp_108_sva_4;
      tmp_110_sva_5 <= tmp_110_sva_4;
      tmp_112_sva_5 <= tmp_112_sva_4;
      tmp_114_sva_5 <= tmp_114_sva_4;
      tmp_116_sva_5 <= tmp_116_sva_4;
      tmp_118_sva_5 <= tmp_118_sva_4;
      tmp_120_sva_5 <= tmp_120_sva_4;
      tmp_122_sva_5 <= tmp_122_sva_4;
      tmp_124_sva_5 <= tmp_124_sva_4;
      tmp_126_sva_5 <= tmp_126_sva_4;
      tmp_60_sva_5 <= tmp_60_sva_4;
      tmp_62_sva_5 <= tmp_62_sva_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_6;
      tmp_10_sva_6 <= tmp_10_sva_5;
      tmp_102_sva_6 <= tmp_102_sva_5;
      tmp_104_sva_6 <= tmp_104_sva_5;
      tmp_106_sva_6 <= tmp_106_sva_5;
      tmp_108_sva_6 <= tmp_108_sva_5;
      tmp_110_sva_6 <= tmp_110_sva_5;
      tmp_112_sva_6 <= tmp_112_sva_5;
      tmp_114_sva_6 <= tmp_114_sva_5;
      tmp_116_sva_6 <= tmp_116_sva_5;
      tmp_118_sva_6 <= tmp_118_sva_5;
      tmp_120_sva_6 <= tmp_120_sva_5;
      tmp_122_sva_6 <= tmp_122_sva_5;
      tmp_124_sva_6 <= tmp_124_sva_5;
      tmp_126_sva_6 <= tmp_126_sva_5;
      tmp_60_sva_6 <= tmp_60_sva_5;
      tmp_62_sva_6 <= tmp_62_sva_5;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_44_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_22 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_64_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_45 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_4;
      tmp_10_sva_4 <= tmp_10_sva_3;
      tmp_102_sva_4 <= tmp_102_sva_3;
      tmp_104_sva_4 <= tmp_104_sva_3;
      tmp_106_sva_4 <= tmp_106_sva_3;
      tmp_108_sva_4 <= tmp_108_sva_3;
      tmp_110_sva_4 <= tmp_110_sva_3;
      tmp_112_sva_4 <= tmp_112_sva_3;
      tmp_114_sva_4 <= tmp_114_sva_3;
      tmp_116_sva_4 <= tmp_116_sva_3;
      tmp_118_sva_4 <= tmp_118_sva_3;
      tmp_120_sva_4 <= tmp_120_sva_3;
      tmp_122_sva_4 <= tmp_122_sva_3;
      tmp_124_sva_4 <= tmp_124_sva_3;
      tmp_126_sva_4 <= tmp_126_sva_3;
      tmp_60_sva_4 <= tmp_60_sva_3;
      tmp_62_sva_4 <= tmp_62_sva_3;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_84_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_65 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_3;
      tmp_10_sva_3 <= tmp_10_sva_2;
      tmp_102_sva_3 <= tmp_102_sva_2;
      tmp_104_sva_3 <= tmp_104_sva_2;
      tmp_106_sva_3 <= tmp_106_sva_2;
      tmp_108_sva_3 <= tmp_108_sva_2;
      tmp_110_sva_3 <= tmp_110_sva_2;
      tmp_112_sva_3 <= tmp_112_sva_2;
      tmp_114_sva_3 <= tmp_114_sva_2;
      tmp_116_sva_3 <= tmp_116_sva_2;
      tmp_118_sva_3 <= tmp_118_sva_2;
      tmp_120_sva_3 <= tmp_120_sva_2;
      tmp_122_sva_3 <= tmp_122_sva_2;
      tmp_124_sva_3 <= tmp_124_sva_2;
      tmp_126_sva_3 <= tmp_126_sva_2;
      tmp_60_sva_3 <= tmp_60_sva_2;
      tmp_62_sva_3 <= tmp_62_sva_2;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_103_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_101 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1074_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_2;
      tmp_10_sva_2 <= tmp_10_sva_1;
      tmp_102_sva_2 <= tmp_102_sva_1;
      tmp_104_sva_2 <= tmp_104_sva_1;
      tmp_106_sva_2 <= tmp_106_sva_1;
      tmp_108_sva_2 <= tmp_108_sva_1;
      tmp_110_sva_2 <= tmp_110_sva_1;
      tmp_112_sva_2 <= tmp_112_sva_1;
      tmp_114_sva_2 <= tmp_114_sva_1;
      tmp_116_sva_2 <= tmp_116_sva_1;
      tmp_118_sva_2 <= tmp_118_sva_1;
      tmp_120_sva_2 <= tmp_120_sva_1;
      tmp_122_sva_2 <= tmp_122_sva_1;
      tmp_124_sva_2 <= tmp_124_sva_1;
      tmp_126_sva_2 <= tmp_126_sva_1;
      tmp_60_sva_2 <= tmp_60_sva_1;
      tmp_62_sva_2 <= tmp_62_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_665_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_123_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( or_dcpl_121 | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1043_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_1011_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_980_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_948_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_917_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_885_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_854_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_822_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_791_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_759_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_728_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_696_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_539_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_507_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( or_142_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_476_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( or_143_cse | INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_444_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      INNER_LOOP2_r_11_4_sva_6_0 <= 7'b0000000;
    end
    else if ( ~ (fsm_output[2]) ) begin
      INNER_LOOP2_r_11_4_sva_6_0 <= MUX_v_7_2_2(7'b0000000, STAGE_LOOP_base_STAGE_LOOP_base_mux_nl,
          INNER_LOOP2_r_or_nl);
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_8;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_8;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_6 ) begin
      reg_mult_31_res_lpi_3_dfm_1_cse <= mult_15_res_lpi_3_dfm_1_mx0;
      reg_mult_30_res_lpi_3_dfm_1_cse <= mult_14_res_lpi_3_dfm_1_mx0;
      reg_mult_29_res_lpi_3_dfm_1_cse <= mult_13_res_lpi_3_dfm_1_mx0;
      reg_mult_28_res_lpi_3_dfm_1_cse <= mult_12_res_lpi_3_dfm_1_mx0;
      reg_mult_27_res_lpi_3_dfm_1_cse <= mult_11_res_lpi_3_dfm_1_mx0;
      reg_mult_26_res_lpi_3_dfm_1_cse <= mult_10_res_lpi_3_dfm_1_mx0;
      reg_mult_25_res_lpi_3_dfm_1_cse <= mult_9_res_lpi_3_dfm_1_mx0;
      reg_mult_24_res_lpi_3_dfm_1_cse <= mult_8_res_lpi_3_dfm_1_mx0;
      reg_mult_23_res_lpi_3_dfm_1_cse <= mult_7_res_lpi_3_dfm_1_mx0;
      reg_mult_22_res_lpi_3_dfm_1_cse <= mult_6_res_lpi_3_dfm_1_mx0;
      reg_mult_21_res_lpi_3_dfm_1_cse <= mult_5_res_lpi_3_dfm_1_mx0;
      reg_mult_20_res_lpi_3_dfm_1_cse <= mult_4_res_lpi_3_dfm_1_mx0;
      reg_mult_19_res_lpi_3_dfm_1_cse <= mult_3_res_lpi_3_dfm_1_mx0;
      reg_mult_18_res_lpi_3_dfm_1_cse <= mult_2_res_lpi_3_dfm_1_mx0;
      reg_mult_17_res_lpi_3_dfm_1_cse <= mult_1_res_lpi_3_dfm_1_mx0;
      reg_mult_16_res_lpi_3_dfm_1_cse <= mult_res_lpi_3_dfm_1_mx0;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_7;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_7;
    end
  end
  always @(posedge clk) begin
    if ( ~ (fsm_output[4]) ) begin
      operator_33_true_1_lshift_psp_9_4_sva <= z_out[9:4];
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_5 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_6;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_6;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_4 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_5;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_5;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_3 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_4;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_4;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_2 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_3;
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_948_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_1 ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm ) begin
      INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_11_4_6_0_980_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      butterFly2_15_tw_equal_tmp_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_3_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_5_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_6_1 <= 1'b0;
      butterFly2_15_tw_equal_tmp_7_1 <= 1'b0;
    end
    else if ( INNER_LOOP1_stage_0 ) begin
      butterFly2_15_tw_equal_tmp_1 <= ~((operator_20_false_acc_cse_sva!=3'b000));
      butterFly2_15_tw_equal_tmp_3_1 <= (operator_20_false_acc_cse_sva==3'b011);
      butterFly2_15_tw_equal_tmp_5_1 <= (operator_20_false_acc_cse_sva==3'b101);
      butterFly2_15_tw_equal_tmp_6_1 <= (operator_20_false_acc_cse_sva==3'b110);
      butterFly2_15_tw_equal_tmp_7_1 <= (operator_20_false_acc_cse_sva==3'b111);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_33_true_3_lshift_psp_1_0_sva <= 2'b00;
    end
    else if ( ~ (fsm_output[9]) ) begin
      operator_33_true_3_lshift_psp_1_0_sva <= operator_33_true_3_lshift_psp_1_0_sva_mx0w3;
    end
  end
  assign butterFly2_21_tw_butterFly2_21_tw_or_nl = c_1_sva | INNER_LOOP4_nor_tmp;
  assign c_mux_nl = MUX_s_1_2_2((operator_20_false_acc_cse_sva[0]), butterFly2_21_tw_butterFly2_21_tw_or_nl,
      fsm_output[9]);
  assign STAGE_LOOP_and_nl = (~ (fsm_output[7])) & or_tmp_1134;
  assign STAGE_LOOP_mux1h_nl = MUX1HOT_v_2_5_2((operator_20_false_acc_cse_sva[2:1]),
      (z_out[1:0]), (operator_20_false_acc_cse_sva[1:0]), operator_33_true_3_lshift_psp_1_0_sva_mx0w3,
      operator_33_true_3_lshift_psp_1_0_sva, {(fsm_output[5]) , STAGE_LOOP_and_nl
      , (fsm_output[7]) , (fsm_output[8]) , (fsm_output[9])});
  assign nor_4_nl = ~((fsm_output[8]) | (fsm_output[5]) | (fsm_output[6]) | (~ and_dcpl_90));
  assign INNER_LOOP1_r_mux_44_nl = MUX_s_1_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7, or_dcpl_218);
  assign modulo_add_1_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_81, z_out_78, z_out_76,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_2_nl = ({modulo_add_1_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_2_nl = nl_acc_2_nl[32:0];
  assign modulo_add_1_qelse_and_nl = (~ z_out_83_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_1_qelse_or_1_nl = (z_out_83_32 & modulo_add_1_qelse_or_m1c) |
      (z_out_83_32 & (fsm_output[7])) | (z_out_85_32 & (fsm_output[9]));
  assign modulo_add_1_qelse_and_4_nl = (~ z_out_83_32) & (fsm_output[7]);
  assign modulo_add_1_qelse_and_5_nl = (~ z_out_85_32) & (fsm_output[9]);
  assign modulo_add_10_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_72, z_out_67, z_out_68,
      z_out_82, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_6_nl = ({modulo_add_10_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[32:0];
  assign modulo_add_10_qelse_and_nl = (~ z_out_84_32) & (fsm_output[2]);
  assign modulo_add_10_qelse_or_nl = (z_out_84_32 & (fsm_output[2])) | (z_out_84_32
      & (fsm_output[4])) | (z_out_84_32 & (fsm_output[7])) | (z_out_86_32 & (fsm_output[9]));
  assign modulo_add_10_qelse_and_5_nl = (~ z_out_84_32) & (fsm_output[4]);
  assign modulo_add_10_qelse_and_6_nl = (~ z_out_84_32) & (fsm_output[7]);
  assign modulo_add_10_qelse_and_7_nl = (~ z_out_86_32) & (fsm_output[9]);
  assign modulo_add_11_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_71, z_out_77, z_out_67,
      z_out_81, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_10_nl = ({modulo_add_11_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[32:0];
  assign modulo_add_11_qelse_and_nl = (~ z_out_86_32) & (fsm_output[2]);
  assign modulo_add_11_qelse_or_nl = (z_out_86_32 & (fsm_output[2])) | (z_out_86_32
      & (fsm_output[4])) | (z_out_87_32 & (fsm_output[7])) | (z_out_87_32 & (fsm_output[9]));
  assign modulo_add_11_qelse_and_5_nl = (~ z_out_86_32) & (fsm_output[4]);
  assign modulo_add_11_qelse_and_6_nl = (~ z_out_87_32) & (fsm_output[7]);
  assign modulo_add_11_qelse_and_7_nl = (~ z_out_87_32) & (fsm_output[9]);
  assign modulo_add_12_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_70, z_out_82, z_out_80,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_14_nl = ({modulo_add_12_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[32:0];
  assign modulo_add_12_qelse_and_nl = (~ z_out_87_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_12_qelse_or_1_nl = (z_out_87_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_88_32 & (fsm_output[7])) | (z_out_90_32 & (fsm_output[9]));
  assign modulo_add_12_qelse_and_4_nl = (~ z_out_88_32) & (fsm_output[7]);
  assign modulo_add_12_qelse_and_5_nl = (~ z_out_90_32) & (fsm_output[9]);
  assign modulo_add_13_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_69, z_out_81, z_out_79,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_18_nl = ({modulo_add_13_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[32:0];
  assign modulo_add_13_qelse_and_nl = (~ z_out_90_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_13_qelse_or_1_nl = (z_out_90_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_90_32 & (fsm_output[7])) | (z_out_91_32 & (fsm_output[9]));
  assign modulo_add_13_qelse_and_4_nl = (~ z_out_90_32) & (fsm_output[7]);
  assign modulo_add_13_qelse_and_5_nl = (~ z_out_91_32) & (fsm_output[9]);
  assign modulo_add_14_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_68, z_out_80, z_out_78,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_22_nl = ({modulo_add_14_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[32:0];
  assign modulo_add_14_qelse_and_nl = (~ z_out_92_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_14_qelse_or_1_nl = (z_out_92_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_93_32 & (fsm_output[7])) | (z_out_94_32 & (fsm_output[9]));
  assign modulo_add_14_qelse_and_4_nl = (~ z_out_93_32) & (fsm_output[7]);
  assign modulo_add_14_qelse_and_5_nl = (~ z_out_94_32) & (fsm_output[9]);
  assign modulo_add_15_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_67, z_out_82, z_out_79,
      z_out_77, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_26_nl = ({modulo_add_15_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_26_nl = nl_acc_26_nl[32:0];
  assign modulo_add_15_qelse_and_nl = (~ z_out_93_32) & (fsm_output[2]);
  assign modulo_add_15_qelse_or_nl = (z_out_93_32 & (fsm_output[2])) | (z_out_93_32
      & (fsm_output[4])) | (z_out_94_32 & (fsm_output[7])) | (z_out_97_32 & (fsm_output[9]));
  assign modulo_add_15_qelse_and_5_nl = (~ z_out_93_32) & (fsm_output[4]);
  assign modulo_add_15_qelse_and_6_nl = (~ z_out_94_32) & (fsm_output[7]);
  assign modulo_add_15_qelse_and_7_nl = (~ z_out_97_32) & (fsm_output[9]);
  assign INNER_LOOP1_r_mux_45_nl = MUX_s_1_2_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_7,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_96_itm_10, fsm_output[7]);
  assign INNER_LOOP1_mux_nl = MUX_s_1_2_2(INNER_LOOP1_stage_0, INNER_LOOP1_stage_0_11,
      or_dcpl_218);
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_1_nl = (z_out_2[0]) & (fsm_output[4]);
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_3_nl = (z_out_2[0]) & (fsm_output[9]);
  assign or_1465_nl = (fsm_output[9:8]!=2'b00);
  assign INNER_LOOP1_r_mux1h_46_nl = MUX1HOT_s_1_4_2(INNER_LOOP1_stage_0_9, INNER_LOOP1_r_INNER_LOOP1_r_and_1_nl,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_11_4_6_0_97_itm_9, INNER_LOOP1_r_INNER_LOOP1_r_and_3_nl,
      {(fsm_output[2]) , or_dcpl_233 , (fsm_output[7]) , or_1465_nl});
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_2_nl = (z_out_2[0]) & (fsm_output[7]);
  assign INNER_LOOP1_mux_11_nl = MUX_s_1_2_2(INNER_LOOP1_stage_0_10, INNER_LOOP1_r_INNER_LOOP1_r_and_2_nl,
      or_tmp_1134);
  assign INNER_LOOP1_r_INNER_LOOP1_r_and_nl = (z_out_2[0]) & (fsm_output[2]);
  assign modulo_add_2_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_80, z_out_77, z_out_75,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_29_nl = ({modulo_add_2_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_29_nl = nl_acc_29_nl[32:0];
  assign modulo_add_23_qelse_and_nl = (~ z_out_96_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_23_qelse_or_1_nl = (z_out_96_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_96_32 & (fsm_output[7])) | (z_out_98_32 & (fsm_output[9]));
  assign modulo_add_23_qelse_and_4_nl = (~ z_out_96_32) & (fsm_output[7]);
  assign modulo_add_23_qelse_and_5_nl = (~ z_out_98_32) & (fsm_output[9]);
  assign modulo_add_3_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_79, z_out_76, z_out_74,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_32_nl = ({modulo_add_3_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_32_nl = nl_acc_32_nl[32:0];
  assign modulo_add_24_qelse_and_nl = (~ z_out_98_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_24_qelse_or_1_nl = (z_out_98_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_97_32 & (fsm_output[7])) | (z_out_96_32 & (fsm_output[9]));
  assign modulo_add_24_qelse_and_4_nl = (~ z_out_97_32) & (fsm_output[7]);
  assign modulo_add_24_qelse_and_5_nl = (~ z_out_96_32) & (fsm_output[9]);
  assign modulo_add_4_qif_mux1h_2_nl = MUX1HOT_v_32_3_2(z_out_78, z_out_75, z_out_73,
      {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_34_nl = ({modulo_add_4_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_34_nl = nl_acc_34_nl[32:0];
  assign modulo_add_25_qelse_and_nl = (~ z_out_97_32) & modulo_add_1_qelse_or_m1c;
  assign modulo_add_25_qelse_or_1_nl = (z_out_97_32 & modulo_add_1_qelse_or_m1c)
      | (z_out_95_32 & (fsm_output[7])) | (z_out_92_32 & (fsm_output[9]));
  assign modulo_add_25_qelse_and_4_nl = (~ z_out_95_32) & (fsm_output[7]);
  assign modulo_add_25_qelse_and_5_nl = (~ z_out_92_32) & (fsm_output[9]);
  assign modulo_add_5_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_77, z_out_76, z_out_74,
      z_out_72, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_37_nl = ({modulo_add_5_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_37_nl = nl_acc_37_nl[32:0];
  assign modulo_add_26_qelse_and_nl = (~ z_out_91_32) & (fsm_output[2]);
  assign modulo_add_26_qelse_or_nl = (z_out_91_32 & (fsm_output[2])) | (z_out_91_32
      & (fsm_output[4])) | (z_out_91_32 & (fsm_output[7])) | (z_out_88_32 & (fsm_output[9]));
  assign modulo_add_26_qelse_and_5_nl = (~ z_out_91_32) & (fsm_output[4]);
  assign modulo_add_26_qelse_and_6_nl = (~ z_out_91_32) & (fsm_output[7]);
  assign modulo_add_26_qelse_and_7_nl = (~ z_out_88_32) & (fsm_output[9]);
  assign modulo_add_6_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_76, z_out_75, z_out_73,
      z_out_71, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_39_nl = ({modulo_add_6_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_39_nl = nl_acc_39_nl[32:0];
  assign modulo_add_27_qelse_and_nl = (~ z_out_89_32) & (fsm_output[2]);
  assign modulo_add_27_qelse_or_nl = (z_out_89_32 & (fsm_output[2])) | (z_out_89_32
      & (fsm_output[4])) | (z_out_85_32 & (fsm_output[7])) | (z_out_84_32 & (fsm_output[9]));
  assign modulo_add_27_qelse_and_5_nl = (~ z_out_89_32) & (fsm_output[4]);
  assign modulo_add_27_qelse_and_6_nl = (~ z_out_85_32) & (fsm_output[7]);
  assign modulo_add_27_qelse_and_7_nl = (~ z_out_84_32) & (fsm_output[9]);
  assign modulo_add_7_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_75, z_out_74, z_out_72,
      z_out_70, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_42_nl = ({modulo_add_7_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_42_nl = nl_acc_42_nl[32:0];
  assign modulo_add_28_qelse_and_nl = (~ z_out_85_32) & (fsm_output[2]);
  assign modulo_add_28_qelse_or_nl = (z_out_85_32 & (fsm_output[2])) | (z_out_85_32
      & (fsm_output[4])) | (z_out_89_32 & (fsm_output[7])) | (z_out_93_32 & (fsm_output[9]));
  assign modulo_add_28_qelse_and_5_nl = (~ z_out_85_32) & (fsm_output[4]);
  assign modulo_add_28_qelse_and_6_nl = (~ z_out_89_32) & (fsm_output[7]);
  assign modulo_add_28_qelse_and_7_nl = (~ z_out_93_32) & (fsm_output[9]);
  assign modulo_add_8_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_74, z_out_73, z_out_71,
      z_out_69, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_44_nl = ({modulo_add_8_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_44_nl = nl_acc_44_nl[32:0];
  assign modulo_add_29_qelse_and_nl = (~ z_out_95_32) & (fsm_output[2]);
  assign modulo_add_29_qelse_or_nl = (z_out_95_32 & (fsm_output[2])) | (z_out_95_32
      & (fsm_output[4])) | (z_out_98_32 & (fsm_output[7])) | (z_out_95_32 & (fsm_output[9]));
  assign modulo_add_29_qelse_and_5_nl = (~ z_out_95_32) & (fsm_output[4]);
  assign modulo_add_29_qelse_and_6_nl = (~ z_out_98_32) & (fsm_output[7]);
  assign modulo_add_29_qelse_and_7_nl = (~ z_out_95_32) & (fsm_output[9]);
  assign modulo_add_9_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_73, z_out_72, z_out_70,
      z_out_68, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_47_nl = ({modulo_add_9_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_47_nl = nl_acc_47_nl[32:0];
  assign modulo_add_30_qelse_and_nl = (~ z_out_94_32) & (fsm_output[2]);
  assign modulo_add_30_qelse_or_nl = (z_out_94_32 & (fsm_output[2])) | (z_out_94_32
      & (fsm_output[4])) | (z_out_92_32 & (fsm_output[7])) | (z_out_89_32 & (fsm_output[9]));
  assign modulo_add_30_qelse_and_5_nl = (~ z_out_94_32) & (fsm_output[4]);
  assign modulo_add_30_qelse_and_6_nl = (~ z_out_92_32) & (fsm_output[7]);
  assign modulo_add_30_qelse_and_7_nl = (~ z_out_89_32) & (fsm_output[9]);
  assign modulo_add_qif_mux1h_2_nl = MUX1HOT_v_32_4_2(z_out_82, z_out_71, z_out_69,
      z_out_67, {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_49_nl = ({modulo_add_qif_mux1h_2_nl , 1'b1}) + ({(~ p_sva) , 1'b1});
  assign acc_49_nl = nl_acc_49_nl[32:0];
  assign modulo_add_31_qelse_and_nl = (~ z_out_88_32) & (fsm_output[2]);
  assign modulo_add_31_qelse_or_nl = (z_out_88_32 & (fsm_output[2])) | (z_out_88_32
      & (fsm_output[4])) | (z_out_86_32 & (fsm_output[7])) | (z_out_83_32 & (fsm_output[9]));
  assign modulo_add_31_qelse_and_5_nl = (~ z_out_88_32) & (fsm_output[4]);
  assign modulo_add_31_qelse_and_6_nl = (~ z_out_86_32) & (fsm_output[7]);
  assign modulo_add_31_qelse_and_7_nl = (~ z_out_83_32) & (fsm_output[9]);
  assign modulo_sub_16_qelse_or_nl = ((z_out_66[31]) & (~ (fsm_output[9]))) | ((z_out_51[31])
      & (fsm_output[9]));
  assign modulo_sub_17_qelse_or_nl = ((z_out_56[31]) & (~ (fsm_output[9]))) | ((z_out_52[31])
      & (fsm_output[9]));
  assign modulo_sub_18_qelse_or_nl = ((z_out_63[31]) & (~ (fsm_output[9]))) | ((z_out_53[31])
      & (fsm_output[9]));
  assign modulo_sub_19_qelse_or_nl = ((z_out_64[31]) & (~ (fsm_output[9]))) | ((z_out_54[31])
      & (fsm_output[9]));
  assign modulo_sub_20_qelse_or_nl = ((z_out_65[31]) & (~ (fsm_output[9]))) | ((z_out_55[31])
      & (fsm_output[9]));
  assign modulo_sub_21_qelse_or_nl = ((z_out_51[31]) & (~ (fsm_output[9]))) | ((z_out_56[31])
      & (fsm_output[9]));
  assign modulo_sub_22_qelse_or_nl = ((z_out_52[31]) & (~ (fsm_output[9]))) | ((z_out_57[31])
      & (fsm_output[9]));
  assign modulo_sub_23_qelse_or_nl = ((z_out_53[31]) & (~ (fsm_output[9]))) | ((z_out_58[31])
      & (fsm_output[9]));
  assign modulo_sub_24_qelse_or_nl = ((z_out_54[31]) & (~ (fsm_output[9]))) | ((z_out_59[31])
      & (fsm_output[9]));
  assign modulo_sub_25_qelse_or_nl = ((z_out_55[31]) & (~ (fsm_output[9]))) | ((z_out_60[31])
      & (fsm_output[9]));
  assign modulo_sub_26_qelse_or_nl = ((z_out_57[31]) & (~ (fsm_output[9]))) | ((z_out_61[31])
      & (fsm_output[9]));
  assign modulo_sub_27_qelse_or_nl = ((z_out_58[31]) & (~ (fsm_output[9]))) | ((z_out_62[31])
      & (fsm_output[9]));
  assign modulo_sub_28_qelse_or_nl = ((z_out_59[31]) & (~ (fsm_output[9]))) | ((z_out_63[31])
      & (fsm_output[9]));
  assign modulo_sub_29_qelse_or_nl = ((z_out_60[31]) & (~ (fsm_output[9]))) | ((z_out_64[31])
      & (fsm_output[9]));
  assign modulo_sub_30_qelse_or_nl = ((z_out_61[31]) & (~ (fsm_output[9]))) | ((z_out_65[31])
      & (fsm_output[9]));
  assign modulo_sub_31_qelse_or_nl = ((z_out_62[31]) & (~ (fsm_output[9]))) | ((z_out_66[31])
      & (fsm_output[9]));
  assign STAGE_LOOP_base_STAGE_LOOP_base_mux_nl = MUX_v_7_2_2((z_out[10:4]), (z_out_2[6:0]),
      fsm_output[4]);
  assign INNER_LOOP2_r_or_nl = (fsm_output[4]) | (fsm_output[1]) | (fsm_output[2]);
  assign operator_20_false_mux_2_nl = MUX_v_3_2_2(({butterFly2_11_tw_h_slc_operator_33_true_2_lshift_psp_2_0_1_0_itm
      , c_1_sva}), operator_20_false_acc_cse_sva, fsm_output[5]);
  assign nl_z_out_1 = operator_20_false_mux_2_nl + ({1'b1 , (~ (fsm_output[5])) ,
      1'b1});
  assign z_out_1 = nl_z_out_1[2:0];
  assign operator_20_false_mux1h_2_nl = MUX1HOT_v_7_4_2(INNER_LOOP1_r_11_4_sva_6_0,
      INNER_LOOP2_r_11_4_sva_6_0, INNER_LOOP3_r_11_4_sva_6_0, INNER_LOOP4_r_11_4_sva_6_0,
      {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_2 = conv_u2u_7_8(operator_20_false_mux1h_2_nl) + 8'b00000001;
  assign z_out_2 = nl_z_out_2[7:0];
  assign modulo_sub_6_qif_mux_2_nl = MUX_v_31_2_2((z_out_57[30:0]), (z_out_55[30:0]),
      fsm_output[7]);
  assign nl_z_out_4 = ({1'b1 , modulo_sub_6_qif_mux_2_nl}) + p_sva;
  assign z_out_4 = nl_z_out_4[31:0];
  assign modulo_sub_37_qif_mux_2_nl = MUX_v_31_2_2((z_out_54[30:0]), (z_out_58[30:0]),
      fsm_output[2]);
  assign nl_z_out_5 = ({1'b1 , modulo_sub_37_qif_mux_2_nl}) + p_sva;
  assign z_out_5 = nl_z_out_5[31:0];
  assign modulo_sub_36_qif_mux_2_nl = MUX_v_31_2_2((z_out_53[30:0]), (z_out_59[30:0]),
      fsm_output[2]);
  assign nl_z_out_8 = ({1'b1 , modulo_sub_36_qif_mux_2_nl}) + p_sva;
  assign z_out_8 = nl_z_out_8[31:0];
  assign modulo_sub_4_qif_mux_2_nl = MUX_v_31_2_2((z_out_55[30:0]), (z_out_57[30:0]),
      fsm_output[7]);
  assign nl_z_out_9 = ({1'b1 , modulo_sub_4_qif_mux_2_nl}) + p_sva;
  assign z_out_9 = nl_z_out_9[31:0];
  assign modulo_sub_35_qif_mux_2_nl = MUX_v_31_2_2((z_out_52[30:0]), (z_out_60[30:0]),
      fsm_output[2]);
  assign nl_z_out_10 = ({1'b1 , modulo_sub_35_qif_mux_2_nl}) + p_sva;
  assign z_out_10 = nl_z_out_10[31:0];
  assign modulo_sub_3_qif_mux_2_nl = MUX_v_31_2_2((z_out_54[30:0]), (z_out_58[30:0]),
      fsm_output[7]);
  assign nl_z_out_12 = ({1'b1 , modulo_sub_3_qif_mux_2_nl}) + p_sva;
  assign z_out_12 = nl_z_out_12[31:0];
  assign modulo_sub_34_qif_mux_2_nl = MUX_v_31_2_2((z_out_51[30:0]), (z_out_61[30:0]),
      fsm_output[2]);
  assign nl_z_out_13 = ({1'b1 , modulo_sub_34_qif_mux_2_nl}) + p_sva;
  assign z_out_13 = nl_z_out_13[31:0];
  assign modulo_sub_2_qif_mux_2_nl = MUX_v_31_2_2((z_out_53[30:0]), (z_out_59[30:0]),
      fsm_output[7]);
  assign nl_z_out_14 = ({1'b1 , modulo_sub_2_qif_mux_2_nl}) + p_sva;
  assign z_out_14 = nl_z_out_14[31:0];
  assign modulo_sub_33_qif_mux_2_nl = MUX_v_31_2_2((z_out_66[30:0]), (z_out_62[30:0]),
      fsm_output[2]);
  assign nl_z_out_16 = ({1'b1 , modulo_sub_33_qif_mux_2_nl}) + p_sva;
  assign z_out_16 = nl_z_out_16[31:0];
  assign modulo_sub_1_qif_mux_2_nl = MUX_v_31_2_2((z_out_52[30:0]), (z_out_60[30:0]),
      fsm_output[7]);
  assign nl_z_out_17 = ({1'b1 , modulo_sub_1_qif_mux_2_nl}) + p_sva;
  assign z_out_17 = nl_z_out_17[31:0];
  assign modulo_sub_32_qif_mux_2_nl = MUX_v_31_2_2((z_out_65[30:0]), (z_out_63[30:0]),
      fsm_output[2]);
  assign nl_z_out_18 = ({1'b1 , modulo_sub_32_qif_mux_2_nl}) + p_sva;
  assign z_out_18 = nl_z_out_18[31:0];
  assign modulo_sub_qif_mux_2_nl = MUX_v_31_2_2((z_out_51[30:0]), (z_out_61[30:0]),
      fsm_output[7]);
  assign nl_z_out_20 = ({1'b1 , modulo_sub_qif_mux_2_nl}) + p_sva;
  assign z_out_20 = nl_z_out_20[31:0];
  assign modulo_sub_31_qif_mux_2_nl = MUX_v_31_2_2((z_out_62[30:0]), (z_out_66[30:0]),
      fsm_output[9]);
  assign nl_z_out_21 = ({1'b1 , modulo_sub_31_qif_mux_2_nl}) + p_sva;
  assign z_out_21 = nl_z_out_21[31:0];
  assign modulo_sub_13_qif_mux_2_nl = MUX_v_31_2_2((z_out_64[30:0]), (z_out_63[30:0]),
      fsm_output[7]);
  assign nl_z_out_22 = ({1'b1 , modulo_sub_13_qif_mux_2_nl}) + p_sva;
  assign z_out_22 = nl_z_out_22[31:0];
  assign modulo_sub_30_qif_mux_2_nl = MUX_v_31_2_2((z_out_61[30:0]), (z_out_65[30:0]),
      fsm_output[9]);
  assign nl_z_out_24 = ({1'b1 , modulo_sub_30_qif_mux_2_nl}) + p_sva;
  assign z_out_24 = nl_z_out_24[31:0];
  assign modulo_sub_45_qif_mux_2_nl = MUX_v_31_2_2((z_out_62[30:0]), (z_out_65[30:0]),
      fsm_output[2]);
  assign nl_z_out_25 = ({1'b1 , modulo_sub_45_qif_mux_2_nl}) + p_sva;
  assign z_out_25 = nl_z_out_25[31:0];
  assign modulo_sub_29_qif_mux_2_nl = MUX_v_31_2_2((z_out_60[30:0]), (z_out_64[30:0]),
      fsm_output[9]);
  assign nl_z_out_26 = ({1'b1 , modulo_sub_29_qif_mux_2_nl}) + p_sva;
  assign z_out_26 = nl_z_out_26[31:0];
  assign modulo_sub_15_qif_mux_2_nl = MUX_v_31_2_2((z_out_66[30:0]), (z_out_64[30:0]),
      fsm_output[7]);
  assign nl_z_out_28 = ({1'b1 , modulo_sub_15_qif_mux_2_nl}) + p_sva;
  assign z_out_28 = nl_z_out_28[31:0];
  assign modulo_sub_28_qif_mux_2_nl = MUX_v_31_2_2((z_out_59[30:0]), (z_out_63[30:0]),
      fsm_output[9]);
  assign nl_z_out_29 = ({1'b1 , modulo_sub_28_qif_mux_2_nl}) + p_sva;
  assign z_out_29 = nl_z_out_29[31:0];
  assign modulo_sub_27_qif_mux_2_nl = MUX_v_31_2_2((z_out_58[30:0]), (z_out_62[30:0]),
      fsm_output[9]);
  assign nl_z_out_31 = ({1'b1 , modulo_sub_27_qif_mux_2_nl}) + p_sva;
  assign z_out_31 = nl_z_out_31[31:0];
  assign modulo_sub_26_qif_mux_2_nl = MUX_v_31_2_2((z_out_57[30:0]), (z_out_61[30:0]),
      fsm_output[9]);
  assign nl_z_out_32 = ({1'b1 , modulo_sub_26_qif_mux_2_nl}) + p_sva;
  assign z_out_32 = nl_z_out_32[31:0];
  assign modulo_sub_25_qif_mux_2_nl = MUX_v_31_2_2((z_out_55[30:0]), (z_out_60[30:0]),
      fsm_output[9]);
  assign nl_z_out_34 = ({1'b1 , modulo_sub_25_qif_mux_2_nl}) + p_sva;
  assign z_out_34 = nl_z_out_34[31:0];
  assign modulo_sub_24_qif_mux_2_nl = MUX_v_31_2_2((z_out_54[30:0]), (z_out_59[30:0]),
      fsm_output[9]);
  assign nl_z_out_36 = ({1'b1 , modulo_sub_24_qif_mux_2_nl}) + p_sva;
  assign z_out_36 = nl_z_out_36[31:0];
  assign modulo_sub_23_qif_mux_2_nl = MUX_v_31_2_2((z_out_53[30:0]), (z_out_58[30:0]),
      fsm_output[9]);
  assign nl_z_out_37 = ({1'b1 , modulo_sub_23_qif_mux_2_nl}) + p_sva;
  assign z_out_37 = nl_z_out_37[31:0];
  assign modulo_sub_22_qif_mux_2_nl = MUX_v_31_2_2((z_out_52[30:0]), (z_out_57[30:0]),
      fsm_output[9]);
  assign nl_z_out_39 = ({1'b1 , modulo_sub_22_qif_mux_2_nl}) + p_sva;
  assign z_out_39 = nl_z_out_39[31:0];
  assign modulo_sub_21_qif_mux_2_nl = MUX_v_31_2_2((z_out_51[30:0]), (z_out_56[30:0]),
      fsm_output[9]);
  assign nl_z_out_41 = ({1'b1 , modulo_sub_21_qif_mux_2_nl}) + p_sva;
  assign z_out_41 = nl_z_out_41[31:0];
  assign modulo_sub_20_qif_mux_2_nl = MUX_v_31_2_2((z_out_65[30:0]), (z_out_55[30:0]),
      fsm_output[9]);
  assign nl_z_out_42 = ({1'b1 , modulo_sub_20_qif_mux_2_nl}) + p_sva;
  assign z_out_42 = nl_z_out_42[31:0];
  assign modulo_sub_19_qif_mux_2_nl = MUX_v_31_2_2((z_out_64[30:0]), (z_out_54[30:0]),
      fsm_output[9]);
  assign nl_z_out_44 = ({1'b1 , modulo_sub_19_qif_mux_2_nl}) + p_sva;
  assign z_out_44 = nl_z_out_44[31:0];
  assign modulo_sub_18_qif_mux_2_nl = MUX_v_31_2_2((z_out_63[30:0]), (z_out_53[30:0]),
      fsm_output[9]);
  assign nl_z_out_46 = ({1'b1 , modulo_sub_18_qif_mux_2_nl}) + p_sva;
  assign z_out_46 = nl_z_out_46[31:0];
  assign modulo_sub_17_qif_mux_2_nl = MUX_v_31_2_2((z_out_56[30:0]), (z_out_52[30:0]),
      fsm_output[9]);
  assign nl_z_out_47 = ({1'b1 , modulo_sub_17_qif_mux_2_nl}) + p_sva;
  assign z_out_47 = nl_z_out_47[31:0];
  assign modulo_sub_16_qif_mux_2_nl = MUX_v_31_2_2((z_out_66[30:0]), (z_out_51[30:0]),
      fsm_output[9]);
  assign nl_z_out_49 = ({1'b1 , modulo_sub_16_qif_mux_2_nl}) + p_sva;
  assign z_out_49 = nl_z_out_49[31:0];
  assign butterFly1_mux1h_17_nl = MUX1HOT_v_32_4_2((~ mult_res_lpi_3_dfm_1), (~ reg_mult_21_res_lpi_3_dfm_1_cse),
      (~ reg_mult_24_res_lpi_3_dfm_1_cse), (~ reg_mult_17_res_lpi_3_dfm_1_cse), {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_50_nl = ({tmp_10_sva_7 , 1'b1}) + ({butterFly1_mux1h_17_nl , 1'b1});
  assign acc_50_nl = nl_acc_50_nl[32:0];
  assign z_out_51 = readslicef_33_32_1(acc_50_nl);
  assign butterFly1_1_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_1_res_lpi_3_dfm_1),
      (~ reg_mult_22_res_lpi_3_dfm_1_cse), (~ reg_mult_29_res_lpi_3_dfm_1_cse), (~
      reg_mult_25_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_51_nl = ({tmp_102_sva_7 , 1'b1}) + ({butterFly1_1_mux1h_13_nl , 1'b1});
  assign acc_51_nl = nl_acc_51_nl[32:0];
  assign z_out_52 = readslicef_33_32_1(acc_51_nl);
  assign butterFly1_2_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_2_res_lpi_3_dfm_1),
      (~ reg_mult_23_res_lpi_3_dfm_1_cse), (~ reg_mult_31_res_lpi_3_dfm_1_cse), (~
      reg_mult_28_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_52_nl = ({tmp_104_sva_7 , 1'b1}) + ({butterFly1_2_mux1h_13_nl , 1'b1});
  assign acc_52_nl = nl_acc_52_nl[32:0];
  assign z_out_53 = readslicef_33_32_1(acc_52_nl);
  assign butterFly1_3_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_3_res_lpi_3_dfm_1),
      (~ reg_mult_24_res_lpi_3_dfm_1_cse), (~ reg_mult_27_res_lpi_3_dfm_1_cse), (~
      reg_mult_20_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_53_nl = ({tmp_106_sva_7 , 1'b1}) + ({butterFly1_3_mux1h_13_nl , 1'b1});
  assign acc_53_nl = nl_acc_53_nl[32:0];
  assign z_out_54 = readslicef_33_32_1(acc_53_nl);
  assign butterFly1_4_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_4_res_lpi_3_dfm_1),
      (~ reg_mult_25_res_lpi_3_dfm_1_cse), (~ reg_mult_23_res_lpi_3_dfm_1_cse), (~
      reg_mult_22_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_54_nl = ({tmp_108_sva_7 , 1'b1}) + ({butterFly1_4_mux1h_13_nl , 1'b1});
  assign acc_54_nl = nl_acc_54_nl[32:0];
  assign z_out_55 = readslicef_33_32_1(acc_54_nl);
  assign butterFly1_5_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_5_res_lpi_3_dfm_1),
      (~ reg_mult_17_res_lpi_3_dfm_1_cse), (~ reg_mult_19_res_lpi_3_dfm_1_cse), (~
      reg_mult_30_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_55_nl = ({tmp_110_sva_7 , 1'b1}) + ({butterFly1_5_mux1h_13_nl , 1'b1});
  assign acc_55_nl = nl_acc_55_nl[32:0];
  assign z_out_56 = readslicef_33_32_1(acc_55_nl);
  assign butterFly1_6_mux1h_13_nl = MUX1HOT_v_32_3_2((~ mult_6_res_lpi_3_dfm_1),
      (~ reg_mult_26_res_lpi_3_dfm_1_cse), (~ reg_mult_18_res_lpi_3_dfm_1_cse), {(fsm_output[2])
      , or_dcpl_194 , (fsm_output[7])});
  assign nl_acc_56_nl = ({tmp_112_sva_7 , 1'b1}) + ({butterFly1_6_mux1h_13_nl , 1'b1});
  assign acc_56_nl = nl_acc_56_nl[32:0];
  assign z_out_57 = readslicef_33_32_1(acc_56_nl);
  assign butterFly1_7_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_7_res_lpi_3_dfm_1),
      (~ reg_mult_27_res_lpi_3_dfm_1_cse), (~ reg_mult_26_res_lpi_3_dfm_1_cse), (~
      reg_mult_18_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_57_nl = ({tmp_114_sva_7 , 1'b1}) + ({butterFly1_7_mux1h_13_nl , 1'b1});
  assign acc_57_nl = nl_acc_57_nl[32:0];
  assign z_out_58 = readslicef_33_32_1(acc_57_nl);
  assign butterFly1_8_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_8_res_lpi_3_dfm_1),
      (~ reg_mult_28_res_lpi_3_dfm_1_cse), (~ reg_mult_30_res_lpi_3_dfm_1_cse), (~
      reg_mult_19_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_58_nl = ({tmp_116_sva_7 , 1'b1}) + ({butterFly1_8_mux1h_13_nl , 1'b1});
  assign acc_58_nl = nl_acc_58_nl[32:0];
  assign z_out_59 = readslicef_33_32_1(acc_58_nl);
  assign butterFly1_9_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_9_res_lpi_3_dfm_1),
      (~ reg_mult_29_res_lpi_3_dfm_1_cse), (~ reg_mult_22_res_lpi_3_dfm_1_cse), (~
      reg_mult_23_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_59_nl = ({tmp_118_sva_7 , 1'b1}) + ({butterFly1_9_mux1h_13_nl , 1'b1});
  assign acc_59_nl = nl_acc_59_nl[32:0];
  assign z_out_60 = readslicef_33_32_1(acc_59_nl);
  assign butterFly1_10_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_10_res_lpi_3_dfm_1),
      (~ reg_mult_30_res_lpi_3_dfm_1_cse), (~ reg_mult_20_res_lpi_3_dfm_1_cse), (~
      reg_mult_27_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_60_nl = ({tmp_120_sva_7 , 1'b1}) + ({butterFly1_10_mux1h_13_nl ,
      1'b1});
  assign acc_60_nl = nl_acc_60_nl[32:0];
  assign z_out_61 = readslicef_33_32_1(acc_60_nl);
  assign butterFly1_11_mux1h_13_nl = MUX1HOT_v_32_3_2((~ mult_11_res_lpi_3_dfm_1),
      (~ reg_mult_31_res_lpi_3_dfm_1_cse), (~ reg_mult_28_res_lpi_3_dfm_1_cse), {(fsm_output[2])
      , or_dcpl_194 , (fsm_output[7])});
  assign nl_acc_61_nl = ({tmp_122_sva_7 , 1'b1}) + ({butterFly1_11_mux1h_13_nl ,
      1'b1});
  assign acc_61_nl = nl_acc_61_nl[32:0];
  assign z_out_62 = readslicef_33_32_1(acc_61_nl);
  assign butterFly1_12_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_12_res_lpi_3_dfm_1),
      (~ reg_mult_18_res_lpi_3_dfm_1_cse), (~ reg_mult_25_res_lpi_3_dfm_1_cse), (~
      reg_mult_29_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_62_nl = ({tmp_124_sva_7 , 1'b1}) + ({butterFly1_12_mux1h_13_nl ,
      1'b1});
  assign acc_62_nl = nl_acc_62_nl[32:0];
  assign z_out_63 = readslicef_33_32_1(acc_62_nl);
  assign butterFly1_13_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_13_res_lpi_3_dfm_1),
      (~ reg_mult_19_res_lpi_3_dfm_1_cse), (~ reg_mult_17_res_lpi_3_dfm_1_cse), (~
      reg_mult_24_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_63_nl = ({tmp_126_sva_7 , 1'b1}) + ({butterFly1_13_mux1h_13_nl ,
      1'b1});
  assign acc_63_nl = nl_acc_63_nl[32:0];
  assign z_out_64 = readslicef_33_32_1(acc_63_nl);
  assign butterFly1_14_mux1h_13_nl = MUX1HOT_v_32_4_2((~ mult_14_res_lpi_3_dfm_1),
      (~ reg_mult_20_res_lpi_3_dfm_1_cse), (~ reg_mult_16_res_lpi_3_dfm_1_cse), (~
      reg_mult_21_res_lpi_3_dfm_1_cse), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_64_nl = ({tmp_60_sva_7 , 1'b1}) + ({butterFly1_14_mux1h_13_nl , 1'b1});
  assign acc_64_nl = nl_acc_64_nl[32:0];
  assign z_out_65 = readslicef_33_32_1(acc_64_nl);
  assign butterFly1_15_mux1h_13_nl = MUX1HOT_v_32_3_2((~ mult_15_res_lpi_3_dfm_1),
      (~ reg_mult_16_res_lpi_3_dfm_1_cse), (~ reg_mult_21_res_lpi_3_dfm_1_cse), {(fsm_output[2])
      , or_dcpl_194 , (fsm_output[7])});
  assign nl_acc_65_nl = ({tmp_62_sva_7 , 1'b1}) + ({butterFly1_15_mux1h_13_nl , 1'b1});
  assign acc_65_nl = nl_acc_65_nl[32:0];
  assign z_out_66 = readslicef_33_32_1(acc_65_nl);
  assign butterFly1_15_mux1h_14_nl = MUX1HOT_v_32_3_2(mult_15_res_lpi_3_dfm_1, reg_mult_16_res_lpi_3_dfm_1_cse,
      reg_mult_21_res_lpi_3_dfm_1_cse, {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
  assign nl_z_out_67 = tmp_62_sva_7 + butterFly1_15_mux1h_14_nl;
  assign z_out_67 = nl_z_out_67[31:0];
  assign butterFly1_14_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_14_res_lpi_3_dfm_1, reg_mult_20_res_lpi_3_dfm_1_cse,
      reg_mult_16_res_lpi_3_dfm_1_cse, reg_mult_21_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_68 = tmp_60_sva_7 + butterFly1_14_mux1h_14_nl;
  assign z_out_68 = nl_z_out_68[31:0];
  assign butterFly1_13_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_13_res_lpi_3_dfm_1, reg_mult_19_res_lpi_3_dfm_1_cse,
      reg_mult_17_res_lpi_3_dfm_1_cse, reg_mult_24_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_69 = tmp_126_sva_7 + butterFly1_13_mux1h_14_nl;
  assign z_out_69 = nl_z_out_69[31:0];
  assign butterFly1_12_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_12_res_lpi_3_dfm_1, reg_mult_18_res_lpi_3_dfm_1_cse,
      reg_mult_25_res_lpi_3_dfm_1_cse, reg_mult_29_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_70 = tmp_124_sva_7 + butterFly1_12_mux1h_14_nl;
  assign z_out_70 = nl_z_out_70[31:0];
  assign butterFly1_11_mux1h_14_nl = MUX1HOT_v_32_3_2(mult_11_res_lpi_3_dfm_1, reg_mult_31_res_lpi_3_dfm_1_cse,
      reg_mult_28_res_lpi_3_dfm_1_cse, {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
  assign nl_z_out_71 = tmp_122_sva_7 + butterFly1_11_mux1h_14_nl;
  assign z_out_71 = nl_z_out_71[31:0];
  assign butterFly1_10_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_10_res_lpi_3_dfm_1, reg_mult_30_res_lpi_3_dfm_1_cse,
      reg_mult_20_res_lpi_3_dfm_1_cse, reg_mult_27_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_72 = tmp_120_sva_7 + butterFly1_10_mux1h_14_nl;
  assign z_out_72 = nl_z_out_72[31:0];
  assign butterFly1_9_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_9_res_lpi_3_dfm_1, reg_mult_29_res_lpi_3_dfm_1_cse,
      reg_mult_22_res_lpi_3_dfm_1_cse, reg_mult_23_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_73 = tmp_118_sva_7 + butterFly1_9_mux1h_14_nl;
  assign z_out_73 = nl_z_out_73[31:0];
  assign butterFly1_8_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_8_res_lpi_3_dfm_1, reg_mult_28_res_lpi_3_dfm_1_cse,
      reg_mult_30_res_lpi_3_dfm_1_cse, reg_mult_19_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_74 = tmp_116_sva_7 + butterFly1_8_mux1h_14_nl;
  assign z_out_74 = nl_z_out_74[31:0];
  assign butterFly1_7_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_7_res_lpi_3_dfm_1, reg_mult_27_res_lpi_3_dfm_1_cse,
      reg_mult_26_res_lpi_3_dfm_1_cse, reg_mult_18_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_75 = tmp_114_sva_7 + butterFly1_7_mux1h_14_nl;
  assign z_out_75 = nl_z_out_75[31:0];
  assign butterFly1_6_mux1h_14_nl = MUX1HOT_v_32_3_2(mult_6_res_lpi_3_dfm_1, reg_mult_26_res_lpi_3_dfm_1_cse,
      reg_mult_18_res_lpi_3_dfm_1_cse, {(fsm_output[2]) , or_dcpl_194 , (fsm_output[7])});
  assign nl_z_out_76 = tmp_112_sva_7 + butterFly1_6_mux1h_14_nl;
  assign z_out_76 = nl_z_out_76[31:0];
  assign butterFly1_5_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_5_res_lpi_3_dfm_1, reg_mult_17_res_lpi_3_dfm_1_cse,
      reg_mult_19_res_lpi_3_dfm_1_cse, reg_mult_30_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_77 = tmp_110_sva_7 + butterFly1_5_mux1h_14_nl;
  assign z_out_77 = nl_z_out_77[31:0];
  assign butterFly1_4_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_4_res_lpi_3_dfm_1, reg_mult_25_res_lpi_3_dfm_1_cse,
      reg_mult_23_res_lpi_3_dfm_1_cse, reg_mult_22_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_78 = tmp_108_sva_7 + butterFly1_4_mux1h_14_nl;
  assign z_out_78 = nl_z_out_78[31:0];
  assign butterFly1_3_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_3_res_lpi_3_dfm_1, reg_mult_24_res_lpi_3_dfm_1_cse,
      reg_mult_27_res_lpi_3_dfm_1_cse, reg_mult_20_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_79 = tmp_106_sva_7 + butterFly1_3_mux1h_14_nl;
  assign z_out_79 = nl_z_out_79[31:0];
  assign butterFly1_2_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_2_res_lpi_3_dfm_1, reg_mult_23_res_lpi_3_dfm_1_cse,
      reg_mult_31_res_lpi_3_dfm_1_cse, reg_mult_28_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_80 = tmp_104_sva_7 + butterFly1_2_mux1h_14_nl;
  assign z_out_80 = nl_z_out_80[31:0];
  assign butterFly1_1_mux1h_14_nl = MUX1HOT_v_32_4_2(mult_1_res_lpi_3_dfm_1, reg_mult_22_res_lpi_3_dfm_1_cse,
      reg_mult_29_res_lpi_3_dfm_1_cse, reg_mult_25_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_81 = tmp_102_sva_7 + butterFly1_1_mux1h_14_nl;
  assign z_out_81 = nl_z_out_81[31:0];
  assign butterFly1_mux1h_18_nl = MUX1HOT_v_32_4_2(mult_res_lpi_3_dfm_1, reg_mult_21_res_lpi_3_dfm_1_cse,
      reg_mult_24_res_lpi_3_dfm_1_cse, reg_mult_17_res_lpi_3_dfm_1_cse, {(fsm_output[2])
      , (fsm_output[4]) , (fsm_output[7]) , (fsm_output[9])});
  assign nl_z_out_82 = tmp_10_sva_7 + butterFly1_mux1h_18_nl;
  assign z_out_82 = nl_z_out_82[31:0];
  assign modulo_add_1_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_81), (~ z_out_78), (~
      z_out_67), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_82_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_1_mux1h_3_nl
      , 1'b1});
  assign acc_82_nl = nl_acc_82_nl[33:0];
  assign z_out_83_32 = readslicef_34_1_33(acc_82_nl);
  assign modulo_add_10_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_72), (~ z_out_67),
      (~ z_out_68), (~ z_out_71), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_83_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_10_mux1h_3_nl
      , 1'b1});
  assign acc_83_nl = nl_acc_83_nl[33:0];
  assign z_out_84_32 = readslicef_34_1_33(acc_83_nl);
  assign modulo_add_54_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_76), (~ z_out_73),
      (~ z_out_75), (~ z_out_74), {(fsm_output[9]) , (fsm_output[7]) , (fsm_output[2])
      , (fsm_output[4])});
  assign nl_acc_84_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_54_mux1h_3_nl
      , 1'b1});
  assign acc_84_nl = nl_acc_84_nl[33:0];
  assign z_out_85_32 = readslicef_34_1_33(acc_84_nl);
  assign modulo_add_48_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_82), (~ z_out_71),
      (~ z_out_77), (~ z_out_69), {(fsm_output[9]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7])});
  assign nl_acc_85_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_48_mux1h_3_nl
      , 1'b1});
  assign acc_85_nl = nl_acc_85_nl[33:0];
  assign z_out_86_32 = readslicef_34_1_33(acc_85_nl);
  assign modulo_add_33_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_67), (~ z_out_81),
      (~ z_out_70), {(fsm_output[7]) , (fsm_output[9]) , modulo_add_1_qelse_or_m1c});
  assign nl_acc_86_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_33_mux1h_3_nl
      , 1'b1});
  assign acc_86_nl = nl_acc_86_nl[33:0];
  assign z_out_87_32 = readslicef_34_1_33(acc_86_nl);
  assign modulo_add_34_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_82), (~ z_out_72),
      (~ z_out_71), {or_dcpl_210 , (fsm_output[9]) , (fsm_output[4])});
  assign nl_acc_87_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_34_mux1h_3_nl
      , 1'b1});
  assign acc_87_nl = nl_acc_87_nl[33:0];
  assign z_out_88_32 = readslicef_34_1_33(acc_87_nl);
  assign modulo_add_6_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_76), (~ z_out_75), (~
      z_out_72), (~ z_out_68), {(fsm_output[2]) , (fsm_output[4]) , (fsm_output[7])
      , (fsm_output[9])});
  assign nl_acc_88_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_6_mux1h_3_nl
      , 1'b1});
  assign acc_88_nl = nl_acc_88_nl[33:0];
  assign z_out_89_32 = readslicef_34_1_33(acc_88_nl);
  assign modulo_add_50_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_80), (~ z_out_69),
      (~ z_out_81), {(fsm_output[9]) , modulo_add_1_qelse_or_m1c , (fsm_output[7])});
  assign nl_acc_89_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_50_mux1h_3_nl
      , 1'b1});
  assign acc_89_nl = nl_acc_89_nl[33:0];
  assign z_out_90_32 = readslicef_34_1_33(acc_89_nl);
  assign modulo_add_51_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_79), (~ z_out_77),
      (~ z_out_76), (~ z_out_74), {(fsm_output[9]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[7])});
  assign nl_acc_90_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_51_mux1h_3_nl
      , 1'b1});
  assign acc_90_nl = nl_acc_90_nl[33:0];
  assign z_out_91_32 = readslicef_34_1_33(acc_90_nl);
  assign modulo_add_14_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_68), (~ z_out_73),
      (~ z_out_70), {modulo_add_1_qelse_or_m1c , (fsm_output[9]) , (fsm_output[7])});
  assign nl_acc_91_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_14_mux1h_3_nl
      , 1'b1});
  assign acc_91_nl = nl_acc_91_nl[33:0];
  assign z_out_92_32 = readslicef_34_1_33(acc_91_nl);
  assign modulo_add_36_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_80), (~ z_out_67),
      (~ z_out_82), (~ z_out_70), {(fsm_output[7]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[9])});
  assign nl_acc_92_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_36_mux1h_3_nl
      , 1'b1});
  assign acc_92_nl = nl_acc_92_nl[33:0];
  assign z_out_93_32 = readslicef_34_1_33(acc_92_nl);
  assign modulo_add_52_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_78), (~ z_out_79),
      (~ z_out_73), (~ z_out_72), {(fsm_output[9]) , (fsm_output[7]) , (fsm_output[2])
      , (fsm_output[4])});
  assign nl_acc_93_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_52_mux1h_3_nl
      , 1'b1});
  assign acc_93_nl = nl_acc_93_nl[33:0];
  assign z_out_94_32 = readslicef_34_1_33(acc_93_nl);
  assign modulo_add_41_mux1h_3_nl = MUX1HOT_v_32_4_2((~ z_out_75), (~ z_out_74),
      (~ z_out_73), (~ z_out_69), {(fsm_output[7]) , (fsm_output[2]) , (fsm_output[4])
      , (fsm_output[9])});
  assign nl_acc_94_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_41_mux1h_3_nl
      , 1'b1});
  assign acc_94_nl = nl_acc_94_nl[33:0];
  assign z_out_95_32 = readslicef_34_1_33(acc_94_nl);
  assign modulo_add_2_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_80), (~ z_out_77), (~
      z_out_74), {modulo_add_1_qelse_or_m1c , (fsm_output[7]) , (fsm_output[9])});
  assign nl_acc_95_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_2_mux1h_3_nl
      , 1'b1});
  assign acc_95_nl = nl_acc_95_nl[33:0];
  assign z_out_96_32 = readslicef_34_1_33(acc_95_nl);
  assign modulo_add_53_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_77), (~ z_out_76),
      (~ z_out_78), {(fsm_output[9]) , (fsm_output[7]) , modulo_add_1_qelse_or_m1c});
  assign nl_acc_96_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_53_mux1h_3_nl
      , 1'b1});
  assign acc_96_nl = nl_acc_96_nl[33:0];
  assign z_out_97_32 = readslicef_34_1_33(acc_96_nl);
  assign modulo_add_55_mux1h_3_nl = MUX1HOT_v_32_3_2((~ z_out_75), (~ z_out_79),
      (~ z_out_71), {(fsm_output[9]) , modulo_add_1_qelse_or_m1c , (fsm_output[7])});
  assign nl_acc_97_nl = ({1'b1 , p_sva , 1'b1}) + conv_u2u_33_34({modulo_add_55_mux1h_3_nl
      , 1'b1});
  assign acc_97_nl = nl_acc_97_nl[33:0];
  assign z_out_98_32 = readslicef_34_1_33(acc_97_nl);

  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    result = result | ( input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [30:0] MUX1HOT_v_31_3_2;
    input [30:0] input_2;
    input [30:0] input_1;
    input [30:0] input_0;
    input [2:0] sel;
    reg [30:0] result;
  begin
    result = input_0 & {31{sel[0]}};
    result = result | ( input_1 & {31{sel[1]}});
    result = result | ( input_2 & {31{sel[2]}});
    MUX1HOT_v_31_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_12_2;
    input [31:0] input_11;
    input [31:0] input_10;
    input [31:0] input_9;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [11:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    result = result | ( input_9 & {32{sel[9]}});
    result = result | ( input_10 & {32{sel[10]}});
    result = result | ( input_11 & {32{sel[11]}});
    MUX1HOT_v_32_12_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_3_2;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [2:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    MUX1HOT_v_32_3_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_4_2;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [3:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    MUX1HOT_v_32_4_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_5_2;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [4:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    MUX1HOT_v_32_5_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_6_2;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [5:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    MUX1HOT_v_32_6_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_8_2;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [7:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    MUX1HOT_v_32_8_2 = result;
  end
  endfunction


  function automatic [31:0] MUX1HOT_v_32_9_2;
    input [31:0] input_8;
    input [31:0] input_7;
    input [31:0] input_6;
    input [31:0] input_5;
    input [31:0] input_4;
    input [31:0] input_3;
    input [31:0] input_2;
    input [31:0] input_1;
    input [31:0] input_0;
    input [8:0] sel;
    reg [31:0] result;
  begin
    result = input_0 & {32{sel[0]}};
    result = result | ( input_1 & {32{sel[1]}});
    result = result | ( input_2 & {32{sel[2]}});
    result = result | ( input_3 & {32{sel[3]}});
    result = result | ( input_4 & {32{sel[4]}});
    result = result | ( input_5 & {32{sel[5]}});
    result = result | ( input_6 & {32{sel[6]}});
    result = result | ( input_7 & {32{sel[7]}});
    result = result | ( input_8 & {32{sel[8]}});
    MUX1HOT_v_32_9_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | ( input_1 & {6{sel[1]}});
    result = result | ( input_2 & {6{sel[2]}});
    result = result | ( input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_4_2;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [3:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | ( input_1 & {7{sel[1]}});
    result = result | ( input_2 & {7{sel[2]}});
    result = result | ( input_3 & {7{sel[3]}});
    MUX1HOT_v_7_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_33_1_32;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 32;
    readslicef_33_1_32 = tmp[0:0];
  end
  endfunction


  function automatic [31:0] readslicef_33_32_1;
    input [32:0] vector;
    reg [32:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_33_32_1 = tmp[31:0];
  end
  endfunction


  function automatic [0:0] readslicef_34_1_33;
    input [33:0] vector;
    reg [33:0] tmp;
  begin
    tmp = vector >> 33;
    readslicef_34_1_33 = tmp[0:0];
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [32:0] conv_u2u_32_33 ;
    input [31:0]  vector ;
  begin
    conv_u2u_32_33 = {1'b0, vector};
  end
  endfunction


  function automatic [33:0] conv_u2u_33_34 ;
    input [32:0]  vector ;
  begin
    conv_u2u_33_34 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    peaseNTT
// ------------------------------------------------------------------


module peaseNTT (
  clk, rst, xt_rsc_0_0_adra, xt_rsc_0_0_da, xt_rsc_0_0_wea, xt_rsc_0_0_qa, xt_rsc_0_0_adrb,
      xt_rsc_0_0_db, xt_rsc_0_0_web, xt_rsc_0_0_qb, xt_rsc_triosy_0_0_lz, xt_rsc_0_1_adra,
      xt_rsc_0_1_da, xt_rsc_0_1_wea, xt_rsc_0_1_qa, xt_rsc_0_1_adrb, xt_rsc_0_1_db,
      xt_rsc_0_1_web, xt_rsc_0_1_qb, xt_rsc_triosy_0_1_lz, xt_rsc_0_2_adra, xt_rsc_0_2_da,
      xt_rsc_0_2_wea, xt_rsc_0_2_qa, xt_rsc_0_2_adrb, xt_rsc_0_2_db, xt_rsc_0_2_web,
      xt_rsc_0_2_qb, xt_rsc_triosy_0_2_lz, xt_rsc_0_3_adra, xt_rsc_0_3_da, xt_rsc_0_3_wea,
      xt_rsc_0_3_qa, xt_rsc_0_3_adrb, xt_rsc_0_3_db, xt_rsc_0_3_web, xt_rsc_0_3_qb,
      xt_rsc_triosy_0_3_lz, xt_rsc_0_4_adra, xt_rsc_0_4_da, xt_rsc_0_4_wea, xt_rsc_0_4_qa,
      xt_rsc_0_4_adrb, xt_rsc_0_4_db, xt_rsc_0_4_web, xt_rsc_0_4_qb, xt_rsc_triosy_0_4_lz,
      xt_rsc_0_5_adra, xt_rsc_0_5_da, xt_rsc_0_5_wea, xt_rsc_0_5_qa, xt_rsc_0_5_adrb,
      xt_rsc_0_5_db, xt_rsc_0_5_web, xt_rsc_0_5_qb, xt_rsc_triosy_0_5_lz, xt_rsc_0_6_adra,
      xt_rsc_0_6_da, xt_rsc_0_6_wea, xt_rsc_0_6_qa, xt_rsc_0_6_adrb, xt_rsc_0_6_db,
      xt_rsc_0_6_web, xt_rsc_0_6_qb, xt_rsc_triosy_0_6_lz, xt_rsc_0_7_adra, xt_rsc_0_7_da,
      xt_rsc_0_7_wea, xt_rsc_0_7_qa, xt_rsc_0_7_adrb, xt_rsc_0_7_db, xt_rsc_0_7_web,
      xt_rsc_0_7_qb, xt_rsc_triosy_0_7_lz, xt_rsc_0_8_adra, xt_rsc_0_8_da, xt_rsc_0_8_wea,
      xt_rsc_0_8_qa, xt_rsc_0_8_adrb, xt_rsc_0_8_db, xt_rsc_0_8_web, xt_rsc_0_8_qb,
      xt_rsc_triosy_0_8_lz, xt_rsc_0_9_adra, xt_rsc_0_9_da, xt_rsc_0_9_wea, xt_rsc_0_9_qa,
      xt_rsc_0_9_adrb, xt_rsc_0_9_db, xt_rsc_0_9_web, xt_rsc_0_9_qb, xt_rsc_triosy_0_9_lz,
      xt_rsc_0_10_adra, xt_rsc_0_10_da, xt_rsc_0_10_wea, xt_rsc_0_10_qa, xt_rsc_0_10_adrb,
      xt_rsc_0_10_db, xt_rsc_0_10_web, xt_rsc_0_10_qb, xt_rsc_triosy_0_10_lz, xt_rsc_0_11_adra,
      xt_rsc_0_11_da, xt_rsc_0_11_wea, xt_rsc_0_11_qa, xt_rsc_0_11_adrb, xt_rsc_0_11_db,
      xt_rsc_0_11_web, xt_rsc_0_11_qb, xt_rsc_triosy_0_11_lz, xt_rsc_0_12_adra, xt_rsc_0_12_da,
      xt_rsc_0_12_wea, xt_rsc_0_12_qa, xt_rsc_0_12_adrb, xt_rsc_0_12_db, xt_rsc_0_12_web,
      xt_rsc_0_12_qb, xt_rsc_triosy_0_12_lz, xt_rsc_0_13_adra, xt_rsc_0_13_da, xt_rsc_0_13_wea,
      xt_rsc_0_13_qa, xt_rsc_0_13_adrb, xt_rsc_0_13_db, xt_rsc_0_13_web, xt_rsc_0_13_qb,
      xt_rsc_triosy_0_13_lz, xt_rsc_0_14_adra, xt_rsc_0_14_da, xt_rsc_0_14_wea, xt_rsc_0_14_qa,
      xt_rsc_0_14_adrb, xt_rsc_0_14_db, xt_rsc_0_14_web, xt_rsc_0_14_qb, xt_rsc_triosy_0_14_lz,
      xt_rsc_0_15_adra, xt_rsc_0_15_da, xt_rsc_0_15_wea, xt_rsc_0_15_qa, xt_rsc_0_15_adrb,
      xt_rsc_0_15_db, xt_rsc_0_15_web, xt_rsc_0_15_qb, xt_rsc_triosy_0_15_lz, xt_rsc_0_16_adra,
      xt_rsc_0_16_da, xt_rsc_0_16_wea, xt_rsc_0_16_qa, xt_rsc_0_16_adrb, xt_rsc_0_16_db,
      xt_rsc_0_16_web, xt_rsc_0_16_qb, xt_rsc_triosy_0_16_lz, xt_rsc_0_17_adra, xt_rsc_0_17_da,
      xt_rsc_0_17_wea, xt_rsc_0_17_qa, xt_rsc_0_17_adrb, xt_rsc_0_17_db, xt_rsc_0_17_web,
      xt_rsc_0_17_qb, xt_rsc_triosy_0_17_lz, xt_rsc_0_18_adra, xt_rsc_0_18_da, xt_rsc_0_18_wea,
      xt_rsc_0_18_qa, xt_rsc_0_18_adrb, xt_rsc_0_18_db, xt_rsc_0_18_web, xt_rsc_0_18_qb,
      xt_rsc_triosy_0_18_lz, xt_rsc_0_19_adra, xt_rsc_0_19_da, xt_rsc_0_19_wea, xt_rsc_0_19_qa,
      xt_rsc_0_19_adrb, xt_rsc_0_19_db, xt_rsc_0_19_web, xt_rsc_0_19_qb, xt_rsc_triosy_0_19_lz,
      xt_rsc_0_20_adra, xt_rsc_0_20_da, xt_rsc_0_20_wea, xt_rsc_0_20_qa, xt_rsc_0_20_adrb,
      xt_rsc_0_20_db, xt_rsc_0_20_web, xt_rsc_0_20_qb, xt_rsc_triosy_0_20_lz, xt_rsc_0_21_adra,
      xt_rsc_0_21_da, xt_rsc_0_21_wea, xt_rsc_0_21_qa, xt_rsc_0_21_adrb, xt_rsc_0_21_db,
      xt_rsc_0_21_web, xt_rsc_0_21_qb, xt_rsc_triosy_0_21_lz, xt_rsc_0_22_adra, xt_rsc_0_22_da,
      xt_rsc_0_22_wea, xt_rsc_0_22_qa, xt_rsc_0_22_adrb, xt_rsc_0_22_db, xt_rsc_0_22_web,
      xt_rsc_0_22_qb, xt_rsc_triosy_0_22_lz, xt_rsc_0_23_adra, xt_rsc_0_23_da, xt_rsc_0_23_wea,
      xt_rsc_0_23_qa, xt_rsc_0_23_adrb, xt_rsc_0_23_db, xt_rsc_0_23_web, xt_rsc_0_23_qb,
      xt_rsc_triosy_0_23_lz, xt_rsc_0_24_adra, xt_rsc_0_24_da, xt_rsc_0_24_wea, xt_rsc_0_24_qa,
      xt_rsc_0_24_adrb, xt_rsc_0_24_db, xt_rsc_0_24_web, xt_rsc_0_24_qb, xt_rsc_triosy_0_24_lz,
      xt_rsc_0_25_adra, xt_rsc_0_25_da, xt_rsc_0_25_wea, xt_rsc_0_25_qa, xt_rsc_0_25_adrb,
      xt_rsc_0_25_db, xt_rsc_0_25_web, xt_rsc_0_25_qb, xt_rsc_triosy_0_25_lz, xt_rsc_0_26_adra,
      xt_rsc_0_26_da, xt_rsc_0_26_wea, xt_rsc_0_26_qa, xt_rsc_0_26_adrb, xt_rsc_0_26_db,
      xt_rsc_0_26_web, xt_rsc_0_26_qb, xt_rsc_triosy_0_26_lz, xt_rsc_0_27_adra, xt_rsc_0_27_da,
      xt_rsc_0_27_wea, xt_rsc_0_27_qa, xt_rsc_0_27_adrb, xt_rsc_0_27_db, xt_rsc_0_27_web,
      xt_rsc_0_27_qb, xt_rsc_triosy_0_27_lz, xt_rsc_0_28_adra, xt_rsc_0_28_da, xt_rsc_0_28_wea,
      xt_rsc_0_28_qa, xt_rsc_0_28_adrb, xt_rsc_0_28_db, xt_rsc_0_28_web, xt_rsc_0_28_qb,
      xt_rsc_triosy_0_28_lz, xt_rsc_0_29_adra, xt_rsc_0_29_da, xt_rsc_0_29_wea, xt_rsc_0_29_qa,
      xt_rsc_0_29_adrb, xt_rsc_0_29_db, xt_rsc_0_29_web, xt_rsc_0_29_qb, xt_rsc_triosy_0_29_lz,
      xt_rsc_0_30_adra, xt_rsc_0_30_da, xt_rsc_0_30_wea, xt_rsc_0_30_qa, xt_rsc_0_30_adrb,
      xt_rsc_0_30_db, xt_rsc_0_30_web, xt_rsc_0_30_qb, xt_rsc_triosy_0_30_lz, xt_rsc_0_31_adra,
      xt_rsc_0_31_da, xt_rsc_0_31_wea, xt_rsc_0_31_qa, xt_rsc_0_31_adrb, xt_rsc_0_31_db,
      xt_rsc_0_31_web, xt_rsc_0_31_qb, xt_rsc_triosy_0_31_lz, p_rsc_dat, p_rsc_triosy_lz,
      r_rsc_dat, r_rsc_triosy_lz, twiddle_rsc_0_0_adra, twiddle_rsc_0_0_da, twiddle_rsc_0_0_wea,
      twiddle_rsc_0_0_qa, twiddle_rsc_0_0_adrb, twiddle_rsc_0_0_db, twiddle_rsc_0_0_web,
      twiddle_rsc_0_0_qb, twiddle_rsc_triosy_0_0_lz, twiddle_rsc_0_1_adra, twiddle_rsc_0_1_da,
      twiddle_rsc_0_1_wea, twiddle_rsc_0_1_qa, twiddle_rsc_0_1_adrb, twiddle_rsc_0_1_db,
      twiddle_rsc_0_1_web, twiddle_rsc_0_1_qb, twiddle_rsc_triosy_0_1_lz, twiddle_rsc_0_2_adra,
      twiddle_rsc_0_2_da, twiddle_rsc_0_2_wea, twiddle_rsc_0_2_qa, twiddle_rsc_0_2_adrb,
      twiddle_rsc_0_2_db, twiddle_rsc_0_2_web, twiddle_rsc_0_2_qb, twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_0_3_adra, twiddle_rsc_0_3_da, twiddle_rsc_0_3_wea, twiddle_rsc_0_3_qa,
      twiddle_rsc_0_3_adrb, twiddle_rsc_0_3_db, twiddle_rsc_0_3_web, twiddle_rsc_0_3_qb,
      twiddle_rsc_triosy_0_3_lz, twiddle_rsc_0_4_adra, twiddle_rsc_0_4_da, twiddle_rsc_0_4_wea,
      twiddle_rsc_0_4_qa, twiddle_rsc_0_4_adrb, twiddle_rsc_0_4_db, twiddle_rsc_0_4_web,
      twiddle_rsc_0_4_qb, twiddle_rsc_triosy_0_4_lz, twiddle_rsc_0_5_adra, twiddle_rsc_0_5_da,
      twiddle_rsc_0_5_wea, twiddle_rsc_0_5_qa, twiddle_rsc_0_5_adrb, twiddle_rsc_0_5_db,
      twiddle_rsc_0_5_web, twiddle_rsc_0_5_qb, twiddle_rsc_triosy_0_5_lz, twiddle_rsc_0_6_adra,
      twiddle_rsc_0_6_da, twiddle_rsc_0_6_wea, twiddle_rsc_0_6_qa, twiddle_rsc_0_6_adrb,
      twiddle_rsc_0_6_db, twiddle_rsc_0_6_web, twiddle_rsc_0_6_qb, twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_0_7_adra, twiddle_rsc_0_7_da, twiddle_rsc_0_7_wea, twiddle_rsc_0_7_qa,
      twiddle_rsc_0_7_adrb, twiddle_rsc_0_7_db, twiddle_rsc_0_7_web, twiddle_rsc_0_7_qb,
      twiddle_rsc_triosy_0_7_lz, twiddle_rsc_0_8_adra, twiddle_rsc_0_8_da, twiddle_rsc_0_8_wea,
      twiddle_rsc_0_8_qa, twiddle_rsc_0_8_adrb, twiddle_rsc_0_8_db, twiddle_rsc_0_8_web,
      twiddle_rsc_0_8_qb, twiddle_rsc_triosy_0_8_lz, twiddle_rsc_0_9_adra, twiddle_rsc_0_9_da,
      twiddle_rsc_0_9_wea, twiddle_rsc_0_9_qa, twiddle_rsc_0_9_adrb, twiddle_rsc_0_9_db,
      twiddle_rsc_0_9_web, twiddle_rsc_0_9_qb, twiddle_rsc_triosy_0_9_lz, twiddle_rsc_0_10_adra,
      twiddle_rsc_0_10_da, twiddle_rsc_0_10_wea, twiddle_rsc_0_10_qa, twiddle_rsc_0_10_adrb,
      twiddle_rsc_0_10_db, twiddle_rsc_0_10_web, twiddle_rsc_0_10_qb, twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_0_11_adra, twiddle_rsc_0_11_da, twiddle_rsc_0_11_wea, twiddle_rsc_0_11_qa,
      twiddle_rsc_0_11_adrb, twiddle_rsc_0_11_db, twiddle_rsc_0_11_web, twiddle_rsc_0_11_qb,
      twiddle_rsc_triosy_0_11_lz, twiddle_rsc_0_12_adra, twiddle_rsc_0_12_da, twiddle_rsc_0_12_wea,
      twiddle_rsc_0_12_qa, twiddle_rsc_0_12_adrb, twiddle_rsc_0_12_db, twiddle_rsc_0_12_web,
      twiddle_rsc_0_12_qb, twiddle_rsc_triosy_0_12_lz, twiddle_rsc_0_13_adra, twiddle_rsc_0_13_da,
      twiddle_rsc_0_13_wea, twiddle_rsc_0_13_qa, twiddle_rsc_0_13_adrb, twiddle_rsc_0_13_db,
      twiddle_rsc_0_13_web, twiddle_rsc_0_13_qb, twiddle_rsc_triosy_0_13_lz, twiddle_rsc_0_14_adra,
      twiddle_rsc_0_14_da, twiddle_rsc_0_14_wea, twiddle_rsc_0_14_qa, twiddle_rsc_0_14_adrb,
      twiddle_rsc_0_14_db, twiddle_rsc_0_14_web, twiddle_rsc_0_14_qb, twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_0_15_adra, twiddle_rsc_0_15_da, twiddle_rsc_0_15_wea, twiddle_rsc_0_15_qa,
      twiddle_rsc_0_15_adrb, twiddle_rsc_0_15_db, twiddle_rsc_0_15_web, twiddle_rsc_0_15_qb,
      twiddle_rsc_triosy_0_15_lz, twiddle_h_rsc_0_0_adra, twiddle_h_rsc_0_0_da, twiddle_h_rsc_0_0_wea,
      twiddle_h_rsc_0_0_qa, twiddle_h_rsc_0_0_adrb, twiddle_h_rsc_0_0_db, twiddle_h_rsc_0_0_web,
      twiddle_h_rsc_0_0_qb, twiddle_h_rsc_triosy_0_0_lz, twiddle_h_rsc_0_1_adra,
      twiddle_h_rsc_0_1_da, twiddle_h_rsc_0_1_wea, twiddle_h_rsc_0_1_qa, twiddle_h_rsc_0_1_adrb,
      twiddle_h_rsc_0_1_db, twiddle_h_rsc_0_1_web, twiddle_h_rsc_0_1_qb, twiddle_h_rsc_triosy_0_1_lz,
      twiddle_h_rsc_0_2_adra, twiddle_h_rsc_0_2_da, twiddle_h_rsc_0_2_wea, twiddle_h_rsc_0_2_qa,
      twiddle_h_rsc_0_2_adrb, twiddle_h_rsc_0_2_db, twiddle_h_rsc_0_2_web, twiddle_h_rsc_0_2_qb,
      twiddle_h_rsc_triosy_0_2_lz, twiddle_h_rsc_0_3_adra, twiddle_h_rsc_0_3_da,
      twiddle_h_rsc_0_3_wea, twiddle_h_rsc_0_3_qa, twiddle_h_rsc_0_3_adrb, twiddle_h_rsc_0_3_db,
      twiddle_h_rsc_0_3_web, twiddle_h_rsc_0_3_qb, twiddle_h_rsc_triosy_0_3_lz, twiddle_h_rsc_0_4_adra,
      twiddle_h_rsc_0_4_da, twiddle_h_rsc_0_4_wea, twiddle_h_rsc_0_4_qa, twiddle_h_rsc_0_4_adrb,
      twiddle_h_rsc_0_4_db, twiddle_h_rsc_0_4_web, twiddle_h_rsc_0_4_qb, twiddle_h_rsc_triosy_0_4_lz,
      twiddle_h_rsc_0_5_adra, twiddle_h_rsc_0_5_da, twiddle_h_rsc_0_5_wea, twiddle_h_rsc_0_5_qa,
      twiddle_h_rsc_0_5_adrb, twiddle_h_rsc_0_5_db, twiddle_h_rsc_0_5_web, twiddle_h_rsc_0_5_qb,
      twiddle_h_rsc_triosy_0_5_lz, twiddle_h_rsc_0_6_adra, twiddle_h_rsc_0_6_da,
      twiddle_h_rsc_0_6_wea, twiddle_h_rsc_0_6_qa, twiddle_h_rsc_0_6_adrb, twiddle_h_rsc_0_6_db,
      twiddle_h_rsc_0_6_web, twiddle_h_rsc_0_6_qb, twiddle_h_rsc_triosy_0_6_lz, twiddle_h_rsc_0_7_adra,
      twiddle_h_rsc_0_7_da, twiddle_h_rsc_0_7_wea, twiddle_h_rsc_0_7_qa, twiddle_h_rsc_0_7_adrb,
      twiddle_h_rsc_0_7_db, twiddle_h_rsc_0_7_web, twiddle_h_rsc_0_7_qb, twiddle_h_rsc_triosy_0_7_lz,
      twiddle_h_rsc_0_8_adra, twiddle_h_rsc_0_8_da, twiddle_h_rsc_0_8_wea, twiddle_h_rsc_0_8_qa,
      twiddle_h_rsc_0_8_adrb, twiddle_h_rsc_0_8_db, twiddle_h_rsc_0_8_web, twiddle_h_rsc_0_8_qb,
      twiddle_h_rsc_triosy_0_8_lz, twiddle_h_rsc_0_9_adra, twiddle_h_rsc_0_9_da,
      twiddle_h_rsc_0_9_wea, twiddle_h_rsc_0_9_qa, twiddle_h_rsc_0_9_adrb, twiddle_h_rsc_0_9_db,
      twiddle_h_rsc_0_9_web, twiddle_h_rsc_0_9_qb, twiddle_h_rsc_triosy_0_9_lz, twiddle_h_rsc_0_10_adra,
      twiddle_h_rsc_0_10_da, twiddle_h_rsc_0_10_wea, twiddle_h_rsc_0_10_qa, twiddle_h_rsc_0_10_adrb,
      twiddle_h_rsc_0_10_db, twiddle_h_rsc_0_10_web, twiddle_h_rsc_0_10_qb, twiddle_h_rsc_triosy_0_10_lz,
      twiddle_h_rsc_0_11_adra, twiddle_h_rsc_0_11_da, twiddle_h_rsc_0_11_wea, twiddle_h_rsc_0_11_qa,
      twiddle_h_rsc_0_11_adrb, twiddle_h_rsc_0_11_db, twiddle_h_rsc_0_11_web, twiddle_h_rsc_0_11_qb,
      twiddle_h_rsc_triosy_0_11_lz, twiddle_h_rsc_0_12_adra, twiddle_h_rsc_0_12_da,
      twiddle_h_rsc_0_12_wea, twiddle_h_rsc_0_12_qa, twiddle_h_rsc_0_12_adrb, twiddle_h_rsc_0_12_db,
      twiddle_h_rsc_0_12_web, twiddle_h_rsc_0_12_qb, twiddle_h_rsc_triosy_0_12_lz,
      twiddle_h_rsc_0_13_adra, twiddle_h_rsc_0_13_da, twiddle_h_rsc_0_13_wea, twiddle_h_rsc_0_13_qa,
      twiddle_h_rsc_0_13_adrb, twiddle_h_rsc_0_13_db, twiddle_h_rsc_0_13_web, twiddle_h_rsc_0_13_qb,
      twiddle_h_rsc_triosy_0_13_lz, twiddle_h_rsc_0_14_adra, twiddle_h_rsc_0_14_da,
      twiddle_h_rsc_0_14_wea, twiddle_h_rsc_0_14_qa, twiddle_h_rsc_0_14_adrb, twiddle_h_rsc_0_14_db,
      twiddle_h_rsc_0_14_web, twiddle_h_rsc_0_14_qb, twiddle_h_rsc_triosy_0_14_lz,
      twiddle_h_rsc_0_15_adra, twiddle_h_rsc_0_15_da, twiddle_h_rsc_0_15_wea, twiddle_h_rsc_0_15_qa,
      twiddle_h_rsc_0_15_adrb, twiddle_h_rsc_0_15_db, twiddle_h_rsc_0_15_web, twiddle_h_rsc_0_15_qb,
      twiddle_h_rsc_triosy_0_15_lz
);
  input clk;
  input rst;
  output [7:0] xt_rsc_0_0_adra;
  output [31:0] xt_rsc_0_0_da;
  output xt_rsc_0_0_wea;
  input [31:0] xt_rsc_0_0_qa;
  output [7:0] xt_rsc_0_0_adrb;
  output [31:0] xt_rsc_0_0_db;
  output xt_rsc_0_0_web;
  input [31:0] xt_rsc_0_0_qb;
  output xt_rsc_triosy_0_0_lz;
  output [7:0] xt_rsc_0_1_adra;
  output [31:0] xt_rsc_0_1_da;
  output xt_rsc_0_1_wea;
  input [31:0] xt_rsc_0_1_qa;
  output [7:0] xt_rsc_0_1_adrb;
  output [31:0] xt_rsc_0_1_db;
  output xt_rsc_0_1_web;
  input [31:0] xt_rsc_0_1_qb;
  output xt_rsc_triosy_0_1_lz;
  output [7:0] xt_rsc_0_2_adra;
  output [31:0] xt_rsc_0_2_da;
  output xt_rsc_0_2_wea;
  input [31:0] xt_rsc_0_2_qa;
  output [7:0] xt_rsc_0_2_adrb;
  output [31:0] xt_rsc_0_2_db;
  output xt_rsc_0_2_web;
  input [31:0] xt_rsc_0_2_qb;
  output xt_rsc_triosy_0_2_lz;
  output [7:0] xt_rsc_0_3_adra;
  output [31:0] xt_rsc_0_3_da;
  output xt_rsc_0_3_wea;
  input [31:0] xt_rsc_0_3_qa;
  output [7:0] xt_rsc_0_3_adrb;
  output [31:0] xt_rsc_0_3_db;
  output xt_rsc_0_3_web;
  input [31:0] xt_rsc_0_3_qb;
  output xt_rsc_triosy_0_3_lz;
  output [7:0] xt_rsc_0_4_adra;
  output [31:0] xt_rsc_0_4_da;
  output xt_rsc_0_4_wea;
  input [31:0] xt_rsc_0_4_qa;
  output [7:0] xt_rsc_0_4_adrb;
  output [31:0] xt_rsc_0_4_db;
  output xt_rsc_0_4_web;
  input [31:0] xt_rsc_0_4_qb;
  output xt_rsc_triosy_0_4_lz;
  output [7:0] xt_rsc_0_5_adra;
  output [31:0] xt_rsc_0_5_da;
  output xt_rsc_0_5_wea;
  input [31:0] xt_rsc_0_5_qa;
  output [7:0] xt_rsc_0_5_adrb;
  output [31:0] xt_rsc_0_5_db;
  output xt_rsc_0_5_web;
  input [31:0] xt_rsc_0_5_qb;
  output xt_rsc_triosy_0_5_lz;
  output [7:0] xt_rsc_0_6_adra;
  output [31:0] xt_rsc_0_6_da;
  output xt_rsc_0_6_wea;
  input [31:0] xt_rsc_0_6_qa;
  output [7:0] xt_rsc_0_6_adrb;
  output [31:0] xt_rsc_0_6_db;
  output xt_rsc_0_6_web;
  input [31:0] xt_rsc_0_6_qb;
  output xt_rsc_triosy_0_6_lz;
  output [7:0] xt_rsc_0_7_adra;
  output [31:0] xt_rsc_0_7_da;
  output xt_rsc_0_7_wea;
  input [31:0] xt_rsc_0_7_qa;
  output [7:0] xt_rsc_0_7_adrb;
  output [31:0] xt_rsc_0_7_db;
  output xt_rsc_0_7_web;
  input [31:0] xt_rsc_0_7_qb;
  output xt_rsc_triosy_0_7_lz;
  output [7:0] xt_rsc_0_8_adra;
  output [31:0] xt_rsc_0_8_da;
  output xt_rsc_0_8_wea;
  input [31:0] xt_rsc_0_8_qa;
  output [7:0] xt_rsc_0_8_adrb;
  output [31:0] xt_rsc_0_8_db;
  output xt_rsc_0_8_web;
  input [31:0] xt_rsc_0_8_qb;
  output xt_rsc_triosy_0_8_lz;
  output [7:0] xt_rsc_0_9_adra;
  output [31:0] xt_rsc_0_9_da;
  output xt_rsc_0_9_wea;
  input [31:0] xt_rsc_0_9_qa;
  output [7:0] xt_rsc_0_9_adrb;
  output [31:0] xt_rsc_0_9_db;
  output xt_rsc_0_9_web;
  input [31:0] xt_rsc_0_9_qb;
  output xt_rsc_triosy_0_9_lz;
  output [7:0] xt_rsc_0_10_adra;
  output [31:0] xt_rsc_0_10_da;
  output xt_rsc_0_10_wea;
  input [31:0] xt_rsc_0_10_qa;
  output [7:0] xt_rsc_0_10_adrb;
  output [31:0] xt_rsc_0_10_db;
  output xt_rsc_0_10_web;
  input [31:0] xt_rsc_0_10_qb;
  output xt_rsc_triosy_0_10_lz;
  output [7:0] xt_rsc_0_11_adra;
  output [31:0] xt_rsc_0_11_da;
  output xt_rsc_0_11_wea;
  input [31:0] xt_rsc_0_11_qa;
  output [7:0] xt_rsc_0_11_adrb;
  output [31:0] xt_rsc_0_11_db;
  output xt_rsc_0_11_web;
  input [31:0] xt_rsc_0_11_qb;
  output xt_rsc_triosy_0_11_lz;
  output [7:0] xt_rsc_0_12_adra;
  output [31:0] xt_rsc_0_12_da;
  output xt_rsc_0_12_wea;
  input [31:0] xt_rsc_0_12_qa;
  output [7:0] xt_rsc_0_12_adrb;
  output [31:0] xt_rsc_0_12_db;
  output xt_rsc_0_12_web;
  input [31:0] xt_rsc_0_12_qb;
  output xt_rsc_triosy_0_12_lz;
  output [7:0] xt_rsc_0_13_adra;
  output [31:0] xt_rsc_0_13_da;
  output xt_rsc_0_13_wea;
  input [31:0] xt_rsc_0_13_qa;
  output [7:0] xt_rsc_0_13_adrb;
  output [31:0] xt_rsc_0_13_db;
  output xt_rsc_0_13_web;
  input [31:0] xt_rsc_0_13_qb;
  output xt_rsc_triosy_0_13_lz;
  output [7:0] xt_rsc_0_14_adra;
  output [31:0] xt_rsc_0_14_da;
  output xt_rsc_0_14_wea;
  input [31:0] xt_rsc_0_14_qa;
  output [7:0] xt_rsc_0_14_adrb;
  output [31:0] xt_rsc_0_14_db;
  output xt_rsc_0_14_web;
  input [31:0] xt_rsc_0_14_qb;
  output xt_rsc_triosy_0_14_lz;
  output [7:0] xt_rsc_0_15_adra;
  output [31:0] xt_rsc_0_15_da;
  output xt_rsc_0_15_wea;
  input [31:0] xt_rsc_0_15_qa;
  output [7:0] xt_rsc_0_15_adrb;
  output [31:0] xt_rsc_0_15_db;
  output xt_rsc_0_15_web;
  input [31:0] xt_rsc_0_15_qb;
  output xt_rsc_triosy_0_15_lz;
  output [7:0] xt_rsc_0_16_adra;
  output [31:0] xt_rsc_0_16_da;
  output xt_rsc_0_16_wea;
  input [31:0] xt_rsc_0_16_qa;
  output [7:0] xt_rsc_0_16_adrb;
  output [31:0] xt_rsc_0_16_db;
  output xt_rsc_0_16_web;
  input [31:0] xt_rsc_0_16_qb;
  output xt_rsc_triosy_0_16_lz;
  output [7:0] xt_rsc_0_17_adra;
  output [31:0] xt_rsc_0_17_da;
  output xt_rsc_0_17_wea;
  input [31:0] xt_rsc_0_17_qa;
  output [7:0] xt_rsc_0_17_adrb;
  output [31:0] xt_rsc_0_17_db;
  output xt_rsc_0_17_web;
  input [31:0] xt_rsc_0_17_qb;
  output xt_rsc_triosy_0_17_lz;
  output [7:0] xt_rsc_0_18_adra;
  output [31:0] xt_rsc_0_18_da;
  output xt_rsc_0_18_wea;
  input [31:0] xt_rsc_0_18_qa;
  output [7:0] xt_rsc_0_18_adrb;
  output [31:0] xt_rsc_0_18_db;
  output xt_rsc_0_18_web;
  input [31:0] xt_rsc_0_18_qb;
  output xt_rsc_triosy_0_18_lz;
  output [7:0] xt_rsc_0_19_adra;
  output [31:0] xt_rsc_0_19_da;
  output xt_rsc_0_19_wea;
  input [31:0] xt_rsc_0_19_qa;
  output [7:0] xt_rsc_0_19_adrb;
  output [31:0] xt_rsc_0_19_db;
  output xt_rsc_0_19_web;
  input [31:0] xt_rsc_0_19_qb;
  output xt_rsc_triosy_0_19_lz;
  output [7:0] xt_rsc_0_20_adra;
  output [31:0] xt_rsc_0_20_da;
  output xt_rsc_0_20_wea;
  input [31:0] xt_rsc_0_20_qa;
  output [7:0] xt_rsc_0_20_adrb;
  output [31:0] xt_rsc_0_20_db;
  output xt_rsc_0_20_web;
  input [31:0] xt_rsc_0_20_qb;
  output xt_rsc_triosy_0_20_lz;
  output [7:0] xt_rsc_0_21_adra;
  output [31:0] xt_rsc_0_21_da;
  output xt_rsc_0_21_wea;
  input [31:0] xt_rsc_0_21_qa;
  output [7:0] xt_rsc_0_21_adrb;
  output [31:0] xt_rsc_0_21_db;
  output xt_rsc_0_21_web;
  input [31:0] xt_rsc_0_21_qb;
  output xt_rsc_triosy_0_21_lz;
  output [7:0] xt_rsc_0_22_adra;
  output [31:0] xt_rsc_0_22_da;
  output xt_rsc_0_22_wea;
  input [31:0] xt_rsc_0_22_qa;
  output [7:0] xt_rsc_0_22_adrb;
  output [31:0] xt_rsc_0_22_db;
  output xt_rsc_0_22_web;
  input [31:0] xt_rsc_0_22_qb;
  output xt_rsc_triosy_0_22_lz;
  output [7:0] xt_rsc_0_23_adra;
  output [31:0] xt_rsc_0_23_da;
  output xt_rsc_0_23_wea;
  input [31:0] xt_rsc_0_23_qa;
  output [7:0] xt_rsc_0_23_adrb;
  output [31:0] xt_rsc_0_23_db;
  output xt_rsc_0_23_web;
  input [31:0] xt_rsc_0_23_qb;
  output xt_rsc_triosy_0_23_lz;
  output [7:0] xt_rsc_0_24_adra;
  output [31:0] xt_rsc_0_24_da;
  output xt_rsc_0_24_wea;
  input [31:0] xt_rsc_0_24_qa;
  output [7:0] xt_rsc_0_24_adrb;
  output [31:0] xt_rsc_0_24_db;
  output xt_rsc_0_24_web;
  input [31:0] xt_rsc_0_24_qb;
  output xt_rsc_triosy_0_24_lz;
  output [7:0] xt_rsc_0_25_adra;
  output [31:0] xt_rsc_0_25_da;
  output xt_rsc_0_25_wea;
  input [31:0] xt_rsc_0_25_qa;
  output [7:0] xt_rsc_0_25_adrb;
  output [31:0] xt_rsc_0_25_db;
  output xt_rsc_0_25_web;
  input [31:0] xt_rsc_0_25_qb;
  output xt_rsc_triosy_0_25_lz;
  output [7:0] xt_rsc_0_26_adra;
  output [31:0] xt_rsc_0_26_da;
  output xt_rsc_0_26_wea;
  input [31:0] xt_rsc_0_26_qa;
  output [7:0] xt_rsc_0_26_adrb;
  output [31:0] xt_rsc_0_26_db;
  output xt_rsc_0_26_web;
  input [31:0] xt_rsc_0_26_qb;
  output xt_rsc_triosy_0_26_lz;
  output [7:0] xt_rsc_0_27_adra;
  output [31:0] xt_rsc_0_27_da;
  output xt_rsc_0_27_wea;
  input [31:0] xt_rsc_0_27_qa;
  output [7:0] xt_rsc_0_27_adrb;
  output [31:0] xt_rsc_0_27_db;
  output xt_rsc_0_27_web;
  input [31:0] xt_rsc_0_27_qb;
  output xt_rsc_triosy_0_27_lz;
  output [7:0] xt_rsc_0_28_adra;
  output [31:0] xt_rsc_0_28_da;
  output xt_rsc_0_28_wea;
  input [31:0] xt_rsc_0_28_qa;
  output [7:0] xt_rsc_0_28_adrb;
  output [31:0] xt_rsc_0_28_db;
  output xt_rsc_0_28_web;
  input [31:0] xt_rsc_0_28_qb;
  output xt_rsc_triosy_0_28_lz;
  output [7:0] xt_rsc_0_29_adra;
  output [31:0] xt_rsc_0_29_da;
  output xt_rsc_0_29_wea;
  input [31:0] xt_rsc_0_29_qa;
  output [7:0] xt_rsc_0_29_adrb;
  output [31:0] xt_rsc_0_29_db;
  output xt_rsc_0_29_web;
  input [31:0] xt_rsc_0_29_qb;
  output xt_rsc_triosy_0_29_lz;
  output [7:0] xt_rsc_0_30_adra;
  output [31:0] xt_rsc_0_30_da;
  output xt_rsc_0_30_wea;
  input [31:0] xt_rsc_0_30_qa;
  output [7:0] xt_rsc_0_30_adrb;
  output [31:0] xt_rsc_0_30_db;
  output xt_rsc_0_30_web;
  input [31:0] xt_rsc_0_30_qb;
  output xt_rsc_triosy_0_30_lz;
  output [7:0] xt_rsc_0_31_adra;
  output [31:0] xt_rsc_0_31_da;
  output xt_rsc_0_31_wea;
  input [31:0] xt_rsc_0_31_qa;
  output [7:0] xt_rsc_0_31_adrb;
  output [31:0] xt_rsc_0_31_db;
  output xt_rsc_0_31_web;
  input [31:0] xt_rsc_0_31_qb;
  output xt_rsc_triosy_0_31_lz;
  input [31:0] p_rsc_dat;
  output p_rsc_triosy_lz;
  input [31:0] r_rsc_dat;
  output r_rsc_triosy_lz;
  output [7:0] twiddle_rsc_0_0_adra;
  output [31:0] twiddle_rsc_0_0_da;
  output twiddle_rsc_0_0_wea;
  input [31:0] twiddle_rsc_0_0_qa;
  output [7:0] twiddle_rsc_0_0_adrb;
  output [31:0] twiddle_rsc_0_0_db;
  output twiddle_rsc_0_0_web;
  input [31:0] twiddle_rsc_0_0_qb;
  output twiddle_rsc_triosy_0_0_lz;
  output [7:0] twiddle_rsc_0_1_adra;
  output [31:0] twiddle_rsc_0_1_da;
  output twiddle_rsc_0_1_wea;
  input [31:0] twiddle_rsc_0_1_qa;
  output [7:0] twiddle_rsc_0_1_adrb;
  output [31:0] twiddle_rsc_0_1_db;
  output twiddle_rsc_0_1_web;
  input [31:0] twiddle_rsc_0_1_qb;
  output twiddle_rsc_triosy_0_1_lz;
  output [7:0] twiddle_rsc_0_2_adra;
  output [31:0] twiddle_rsc_0_2_da;
  output twiddle_rsc_0_2_wea;
  input [31:0] twiddle_rsc_0_2_qa;
  output [7:0] twiddle_rsc_0_2_adrb;
  output [31:0] twiddle_rsc_0_2_db;
  output twiddle_rsc_0_2_web;
  input [31:0] twiddle_rsc_0_2_qb;
  output twiddle_rsc_triosy_0_2_lz;
  output [7:0] twiddle_rsc_0_3_adra;
  output [31:0] twiddle_rsc_0_3_da;
  output twiddle_rsc_0_3_wea;
  input [31:0] twiddle_rsc_0_3_qa;
  output [7:0] twiddle_rsc_0_3_adrb;
  output [31:0] twiddle_rsc_0_3_db;
  output twiddle_rsc_0_3_web;
  input [31:0] twiddle_rsc_0_3_qb;
  output twiddle_rsc_triosy_0_3_lz;
  output [7:0] twiddle_rsc_0_4_adra;
  output [31:0] twiddle_rsc_0_4_da;
  output twiddle_rsc_0_4_wea;
  input [31:0] twiddle_rsc_0_4_qa;
  output [7:0] twiddle_rsc_0_4_adrb;
  output [31:0] twiddle_rsc_0_4_db;
  output twiddle_rsc_0_4_web;
  input [31:0] twiddle_rsc_0_4_qb;
  output twiddle_rsc_triosy_0_4_lz;
  output [7:0] twiddle_rsc_0_5_adra;
  output [31:0] twiddle_rsc_0_5_da;
  output twiddle_rsc_0_5_wea;
  input [31:0] twiddle_rsc_0_5_qa;
  output [7:0] twiddle_rsc_0_5_adrb;
  output [31:0] twiddle_rsc_0_5_db;
  output twiddle_rsc_0_5_web;
  input [31:0] twiddle_rsc_0_5_qb;
  output twiddle_rsc_triosy_0_5_lz;
  output [7:0] twiddle_rsc_0_6_adra;
  output [31:0] twiddle_rsc_0_6_da;
  output twiddle_rsc_0_6_wea;
  input [31:0] twiddle_rsc_0_6_qa;
  output [7:0] twiddle_rsc_0_6_adrb;
  output [31:0] twiddle_rsc_0_6_db;
  output twiddle_rsc_0_6_web;
  input [31:0] twiddle_rsc_0_6_qb;
  output twiddle_rsc_triosy_0_6_lz;
  output [7:0] twiddle_rsc_0_7_adra;
  output [31:0] twiddle_rsc_0_7_da;
  output twiddle_rsc_0_7_wea;
  input [31:0] twiddle_rsc_0_7_qa;
  output [7:0] twiddle_rsc_0_7_adrb;
  output [31:0] twiddle_rsc_0_7_db;
  output twiddle_rsc_0_7_web;
  input [31:0] twiddle_rsc_0_7_qb;
  output twiddle_rsc_triosy_0_7_lz;
  output [7:0] twiddle_rsc_0_8_adra;
  output [31:0] twiddle_rsc_0_8_da;
  output twiddle_rsc_0_8_wea;
  input [31:0] twiddle_rsc_0_8_qa;
  output [7:0] twiddle_rsc_0_8_adrb;
  output [31:0] twiddle_rsc_0_8_db;
  output twiddle_rsc_0_8_web;
  input [31:0] twiddle_rsc_0_8_qb;
  output twiddle_rsc_triosy_0_8_lz;
  output [7:0] twiddle_rsc_0_9_adra;
  output [31:0] twiddle_rsc_0_9_da;
  output twiddle_rsc_0_9_wea;
  input [31:0] twiddle_rsc_0_9_qa;
  output [7:0] twiddle_rsc_0_9_adrb;
  output [31:0] twiddle_rsc_0_9_db;
  output twiddle_rsc_0_9_web;
  input [31:0] twiddle_rsc_0_9_qb;
  output twiddle_rsc_triosy_0_9_lz;
  output [7:0] twiddle_rsc_0_10_adra;
  output [31:0] twiddle_rsc_0_10_da;
  output twiddle_rsc_0_10_wea;
  input [31:0] twiddle_rsc_0_10_qa;
  output [7:0] twiddle_rsc_0_10_adrb;
  output [31:0] twiddle_rsc_0_10_db;
  output twiddle_rsc_0_10_web;
  input [31:0] twiddle_rsc_0_10_qb;
  output twiddle_rsc_triosy_0_10_lz;
  output [7:0] twiddle_rsc_0_11_adra;
  output [31:0] twiddle_rsc_0_11_da;
  output twiddle_rsc_0_11_wea;
  input [31:0] twiddle_rsc_0_11_qa;
  output [7:0] twiddle_rsc_0_11_adrb;
  output [31:0] twiddle_rsc_0_11_db;
  output twiddle_rsc_0_11_web;
  input [31:0] twiddle_rsc_0_11_qb;
  output twiddle_rsc_triosy_0_11_lz;
  output [7:0] twiddle_rsc_0_12_adra;
  output [31:0] twiddle_rsc_0_12_da;
  output twiddle_rsc_0_12_wea;
  input [31:0] twiddle_rsc_0_12_qa;
  output [7:0] twiddle_rsc_0_12_adrb;
  output [31:0] twiddle_rsc_0_12_db;
  output twiddle_rsc_0_12_web;
  input [31:0] twiddle_rsc_0_12_qb;
  output twiddle_rsc_triosy_0_12_lz;
  output [7:0] twiddle_rsc_0_13_adra;
  output [31:0] twiddle_rsc_0_13_da;
  output twiddle_rsc_0_13_wea;
  input [31:0] twiddle_rsc_0_13_qa;
  output [7:0] twiddle_rsc_0_13_adrb;
  output [31:0] twiddle_rsc_0_13_db;
  output twiddle_rsc_0_13_web;
  input [31:0] twiddle_rsc_0_13_qb;
  output twiddle_rsc_triosy_0_13_lz;
  output [7:0] twiddle_rsc_0_14_adra;
  output [31:0] twiddle_rsc_0_14_da;
  output twiddle_rsc_0_14_wea;
  input [31:0] twiddle_rsc_0_14_qa;
  output [7:0] twiddle_rsc_0_14_adrb;
  output [31:0] twiddle_rsc_0_14_db;
  output twiddle_rsc_0_14_web;
  input [31:0] twiddle_rsc_0_14_qb;
  output twiddle_rsc_triosy_0_14_lz;
  output [7:0] twiddle_rsc_0_15_adra;
  output [31:0] twiddle_rsc_0_15_da;
  output twiddle_rsc_0_15_wea;
  input [31:0] twiddle_rsc_0_15_qa;
  output [7:0] twiddle_rsc_0_15_adrb;
  output [31:0] twiddle_rsc_0_15_db;
  output twiddle_rsc_0_15_web;
  input [31:0] twiddle_rsc_0_15_qb;
  output twiddle_rsc_triosy_0_15_lz;
  output [7:0] twiddle_h_rsc_0_0_adra;
  output [31:0] twiddle_h_rsc_0_0_da;
  output twiddle_h_rsc_0_0_wea;
  input [31:0] twiddle_h_rsc_0_0_qa;
  output [7:0] twiddle_h_rsc_0_0_adrb;
  output [31:0] twiddle_h_rsc_0_0_db;
  output twiddle_h_rsc_0_0_web;
  input [31:0] twiddle_h_rsc_0_0_qb;
  output twiddle_h_rsc_triosy_0_0_lz;
  output [7:0] twiddle_h_rsc_0_1_adra;
  output [31:0] twiddle_h_rsc_0_1_da;
  output twiddle_h_rsc_0_1_wea;
  input [31:0] twiddle_h_rsc_0_1_qa;
  output [7:0] twiddle_h_rsc_0_1_adrb;
  output [31:0] twiddle_h_rsc_0_1_db;
  output twiddle_h_rsc_0_1_web;
  input [31:0] twiddle_h_rsc_0_1_qb;
  output twiddle_h_rsc_triosy_0_1_lz;
  output [7:0] twiddle_h_rsc_0_2_adra;
  output [31:0] twiddle_h_rsc_0_2_da;
  output twiddle_h_rsc_0_2_wea;
  input [31:0] twiddle_h_rsc_0_2_qa;
  output [7:0] twiddle_h_rsc_0_2_adrb;
  output [31:0] twiddle_h_rsc_0_2_db;
  output twiddle_h_rsc_0_2_web;
  input [31:0] twiddle_h_rsc_0_2_qb;
  output twiddle_h_rsc_triosy_0_2_lz;
  output [7:0] twiddle_h_rsc_0_3_adra;
  output [31:0] twiddle_h_rsc_0_3_da;
  output twiddle_h_rsc_0_3_wea;
  input [31:0] twiddle_h_rsc_0_3_qa;
  output [7:0] twiddle_h_rsc_0_3_adrb;
  output [31:0] twiddle_h_rsc_0_3_db;
  output twiddle_h_rsc_0_3_web;
  input [31:0] twiddle_h_rsc_0_3_qb;
  output twiddle_h_rsc_triosy_0_3_lz;
  output [7:0] twiddle_h_rsc_0_4_adra;
  output [31:0] twiddle_h_rsc_0_4_da;
  output twiddle_h_rsc_0_4_wea;
  input [31:0] twiddle_h_rsc_0_4_qa;
  output [7:0] twiddle_h_rsc_0_4_adrb;
  output [31:0] twiddle_h_rsc_0_4_db;
  output twiddle_h_rsc_0_4_web;
  input [31:0] twiddle_h_rsc_0_4_qb;
  output twiddle_h_rsc_triosy_0_4_lz;
  output [7:0] twiddle_h_rsc_0_5_adra;
  output [31:0] twiddle_h_rsc_0_5_da;
  output twiddle_h_rsc_0_5_wea;
  input [31:0] twiddle_h_rsc_0_5_qa;
  output [7:0] twiddle_h_rsc_0_5_adrb;
  output [31:0] twiddle_h_rsc_0_5_db;
  output twiddle_h_rsc_0_5_web;
  input [31:0] twiddle_h_rsc_0_5_qb;
  output twiddle_h_rsc_triosy_0_5_lz;
  output [7:0] twiddle_h_rsc_0_6_adra;
  output [31:0] twiddle_h_rsc_0_6_da;
  output twiddle_h_rsc_0_6_wea;
  input [31:0] twiddle_h_rsc_0_6_qa;
  output [7:0] twiddle_h_rsc_0_6_adrb;
  output [31:0] twiddle_h_rsc_0_6_db;
  output twiddle_h_rsc_0_6_web;
  input [31:0] twiddle_h_rsc_0_6_qb;
  output twiddle_h_rsc_triosy_0_6_lz;
  output [7:0] twiddle_h_rsc_0_7_adra;
  output [31:0] twiddle_h_rsc_0_7_da;
  output twiddle_h_rsc_0_7_wea;
  input [31:0] twiddle_h_rsc_0_7_qa;
  output [7:0] twiddle_h_rsc_0_7_adrb;
  output [31:0] twiddle_h_rsc_0_7_db;
  output twiddle_h_rsc_0_7_web;
  input [31:0] twiddle_h_rsc_0_7_qb;
  output twiddle_h_rsc_triosy_0_7_lz;
  output [7:0] twiddle_h_rsc_0_8_adra;
  output [31:0] twiddle_h_rsc_0_8_da;
  output twiddle_h_rsc_0_8_wea;
  input [31:0] twiddle_h_rsc_0_8_qa;
  output [7:0] twiddle_h_rsc_0_8_adrb;
  output [31:0] twiddle_h_rsc_0_8_db;
  output twiddle_h_rsc_0_8_web;
  input [31:0] twiddle_h_rsc_0_8_qb;
  output twiddle_h_rsc_triosy_0_8_lz;
  output [7:0] twiddle_h_rsc_0_9_adra;
  output [31:0] twiddle_h_rsc_0_9_da;
  output twiddle_h_rsc_0_9_wea;
  input [31:0] twiddle_h_rsc_0_9_qa;
  output [7:0] twiddle_h_rsc_0_9_adrb;
  output [31:0] twiddle_h_rsc_0_9_db;
  output twiddle_h_rsc_0_9_web;
  input [31:0] twiddle_h_rsc_0_9_qb;
  output twiddle_h_rsc_triosy_0_9_lz;
  output [7:0] twiddle_h_rsc_0_10_adra;
  output [31:0] twiddle_h_rsc_0_10_da;
  output twiddle_h_rsc_0_10_wea;
  input [31:0] twiddle_h_rsc_0_10_qa;
  output [7:0] twiddle_h_rsc_0_10_adrb;
  output [31:0] twiddle_h_rsc_0_10_db;
  output twiddle_h_rsc_0_10_web;
  input [31:0] twiddle_h_rsc_0_10_qb;
  output twiddle_h_rsc_triosy_0_10_lz;
  output [7:0] twiddle_h_rsc_0_11_adra;
  output [31:0] twiddle_h_rsc_0_11_da;
  output twiddle_h_rsc_0_11_wea;
  input [31:0] twiddle_h_rsc_0_11_qa;
  output [7:0] twiddle_h_rsc_0_11_adrb;
  output [31:0] twiddle_h_rsc_0_11_db;
  output twiddle_h_rsc_0_11_web;
  input [31:0] twiddle_h_rsc_0_11_qb;
  output twiddle_h_rsc_triosy_0_11_lz;
  output [7:0] twiddle_h_rsc_0_12_adra;
  output [31:0] twiddle_h_rsc_0_12_da;
  output twiddle_h_rsc_0_12_wea;
  input [31:0] twiddle_h_rsc_0_12_qa;
  output [7:0] twiddle_h_rsc_0_12_adrb;
  output [31:0] twiddle_h_rsc_0_12_db;
  output twiddle_h_rsc_0_12_web;
  input [31:0] twiddle_h_rsc_0_12_qb;
  output twiddle_h_rsc_triosy_0_12_lz;
  output [7:0] twiddle_h_rsc_0_13_adra;
  output [31:0] twiddle_h_rsc_0_13_da;
  output twiddle_h_rsc_0_13_wea;
  input [31:0] twiddle_h_rsc_0_13_qa;
  output [7:0] twiddle_h_rsc_0_13_adrb;
  output [31:0] twiddle_h_rsc_0_13_db;
  output twiddle_h_rsc_0_13_web;
  input [31:0] twiddle_h_rsc_0_13_qb;
  output twiddle_h_rsc_triosy_0_13_lz;
  output [7:0] twiddle_h_rsc_0_14_adra;
  output [31:0] twiddle_h_rsc_0_14_da;
  output twiddle_h_rsc_0_14_wea;
  input [31:0] twiddle_h_rsc_0_14_qa;
  output [7:0] twiddle_h_rsc_0_14_adrb;
  output [31:0] twiddle_h_rsc_0_14_db;
  output twiddle_h_rsc_0_14_web;
  input [31:0] twiddle_h_rsc_0_14_qb;
  output twiddle_h_rsc_triosy_0_14_lz;
  output [7:0] twiddle_h_rsc_0_15_adra;
  output [31:0] twiddle_h_rsc_0_15_da;
  output twiddle_h_rsc_0_15_wea;
  input [31:0] twiddle_h_rsc_0_15_qa;
  output [7:0] twiddle_h_rsc_0_15_adrb;
  output [31:0] twiddle_h_rsc_0_15_db;
  output twiddle_h_rsc_0_15_web;
  input [31:0] twiddle_h_rsc_0_15_qb;
  output twiddle_h_rsc_triosy_0_15_lz;


  // Interconnect Declarations
  wire [15:0] yt_rsc_0_0_i_adra_d;
  wire yt_rsc_0_0_i_clka_en_d;
  wire [63:0] yt_rsc_0_0_i_da_d;
  wire [63:0] yt_rsc_0_0_i_qa_d;
  wire [1:0] yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_1_i_adra_d;
  wire [63:0] yt_rsc_0_1_i_da_d;
  wire [63:0] yt_rsc_0_1_i_qa_d;
  wire [1:0] yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_2_i_adra_d;
  wire [63:0] yt_rsc_0_2_i_da_d;
  wire [63:0] yt_rsc_0_2_i_qa_d;
  wire [1:0] yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_3_i_adra_d;
  wire [63:0] yt_rsc_0_3_i_da_d;
  wire [63:0] yt_rsc_0_3_i_qa_d;
  wire [1:0] yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_4_i_adra_d;
  wire [63:0] yt_rsc_0_4_i_da_d;
  wire [63:0] yt_rsc_0_4_i_qa_d;
  wire [1:0] yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_5_i_adra_d;
  wire [63:0] yt_rsc_0_5_i_da_d;
  wire [63:0] yt_rsc_0_5_i_qa_d;
  wire [1:0] yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_6_i_adra_d;
  wire [63:0] yt_rsc_0_6_i_da_d;
  wire [63:0] yt_rsc_0_6_i_qa_d;
  wire [1:0] yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_7_i_adra_d;
  wire [63:0] yt_rsc_0_7_i_da_d;
  wire [63:0] yt_rsc_0_7_i_qa_d;
  wire [1:0] yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_8_i_adra_d;
  wire [63:0] yt_rsc_0_8_i_da_d;
  wire [63:0] yt_rsc_0_8_i_qa_d;
  wire [1:0] yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_9_i_adra_d;
  wire [63:0] yt_rsc_0_9_i_da_d;
  wire [63:0] yt_rsc_0_9_i_qa_d;
  wire [1:0] yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_10_i_adra_d;
  wire [63:0] yt_rsc_0_10_i_da_d;
  wire [63:0] yt_rsc_0_10_i_qa_d;
  wire [1:0] yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_11_i_adra_d;
  wire [63:0] yt_rsc_0_11_i_da_d;
  wire [63:0] yt_rsc_0_11_i_qa_d;
  wire [1:0] yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_12_i_adra_d;
  wire [63:0] yt_rsc_0_12_i_da_d;
  wire [63:0] yt_rsc_0_12_i_qa_d;
  wire [1:0] yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_13_i_adra_d;
  wire [63:0] yt_rsc_0_13_i_da_d;
  wire [63:0] yt_rsc_0_13_i_qa_d;
  wire [1:0] yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_14_i_adra_d;
  wire [63:0] yt_rsc_0_14_i_da_d;
  wire [63:0] yt_rsc_0_14_i_qa_d;
  wire [1:0] yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_15_i_adra_d;
  wire [63:0] yt_rsc_0_15_i_da_d;
  wire [63:0] yt_rsc_0_15_i_qa_d;
  wire [1:0] yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_16_i_adra_d;
  wire yt_rsc_0_16_i_clka_en_d;
  wire [63:0] yt_rsc_0_16_i_da_d;
  wire [63:0] yt_rsc_0_16_i_qa_d;
  wire [1:0] yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_17_i_adra_d;
  wire [63:0] yt_rsc_0_17_i_da_d;
  wire [63:0] yt_rsc_0_17_i_qa_d;
  wire [1:0] yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_18_i_adra_d;
  wire [63:0] yt_rsc_0_18_i_da_d;
  wire [63:0] yt_rsc_0_18_i_qa_d;
  wire [1:0] yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_19_i_adra_d;
  wire [63:0] yt_rsc_0_19_i_da_d;
  wire [63:0] yt_rsc_0_19_i_qa_d;
  wire [1:0] yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_20_i_adra_d;
  wire [63:0] yt_rsc_0_20_i_da_d;
  wire [63:0] yt_rsc_0_20_i_qa_d;
  wire [1:0] yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_21_i_adra_d;
  wire [63:0] yt_rsc_0_21_i_da_d;
  wire [63:0] yt_rsc_0_21_i_qa_d;
  wire [1:0] yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_22_i_adra_d;
  wire [63:0] yt_rsc_0_22_i_da_d;
  wire [63:0] yt_rsc_0_22_i_qa_d;
  wire [1:0] yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_23_i_adra_d;
  wire [63:0] yt_rsc_0_23_i_da_d;
  wire [63:0] yt_rsc_0_23_i_qa_d;
  wire [1:0] yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_24_i_adra_d;
  wire [63:0] yt_rsc_0_24_i_da_d;
  wire [63:0] yt_rsc_0_24_i_qa_d;
  wire [1:0] yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_25_i_adra_d;
  wire [63:0] yt_rsc_0_25_i_da_d;
  wire [63:0] yt_rsc_0_25_i_qa_d;
  wire [1:0] yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_26_i_adra_d;
  wire [63:0] yt_rsc_0_26_i_da_d;
  wire [63:0] yt_rsc_0_26_i_qa_d;
  wire [1:0] yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_27_i_adra_d;
  wire [63:0] yt_rsc_0_27_i_da_d;
  wire [63:0] yt_rsc_0_27_i_qa_d;
  wire [1:0] yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_28_i_adra_d;
  wire [63:0] yt_rsc_0_28_i_da_d;
  wire [63:0] yt_rsc_0_28_i_qa_d;
  wire [1:0] yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_29_i_adra_d;
  wire [63:0] yt_rsc_0_29_i_da_d;
  wire [63:0] yt_rsc_0_29_i_qa_d;
  wire [1:0] yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_30_i_adra_d;
  wire [63:0] yt_rsc_0_30_i_da_d;
  wire [63:0] yt_rsc_0_30_i_qa_d;
  wire [1:0] yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] yt_rsc_0_31_i_adra_d;
  wire [63:0] yt_rsc_0_31_i_da_d;
  wire [63:0] yt_rsc_0_31_i_qa_d;
  wire [1:0] yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_0_i_adra_d;
  wire [63:0] xt_rsc_0_0_i_da_d;
  wire [63:0] xt_rsc_0_0_i_qa_d;
  wire [1:0] xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_1_i_adra_d;
  wire [63:0] xt_rsc_0_1_i_da_d;
  wire [63:0] xt_rsc_0_1_i_qa_d;
  wire [1:0] xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_2_i_adra_d;
  wire [63:0] xt_rsc_0_2_i_da_d;
  wire [63:0] xt_rsc_0_2_i_qa_d;
  wire [1:0] xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_3_i_adra_d;
  wire [63:0] xt_rsc_0_3_i_da_d;
  wire [63:0] xt_rsc_0_3_i_qa_d;
  wire [1:0] xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_4_i_adra_d;
  wire [63:0] xt_rsc_0_4_i_da_d;
  wire [63:0] xt_rsc_0_4_i_qa_d;
  wire [1:0] xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_5_i_adra_d;
  wire [63:0] xt_rsc_0_5_i_da_d;
  wire [63:0] xt_rsc_0_5_i_qa_d;
  wire [1:0] xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_6_i_adra_d;
  wire [63:0] xt_rsc_0_6_i_da_d;
  wire [63:0] xt_rsc_0_6_i_qa_d;
  wire [1:0] xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_7_i_adra_d;
  wire [63:0] xt_rsc_0_7_i_da_d;
  wire [63:0] xt_rsc_0_7_i_qa_d;
  wire [1:0] xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_8_i_adra_d;
  wire [63:0] xt_rsc_0_8_i_da_d;
  wire [63:0] xt_rsc_0_8_i_qa_d;
  wire [1:0] xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_9_i_adra_d;
  wire [63:0] xt_rsc_0_9_i_da_d;
  wire [63:0] xt_rsc_0_9_i_qa_d;
  wire [1:0] xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_10_i_adra_d;
  wire [63:0] xt_rsc_0_10_i_da_d;
  wire [63:0] xt_rsc_0_10_i_qa_d;
  wire [1:0] xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_11_i_adra_d;
  wire [63:0] xt_rsc_0_11_i_da_d;
  wire [63:0] xt_rsc_0_11_i_qa_d;
  wire [1:0] xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_12_i_adra_d;
  wire [63:0] xt_rsc_0_12_i_da_d;
  wire [63:0] xt_rsc_0_12_i_qa_d;
  wire [1:0] xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_13_i_adra_d;
  wire [63:0] xt_rsc_0_13_i_da_d;
  wire [63:0] xt_rsc_0_13_i_qa_d;
  wire [1:0] xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_14_i_adra_d;
  wire [63:0] xt_rsc_0_14_i_da_d;
  wire [63:0] xt_rsc_0_14_i_qa_d;
  wire [1:0] xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_15_i_adra_d;
  wire [63:0] xt_rsc_0_15_i_da_d;
  wire [63:0] xt_rsc_0_15_i_qa_d;
  wire [1:0] xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_16_i_adra_d;
  wire [63:0] xt_rsc_0_16_i_da_d;
  wire [63:0] xt_rsc_0_16_i_qa_d;
  wire [1:0] xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_17_i_adra_d;
  wire [63:0] xt_rsc_0_17_i_da_d;
  wire [63:0] xt_rsc_0_17_i_qa_d;
  wire [1:0] xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_18_i_adra_d;
  wire [63:0] xt_rsc_0_18_i_da_d;
  wire [63:0] xt_rsc_0_18_i_qa_d;
  wire [1:0] xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_19_i_adra_d;
  wire [63:0] xt_rsc_0_19_i_da_d;
  wire [63:0] xt_rsc_0_19_i_qa_d;
  wire [1:0] xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_20_i_adra_d;
  wire [63:0] xt_rsc_0_20_i_da_d;
  wire [63:0] xt_rsc_0_20_i_qa_d;
  wire [1:0] xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_21_i_adra_d;
  wire [63:0] xt_rsc_0_21_i_da_d;
  wire [63:0] xt_rsc_0_21_i_qa_d;
  wire [1:0] xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_22_i_adra_d;
  wire [63:0] xt_rsc_0_22_i_da_d;
  wire [63:0] xt_rsc_0_22_i_qa_d;
  wire [1:0] xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_23_i_adra_d;
  wire [63:0] xt_rsc_0_23_i_da_d;
  wire [63:0] xt_rsc_0_23_i_qa_d;
  wire [1:0] xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_24_i_adra_d;
  wire [63:0] xt_rsc_0_24_i_da_d;
  wire [63:0] xt_rsc_0_24_i_qa_d;
  wire [1:0] xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_25_i_adra_d;
  wire [63:0] xt_rsc_0_25_i_da_d;
  wire [63:0] xt_rsc_0_25_i_qa_d;
  wire [1:0] xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_26_i_adra_d;
  wire [63:0] xt_rsc_0_26_i_da_d;
  wire [63:0] xt_rsc_0_26_i_qa_d;
  wire [1:0] xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_27_i_adra_d;
  wire [63:0] xt_rsc_0_27_i_da_d;
  wire [63:0] xt_rsc_0_27_i_qa_d;
  wire [1:0] xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_28_i_adra_d;
  wire [63:0] xt_rsc_0_28_i_da_d;
  wire [63:0] xt_rsc_0_28_i_qa_d;
  wire [1:0] xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_29_i_adra_d;
  wire [63:0] xt_rsc_0_29_i_da_d;
  wire [63:0] xt_rsc_0_29_i_qa_d;
  wire [1:0] xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_30_i_adra_d;
  wire [63:0] xt_rsc_0_30_i_da_d;
  wire [63:0] xt_rsc_0_30_i_qa_d;
  wire [1:0] xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [15:0] xt_rsc_0_31_i_adra_d;
  wire [63:0] xt_rsc_0_31_i_da_d;
  wire [63:0] xt_rsc_0_31_i_qa_d;
  wire [1:0] xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_0_i_adra_d;
  wire [63:0] twiddle_rsc_0_0_i_qa_d;
  wire [1:0] twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_1_i_adra_d;
  wire [63:0] twiddle_rsc_0_1_i_qa_d;
  wire [1:0] twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_2_i_adra_d;
  wire [63:0] twiddle_rsc_0_2_i_qa_d;
  wire [1:0] twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_3_i_adra_d;
  wire [63:0] twiddle_rsc_0_3_i_qa_d;
  wire [1:0] twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_4_i_adra_d;
  wire [63:0] twiddle_rsc_0_4_i_qa_d;
  wire [1:0] twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_5_i_adra_d;
  wire [63:0] twiddle_rsc_0_5_i_qa_d;
  wire [1:0] twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_6_i_adra_d;
  wire [63:0] twiddle_rsc_0_6_i_qa_d;
  wire [1:0] twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_7_i_adra_d;
  wire [63:0] twiddle_rsc_0_7_i_qa_d;
  wire [1:0] twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_8_i_adra_d;
  wire [63:0] twiddle_rsc_0_8_i_qa_d;
  wire [1:0] twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_9_i_adra_d;
  wire [63:0] twiddle_rsc_0_9_i_qa_d;
  wire [1:0] twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_10_i_adra_d;
  wire [63:0] twiddle_rsc_0_10_i_qa_d;
  wire [1:0] twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_11_i_adra_d;
  wire [63:0] twiddle_rsc_0_11_i_qa_d;
  wire [1:0] twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_12_i_adra_d;
  wire [63:0] twiddle_rsc_0_12_i_qa_d;
  wire [1:0] twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_13_i_adra_d;
  wire [63:0] twiddle_rsc_0_13_i_qa_d;
  wire [1:0] twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_14_i_adra_d;
  wire [63:0] twiddle_rsc_0_14_i_qa_d;
  wire [1:0] twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_rsc_0_15_i_adra_d;
  wire [63:0] twiddle_rsc_0_15_i_qa_d;
  wire [1:0] twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_0_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_0_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_1_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_1_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_2_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_2_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_3_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_3_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_4_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_4_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_5_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_5_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_6_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_6_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_7_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_7_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_8_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_8_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_9_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_9_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_10_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_10_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_11_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_11_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_12_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_12_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_13_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_13_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_14_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_14_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire [7:0] twiddle_h_rsc_0_15_i_adra_d;
  wire [63:0] twiddle_h_rsc_0_15_i_qa_d;
  wire [1:0] twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d;
  wire yt_rsc_0_0_clkb_en;
  wire yt_rsc_0_0_clka_en;
  wire [31:0] yt_rsc_0_0_qb;
  wire yt_rsc_0_0_web;
  wire [31:0] yt_rsc_0_0_db;
  wire [7:0] yt_rsc_0_0_adrb;
  wire [31:0] yt_rsc_0_0_qa;
  wire yt_rsc_0_0_wea;
  wire [31:0] yt_rsc_0_0_da;
  wire [7:0] yt_rsc_0_0_adra;
  wire yt_rsc_0_1_clkb_en;
  wire yt_rsc_0_1_clka_en;
  wire [31:0] yt_rsc_0_1_qb;
  wire yt_rsc_0_1_web;
  wire [31:0] yt_rsc_0_1_db;
  wire [7:0] yt_rsc_0_1_adrb;
  wire [31:0] yt_rsc_0_1_qa;
  wire yt_rsc_0_1_wea;
  wire [31:0] yt_rsc_0_1_da;
  wire [7:0] yt_rsc_0_1_adra;
  wire yt_rsc_0_2_clkb_en;
  wire yt_rsc_0_2_clka_en;
  wire [31:0] yt_rsc_0_2_qb;
  wire yt_rsc_0_2_web;
  wire [31:0] yt_rsc_0_2_db;
  wire [7:0] yt_rsc_0_2_adrb;
  wire [31:0] yt_rsc_0_2_qa;
  wire yt_rsc_0_2_wea;
  wire [31:0] yt_rsc_0_2_da;
  wire [7:0] yt_rsc_0_2_adra;
  wire yt_rsc_0_3_clkb_en;
  wire yt_rsc_0_3_clka_en;
  wire [31:0] yt_rsc_0_3_qb;
  wire yt_rsc_0_3_web;
  wire [31:0] yt_rsc_0_3_db;
  wire [7:0] yt_rsc_0_3_adrb;
  wire [31:0] yt_rsc_0_3_qa;
  wire yt_rsc_0_3_wea;
  wire [31:0] yt_rsc_0_3_da;
  wire [7:0] yt_rsc_0_3_adra;
  wire yt_rsc_0_4_clkb_en;
  wire yt_rsc_0_4_clka_en;
  wire [31:0] yt_rsc_0_4_qb;
  wire yt_rsc_0_4_web;
  wire [31:0] yt_rsc_0_4_db;
  wire [7:0] yt_rsc_0_4_adrb;
  wire [31:0] yt_rsc_0_4_qa;
  wire yt_rsc_0_4_wea;
  wire [31:0] yt_rsc_0_4_da;
  wire [7:0] yt_rsc_0_4_adra;
  wire yt_rsc_0_5_clkb_en;
  wire yt_rsc_0_5_clka_en;
  wire [31:0] yt_rsc_0_5_qb;
  wire yt_rsc_0_5_web;
  wire [31:0] yt_rsc_0_5_db;
  wire [7:0] yt_rsc_0_5_adrb;
  wire [31:0] yt_rsc_0_5_qa;
  wire yt_rsc_0_5_wea;
  wire [31:0] yt_rsc_0_5_da;
  wire [7:0] yt_rsc_0_5_adra;
  wire yt_rsc_0_6_clkb_en;
  wire yt_rsc_0_6_clka_en;
  wire [31:0] yt_rsc_0_6_qb;
  wire yt_rsc_0_6_web;
  wire [31:0] yt_rsc_0_6_db;
  wire [7:0] yt_rsc_0_6_adrb;
  wire [31:0] yt_rsc_0_6_qa;
  wire yt_rsc_0_6_wea;
  wire [31:0] yt_rsc_0_6_da;
  wire [7:0] yt_rsc_0_6_adra;
  wire yt_rsc_0_7_clkb_en;
  wire yt_rsc_0_7_clka_en;
  wire [31:0] yt_rsc_0_7_qb;
  wire yt_rsc_0_7_web;
  wire [31:0] yt_rsc_0_7_db;
  wire [7:0] yt_rsc_0_7_adrb;
  wire [31:0] yt_rsc_0_7_qa;
  wire yt_rsc_0_7_wea;
  wire [31:0] yt_rsc_0_7_da;
  wire [7:0] yt_rsc_0_7_adra;
  wire yt_rsc_0_8_clkb_en;
  wire yt_rsc_0_8_clka_en;
  wire [31:0] yt_rsc_0_8_qb;
  wire yt_rsc_0_8_web;
  wire [31:0] yt_rsc_0_8_db;
  wire [7:0] yt_rsc_0_8_adrb;
  wire [31:0] yt_rsc_0_8_qa;
  wire yt_rsc_0_8_wea;
  wire [31:0] yt_rsc_0_8_da;
  wire [7:0] yt_rsc_0_8_adra;
  wire yt_rsc_0_9_clkb_en;
  wire yt_rsc_0_9_clka_en;
  wire [31:0] yt_rsc_0_9_qb;
  wire yt_rsc_0_9_web;
  wire [31:0] yt_rsc_0_9_db;
  wire [7:0] yt_rsc_0_9_adrb;
  wire [31:0] yt_rsc_0_9_qa;
  wire yt_rsc_0_9_wea;
  wire [31:0] yt_rsc_0_9_da;
  wire [7:0] yt_rsc_0_9_adra;
  wire yt_rsc_0_10_clkb_en;
  wire yt_rsc_0_10_clka_en;
  wire [31:0] yt_rsc_0_10_qb;
  wire yt_rsc_0_10_web;
  wire [31:0] yt_rsc_0_10_db;
  wire [7:0] yt_rsc_0_10_adrb;
  wire [31:0] yt_rsc_0_10_qa;
  wire yt_rsc_0_10_wea;
  wire [31:0] yt_rsc_0_10_da;
  wire [7:0] yt_rsc_0_10_adra;
  wire yt_rsc_0_11_clkb_en;
  wire yt_rsc_0_11_clka_en;
  wire [31:0] yt_rsc_0_11_qb;
  wire yt_rsc_0_11_web;
  wire [31:0] yt_rsc_0_11_db;
  wire [7:0] yt_rsc_0_11_adrb;
  wire [31:0] yt_rsc_0_11_qa;
  wire yt_rsc_0_11_wea;
  wire [31:0] yt_rsc_0_11_da;
  wire [7:0] yt_rsc_0_11_adra;
  wire yt_rsc_0_12_clkb_en;
  wire yt_rsc_0_12_clka_en;
  wire [31:0] yt_rsc_0_12_qb;
  wire yt_rsc_0_12_web;
  wire [31:0] yt_rsc_0_12_db;
  wire [7:0] yt_rsc_0_12_adrb;
  wire [31:0] yt_rsc_0_12_qa;
  wire yt_rsc_0_12_wea;
  wire [31:0] yt_rsc_0_12_da;
  wire [7:0] yt_rsc_0_12_adra;
  wire yt_rsc_0_13_clkb_en;
  wire yt_rsc_0_13_clka_en;
  wire [31:0] yt_rsc_0_13_qb;
  wire yt_rsc_0_13_web;
  wire [31:0] yt_rsc_0_13_db;
  wire [7:0] yt_rsc_0_13_adrb;
  wire [31:0] yt_rsc_0_13_qa;
  wire yt_rsc_0_13_wea;
  wire [31:0] yt_rsc_0_13_da;
  wire [7:0] yt_rsc_0_13_adra;
  wire yt_rsc_0_14_clkb_en;
  wire yt_rsc_0_14_clka_en;
  wire [31:0] yt_rsc_0_14_qb;
  wire yt_rsc_0_14_web;
  wire [31:0] yt_rsc_0_14_db;
  wire [7:0] yt_rsc_0_14_adrb;
  wire [31:0] yt_rsc_0_14_qa;
  wire yt_rsc_0_14_wea;
  wire [31:0] yt_rsc_0_14_da;
  wire [7:0] yt_rsc_0_14_adra;
  wire yt_rsc_0_15_clkb_en;
  wire yt_rsc_0_15_clka_en;
  wire [31:0] yt_rsc_0_15_qb;
  wire yt_rsc_0_15_web;
  wire [31:0] yt_rsc_0_15_db;
  wire [7:0] yt_rsc_0_15_adrb;
  wire [31:0] yt_rsc_0_15_qa;
  wire yt_rsc_0_15_wea;
  wire [31:0] yt_rsc_0_15_da;
  wire [7:0] yt_rsc_0_15_adra;
  wire yt_rsc_0_16_clkb_en;
  wire yt_rsc_0_16_clka_en;
  wire [31:0] yt_rsc_0_16_qb;
  wire yt_rsc_0_16_web;
  wire [31:0] yt_rsc_0_16_db;
  wire [7:0] yt_rsc_0_16_adrb;
  wire [31:0] yt_rsc_0_16_qa;
  wire yt_rsc_0_16_wea;
  wire [31:0] yt_rsc_0_16_da;
  wire [7:0] yt_rsc_0_16_adra;
  wire yt_rsc_0_17_clkb_en;
  wire yt_rsc_0_17_clka_en;
  wire [31:0] yt_rsc_0_17_qb;
  wire yt_rsc_0_17_web;
  wire [31:0] yt_rsc_0_17_db;
  wire [7:0] yt_rsc_0_17_adrb;
  wire [31:0] yt_rsc_0_17_qa;
  wire yt_rsc_0_17_wea;
  wire [31:0] yt_rsc_0_17_da;
  wire [7:0] yt_rsc_0_17_adra;
  wire yt_rsc_0_18_clkb_en;
  wire yt_rsc_0_18_clka_en;
  wire [31:0] yt_rsc_0_18_qb;
  wire yt_rsc_0_18_web;
  wire [31:0] yt_rsc_0_18_db;
  wire [7:0] yt_rsc_0_18_adrb;
  wire [31:0] yt_rsc_0_18_qa;
  wire yt_rsc_0_18_wea;
  wire [31:0] yt_rsc_0_18_da;
  wire [7:0] yt_rsc_0_18_adra;
  wire yt_rsc_0_19_clkb_en;
  wire yt_rsc_0_19_clka_en;
  wire [31:0] yt_rsc_0_19_qb;
  wire yt_rsc_0_19_web;
  wire [31:0] yt_rsc_0_19_db;
  wire [7:0] yt_rsc_0_19_adrb;
  wire [31:0] yt_rsc_0_19_qa;
  wire yt_rsc_0_19_wea;
  wire [31:0] yt_rsc_0_19_da;
  wire [7:0] yt_rsc_0_19_adra;
  wire yt_rsc_0_20_clkb_en;
  wire yt_rsc_0_20_clka_en;
  wire [31:0] yt_rsc_0_20_qb;
  wire yt_rsc_0_20_web;
  wire [31:0] yt_rsc_0_20_db;
  wire [7:0] yt_rsc_0_20_adrb;
  wire [31:0] yt_rsc_0_20_qa;
  wire yt_rsc_0_20_wea;
  wire [31:0] yt_rsc_0_20_da;
  wire [7:0] yt_rsc_0_20_adra;
  wire yt_rsc_0_21_clkb_en;
  wire yt_rsc_0_21_clka_en;
  wire [31:0] yt_rsc_0_21_qb;
  wire yt_rsc_0_21_web;
  wire [31:0] yt_rsc_0_21_db;
  wire [7:0] yt_rsc_0_21_adrb;
  wire [31:0] yt_rsc_0_21_qa;
  wire yt_rsc_0_21_wea;
  wire [31:0] yt_rsc_0_21_da;
  wire [7:0] yt_rsc_0_21_adra;
  wire yt_rsc_0_22_clkb_en;
  wire yt_rsc_0_22_clka_en;
  wire [31:0] yt_rsc_0_22_qb;
  wire yt_rsc_0_22_web;
  wire [31:0] yt_rsc_0_22_db;
  wire [7:0] yt_rsc_0_22_adrb;
  wire [31:0] yt_rsc_0_22_qa;
  wire yt_rsc_0_22_wea;
  wire [31:0] yt_rsc_0_22_da;
  wire [7:0] yt_rsc_0_22_adra;
  wire yt_rsc_0_23_clkb_en;
  wire yt_rsc_0_23_clka_en;
  wire [31:0] yt_rsc_0_23_qb;
  wire yt_rsc_0_23_web;
  wire [31:0] yt_rsc_0_23_db;
  wire [7:0] yt_rsc_0_23_adrb;
  wire [31:0] yt_rsc_0_23_qa;
  wire yt_rsc_0_23_wea;
  wire [31:0] yt_rsc_0_23_da;
  wire [7:0] yt_rsc_0_23_adra;
  wire yt_rsc_0_24_clkb_en;
  wire yt_rsc_0_24_clka_en;
  wire [31:0] yt_rsc_0_24_qb;
  wire yt_rsc_0_24_web;
  wire [31:0] yt_rsc_0_24_db;
  wire [7:0] yt_rsc_0_24_adrb;
  wire [31:0] yt_rsc_0_24_qa;
  wire yt_rsc_0_24_wea;
  wire [31:0] yt_rsc_0_24_da;
  wire [7:0] yt_rsc_0_24_adra;
  wire yt_rsc_0_25_clkb_en;
  wire yt_rsc_0_25_clka_en;
  wire [31:0] yt_rsc_0_25_qb;
  wire yt_rsc_0_25_web;
  wire [31:0] yt_rsc_0_25_db;
  wire [7:0] yt_rsc_0_25_adrb;
  wire [31:0] yt_rsc_0_25_qa;
  wire yt_rsc_0_25_wea;
  wire [31:0] yt_rsc_0_25_da;
  wire [7:0] yt_rsc_0_25_adra;
  wire yt_rsc_0_26_clkb_en;
  wire yt_rsc_0_26_clka_en;
  wire [31:0] yt_rsc_0_26_qb;
  wire yt_rsc_0_26_web;
  wire [31:0] yt_rsc_0_26_db;
  wire [7:0] yt_rsc_0_26_adrb;
  wire [31:0] yt_rsc_0_26_qa;
  wire yt_rsc_0_26_wea;
  wire [31:0] yt_rsc_0_26_da;
  wire [7:0] yt_rsc_0_26_adra;
  wire yt_rsc_0_27_clkb_en;
  wire yt_rsc_0_27_clka_en;
  wire [31:0] yt_rsc_0_27_qb;
  wire yt_rsc_0_27_web;
  wire [31:0] yt_rsc_0_27_db;
  wire [7:0] yt_rsc_0_27_adrb;
  wire [31:0] yt_rsc_0_27_qa;
  wire yt_rsc_0_27_wea;
  wire [31:0] yt_rsc_0_27_da;
  wire [7:0] yt_rsc_0_27_adra;
  wire yt_rsc_0_28_clkb_en;
  wire yt_rsc_0_28_clka_en;
  wire [31:0] yt_rsc_0_28_qb;
  wire yt_rsc_0_28_web;
  wire [31:0] yt_rsc_0_28_db;
  wire [7:0] yt_rsc_0_28_adrb;
  wire [31:0] yt_rsc_0_28_qa;
  wire yt_rsc_0_28_wea;
  wire [31:0] yt_rsc_0_28_da;
  wire [7:0] yt_rsc_0_28_adra;
  wire yt_rsc_0_29_clkb_en;
  wire yt_rsc_0_29_clka_en;
  wire [31:0] yt_rsc_0_29_qb;
  wire yt_rsc_0_29_web;
  wire [31:0] yt_rsc_0_29_db;
  wire [7:0] yt_rsc_0_29_adrb;
  wire [31:0] yt_rsc_0_29_qa;
  wire yt_rsc_0_29_wea;
  wire [31:0] yt_rsc_0_29_da;
  wire [7:0] yt_rsc_0_29_adra;
  wire yt_rsc_0_30_clkb_en;
  wire yt_rsc_0_30_clka_en;
  wire [31:0] yt_rsc_0_30_qb;
  wire yt_rsc_0_30_web;
  wire [31:0] yt_rsc_0_30_db;
  wire [7:0] yt_rsc_0_30_adrb;
  wire [31:0] yt_rsc_0_30_qa;
  wire yt_rsc_0_30_wea;
  wire [31:0] yt_rsc_0_30_da;
  wire [7:0] yt_rsc_0_30_adra;
  wire yt_rsc_0_31_clkb_en;
  wire yt_rsc_0_31_clka_en;
  wire [31:0] yt_rsc_0_31_qb;
  wire yt_rsc_0_31_web;
  wire [31:0] yt_rsc_0_31_db;
  wire [7:0] yt_rsc_0_31_adrb;
  wire [31:0] yt_rsc_0_31_qa;
  wire yt_rsc_0_31_wea;
  wire [31:0] yt_rsc_0_31_da;
  wire [7:0] yt_rsc_0_31_adra;
  wire [1:0] yt_rsc_0_0_i_wea_d_iff;
  wire [1:0] yt_rsc_0_16_i_wea_d_iff;
  wire [1:0] xt_rsc_0_0_i_wea_d_iff;
  wire [1:0] xt_rsc_0_16_i_wea_d_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [15:0] nl_twiddle_rsc_0_0_i_adra_d;
  assign nl_twiddle_rsc_0_0_i_adra_d = {8'b00000000 , twiddle_rsc_0_0_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_1_i_adra_d;
  assign nl_twiddle_rsc_0_1_i_adra_d = {8'b00000000 , twiddle_rsc_0_1_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_2_i_adra_d;
  assign nl_twiddle_rsc_0_2_i_adra_d = {8'b00000000 , twiddle_rsc_0_2_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_3_i_adra_d;
  assign nl_twiddle_rsc_0_3_i_adra_d = {8'b00000000 , twiddle_rsc_0_3_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_4_i_adra_d;
  assign nl_twiddle_rsc_0_4_i_adra_d = {8'b00000000 , twiddle_rsc_0_4_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_5_i_adra_d;
  assign nl_twiddle_rsc_0_5_i_adra_d = {8'b00000000 , twiddle_rsc_0_5_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_6_i_adra_d;
  assign nl_twiddle_rsc_0_6_i_adra_d = {8'b00000000 , twiddle_rsc_0_6_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_7_i_adra_d;
  assign nl_twiddle_rsc_0_7_i_adra_d = {8'b00000000 , twiddle_rsc_0_7_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_8_i_adra_d;
  assign nl_twiddle_rsc_0_8_i_adra_d = {8'b00000000 , twiddle_rsc_0_8_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_9_i_adra_d;
  assign nl_twiddle_rsc_0_9_i_adra_d = {8'b00000000 , twiddle_rsc_0_9_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_10_i_adra_d;
  assign nl_twiddle_rsc_0_10_i_adra_d = {8'b00000000 , twiddle_rsc_0_10_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_11_i_adra_d;
  assign nl_twiddle_rsc_0_11_i_adra_d = {8'b00000000 , twiddle_rsc_0_11_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_12_i_adra_d;
  assign nl_twiddle_rsc_0_12_i_adra_d = {8'b00000000 , twiddle_rsc_0_12_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_13_i_adra_d;
  assign nl_twiddle_rsc_0_13_i_adra_d = {8'b00000000 , twiddle_rsc_0_13_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_14_i_adra_d;
  assign nl_twiddle_rsc_0_14_i_adra_d = {8'b00000000 , twiddle_rsc_0_14_i_adra_d};
  wire [15:0] nl_twiddle_rsc_0_15_i_adra_d;
  assign nl_twiddle_rsc_0_15_i_adra_d = {8'b00000000 , twiddle_rsc_0_15_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_0_i_adra_d;
  assign nl_twiddle_h_rsc_0_0_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_0_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_1_i_adra_d;
  assign nl_twiddle_h_rsc_0_1_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_1_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_2_i_adra_d;
  assign nl_twiddle_h_rsc_0_2_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_2_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_3_i_adra_d;
  assign nl_twiddle_h_rsc_0_3_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_3_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_4_i_adra_d;
  assign nl_twiddle_h_rsc_0_4_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_4_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_5_i_adra_d;
  assign nl_twiddle_h_rsc_0_5_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_5_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_6_i_adra_d;
  assign nl_twiddle_h_rsc_0_6_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_6_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_7_i_adra_d;
  assign nl_twiddle_h_rsc_0_7_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_7_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_8_i_adra_d;
  assign nl_twiddle_h_rsc_0_8_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_8_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_9_i_adra_d;
  assign nl_twiddle_h_rsc_0_9_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_9_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_10_i_adra_d;
  assign nl_twiddle_h_rsc_0_10_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_10_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_11_i_adra_d;
  assign nl_twiddle_h_rsc_0_11_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_11_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_12_i_adra_d;
  assign nl_twiddle_h_rsc_0_12_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_12_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_13_i_adra_d;
  assign nl_twiddle_h_rsc_0_13_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_13_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_14_i_adra_d;
  assign nl_twiddle_h_rsc_0_14_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_14_i_adra_d};
  wire [15:0] nl_twiddle_h_rsc_0_15_i_adra_d;
  assign nl_twiddle_h_rsc_0_15_i_adra_d = {8'b00000000 , twiddle_h_rsc_0_15_i_adra_d};
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_0_comp (
      .adra(yt_rsc_0_0_adra),
      .adrb(yt_rsc_0_0_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_0_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_0_clkb_en),
      .da(yt_rsc_0_0_da),
      .db(yt_rsc_0_0_db),
      .qa(yt_rsc_0_0_qa),
      .qb(yt_rsc_0_0_qb),
      .wea(yt_rsc_0_0_wea),
      .web(yt_rsc_0_0_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_1_comp (
      .adra(yt_rsc_0_1_adra),
      .adrb(yt_rsc_0_1_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_1_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_1_clkb_en),
      .da(yt_rsc_0_1_da),
      .db(yt_rsc_0_1_db),
      .qa(yt_rsc_0_1_qa),
      .qb(yt_rsc_0_1_qb),
      .wea(yt_rsc_0_1_wea),
      .web(yt_rsc_0_1_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_2_comp (
      .adra(yt_rsc_0_2_adra),
      .adrb(yt_rsc_0_2_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_2_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_2_clkb_en),
      .da(yt_rsc_0_2_da),
      .db(yt_rsc_0_2_db),
      .qa(yt_rsc_0_2_qa),
      .qb(yt_rsc_0_2_qb),
      .wea(yt_rsc_0_2_wea),
      .web(yt_rsc_0_2_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_3_comp (
      .adra(yt_rsc_0_3_adra),
      .adrb(yt_rsc_0_3_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_3_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_3_clkb_en),
      .da(yt_rsc_0_3_da),
      .db(yt_rsc_0_3_db),
      .qa(yt_rsc_0_3_qa),
      .qb(yt_rsc_0_3_qb),
      .wea(yt_rsc_0_3_wea),
      .web(yt_rsc_0_3_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_4_comp (
      .adra(yt_rsc_0_4_adra),
      .adrb(yt_rsc_0_4_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_4_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_4_clkb_en),
      .da(yt_rsc_0_4_da),
      .db(yt_rsc_0_4_db),
      .qa(yt_rsc_0_4_qa),
      .qb(yt_rsc_0_4_qb),
      .wea(yt_rsc_0_4_wea),
      .web(yt_rsc_0_4_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_5_comp (
      .adra(yt_rsc_0_5_adra),
      .adrb(yt_rsc_0_5_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_5_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_5_clkb_en),
      .da(yt_rsc_0_5_da),
      .db(yt_rsc_0_5_db),
      .qa(yt_rsc_0_5_qa),
      .qb(yt_rsc_0_5_qb),
      .wea(yt_rsc_0_5_wea),
      .web(yt_rsc_0_5_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_6_comp (
      .adra(yt_rsc_0_6_adra),
      .adrb(yt_rsc_0_6_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_6_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_6_clkb_en),
      .da(yt_rsc_0_6_da),
      .db(yt_rsc_0_6_db),
      .qa(yt_rsc_0_6_qa),
      .qb(yt_rsc_0_6_qb),
      .wea(yt_rsc_0_6_wea),
      .web(yt_rsc_0_6_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_7_comp (
      .adra(yt_rsc_0_7_adra),
      .adrb(yt_rsc_0_7_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_7_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_7_clkb_en),
      .da(yt_rsc_0_7_da),
      .db(yt_rsc_0_7_db),
      .qa(yt_rsc_0_7_qa),
      .qb(yt_rsc_0_7_qb),
      .wea(yt_rsc_0_7_wea),
      .web(yt_rsc_0_7_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_8_comp (
      .adra(yt_rsc_0_8_adra),
      .adrb(yt_rsc_0_8_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_8_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_8_clkb_en),
      .da(yt_rsc_0_8_da),
      .db(yt_rsc_0_8_db),
      .qa(yt_rsc_0_8_qa),
      .qb(yt_rsc_0_8_qb),
      .wea(yt_rsc_0_8_wea),
      .web(yt_rsc_0_8_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_9_comp (
      .adra(yt_rsc_0_9_adra),
      .adrb(yt_rsc_0_9_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_9_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_9_clkb_en),
      .da(yt_rsc_0_9_da),
      .db(yt_rsc_0_9_db),
      .qa(yt_rsc_0_9_qa),
      .qb(yt_rsc_0_9_qb),
      .wea(yt_rsc_0_9_wea),
      .web(yt_rsc_0_9_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_10_comp (
      .adra(yt_rsc_0_10_adra),
      .adrb(yt_rsc_0_10_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_10_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_10_clkb_en),
      .da(yt_rsc_0_10_da),
      .db(yt_rsc_0_10_db),
      .qa(yt_rsc_0_10_qa),
      .qb(yt_rsc_0_10_qb),
      .wea(yt_rsc_0_10_wea),
      .web(yt_rsc_0_10_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_11_comp (
      .adra(yt_rsc_0_11_adra),
      .adrb(yt_rsc_0_11_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_11_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_11_clkb_en),
      .da(yt_rsc_0_11_da),
      .db(yt_rsc_0_11_db),
      .qa(yt_rsc_0_11_qa),
      .qb(yt_rsc_0_11_qb),
      .wea(yt_rsc_0_11_wea),
      .web(yt_rsc_0_11_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_12_comp (
      .adra(yt_rsc_0_12_adra),
      .adrb(yt_rsc_0_12_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_12_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_12_clkb_en),
      .da(yt_rsc_0_12_da),
      .db(yt_rsc_0_12_db),
      .qa(yt_rsc_0_12_qa),
      .qb(yt_rsc_0_12_qb),
      .wea(yt_rsc_0_12_wea),
      .web(yt_rsc_0_12_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_13_comp (
      .adra(yt_rsc_0_13_adra),
      .adrb(yt_rsc_0_13_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_13_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_13_clkb_en),
      .da(yt_rsc_0_13_da),
      .db(yt_rsc_0_13_db),
      .qa(yt_rsc_0_13_qa),
      .qb(yt_rsc_0_13_qb),
      .wea(yt_rsc_0_13_wea),
      .web(yt_rsc_0_13_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_14_comp (
      .adra(yt_rsc_0_14_adra),
      .adrb(yt_rsc_0_14_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_14_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_14_clkb_en),
      .da(yt_rsc_0_14_da),
      .db(yt_rsc_0_14_db),
      .qa(yt_rsc_0_14_qa),
      .qb(yt_rsc_0_14_qb),
      .wea(yt_rsc_0_14_wea),
      .web(yt_rsc_0_14_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_15_comp (
      .adra(yt_rsc_0_15_adra),
      .adrb(yt_rsc_0_15_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_15_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_15_clkb_en),
      .da(yt_rsc_0_15_da),
      .db(yt_rsc_0_15_db),
      .qa(yt_rsc_0_15_qa),
      .qb(yt_rsc_0_15_qb),
      .wea(yt_rsc_0_15_wea),
      .web(yt_rsc_0_15_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_16_comp (
      .adra(yt_rsc_0_16_adra),
      .adrb(yt_rsc_0_16_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_16_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_16_clkb_en),
      .da(yt_rsc_0_16_da),
      .db(yt_rsc_0_16_db),
      .qa(yt_rsc_0_16_qa),
      .qb(yt_rsc_0_16_qb),
      .wea(yt_rsc_0_16_wea),
      .web(yt_rsc_0_16_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_17_comp (
      .adra(yt_rsc_0_17_adra),
      .adrb(yt_rsc_0_17_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_17_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_17_clkb_en),
      .da(yt_rsc_0_17_da),
      .db(yt_rsc_0_17_db),
      .qa(yt_rsc_0_17_qa),
      .qb(yt_rsc_0_17_qb),
      .wea(yt_rsc_0_17_wea),
      .web(yt_rsc_0_17_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_18_comp (
      .adra(yt_rsc_0_18_adra),
      .adrb(yt_rsc_0_18_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_18_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_18_clkb_en),
      .da(yt_rsc_0_18_da),
      .db(yt_rsc_0_18_db),
      .qa(yt_rsc_0_18_qa),
      .qb(yt_rsc_0_18_qb),
      .wea(yt_rsc_0_18_wea),
      .web(yt_rsc_0_18_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_19_comp (
      .adra(yt_rsc_0_19_adra),
      .adrb(yt_rsc_0_19_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_19_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_19_clkb_en),
      .da(yt_rsc_0_19_da),
      .db(yt_rsc_0_19_db),
      .qa(yt_rsc_0_19_qa),
      .qb(yt_rsc_0_19_qb),
      .wea(yt_rsc_0_19_wea),
      .web(yt_rsc_0_19_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_20_comp (
      .adra(yt_rsc_0_20_adra),
      .adrb(yt_rsc_0_20_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_20_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_20_clkb_en),
      .da(yt_rsc_0_20_da),
      .db(yt_rsc_0_20_db),
      .qa(yt_rsc_0_20_qa),
      .qb(yt_rsc_0_20_qb),
      .wea(yt_rsc_0_20_wea),
      .web(yt_rsc_0_20_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_21_comp (
      .adra(yt_rsc_0_21_adra),
      .adrb(yt_rsc_0_21_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_21_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_21_clkb_en),
      .da(yt_rsc_0_21_da),
      .db(yt_rsc_0_21_db),
      .qa(yt_rsc_0_21_qa),
      .qb(yt_rsc_0_21_qb),
      .wea(yt_rsc_0_21_wea),
      .web(yt_rsc_0_21_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_22_comp (
      .adra(yt_rsc_0_22_adra),
      .adrb(yt_rsc_0_22_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_22_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_22_clkb_en),
      .da(yt_rsc_0_22_da),
      .db(yt_rsc_0_22_db),
      .qa(yt_rsc_0_22_qa),
      .qb(yt_rsc_0_22_qb),
      .wea(yt_rsc_0_22_wea),
      .web(yt_rsc_0_22_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_23_comp (
      .adra(yt_rsc_0_23_adra),
      .adrb(yt_rsc_0_23_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_23_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_23_clkb_en),
      .da(yt_rsc_0_23_da),
      .db(yt_rsc_0_23_db),
      .qa(yt_rsc_0_23_qa),
      .qb(yt_rsc_0_23_qb),
      .wea(yt_rsc_0_23_wea),
      .web(yt_rsc_0_23_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_24_comp (
      .adra(yt_rsc_0_24_adra),
      .adrb(yt_rsc_0_24_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_24_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_24_clkb_en),
      .da(yt_rsc_0_24_da),
      .db(yt_rsc_0_24_db),
      .qa(yt_rsc_0_24_qa),
      .qb(yt_rsc_0_24_qb),
      .wea(yt_rsc_0_24_wea),
      .web(yt_rsc_0_24_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_25_comp (
      .adra(yt_rsc_0_25_adra),
      .adrb(yt_rsc_0_25_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_25_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_25_clkb_en),
      .da(yt_rsc_0_25_da),
      .db(yt_rsc_0_25_db),
      .qa(yt_rsc_0_25_qa),
      .qb(yt_rsc_0_25_qb),
      .wea(yt_rsc_0_25_wea),
      .web(yt_rsc_0_25_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_26_comp (
      .adra(yt_rsc_0_26_adra),
      .adrb(yt_rsc_0_26_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_26_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_26_clkb_en),
      .da(yt_rsc_0_26_da),
      .db(yt_rsc_0_26_db),
      .qa(yt_rsc_0_26_qa),
      .qb(yt_rsc_0_26_qb),
      .wea(yt_rsc_0_26_wea),
      .web(yt_rsc_0_26_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_27_comp (
      .adra(yt_rsc_0_27_adra),
      .adrb(yt_rsc_0_27_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_27_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_27_clkb_en),
      .da(yt_rsc_0_27_da),
      .db(yt_rsc_0_27_db),
      .qa(yt_rsc_0_27_qa),
      .qb(yt_rsc_0_27_qb),
      .wea(yt_rsc_0_27_wea),
      .web(yt_rsc_0_27_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_28_comp (
      .adra(yt_rsc_0_28_adra),
      .adrb(yt_rsc_0_28_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_28_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_28_clkb_en),
      .da(yt_rsc_0_28_da),
      .db(yt_rsc_0_28_db),
      .qa(yt_rsc_0_28_qa),
      .qb(yt_rsc_0_28_qb),
      .wea(yt_rsc_0_28_wea),
      .web(yt_rsc_0_28_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_29_comp (
      .adra(yt_rsc_0_29_adra),
      .adrb(yt_rsc_0_29_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_29_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_29_clkb_en),
      .da(yt_rsc_0_29_da),
      .db(yt_rsc_0_29_db),
      .qa(yt_rsc_0_29_qa),
      .qb(yt_rsc_0_29_qb),
      .wea(yt_rsc_0_29_wea),
      .web(yt_rsc_0_29_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_30_comp (
      .adra(yt_rsc_0_30_adra),
      .adrb(yt_rsc_0_30_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_30_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_30_clkb_en),
      .da(yt_rsc_0_30_da),
      .db(yt_rsc_0_30_db),
      .qa(yt_rsc_0_30_qa),
      .qb(yt_rsc_0_30_qb),
      .wea(yt_rsc_0_30_wea),
      .web(yt_rsc_0_30_web)
    );
  BLOCK_DPRAM_RBW_DUAL #(.addr_width(32'sd8),
  .data_width(32'sd32),
  .depth(32'sd256),
  .latency(32'sd1)) yt_rsc_0_31_comp (
      .adra(yt_rsc_0_31_adra),
      .adrb(yt_rsc_0_31_adrb),
      .clka(clk),
      .clka_en(yt_rsc_0_31_clkb_en),
      .clkb(clk),
      .clkb_en(yt_rsc_0_31_clkb_en),
      .da(yt_rsc_0_31_da),
      .db(yt_rsc_0_31_db),
      .qa(yt_rsc_0_31_qa),
      .qb(yt_rsc_0_31_qb),
      .wea(yt_rsc_0_31_wea),
      .web(yt_rsc_0_31_web)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_7_8_32_256_256_32_1_gen yt_rsc_0_0_i
      (
      .clkb_en(yt_rsc_0_0_clkb_en),
      .clka_en(yt_rsc_0_0_clka_en),
      .qb(yt_rsc_0_0_qb),
      .web(yt_rsc_0_0_web),
      .db(yt_rsc_0_0_db),
      .adrb(yt_rsc_0_0_adrb),
      .qa(yt_rsc_0_0_qa),
      .wea(yt_rsc_0_0_wea),
      .da(yt_rsc_0_0_da),
      .adra(yt_rsc_0_0_adra),
      .adra_d(yt_rsc_0_0_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_0_i_da_d),
      .qa_d(yt_rsc_0_0_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_8_8_32_256_256_32_1_gen yt_rsc_0_1_i
      (
      .clkb_en(yt_rsc_0_1_clkb_en),
      .clka_en(yt_rsc_0_1_clka_en),
      .qb(yt_rsc_0_1_qb),
      .web(yt_rsc_0_1_web),
      .db(yt_rsc_0_1_db),
      .adrb(yt_rsc_0_1_adrb),
      .qa(yt_rsc_0_1_qa),
      .wea(yt_rsc_0_1_wea),
      .da(yt_rsc_0_1_da),
      .adra(yt_rsc_0_1_adra),
      .adra_d(yt_rsc_0_1_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_1_i_da_d),
      .qa_d(yt_rsc_0_1_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_9_8_32_256_256_32_1_gen yt_rsc_0_2_i
      (
      .clkb_en(yt_rsc_0_2_clkb_en),
      .clka_en(yt_rsc_0_2_clka_en),
      .qb(yt_rsc_0_2_qb),
      .web(yt_rsc_0_2_web),
      .db(yt_rsc_0_2_db),
      .adrb(yt_rsc_0_2_adrb),
      .qa(yt_rsc_0_2_qa),
      .wea(yt_rsc_0_2_wea),
      .da(yt_rsc_0_2_da),
      .adra(yt_rsc_0_2_adra),
      .adra_d(yt_rsc_0_2_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_2_i_da_d),
      .qa_d(yt_rsc_0_2_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_10_8_32_256_256_32_1_gen yt_rsc_0_3_i
      (
      .clkb_en(yt_rsc_0_3_clkb_en),
      .clka_en(yt_rsc_0_3_clka_en),
      .qb(yt_rsc_0_3_qb),
      .web(yt_rsc_0_3_web),
      .db(yt_rsc_0_3_db),
      .adrb(yt_rsc_0_3_adrb),
      .qa(yt_rsc_0_3_qa),
      .wea(yt_rsc_0_3_wea),
      .da(yt_rsc_0_3_da),
      .adra(yt_rsc_0_3_adra),
      .adra_d(yt_rsc_0_3_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_3_i_da_d),
      .qa_d(yt_rsc_0_3_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_11_8_32_256_256_32_1_gen yt_rsc_0_4_i
      (
      .clkb_en(yt_rsc_0_4_clkb_en),
      .clka_en(yt_rsc_0_4_clka_en),
      .qb(yt_rsc_0_4_qb),
      .web(yt_rsc_0_4_web),
      .db(yt_rsc_0_4_db),
      .adrb(yt_rsc_0_4_adrb),
      .qa(yt_rsc_0_4_qa),
      .wea(yt_rsc_0_4_wea),
      .da(yt_rsc_0_4_da),
      .adra(yt_rsc_0_4_adra),
      .adra_d(yt_rsc_0_4_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_4_i_da_d),
      .qa_d(yt_rsc_0_4_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_12_8_32_256_256_32_1_gen yt_rsc_0_5_i
      (
      .clkb_en(yt_rsc_0_5_clkb_en),
      .clka_en(yt_rsc_0_5_clka_en),
      .qb(yt_rsc_0_5_qb),
      .web(yt_rsc_0_5_web),
      .db(yt_rsc_0_5_db),
      .adrb(yt_rsc_0_5_adrb),
      .qa(yt_rsc_0_5_qa),
      .wea(yt_rsc_0_5_wea),
      .da(yt_rsc_0_5_da),
      .adra(yt_rsc_0_5_adra),
      .adra_d(yt_rsc_0_5_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_5_i_da_d),
      .qa_d(yt_rsc_0_5_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_13_8_32_256_256_32_1_gen yt_rsc_0_6_i
      (
      .clkb_en(yt_rsc_0_6_clkb_en),
      .clka_en(yt_rsc_0_6_clka_en),
      .qb(yt_rsc_0_6_qb),
      .web(yt_rsc_0_6_web),
      .db(yt_rsc_0_6_db),
      .adrb(yt_rsc_0_6_adrb),
      .qa(yt_rsc_0_6_qa),
      .wea(yt_rsc_0_6_wea),
      .da(yt_rsc_0_6_da),
      .adra(yt_rsc_0_6_adra),
      .adra_d(yt_rsc_0_6_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_6_i_da_d),
      .qa_d(yt_rsc_0_6_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_14_8_32_256_256_32_1_gen yt_rsc_0_7_i
      (
      .clkb_en(yt_rsc_0_7_clkb_en),
      .clka_en(yt_rsc_0_7_clka_en),
      .qb(yt_rsc_0_7_qb),
      .web(yt_rsc_0_7_web),
      .db(yt_rsc_0_7_db),
      .adrb(yt_rsc_0_7_adrb),
      .qa(yt_rsc_0_7_qa),
      .wea(yt_rsc_0_7_wea),
      .da(yt_rsc_0_7_da),
      .adra(yt_rsc_0_7_adra),
      .adra_d(yt_rsc_0_7_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_7_i_da_d),
      .qa_d(yt_rsc_0_7_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_15_8_32_256_256_32_1_gen yt_rsc_0_8_i
      (
      .clkb_en(yt_rsc_0_8_clkb_en),
      .clka_en(yt_rsc_0_8_clka_en),
      .qb(yt_rsc_0_8_qb),
      .web(yt_rsc_0_8_web),
      .db(yt_rsc_0_8_db),
      .adrb(yt_rsc_0_8_adrb),
      .qa(yt_rsc_0_8_qa),
      .wea(yt_rsc_0_8_wea),
      .da(yt_rsc_0_8_da),
      .adra(yt_rsc_0_8_adra),
      .adra_d(yt_rsc_0_8_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_8_i_da_d),
      .qa_d(yt_rsc_0_8_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_16_8_32_256_256_32_1_gen yt_rsc_0_9_i
      (
      .clkb_en(yt_rsc_0_9_clkb_en),
      .clka_en(yt_rsc_0_9_clka_en),
      .qb(yt_rsc_0_9_qb),
      .web(yt_rsc_0_9_web),
      .db(yt_rsc_0_9_db),
      .adrb(yt_rsc_0_9_adrb),
      .qa(yt_rsc_0_9_qa),
      .wea(yt_rsc_0_9_wea),
      .da(yt_rsc_0_9_da),
      .adra(yt_rsc_0_9_adra),
      .adra_d(yt_rsc_0_9_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_9_i_da_d),
      .qa_d(yt_rsc_0_9_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_17_8_32_256_256_32_1_gen yt_rsc_0_10_i
      (
      .clkb_en(yt_rsc_0_10_clkb_en),
      .clka_en(yt_rsc_0_10_clka_en),
      .qb(yt_rsc_0_10_qb),
      .web(yt_rsc_0_10_web),
      .db(yt_rsc_0_10_db),
      .adrb(yt_rsc_0_10_adrb),
      .qa(yt_rsc_0_10_qa),
      .wea(yt_rsc_0_10_wea),
      .da(yt_rsc_0_10_da),
      .adra(yt_rsc_0_10_adra),
      .adra_d(yt_rsc_0_10_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_10_i_da_d),
      .qa_d(yt_rsc_0_10_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_18_8_32_256_256_32_1_gen yt_rsc_0_11_i
      (
      .clkb_en(yt_rsc_0_11_clkb_en),
      .clka_en(yt_rsc_0_11_clka_en),
      .qb(yt_rsc_0_11_qb),
      .web(yt_rsc_0_11_web),
      .db(yt_rsc_0_11_db),
      .adrb(yt_rsc_0_11_adrb),
      .qa(yt_rsc_0_11_qa),
      .wea(yt_rsc_0_11_wea),
      .da(yt_rsc_0_11_da),
      .adra(yt_rsc_0_11_adra),
      .adra_d(yt_rsc_0_11_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_11_i_da_d),
      .qa_d(yt_rsc_0_11_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_19_8_32_256_256_32_1_gen yt_rsc_0_12_i
      (
      .clkb_en(yt_rsc_0_12_clkb_en),
      .clka_en(yt_rsc_0_12_clka_en),
      .qb(yt_rsc_0_12_qb),
      .web(yt_rsc_0_12_web),
      .db(yt_rsc_0_12_db),
      .adrb(yt_rsc_0_12_adrb),
      .qa(yt_rsc_0_12_qa),
      .wea(yt_rsc_0_12_wea),
      .da(yt_rsc_0_12_da),
      .adra(yt_rsc_0_12_adra),
      .adra_d(yt_rsc_0_12_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_12_i_da_d),
      .qa_d(yt_rsc_0_12_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_20_8_32_256_256_32_1_gen yt_rsc_0_13_i
      (
      .clkb_en(yt_rsc_0_13_clkb_en),
      .clka_en(yt_rsc_0_13_clka_en),
      .qb(yt_rsc_0_13_qb),
      .web(yt_rsc_0_13_web),
      .db(yt_rsc_0_13_db),
      .adrb(yt_rsc_0_13_adrb),
      .qa(yt_rsc_0_13_qa),
      .wea(yt_rsc_0_13_wea),
      .da(yt_rsc_0_13_da),
      .adra(yt_rsc_0_13_adra),
      .adra_d(yt_rsc_0_13_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_13_i_da_d),
      .qa_d(yt_rsc_0_13_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_21_8_32_256_256_32_1_gen yt_rsc_0_14_i
      (
      .clkb_en(yt_rsc_0_14_clkb_en),
      .clka_en(yt_rsc_0_14_clka_en),
      .qb(yt_rsc_0_14_qb),
      .web(yt_rsc_0_14_web),
      .db(yt_rsc_0_14_db),
      .adrb(yt_rsc_0_14_adrb),
      .qa(yt_rsc_0_14_qa),
      .wea(yt_rsc_0_14_wea),
      .da(yt_rsc_0_14_da),
      .adra(yt_rsc_0_14_adra),
      .adra_d(yt_rsc_0_14_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_14_i_da_d),
      .qa_d(yt_rsc_0_14_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_22_8_32_256_256_32_1_gen yt_rsc_0_15_i
      (
      .clkb_en(yt_rsc_0_15_clkb_en),
      .clka_en(yt_rsc_0_15_clka_en),
      .qb(yt_rsc_0_15_qb),
      .web(yt_rsc_0_15_web),
      .db(yt_rsc_0_15_db),
      .adrb(yt_rsc_0_15_adrb),
      .qa(yt_rsc_0_15_qa),
      .wea(yt_rsc_0_15_wea),
      .da(yt_rsc_0_15_da),
      .adra(yt_rsc_0_15_adra),
      .adra_d(yt_rsc_0_15_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_0_i_clka_en_d),
      .da_d(yt_rsc_0_15_i_da_d),
      .qa_d(yt_rsc_0_15_i_qa_d),
      .wea_d(yt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_23_8_32_256_256_32_1_gen yt_rsc_0_16_i
      (
      .clkb_en(yt_rsc_0_16_clkb_en),
      .clka_en(yt_rsc_0_16_clka_en),
      .qb(yt_rsc_0_16_qb),
      .web(yt_rsc_0_16_web),
      .db(yt_rsc_0_16_db),
      .adrb(yt_rsc_0_16_adrb),
      .qa(yt_rsc_0_16_qa),
      .wea(yt_rsc_0_16_wea),
      .da(yt_rsc_0_16_da),
      .adra(yt_rsc_0_16_adra),
      .adra_d(yt_rsc_0_16_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_16_i_da_d),
      .qa_d(yt_rsc_0_16_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_24_8_32_256_256_32_1_gen yt_rsc_0_17_i
      (
      .clkb_en(yt_rsc_0_17_clkb_en),
      .clka_en(yt_rsc_0_17_clka_en),
      .qb(yt_rsc_0_17_qb),
      .web(yt_rsc_0_17_web),
      .db(yt_rsc_0_17_db),
      .adrb(yt_rsc_0_17_adrb),
      .qa(yt_rsc_0_17_qa),
      .wea(yt_rsc_0_17_wea),
      .da(yt_rsc_0_17_da),
      .adra(yt_rsc_0_17_adra),
      .adra_d(yt_rsc_0_17_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_17_i_da_d),
      .qa_d(yt_rsc_0_17_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_25_8_32_256_256_32_1_gen yt_rsc_0_18_i
      (
      .clkb_en(yt_rsc_0_18_clkb_en),
      .clka_en(yt_rsc_0_18_clka_en),
      .qb(yt_rsc_0_18_qb),
      .web(yt_rsc_0_18_web),
      .db(yt_rsc_0_18_db),
      .adrb(yt_rsc_0_18_adrb),
      .qa(yt_rsc_0_18_qa),
      .wea(yt_rsc_0_18_wea),
      .da(yt_rsc_0_18_da),
      .adra(yt_rsc_0_18_adra),
      .adra_d(yt_rsc_0_18_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_18_i_da_d),
      .qa_d(yt_rsc_0_18_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_26_8_32_256_256_32_1_gen yt_rsc_0_19_i
      (
      .clkb_en(yt_rsc_0_19_clkb_en),
      .clka_en(yt_rsc_0_19_clka_en),
      .qb(yt_rsc_0_19_qb),
      .web(yt_rsc_0_19_web),
      .db(yt_rsc_0_19_db),
      .adrb(yt_rsc_0_19_adrb),
      .qa(yt_rsc_0_19_qa),
      .wea(yt_rsc_0_19_wea),
      .da(yt_rsc_0_19_da),
      .adra(yt_rsc_0_19_adra),
      .adra_d(yt_rsc_0_19_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_19_i_da_d),
      .qa_d(yt_rsc_0_19_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_27_8_32_256_256_32_1_gen yt_rsc_0_20_i
      (
      .clkb_en(yt_rsc_0_20_clkb_en),
      .clka_en(yt_rsc_0_20_clka_en),
      .qb(yt_rsc_0_20_qb),
      .web(yt_rsc_0_20_web),
      .db(yt_rsc_0_20_db),
      .adrb(yt_rsc_0_20_adrb),
      .qa(yt_rsc_0_20_qa),
      .wea(yt_rsc_0_20_wea),
      .da(yt_rsc_0_20_da),
      .adra(yt_rsc_0_20_adra),
      .adra_d(yt_rsc_0_20_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_20_i_da_d),
      .qa_d(yt_rsc_0_20_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_28_8_32_256_256_32_1_gen yt_rsc_0_21_i
      (
      .clkb_en(yt_rsc_0_21_clkb_en),
      .clka_en(yt_rsc_0_21_clka_en),
      .qb(yt_rsc_0_21_qb),
      .web(yt_rsc_0_21_web),
      .db(yt_rsc_0_21_db),
      .adrb(yt_rsc_0_21_adrb),
      .qa(yt_rsc_0_21_qa),
      .wea(yt_rsc_0_21_wea),
      .da(yt_rsc_0_21_da),
      .adra(yt_rsc_0_21_adra),
      .adra_d(yt_rsc_0_21_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_21_i_da_d),
      .qa_d(yt_rsc_0_21_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_29_8_32_256_256_32_1_gen yt_rsc_0_22_i
      (
      .clkb_en(yt_rsc_0_22_clkb_en),
      .clka_en(yt_rsc_0_22_clka_en),
      .qb(yt_rsc_0_22_qb),
      .web(yt_rsc_0_22_web),
      .db(yt_rsc_0_22_db),
      .adrb(yt_rsc_0_22_adrb),
      .qa(yt_rsc_0_22_qa),
      .wea(yt_rsc_0_22_wea),
      .da(yt_rsc_0_22_da),
      .adra(yt_rsc_0_22_adra),
      .adra_d(yt_rsc_0_22_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_22_i_da_d),
      .qa_d(yt_rsc_0_22_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_30_8_32_256_256_32_1_gen yt_rsc_0_23_i
      (
      .clkb_en(yt_rsc_0_23_clkb_en),
      .clka_en(yt_rsc_0_23_clka_en),
      .qb(yt_rsc_0_23_qb),
      .web(yt_rsc_0_23_web),
      .db(yt_rsc_0_23_db),
      .adrb(yt_rsc_0_23_adrb),
      .qa(yt_rsc_0_23_qa),
      .wea(yt_rsc_0_23_wea),
      .da(yt_rsc_0_23_da),
      .adra(yt_rsc_0_23_adra),
      .adra_d(yt_rsc_0_23_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_23_i_da_d),
      .qa_d(yt_rsc_0_23_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_31_8_32_256_256_32_1_gen yt_rsc_0_24_i
      (
      .clkb_en(yt_rsc_0_24_clkb_en),
      .clka_en(yt_rsc_0_24_clka_en),
      .qb(yt_rsc_0_24_qb),
      .web(yt_rsc_0_24_web),
      .db(yt_rsc_0_24_db),
      .adrb(yt_rsc_0_24_adrb),
      .qa(yt_rsc_0_24_qa),
      .wea(yt_rsc_0_24_wea),
      .da(yt_rsc_0_24_da),
      .adra(yt_rsc_0_24_adra),
      .adra_d(yt_rsc_0_24_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_24_i_da_d),
      .qa_d(yt_rsc_0_24_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_32_8_32_256_256_32_1_gen yt_rsc_0_25_i
      (
      .clkb_en(yt_rsc_0_25_clkb_en),
      .clka_en(yt_rsc_0_25_clka_en),
      .qb(yt_rsc_0_25_qb),
      .web(yt_rsc_0_25_web),
      .db(yt_rsc_0_25_db),
      .adrb(yt_rsc_0_25_adrb),
      .qa(yt_rsc_0_25_qa),
      .wea(yt_rsc_0_25_wea),
      .da(yt_rsc_0_25_da),
      .adra(yt_rsc_0_25_adra),
      .adra_d(yt_rsc_0_25_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_25_i_da_d),
      .qa_d(yt_rsc_0_25_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_33_8_32_256_256_32_1_gen yt_rsc_0_26_i
      (
      .clkb_en(yt_rsc_0_26_clkb_en),
      .clka_en(yt_rsc_0_26_clka_en),
      .qb(yt_rsc_0_26_qb),
      .web(yt_rsc_0_26_web),
      .db(yt_rsc_0_26_db),
      .adrb(yt_rsc_0_26_adrb),
      .qa(yt_rsc_0_26_qa),
      .wea(yt_rsc_0_26_wea),
      .da(yt_rsc_0_26_da),
      .adra(yt_rsc_0_26_adra),
      .adra_d(yt_rsc_0_26_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_26_i_da_d),
      .qa_d(yt_rsc_0_26_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_34_8_32_256_256_32_1_gen yt_rsc_0_27_i
      (
      .clkb_en(yt_rsc_0_27_clkb_en),
      .clka_en(yt_rsc_0_27_clka_en),
      .qb(yt_rsc_0_27_qb),
      .web(yt_rsc_0_27_web),
      .db(yt_rsc_0_27_db),
      .adrb(yt_rsc_0_27_adrb),
      .qa(yt_rsc_0_27_qa),
      .wea(yt_rsc_0_27_wea),
      .da(yt_rsc_0_27_da),
      .adra(yt_rsc_0_27_adra),
      .adra_d(yt_rsc_0_27_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_27_i_da_d),
      .qa_d(yt_rsc_0_27_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_35_8_32_256_256_32_1_gen yt_rsc_0_28_i
      (
      .clkb_en(yt_rsc_0_28_clkb_en),
      .clka_en(yt_rsc_0_28_clka_en),
      .qb(yt_rsc_0_28_qb),
      .web(yt_rsc_0_28_web),
      .db(yt_rsc_0_28_db),
      .adrb(yt_rsc_0_28_adrb),
      .qa(yt_rsc_0_28_qa),
      .wea(yt_rsc_0_28_wea),
      .da(yt_rsc_0_28_da),
      .adra(yt_rsc_0_28_adra),
      .adra_d(yt_rsc_0_28_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_28_i_da_d),
      .qa_d(yt_rsc_0_28_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_36_8_32_256_256_32_1_gen yt_rsc_0_29_i
      (
      .clkb_en(yt_rsc_0_29_clkb_en),
      .clka_en(yt_rsc_0_29_clka_en),
      .qb(yt_rsc_0_29_qb),
      .web(yt_rsc_0_29_web),
      .db(yt_rsc_0_29_db),
      .adrb(yt_rsc_0_29_adrb),
      .qa(yt_rsc_0_29_qa),
      .wea(yt_rsc_0_29_wea),
      .da(yt_rsc_0_29_da),
      .adra(yt_rsc_0_29_adra),
      .adra_d(yt_rsc_0_29_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_29_i_da_d),
      .qa_d(yt_rsc_0_29_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_37_8_32_256_256_32_1_gen yt_rsc_0_30_i
      (
      .clkb_en(yt_rsc_0_30_clkb_en),
      .clka_en(yt_rsc_0_30_clka_en),
      .qb(yt_rsc_0_30_qb),
      .web(yt_rsc_0_30_web),
      .db(yt_rsc_0_30_db),
      .adrb(yt_rsc_0_30_adrb),
      .qa(yt_rsc_0_30_qa),
      .wea(yt_rsc_0_30_wea),
      .da(yt_rsc_0_30_da),
      .adra(yt_rsc_0_30_adra),
      .adra_d(yt_rsc_0_30_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_30_i_da_d),
      .qa_d(yt_rsc_0_30_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_en_38_8_32_256_256_32_1_gen yt_rsc_0_31_i
      (
      .clkb_en(yt_rsc_0_31_clkb_en),
      .clka_en(yt_rsc_0_31_clka_en),
      .qb(yt_rsc_0_31_qb),
      .web(yt_rsc_0_31_web),
      .db(yt_rsc_0_31_db),
      .adrb(yt_rsc_0_31_adrb),
      .qa(yt_rsc_0_31_qa),
      .wea(yt_rsc_0_31_wea),
      .da(yt_rsc_0_31_da),
      .adra(yt_rsc_0_31_adra),
      .adra_d(yt_rsc_0_31_i_adra_d),
      .clka(clk),
      .clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .clkb_en_d(yt_rsc_0_16_i_clka_en_d),
      .da_d(yt_rsc_0_31_i_da_d),
      .qa_d(yt_rsc_0_31_i_qa_d),
      .wea_d(yt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(yt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_39_8_32_256_256_32_1_gen xt_rsc_0_0_i
      (
      .qb(xt_rsc_0_0_qb),
      .web(xt_rsc_0_0_web),
      .db(xt_rsc_0_0_db),
      .adrb(xt_rsc_0_0_adrb),
      .qa(xt_rsc_0_0_qa),
      .wea(xt_rsc_0_0_wea),
      .da(xt_rsc_0_0_da),
      .adra(xt_rsc_0_0_adra),
      .adra_d(xt_rsc_0_0_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_0_i_da_d),
      .qa_d(xt_rsc_0_0_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_40_8_32_256_256_32_1_gen xt_rsc_0_1_i
      (
      .qb(xt_rsc_0_1_qb),
      .web(xt_rsc_0_1_web),
      .db(xt_rsc_0_1_db),
      .adrb(xt_rsc_0_1_adrb),
      .qa(xt_rsc_0_1_qa),
      .wea(xt_rsc_0_1_wea),
      .da(xt_rsc_0_1_da),
      .adra(xt_rsc_0_1_adra),
      .adra_d(xt_rsc_0_1_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_1_i_da_d),
      .qa_d(xt_rsc_0_1_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_41_8_32_256_256_32_1_gen xt_rsc_0_2_i
      (
      .qb(xt_rsc_0_2_qb),
      .web(xt_rsc_0_2_web),
      .db(xt_rsc_0_2_db),
      .adrb(xt_rsc_0_2_adrb),
      .qa(xt_rsc_0_2_qa),
      .wea(xt_rsc_0_2_wea),
      .da(xt_rsc_0_2_da),
      .adra(xt_rsc_0_2_adra),
      .adra_d(xt_rsc_0_2_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_2_i_da_d),
      .qa_d(xt_rsc_0_2_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_42_8_32_256_256_32_1_gen xt_rsc_0_3_i
      (
      .qb(xt_rsc_0_3_qb),
      .web(xt_rsc_0_3_web),
      .db(xt_rsc_0_3_db),
      .adrb(xt_rsc_0_3_adrb),
      .qa(xt_rsc_0_3_qa),
      .wea(xt_rsc_0_3_wea),
      .da(xt_rsc_0_3_da),
      .adra(xt_rsc_0_3_adra),
      .adra_d(xt_rsc_0_3_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_3_i_da_d),
      .qa_d(xt_rsc_0_3_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_43_8_32_256_256_32_1_gen xt_rsc_0_4_i
      (
      .qb(xt_rsc_0_4_qb),
      .web(xt_rsc_0_4_web),
      .db(xt_rsc_0_4_db),
      .adrb(xt_rsc_0_4_adrb),
      .qa(xt_rsc_0_4_qa),
      .wea(xt_rsc_0_4_wea),
      .da(xt_rsc_0_4_da),
      .adra(xt_rsc_0_4_adra),
      .adra_d(xt_rsc_0_4_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_4_i_da_d),
      .qa_d(xt_rsc_0_4_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_44_8_32_256_256_32_1_gen xt_rsc_0_5_i
      (
      .qb(xt_rsc_0_5_qb),
      .web(xt_rsc_0_5_web),
      .db(xt_rsc_0_5_db),
      .adrb(xt_rsc_0_5_adrb),
      .qa(xt_rsc_0_5_qa),
      .wea(xt_rsc_0_5_wea),
      .da(xt_rsc_0_5_da),
      .adra(xt_rsc_0_5_adra),
      .adra_d(xt_rsc_0_5_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_5_i_da_d),
      .qa_d(xt_rsc_0_5_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_45_8_32_256_256_32_1_gen xt_rsc_0_6_i
      (
      .qb(xt_rsc_0_6_qb),
      .web(xt_rsc_0_6_web),
      .db(xt_rsc_0_6_db),
      .adrb(xt_rsc_0_6_adrb),
      .qa(xt_rsc_0_6_qa),
      .wea(xt_rsc_0_6_wea),
      .da(xt_rsc_0_6_da),
      .adra(xt_rsc_0_6_adra),
      .adra_d(xt_rsc_0_6_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_6_i_da_d),
      .qa_d(xt_rsc_0_6_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_46_8_32_256_256_32_1_gen xt_rsc_0_7_i
      (
      .qb(xt_rsc_0_7_qb),
      .web(xt_rsc_0_7_web),
      .db(xt_rsc_0_7_db),
      .adrb(xt_rsc_0_7_adrb),
      .qa(xt_rsc_0_7_qa),
      .wea(xt_rsc_0_7_wea),
      .da(xt_rsc_0_7_da),
      .adra(xt_rsc_0_7_adra),
      .adra_d(xt_rsc_0_7_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_7_i_da_d),
      .qa_d(xt_rsc_0_7_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_47_8_32_256_256_32_1_gen xt_rsc_0_8_i
      (
      .qb(xt_rsc_0_8_qb),
      .web(xt_rsc_0_8_web),
      .db(xt_rsc_0_8_db),
      .adrb(xt_rsc_0_8_adrb),
      .qa(xt_rsc_0_8_qa),
      .wea(xt_rsc_0_8_wea),
      .da(xt_rsc_0_8_da),
      .adra(xt_rsc_0_8_adra),
      .adra_d(xt_rsc_0_8_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_8_i_da_d),
      .qa_d(xt_rsc_0_8_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_48_8_32_256_256_32_1_gen xt_rsc_0_9_i
      (
      .qb(xt_rsc_0_9_qb),
      .web(xt_rsc_0_9_web),
      .db(xt_rsc_0_9_db),
      .adrb(xt_rsc_0_9_adrb),
      .qa(xt_rsc_0_9_qa),
      .wea(xt_rsc_0_9_wea),
      .da(xt_rsc_0_9_da),
      .adra(xt_rsc_0_9_adra),
      .adra_d(xt_rsc_0_9_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_9_i_da_d),
      .qa_d(xt_rsc_0_9_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_49_8_32_256_256_32_1_gen xt_rsc_0_10_i
      (
      .qb(xt_rsc_0_10_qb),
      .web(xt_rsc_0_10_web),
      .db(xt_rsc_0_10_db),
      .adrb(xt_rsc_0_10_adrb),
      .qa(xt_rsc_0_10_qa),
      .wea(xt_rsc_0_10_wea),
      .da(xt_rsc_0_10_da),
      .adra(xt_rsc_0_10_adra),
      .adra_d(xt_rsc_0_10_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_10_i_da_d),
      .qa_d(xt_rsc_0_10_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_50_8_32_256_256_32_1_gen xt_rsc_0_11_i
      (
      .qb(xt_rsc_0_11_qb),
      .web(xt_rsc_0_11_web),
      .db(xt_rsc_0_11_db),
      .adrb(xt_rsc_0_11_adrb),
      .qa(xt_rsc_0_11_qa),
      .wea(xt_rsc_0_11_wea),
      .da(xt_rsc_0_11_da),
      .adra(xt_rsc_0_11_adra),
      .adra_d(xt_rsc_0_11_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_11_i_da_d),
      .qa_d(xt_rsc_0_11_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_51_8_32_256_256_32_1_gen xt_rsc_0_12_i
      (
      .qb(xt_rsc_0_12_qb),
      .web(xt_rsc_0_12_web),
      .db(xt_rsc_0_12_db),
      .adrb(xt_rsc_0_12_adrb),
      .qa(xt_rsc_0_12_qa),
      .wea(xt_rsc_0_12_wea),
      .da(xt_rsc_0_12_da),
      .adra(xt_rsc_0_12_adra),
      .adra_d(xt_rsc_0_12_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_12_i_da_d),
      .qa_d(xt_rsc_0_12_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_52_8_32_256_256_32_1_gen xt_rsc_0_13_i
      (
      .qb(xt_rsc_0_13_qb),
      .web(xt_rsc_0_13_web),
      .db(xt_rsc_0_13_db),
      .adrb(xt_rsc_0_13_adrb),
      .qa(xt_rsc_0_13_qa),
      .wea(xt_rsc_0_13_wea),
      .da(xt_rsc_0_13_da),
      .adra(xt_rsc_0_13_adra),
      .adra_d(xt_rsc_0_13_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_13_i_da_d),
      .qa_d(xt_rsc_0_13_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_53_8_32_256_256_32_1_gen xt_rsc_0_14_i
      (
      .qb(xt_rsc_0_14_qb),
      .web(xt_rsc_0_14_web),
      .db(xt_rsc_0_14_db),
      .adrb(xt_rsc_0_14_adrb),
      .qa(xt_rsc_0_14_qa),
      .wea(xt_rsc_0_14_wea),
      .da(xt_rsc_0_14_da),
      .adra(xt_rsc_0_14_adra),
      .adra_d(xt_rsc_0_14_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_14_i_da_d),
      .qa_d(xt_rsc_0_14_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_54_8_32_256_256_32_1_gen xt_rsc_0_15_i
      (
      .qb(xt_rsc_0_15_qb),
      .web(xt_rsc_0_15_web),
      .db(xt_rsc_0_15_db),
      .adrb(xt_rsc_0_15_adrb),
      .qa(xt_rsc_0_15_qa),
      .wea(xt_rsc_0_15_wea),
      .da(xt_rsc_0_15_da),
      .adra(xt_rsc_0_15_adra),
      .adra_d(xt_rsc_0_15_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_15_i_da_d),
      .qa_d(xt_rsc_0_15_i_qa_d),
      .wea_d(xt_rsc_0_0_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_0_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_55_8_32_256_256_32_1_gen xt_rsc_0_16_i
      (
      .qb(xt_rsc_0_16_qb),
      .web(xt_rsc_0_16_web),
      .db(xt_rsc_0_16_db),
      .adrb(xt_rsc_0_16_adrb),
      .qa(xt_rsc_0_16_qa),
      .wea(xt_rsc_0_16_wea),
      .da(xt_rsc_0_16_da),
      .adra(xt_rsc_0_16_adra),
      .adra_d(xt_rsc_0_16_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_16_i_da_d),
      .qa_d(xt_rsc_0_16_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_56_8_32_256_256_32_1_gen xt_rsc_0_17_i
      (
      .qb(xt_rsc_0_17_qb),
      .web(xt_rsc_0_17_web),
      .db(xt_rsc_0_17_db),
      .adrb(xt_rsc_0_17_adrb),
      .qa(xt_rsc_0_17_qa),
      .wea(xt_rsc_0_17_wea),
      .da(xt_rsc_0_17_da),
      .adra(xt_rsc_0_17_adra),
      .adra_d(xt_rsc_0_17_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_17_i_da_d),
      .qa_d(xt_rsc_0_17_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_57_8_32_256_256_32_1_gen xt_rsc_0_18_i
      (
      .qb(xt_rsc_0_18_qb),
      .web(xt_rsc_0_18_web),
      .db(xt_rsc_0_18_db),
      .adrb(xt_rsc_0_18_adrb),
      .qa(xt_rsc_0_18_qa),
      .wea(xt_rsc_0_18_wea),
      .da(xt_rsc_0_18_da),
      .adra(xt_rsc_0_18_adra),
      .adra_d(xt_rsc_0_18_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_18_i_da_d),
      .qa_d(xt_rsc_0_18_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_58_8_32_256_256_32_1_gen xt_rsc_0_19_i
      (
      .qb(xt_rsc_0_19_qb),
      .web(xt_rsc_0_19_web),
      .db(xt_rsc_0_19_db),
      .adrb(xt_rsc_0_19_adrb),
      .qa(xt_rsc_0_19_qa),
      .wea(xt_rsc_0_19_wea),
      .da(xt_rsc_0_19_da),
      .adra(xt_rsc_0_19_adra),
      .adra_d(xt_rsc_0_19_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_19_i_da_d),
      .qa_d(xt_rsc_0_19_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_59_8_32_256_256_32_1_gen xt_rsc_0_20_i
      (
      .qb(xt_rsc_0_20_qb),
      .web(xt_rsc_0_20_web),
      .db(xt_rsc_0_20_db),
      .adrb(xt_rsc_0_20_adrb),
      .qa(xt_rsc_0_20_qa),
      .wea(xt_rsc_0_20_wea),
      .da(xt_rsc_0_20_da),
      .adra(xt_rsc_0_20_adra),
      .adra_d(xt_rsc_0_20_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_20_i_da_d),
      .qa_d(xt_rsc_0_20_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_60_8_32_256_256_32_1_gen xt_rsc_0_21_i
      (
      .qb(xt_rsc_0_21_qb),
      .web(xt_rsc_0_21_web),
      .db(xt_rsc_0_21_db),
      .adrb(xt_rsc_0_21_adrb),
      .qa(xt_rsc_0_21_qa),
      .wea(xt_rsc_0_21_wea),
      .da(xt_rsc_0_21_da),
      .adra(xt_rsc_0_21_adra),
      .adra_d(xt_rsc_0_21_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_21_i_da_d),
      .qa_d(xt_rsc_0_21_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_61_8_32_256_256_32_1_gen xt_rsc_0_22_i
      (
      .qb(xt_rsc_0_22_qb),
      .web(xt_rsc_0_22_web),
      .db(xt_rsc_0_22_db),
      .adrb(xt_rsc_0_22_adrb),
      .qa(xt_rsc_0_22_qa),
      .wea(xt_rsc_0_22_wea),
      .da(xt_rsc_0_22_da),
      .adra(xt_rsc_0_22_adra),
      .adra_d(xt_rsc_0_22_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_22_i_da_d),
      .qa_d(xt_rsc_0_22_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_62_8_32_256_256_32_1_gen xt_rsc_0_23_i
      (
      .qb(xt_rsc_0_23_qb),
      .web(xt_rsc_0_23_web),
      .db(xt_rsc_0_23_db),
      .adrb(xt_rsc_0_23_adrb),
      .qa(xt_rsc_0_23_qa),
      .wea(xt_rsc_0_23_wea),
      .da(xt_rsc_0_23_da),
      .adra(xt_rsc_0_23_adra),
      .adra_d(xt_rsc_0_23_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_23_i_da_d),
      .qa_d(xt_rsc_0_23_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_63_8_32_256_256_32_1_gen xt_rsc_0_24_i
      (
      .qb(xt_rsc_0_24_qb),
      .web(xt_rsc_0_24_web),
      .db(xt_rsc_0_24_db),
      .adrb(xt_rsc_0_24_adrb),
      .qa(xt_rsc_0_24_qa),
      .wea(xt_rsc_0_24_wea),
      .da(xt_rsc_0_24_da),
      .adra(xt_rsc_0_24_adra),
      .adra_d(xt_rsc_0_24_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_24_i_da_d),
      .qa_d(xt_rsc_0_24_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_64_8_32_256_256_32_1_gen xt_rsc_0_25_i
      (
      .qb(xt_rsc_0_25_qb),
      .web(xt_rsc_0_25_web),
      .db(xt_rsc_0_25_db),
      .adrb(xt_rsc_0_25_adrb),
      .qa(xt_rsc_0_25_qa),
      .wea(xt_rsc_0_25_wea),
      .da(xt_rsc_0_25_da),
      .adra(xt_rsc_0_25_adra),
      .adra_d(xt_rsc_0_25_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_25_i_da_d),
      .qa_d(xt_rsc_0_25_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_65_8_32_256_256_32_1_gen xt_rsc_0_26_i
      (
      .qb(xt_rsc_0_26_qb),
      .web(xt_rsc_0_26_web),
      .db(xt_rsc_0_26_db),
      .adrb(xt_rsc_0_26_adrb),
      .qa(xt_rsc_0_26_qa),
      .wea(xt_rsc_0_26_wea),
      .da(xt_rsc_0_26_da),
      .adra(xt_rsc_0_26_adra),
      .adra_d(xt_rsc_0_26_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_26_i_da_d),
      .qa_d(xt_rsc_0_26_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_66_8_32_256_256_32_1_gen xt_rsc_0_27_i
      (
      .qb(xt_rsc_0_27_qb),
      .web(xt_rsc_0_27_web),
      .db(xt_rsc_0_27_db),
      .adrb(xt_rsc_0_27_adrb),
      .qa(xt_rsc_0_27_qa),
      .wea(xt_rsc_0_27_wea),
      .da(xt_rsc_0_27_da),
      .adra(xt_rsc_0_27_adra),
      .adra_d(xt_rsc_0_27_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_27_i_da_d),
      .qa_d(xt_rsc_0_27_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_67_8_32_256_256_32_1_gen xt_rsc_0_28_i
      (
      .qb(xt_rsc_0_28_qb),
      .web(xt_rsc_0_28_web),
      .db(xt_rsc_0_28_db),
      .adrb(xt_rsc_0_28_adrb),
      .qa(xt_rsc_0_28_qa),
      .wea(xt_rsc_0_28_wea),
      .da(xt_rsc_0_28_da),
      .adra(xt_rsc_0_28_adra),
      .adra_d(xt_rsc_0_28_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_28_i_da_d),
      .qa_d(xt_rsc_0_28_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_68_8_32_256_256_32_1_gen xt_rsc_0_29_i
      (
      .qb(xt_rsc_0_29_qb),
      .web(xt_rsc_0_29_web),
      .db(xt_rsc_0_29_db),
      .adrb(xt_rsc_0_29_adrb),
      .qa(xt_rsc_0_29_qa),
      .wea(xt_rsc_0_29_wea),
      .da(xt_rsc_0_29_da),
      .adra(xt_rsc_0_29_adra),
      .adra_d(xt_rsc_0_29_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_29_i_da_d),
      .qa_d(xt_rsc_0_29_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_69_8_32_256_256_32_1_gen xt_rsc_0_30_i
      (
      .qb(xt_rsc_0_30_qb),
      .web(xt_rsc_0_30_web),
      .db(xt_rsc_0_30_db),
      .adrb(xt_rsc_0_30_adrb),
      .qa(xt_rsc_0_30_qa),
      .wea(xt_rsc_0_30_wea),
      .da(xt_rsc_0_30_da),
      .adra(xt_rsc_0_30_adra),
      .adra_d(xt_rsc_0_30_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_30_i_da_d),
      .qa_d(xt_rsc_0_30_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_70_8_32_256_256_32_1_gen xt_rsc_0_31_i
      (
      .qb(xt_rsc_0_31_qb),
      .web(xt_rsc_0_31_web),
      .db(xt_rsc_0_31_db),
      .adrb(xt_rsc_0_31_adrb),
      .qa(xt_rsc_0_31_qa),
      .wea(xt_rsc_0_31_wea),
      .da(xt_rsc_0_31_da),
      .adra(xt_rsc_0_31_adra),
      .adra_d(xt_rsc_0_31_i_adra_d),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(xt_rsc_0_31_i_da_d),
      .qa_d(xt_rsc_0_31_i_qa_d),
      .wea_d(xt_rsc_0_16_i_wea_d_iff),
      .rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(xt_rsc_0_16_i_wea_d_iff)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_71_8_32_256_256_32_1_gen twiddle_rsc_0_0_i
      (
      .qb(twiddle_rsc_0_0_qb),
      .web(twiddle_rsc_0_0_web),
      .db(twiddle_rsc_0_0_db),
      .adrb(twiddle_rsc_0_0_adrb),
      .qa(twiddle_rsc_0_0_qa),
      .wea(twiddle_rsc_0_0_wea),
      .da(twiddle_rsc_0_0_da),
      .adra(twiddle_rsc_0_0_adra),
      .adra_d(nl_twiddle_rsc_0_0_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_0_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_72_8_32_256_256_32_1_gen twiddle_rsc_0_1_i
      (
      .qb(twiddle_rsc_0_1_qb),
      .web(twiddle_rsc_0_1_web),
      .db(twiddle_rsc_0_1_db),
      .adrb(twiddle_rsc_0_1_adrb),
      .qa(twiddle_rsc_0_1_qa),
      .wea(twiddle_rsc_0_1_wea),
      .da(twiddle_rsc_0_1_da),
      .adra(twiddle_rsc_0_1_adra),
      .adra_d(nl_twiddle_rsc_0_1_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_1_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_73_8_32_256_256_32_1_gen twiddle_rsc_0_2_i
      (
      .qb(twiddle_rsc_0_2_qb),
      .web(twiddle_rsc_0_2_web),
      .db(twiddle_rsc_0_2_db),
      .adrb(twiddle_rsc_0_2_adrb),
      .qa(twiddle_rsc_0_2_qa),
      .wea(twiddle_rsc_0_2_wea),
      .da(twiddle_rsc_0_2_da),
      .adra(twiddle_rsc_0_2_adra),
      .adra_d(nl_twiddle_rsc_0_2_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_2_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_74_8_32_256_256_32_1_gen twiddle_rsc_0_3_i
      (
      .qb(twiddle_rsc_0_3_qb),
      .web(twiddle_rsc_0_3_web),
      .db(twiddle_rsc_0_3_db),
      .adrb(twiddle_rsc_0_3_adrb),
      .qa(twiddle_rsc_0_3_qa),
      .wea(twiddle_rsc_0_3_wea),
      .da(twiddle_rsc_0_3_da),
      .adra(twiddle_rsc_0_3_adra),
      .adra_d(nl_twiddle_rsc_0_3_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_3_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_75_8_32_256_256_32_1_gen twiddle_rsc_0_4_i
      (
      .qb(twiddle_rsc_0_4_qb),
      .web(twiddle_rsc_0_4_web),
      .db(twiddle_rsc_0_4_db),
      .adrb(twiddle_rsc_0_4_adrb),
      .qa(twiddle_rsc_0_4_qa),
      .wea(twiddle_rsc_0_4_wea),
      .da(twiddle_rsc_0_4_da),
      .adra(twiddle_rsc_0_4_adra),
      .adra_d(nl_twiddle_rsc_0_4_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_4_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_76_8_32_256_256_32_1_gen twiddle_rsc_0_5_i
      (
      .qb(twiddle_rsc_0_5_qb),
      .web(twiddle_rsc_0_5_web),
      .db(twiddle_rsc_0_5_db),
      .adrb(twiddle_rsc_0_5_adrb),
      .qa(twiddle_rsc_0_5_qa),
      .wea(twiddle_rsc_0_5_wea),
      .da(twiddle_rsc_0_5_da),
      .adra(twiddle_rsc_0_5_adra),
      .adra_d(nl_twiddle_rsc_0_5_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_5_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_77_8_32_256_256_32_1_gen twiddle_rsc_0_6_i
      (
      .qb(twiddle_rsc_0_6_qb),
      .web(twiddle_rsc_0_6_web),
      .db(twiddle_rsc_0_6_db),
      .adrb(twiddle_rsc_0_6_adrb),
      .qa(twiddle_rsc_0_6_qa),
      .wea(twiddle_rsc_0_6_wea),
      .da(twiddle_rsc_0_6_da),
      .adra(twiddle_rsc_0_6_adra),
      .adra_d(nl_twiddle_rsc_0_6_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_6_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_78_8_32_256_256_32_1_gen twiddle_rsc_0_7_i
      (
      .qb(twiddle_rsc_0_7_qb),
      .web(twiddle_rsc_0_7_web),
      .db(twiddle_rsc_0_7_db),
      .adrb(twiddle_rsc_0_7_adrb),
      .qa(twiddle_rsc_0_7_qa),
      .wea(twiddle_rsc_0_7_wea),
      .da(twiddle_rsc_0_7_da),
      .adra(twiddle_rsc_0_7_adra),
      .adra_d(nl_twiddle_rsc_0_7_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_7_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_79_8_32_256_256_32_1_gen twiddle_rsc_0_8_i
      (
      .qb(twiddle_rsc_0_8_qb),
      .web(twiddle_rsc_0_8_web),
      .db(twiddle_rsc_0_8_db),
      .adrb(twiddle_rsc_0_8_adrb),
      .qa(twiddle_rsc_0_8_qa),
      .wea(twiddle_rsc_0_8_wea),
      .da(twiddle_rsc_0_8_da),
      .adra(twiddle_rsc_0_8_adra),
      .adra_d(nl_twiddle_rsc_0_8_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_8_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_80_8_32_256_256_32_1_gen twiddle_rsc_0_9_i
      (
      .qb(twiddle_rsc_0_9_qb),
      .web(twiddle_rsc_0_9_web),
      .db(twiddle_rsc_0_9_db),
      .adrb(twiddle_rsc_0_9_adrb),
      .qa(twiddle_rsc_0_9_qa),
      .wea(twiddle_rsc_0_9_wea),
      .da(twiddle_rsc_0_9_da),
      .adra(twiddle_rsc_0_9_adra),
      .adra_d(nl_twiddle_rsc_0_9_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_9_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_81_8_32_256_256_32_1_gen twiddle_rsc_0_10_i
      (
      .qb(twiddle_rsc_0_10_qb),
      .web(twiddle_rsc_0_10_web),
      .db(twiddle_rsc_0_10_db),
      .adrb(twiddle_rsc_0_10_adrb),
      .qa(twiddle_rsc_0_10_qa),
      .wea(twiddle_rsc_0_10_wea),
      .da(twiddle_rsc_0_10_da),
      .adra(twiddle_rsc_0_10_adra),
      .adra_d(nl_twiddle_rsc_0_10_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_10_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_82_8_32_256_256_32_1_gen twiddle_rsc_0_11_i
      (
      .qb(twiddle_rsc_0_11_qb),
      .web(twiddle_rsc_0_11_web),
      .db(twiddle_rsc_0_11_db),
      .adrb(twiddle_rsc_0_11_adrb),
      .qa(twiddle_rsc_0_11_qa),
      .wea(twiddle_rsc_0_11_wea),
      .da(twiddle_rsc_0_11_da),
      .adra(twiddle_rsc_0_11_adra),
      .adra_d(nl_twiddle_rsc_0_11_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_11_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_83_8_32_256_256_32_1_gen twiddle_rsc_0_12_i
      (
      .qb(twiddle_rsc_0_12_qb),
      .web(twiddle_rsc_0_12_web),
      .db(twiddle_rsc_0_12_db),
      .adrb(twiddle_rsc_0_12_adrb),
      .qa(twiddle_rsc_0_12_qa),
      .wea(twiddle_rsc_0_12_wea),
      .da(twiddle_rsc_0_12_da),
      .adra(twiddle_rsc_0_12_adra),
      .adra_d(nl_twiddle_rsc_0_12_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_12_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_84_8_32_256_256_32_1_gen twiddle_rsc_0_13_i
      (
      .qb(twiddle_rsc_0_13_qb),
      .web(twiddle_rsc_0_13_web),
      .db(twiddle_rsc_0_13_db),
      .adrb(twiddle_rsc_0_13_adrb),
      .qa(twiddle_rsc_0_13_qa),
      .wea(twiddle_rsc_0_13_wea),
      .da(twiddle_rsc_0_13_da),
      .adra(twiddle_rsc_0_13_adra),
      .adra_d(nl_twiddle_rsc_0_13_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_13_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_85_8_32_256_256_32_1_gen twiddle_rsc_0_14_i
      (
      .qb(twiddle_rsc_0_14_qb),
      .web(twiddle_rsc_0_14_web),
      .db(twiddle_rsc_0_14_db),
      .adrb(twiddle_rsc_0_14_adrb),
      .qa(twiddle_rsc_0_14_qa),
      .wea(twiddle_rsc_0_14_wea),
      .da(twiddle_rsc_0_14_da),
      .adra(twiddle_rsc_0_14_adra),
      .adra_d(nl_twiddle_rsc_0_14_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_14_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_86_8_32_256_256_32_1_gen twiddle_rsc_0_15_i
      (
      .qb(twiddle_rsc_0_15_qb),
      .web(twiddle_rsc_0_15_web),
      .db(twiddle_rsc_0_15_db),
      .adrb(twiddle_rsc_0_15_adrb),
      .qa(twiddle_rsc_0_15_qa),
      .wea(twiddle_rsc_0_15_wea),
      .da(twiddle_rsc_0_15_da),
      .adra(twiddle_rsc_0_15_adra),
      .adra_d(nl_twiddle_rsc_0_15_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_rsc_0_15_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_87_8_32_256_256_32_1_gen twiddle_h_rsc_0_0_i
      (
      .qb(twiddle_h_rsc_0_0_qb),
      .web(twiddle_h_rsc_0_0_web),
      .db(twiddle_h_rsc_0_0_db),
      .adrb(twiddle_h_rsc_0_0_adrb),
      .qa(twiddle_h_rsc_0_0_qa),
      .wea(twiddle_h_rsc_0_0_wea),
      .da(twiddle_h_rsc_0_0_da),
      .adra(twiddle_h_rsc_0_0_adra),
      .adra_d(nl_twiddle_h_rsc_0_0_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_0_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_88_8_32_256_256_32_1_gen twiddle_h_rsc_0_1_i
      (
      .qb(twiddle_h_rsc_0_1_qb),
      .web(twiddle_h_rsc_0_1_web),
      .db(twiddle_h_rsc_0_1_db),
      .adrb(twiddle_h_rsc_0_1_adrb),
      .qa(twiddle_h_rsc_0_1_qa),
      .wea(twiddle_h_rsc_0_1_wea),
      .da(twiddle_h_rsc_0_1_da),
      .adra(twiddle_h_rsc_0_1_adra),
      .adra_d(nl_twiddle_h_rsc_0_1_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_1_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_89_8_32_256_256_32_1_gen twiddle_h_rsc_0_2_i
      (
      .qb(twiddle_h_rsc_0_2_qb),
      .web(twiddle_h_rsc_0_2_web),
      .db(twiddle_h_rsc_0_2_db),
      .adrb(twiddle_h_rsc_0_2_adrb),
      .qa(twiddle_h_rsc_0_2_qa),
      .wea(twiddle_h_rsc_0_2_wea),
      .da(twiddle_h_rsc_0_2_da),
      .adra(twiddle_h_rsc_0_2_adra),
      .adra_d(nl_twiddle_h_rsc_0_2_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_2_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_90_8_32_256_256_32_1_gen twiddle_h_rsc_0_3_i
      (
      .qb(twiddle_h_rsc_0_3_qb),
      .web(twiddle_h_rsc_0_3_web),
      .db(twiddle_h_rsc_0_3_db),
      .adrb(twiddle_h_rsc_0_3_adrb),
      .qa(twiddle_h_rsc_0_3_qa),
      .wea(twiddle_h_rsc_0_3_wea),
      .da(twiddle_h_rsc_0_3_da),
      .adra(twiddle_h_rsc_0_3_adra),
      .adra_d(nl_twiddle_h_rsc_0_3_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_3_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_91_8_32_256_256_32_1_gen twiddle_h_rsc_0_4_i
      (
      .qb(twiddle_h_rsc_0_4_qb),
      .web(twiddle_h_rsc_0_4_web),
      .db(twiddle_h_rsc_0_4_db),
      .adrb(twiddle_h_rsc_0_4_adrb),
      .qa(twiddle_h_rsc_0_4_qa),
      .wea(twiddle_h_rsc_0_4_wea),
      .da(twiddle_h_rsc_0_4_da),
      .adra(twiddle_h_rsc_0_4_adra),
      .adra_d(nl_twiddle_h_rsc_0_4_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_4_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_92_8_32_256_256_32_1_gen twiddle_h_rsc_0_5_i
      (
      .qb(twiddle_h_rsc_0_5_qb),
      .web(twiddle_h_rsc_0_5_web),
      .db(twiddle_h_rsc_0_5_db),
      .adrb(twiddle_h_rsc_0_5_adrb),
      .qa(twiddle_h_rsc_0_5_qa),
      .wea(twiddle_h_rsc_0_5_wea),
      .da(twiddle_h_rsc_0_5_da),
      .adra(twiddle_h_rsc_0_5_adra),
      .adra_d(nl_twiddle_h_rsc_0_5_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_5_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_93_8_32_256_256_32_1_gen twiddle_h_rsc_0_6_i
      (
      .qb(twiddle_h_rsc_0_6_qb),
      .web(twiddle_h_rsc_0_6_web),
      .db(twiddle_h_rsc_0_6_db),
      .adrb(twiddle_h_rsc_0_6_adrb),
      .qa(twiddle_h_rsc_0_6_qa),
      .wea(twiddle_h_rsc_0_6_wea),
      .da(twiddle_h_rsc_0_6_da),
      .adra(twiddle_h_rsc_0_6_adra),
      .adra_d(nl_twiddle_h_rsc_0_6_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_6_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_94_8_32_256_256_32_1_gen twiddle_h_rsc_0_7_i
      (
      .qb(twiddle_h_rsc_0_7_qb),
      .web(twiddle_h_rsc_0_7_web),
      .db(twiddle_h_rsc_0_7_db),
      .adrb(twiddle_h_rsc_0_7_adrb),
      .qa(twiddle_h_rsc_0_7_qa),
      .wea(twiddle_h_rsc_0_7_wea),
      .da(twiddle_h_rsc_0_7_da),
      .adra(twiddle_h_rsc_0_7_adra),
      .adra_d(nl_twiddle_h_rsc_0_7_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_7_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_95_8_32_256_256_32_1_gen twiddle_h_rsc_0_8_i
      (
      .qb(twiddle_h_rsc_0_8_qb),
      .web(twiddle_h_rsc_0_8_web),
      .db(twiddle_h_rsc_0_8_db),
      .adrb(twiddle_h_rsc_0_8_adrb),
      .qa(twiddle_h_rsc_0_8_qa),
      .wea(twiddle_h_rsc_0_8_wea),
      .da(twiddle_h_rsc_0_8_da),
      .adra(twiddle_h_rsc_0_8_adra),
      .adra_d(nl_twiddle_h_rsc_0_8_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_8_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_96_8_32_256_256_32_1_gen twiddle_h_rsc_0_9_i
      (
      .qb(twiddle_h_rsc_0_9_qb),
      .web(twiddle_h_rsc_0_9_web),
      .db(twiddle_h_rsc_0_9_db),
      .adrb(twiddle_h_rsc_0_9_adrb),
      .qa(twiddle_h_rsc_0_9_qa),
      .wea(twiddle_h_rsc_0_9_wea),
      .da(twiddle_h_rsc_0_9_da),
      .adra(twiddle_h_rsc_0_9_adra),
      .adra_d(nl_twiddle_h_rsc_0_9_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_9_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_97_8_32_256_256_32_1_gen twiddle_h_rsc_0_10_i
      (
      .qb(twiddle_h_rsc_0_10_qb),
      .web(twiddle_h_rsc_0_10_web),
      .db(twiddle_h_rsc_0_10_db),
      .adrb(twiddle_h_rsc_0_10_adrb),
      .qa(twiddle_h_rsc_0_10_qa),
      .wea(twiddle_h_rsc_0_10_wea),
      .da(twiddle_h_rsc_0_10_da),
      .adra(twiddle_h_rsc_0_10_adra),
      .adra_d(nl_twiddle_h_rsc_0_10_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_10_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_98_8_32_256_256_32_1_gen twiddle_h_rsc_0_11_i
      (
      .qb(twiddle_h_rsc_0_11_qb),
      .web(twiddle_h_rsc_0_11_web),
      .db(twiddle_h_rsc_0_11_db),
      .adrb(twiddle_h_rsc_0_11_adrb),
      .qa(twiddle_h_rsc_0_11_qa),
      .wea(twiddle_h_rsc_0_11_wea),
      .da(twiddle_h_rsc_0_11_da),
      .adra(twiddle_h_rsc_0_11_adra),
      .adra_d(nl_twiddle_h_rsc_0_11_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_11_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_99_8_32_256_256_32_1_gen twiddle_h_rsc_0_12_i
      (
      .qb(twiddle_h_rsc_0_12_qb),
      .web(twiddle_h_rsc_0_12_web),
      .db(twiddle_h_rsc_0_12_db),
      .adrb(twiddle_h_rsc_0_12_adrb),
      .qa(twiddle_h_rsc_0_12_qa),
      .wea(twiddle_h_rsc_0_12_wea),
      .da(twiddle_h_rsc_0_12_da),
      .adra(twiddle_h_rsc_0_12_adra),
      .adra_d(nl_twiddle_h_rsc_0_12_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_12_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_100_8_32_256_256_32_1_gen twiddle_h_rsc_0_13_i
      (
      .qb(twiddle_h_rsc_0_13_qb),
      .web(twiddle_h_rsc_0_13_web),
      .db(twiddle_h_rsc_0_13_db),
      .adrb(twiddle_h_rsc_0_13_adrb),
      .qa(twiddle_h_rsc_0_13_qa),
      .wea(twiddle_h_rsc_0_13_wea),
      .da(twiddle_h_rsc_0_13_da),
      .adra(twiddle_h_rsc_0_13_adra),
      .adra_d(nl_twiddle_h_rsc_0_13_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_13_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_101_8_32_256_256_32_1_gen twiddle_h_rsc_0_14_i
      (
      .qb(twiddle_h_rsc_0_14_qb),
      .web(twiddle_h_rsc_0_14_web),
      .db(twiddle_h_rsc_0_14_db),
      .adrb(twiddle_h_rsc_0_14_adrb),
      .qa(twiddle_h_rsc_0_14_qa),
      .wea(twiddle_h_rsc_0_14_wea),
      .da(twiddle_h_rsc_0_14_da),
      .adra(twiddle_h_rsc_0_14_adra),
      .adra_d(nl_twiddle_h_rsc_0_14_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_14_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_Xilinx_RAMS_BLOCK_DPRAM_RBW_DUAL_rwport_102_8_32_256_256_32_1_gen twiddle_h_rsc_0_15_i
      (
      .qb(twiddle_h_rsc_0_15_qb),
      .web(twiddle_h_rsc_0_15_web),
      .db(twiddle_h_rsc_0_15_db),
      .adrb(twiddle_h_rsc_0_15_adrb),
      .qa(twiddle_h_rsc_0_15_qa),
      .wea(twiddle_h_rsc_0_15_wea),
      .da(twiddle_h_rsc_0_15_da),
      .adra(twiddle_h_rsc_0_15_adra),
      .adra_d(nl_twiddle_h_rsc_0_15_i_adra_d[15:0]),
      .clka(clk),
      .clka_en(1'b1),
      .da_d(64'b0000000000000000000000000000000000000000000000000000000000000000),
      .qa_d(twiddle_h_rsc_0_15_i_qa_d),
      .wea_d(2'b00),
      .rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .rwA_rw_ram_ir_internal_WMASK_B_d(2'b00)
    );
  peaseNTT_core peaseNTT_core_inst (
      .clk(clk),
      .rst(rst),
      .xt_rsc_triosy_0_0_lz(xt_rsc_triosy_0_0_lz),
      .xt_rsc_triosy_0_1_lz(xt_rsc_triosy_0_1_lz),
      .xt_rsc_triosy_0_2_lz(xt_rsc_triosy_0_2_lz),
      .xt_rsc_triosy_0_3_lz(xt_rsc_triosy_0_3_lz),
      .xt_rsc_triosy_0_4_lz(xt_rsc_triosy_0_4_lz),
      .xt_rsc_triosy_0_5_lz(xt_rsc_triosy_0_5_lz),
      .xt_rsc_triosy_0_6_lz(xt_rsc_triosy_0_6_lz),
      .xt_rsc_triosy_0_7_lz(xt_rsc_triosy_0_7_lz),
      .xt_rsc_triosy_0_8_lz(xt_rsc_triosy_0_8_lz),
      .xt_rsc_triosy_0_9_lz(xt_rsc_triosy_0_9_lz),
      .xt_rsc_triosy_0_10_lz(xt_rsc_triosy_0_10_lz),
      .xt_rsc_triosy_0_11_lz(xt_rsc_triosy_0_11_lz),
      .xt_rsc_triosy_0_12_lz(xt_rsc_triosy_0_12_lz),
      .xt_rsc_triosy_0_13_lz(xt_rsc_triosy_0_13_lz),
      .xt_rsc_triosy_0_14_lz(xt_rsc_triosy_0_14_lz),
      .xt_rsc_triosy_0_15_lz(xt_rsc_triosy_0_15_lz),
      .xt_rsc_triosy_0_16_lz(xt_rsc_triosy_0_16_lz),
      .xt_rsc_triosy_0_17_lz(xt_rsc_triosy_0_17_lz),
      .xt_rsc_triosy_0_18_lz(xt_rsc_triosy_0_18_lz),
      .xt_rsc_triosy_0_19_lz(xt_rsc_triosy_0_19_lz),
      .xt_rsc_triosy_0_20_lz(xt_rsc_triosy_0_20_lz),
      .xt_rsc_triosy_0_21_lz(xt_rsc_triosy_0_21_lz),
      .xt_rsc_triosy_0_22_lz(xt_rsc_triosy_0_22_lz),
      .xt_rsc_triosy_0_23_lz(xt_rsc_triosy_0_23_lz),
      .xt_rsc_triosy_0_24_lz(xt_rsc_triosy_0_24_lz),
      .xt_rsc_triosy_0_25_lz(xt_rsc_triosy_0_25_lz),
      .xt_rsc_triosy_0_26_lz(xt_rsc_triosy_0_26_lz),
      .xt_rsc_triosy_0_27_lz(xt_rsc_triosy_0_27_lz),
      .xt_rsc_triosy_0_28_lz(xt_rsc_triosy_0_28_lz),
      .xt_rsc_triosy_0_29_lz(xt_rsc_triosy_0_29_lz),
      .xt_rsc_triosy_0_30_lz(xt_rsc_triosy_0_30_lz),
      .xt_rsc_triosy_0_31_lz(xt_rsc_triosy_0_31_lz),
      .p_rsc_dat(p_rsc_dat),
      .p_rsc_triosy_lz(p_rsc_triosy_lz),
      .r_rsc_triosy_lz(r_rsc_triosy_lz),
      .twiddle_rsc_triosy_0_0_lz(twiddle_rsc_triosy_0_0_lz),
      .twiddle_rsc_triosy_0_1_lz(twiddle_rsc_triosy_0_1_lz),
      .twiddle_rsc_triosy_0_2_lz(twiddle_rsc_triosy_0_2_lz),
      .twiddle_rsc_triosy_0_3_lz(twiddle_rsc_triosy_0_3_lz),
      .twiddle_rsc_triosy_0_4_lz(twiddle_rsc_triosy_0_4_lz),
      .twiddle_rsc_triosy_0_5_lz(twiddle_rsc_triosy_0_5_lz),
      .twiddle_rsc_triosy_0_6_lz(twiddle_rsc_triosy_0_6_lz),
      .twiddle_rsc_triosy_0_7_lz(twiddle_rsc_triosy_0_7_lz),
      .twiddle_rsc_triosy_0_8_lz(twiddle_rsc_triosy_0_8_lz),
      .twiddle_rsc_triosy_0_9_lz(twiddle_rsc_triosy_0_9_lz),
      .twiddle_rsc_triosy_0_10_lz(twiddle_rsc_triosy_0_10_lz),
      .twiddle_rsc_triosy_0_11_lz(twiddle_rsc_triosy_0_11_lz),
      .twiddle_rsc_triosy_0_12_lz(twiddle_rsc_triosy_0_12_lz),
      .twiddle_rsc_triosy_0_13_lz(twiddle_rsc_triosy_0_13_lz),
      .twiddle_rsc_triosy_0_14_lz(twiddle_rsc_triosy_0_14_lz),
      .twiddle_rsc_triosy_0_15_lz(twiddle_rsc_triosy_0_15_lz),
      .twiddle_h_rsc_triosy_0_0_lz(twiddle_h_rsc_triosy_0_0_lz),
      .twiddle_h_rsc_triosy_0_1_lz(twiddle_h_rsc_triosy_0_1_lz),
      .twiddle_h_rsc_triosy_0_2_lz(twiddle_h_rsc_triosy_0_2_lz),
      .twiddle_h_rsc_triosy_0_3_lz(twiddle_h_rsc_triosy_0_3_lz),
      .twiddle_h_rsc_triosy_0_4_lz(twiddle_h_rsc_triosy_0_4_lz),
      .twiddle_h_rsc_triosy_0_5_lz(twiddle_h_rsc_triosy_0_5_lz),
      .twiddle_h_rsc_triosy_0_6_lz(twiddle_h_rsc_triosy_0_6_lz),
      .twiddle_h_rsc_triosy_0_7_lz(twiddle_h_rsc_triosy_0_7_lz),
      .twiddle_h_rsc_triosy_0_8_lz(twiddle_h_rsc_triosy_0_8_lz),
      .twiddle_h_rsc_triosy_0_9_lz(twiddle_h_rsc_triosy_0_9_lz),
      .twiddle_h_rsc_triosy_0_10_lz(twiddle_h_rsc_triosy_0_10_lz),
      .twiddle_h_rsc_triosy_0_11_lz(twiddle_h_rsc_triosy_0_11_lz),
      .twiddle_h_rsc_triosy_0_12_lz(twiddle_h_rsc_triosy_0_12_lz),
      .twiddle_h_rsc_triosy_0_13_lz(twiddle_h_rsc_triosy_0_13_lz),
      .twiddle_h_rsc_triosy_0_14_lz(twiddle_h_rsc_triosy_0_14_lz),
      .twiddle_h_rsc_triosy_0_15_lz(twiddle_h_rsc_triosy_0_15_lz),
      .yt_rsc_0_0_i_adra_d(yt_rsc_0_0_i_adra_d),
      .yt_rsc_0_0_i_clka_en_d(yt_rsc_0_0_i_clka_en_d),
      .yt_rsc_0_0_i_da_d(yt_rsc_0_0_i_da_d),
      .yt_rsc_0_0_i_qa_d(yt_rsc_0_0_i_qa_d),
      .yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_1_i_adra_d(yt_rsc_0_1_i_adra_d),
      .yt_rsc_0_1_i_da_d(yt_rsc_0_1_i_da_d),
      .yt_rsc_0_1_i_qa_d(yt_rsc_0_1_i_qa_d),
      .yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_2_i_adra_d(yt_rsc_0_2_i_adra_d),
      .yt_rsc_0_2_i_da_d(yt_rsc_0_2_i_da_d),
      .yt_rsc_0_2_i_qa_d(yt_rsc_0_2_i_qa_d),
      .yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_3_i_adra_d(yt_rsc_0_3_i_adra_d),
      .yt_rsc_0_3_i_da_d(yt_rsc_0_3_i_da_d),
      .yt_rsc_0_3_i_qa_d(yt_rsc_0_3_i_qa_d),
      .yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_4_i_adra_d(yt_rsc_0_4_i_adra_d),
      .yt_rsc_0_4_i_da_d(yt_rsc_0_4_i_da_d),
      .yt_rsc_0_4_i_qa_d(yt_rsc_0_4_i_qa_d),
      .yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_5_i_adra_d(yt_rsc_0_5_i_adra_d),
      .yt_rsc_0_5_i_da_d(yt_rsc_0_5_i_da_d),
      .yt_rsc_0_5_i_qa_d(yt_rsc_0_5_i_qa_d),
      .yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_6_i_adra_d(yt_rsc_0_6_i_adra_d),
      .yt_rsc_0_6_i_da_d(yt_rsc_0_6_i_da_d),
      .yt_rsc_0_6_i_qa_d(yt_rsc_0_6_i_qa_d),
      .yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_7_i_adra_d(yt_rsc_0_7_i_adra_d),
      .yt_rsc_0_7_i_da_d(yt_rsc_0_7_i_da_d),
      .yt_rsc_0_7_i_qa_d(yt_rsc_0_7_i_qa_d),
      .yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_8_i_adra_d(yt_rsc_0_8_i_adra_d),
      .yt_rsc_0_8_i_da_d(yt_rsc_0_8_i_da_d),
      .yt_rsc_0_8_i_qa_d(yt_rsc_0_8_i_qa_d),
      .yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_9_i_adra_d(yt_rsc_0_9_i_adra_d),
      .yt_rsc_0_9_i_da_d(yt_rsc_0_9_i_da_d),
      .yt_rsc_0_9_i_qa_d(yt_rsc_0_9_i_qa_d),
      .yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_10_i_adra_d(yt_rsc_0_10_i_adra_d),
      .yt_rsc_0_10_i_da_d(yt_rsc_0_10_i_da_d),
      .yt_rsc_0_10_i_qa_d(yt_rsc_0_10_i_qa_d),
      .yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_11_i_adra_d(yt_rsc_0_11_i_adra_d),
      .yt_rsc_0_11_i_da_d(yt_rsc_0_11_i_da_d),
      .yt_rsc_0_11_i_qa_d(yt_rsc_0_11_i_qa_d),
      .yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_12_i_adra_d(yt_rsc_0_12_i_adra_d),
      .yt_rsc_0_12_i_da_d(yt_rsc_0_12_i_da_d),
      .yt_rsc_0_12_i_qa_d(yt_rsc_0_12_i_qa_d),
      .yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_13_i_adra_d(yt_rsc_0_13_i_adra_d),
      .yt_rsc_0_13_i_da_d(yt_rsc_0_13_i_da_d),
      .yt_rsc_0_13_i_qa_d(yt_rsc_0_13_i_qa_d),
      .yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_14_i_adra_d(yt_rsc_0_14_i_adra_d),
      .yt_rsc_0_14_i_da_d(yt_rsc_0_14_i_da_d),
      .yt_rsc_0_14_i_qa_d(yt_rsc_0_14_i_qa_d),
      .yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_15_i_adra_d(yt_rsc_0_15_i_adra_d),
      .yt_rsc_0_15_i_da_d(yt_rsc_0_15_i_da_d),
      .yt_rsc_0_15_i_qa_d(yt_rsc_0_15_i_qa_d),
      .yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_16_i_adra_d(yt_rsc_0_16_i_adra_d),
      .yt_rsc_0_16_i_clka_en_d(yt_rsc_0_16_i_clka_en_d),
      .yt_rsc_0_16_i_da_d(yt_rsc_0_16_i_da_d),
      .yt_rsc_0_16_i_qa_d(yt_rsc_0_16_i_qa_d),
      .yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_17_i_adra_d(yt_rsc_0_17_i_adra_d),
      .yt_rsc_0_17_i_da_d(yt_rsc_0_17_i_da_d),
      .yt_rsc_0_17_i_qa_d(yt_rsc_0_17_i_qa_d),
      .yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_18_i_adra_d(yt_rsc_0_18_i_adra_d),
      .yt_rsc_0_18_i_da_d(yt_rsc_0_18_i_da_d),
      .yt_rsc_0_18_i_qa_d(yt_rsc_0_18_i_qa_d),
      .yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_19_i_adra_d(yt_rsc_0_19_i_adra_d),
      .yt_rsc_0_19_i_da_d(yt_rsc_0_19_i_da_d),
      .yt_rsc_0_19_i_qa_d(yt_rsc_0_19_i_qa_d),
      .yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_20_i_adra_d(yt_rsc_0_20_i_adra_d),
      .yt_rsc_0_20_i_da_d(yt_rsc_0_20_i_da_d),
      .yt_rsc_0_20_i_qa_d(yt_rsc_0_20_i_qa_d),
      .yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_21_i_adra_d(yt_rsc_0_21_i_adra_d),
      .yt_rsc_0_21_i_da_d(yt_rsc_0_21_i_da_d),
      .yt_rsc_0_21_i_qa_d(yt_rsc_0_21_i_qa_d),
      .yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_22_i_adra_d(yt_rsc_0_22_i_adra_d),
      .yt_rsc_0_22_i_da_d(yt_rsc_0_22_i_da_d),
      .yt_rsc_0_22_i_qa_d(yt_rsc_0_22_i_qa_d),
      .yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_23_i_adra_d(yt_rsc_0_23_i_adra_d),
      .yt_rsc_0_23_i_da_d(yt_rsc_0_23_i_da_d),
      .yt_rsc_0_23_i_qa_d(yt_rsc_0_23_i_qa_d),
      .yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_24_i_adra_d(yt_rsc_0_24_i_adra_d),
      .yt_rsc_0_24_i_da_d(yt_rsc_0_24_i_da_d),
      .yt_rsc_0_24_i_qa_d(yt_rsc_0_24_i_qa_d),
      .yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_25_i_adra_d(yt_rsc_0_25_i_adra_d),
      .yt_rsc_0_25_i_da_d(yt_rsc_0_25_i_da_d),
      .yt_rsc_0_25_i_qa_d(yt_rsc_0_25_i_qa_d),
      .yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_26_i_adra_d(yt_rsc_0_26_i_adra_d),
      .yt_rsc_0_26_i_da_d(yt_rsc_0_26_i_da_d),
      .yt_rsc_0_26_i_qa_d(yt_rsc_0_26_i_qa_d),
      .yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_27_i_adra_d(yt_rsc_0_27_i_adra_d),
      .yt_rsc_0_27_i_da_d(yt_rsc_0_27_i_da_d),
      .yt_rsc_0_27_i_qa_d(yt_rsc_0_27_i_qa_d),
      .yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_28_i_adra_d(yt_rsc_0_28_i_adra_d),
      .yt_rsc_0_28_i_da_d(yt_rsc_0_28_i_da_d),
      .yt_rsc_0_28_i_qa_d(yt_rsc_0_28_i_qa_d),
      .yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_29_i_adra_d(yt_rsc_0_29_i_adra_d),
      .yt_rsc_0_29_i_da_d(yt_rsc_0_29_i_da_d),
      .yt_rsc_0_29_i_qa_d(yt_rsc_0_29_i_qa_d),
      .yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_30_i_adra_d(yt_rsc_0_30_i_adra_d),
      .yt_rsc_0_30_i_da_d(yt_rsc_0_30_i_da_d),
      .yt_rsc_0_30_i_qa_d(yt_rsc_0_30_i_qa_d),
      .yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_31_i_adra_d(yt_rsc_0_31_i_adra_d),
      .yt_rsc_0_31_i_da_d(yt_rsc_0_31_i_da_d),
      .yt_rsc_0_31_i_qa_d(yt_rsc_0_31_i_qa_d),
      .yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d(yt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_0_i_adra_d(xt_rsc_0_0_i_adra_d),
      .xt_rsc_0_0_i_da_d(xt_rsc_0_0_i_da_d),
      .xt_rsc_0_0_i_qa_d(xt_rsc_0_0_i_qa_d),
      .xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_1_i_adra_d(xt_rsc_0_1_i_adra_d),
      .xt_rsc_0_1_i_da_d(xt_rsc_0_1_i_da_d),
      .xt_rsc_0_1_i_qa_d(xt_rsc_0_1_i_qa_d),
      .xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_2_i_adra_d(xt_rsc_0_2_i_adra_d),
      .xt_rsc_0_2_i_da_d(xt_rsc_0_2_i_da_d),
      .xt_rsc_0_2_i_qa_d(xt_rsc_0_2_i_qa_d),
      .xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_3_i_adra_d(xt_rsc_0_3_i_adra_d),
      .xt_rsc_0_3_i_da_d(xt_rsc_0_3_i_da_d),
      .xt_rsc_0_3_i_qa_d(xt_rsc_0_3_i_qa_d),
      .xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_4_i_adra_d(xt_rsc_0_4_i_adra_d),
      .xt_rsc_0_4_i_da_d(xt_rsc_0_4_i_da_d),
      .xt_rsc_0_4_i_qa_d(xt_rsc_0_4_i_qa_d),
      .xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_5_i_adra_d(xt_rsc_0_5_i_adra_d),
      .xt_rsc_0_5_i_da_d(xt_rsc_0_5_i_da_d),
      .xt_rsc_0_5_i_qa_d(xt_rsc_0_5_i_qa_d),
      .xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_6_i_adra_d(xt_rsc_0_6_i_adra_d),
      .xt_rsc_0_6_i_da_d(xt_rsc_0_6_i_da_d),
      .xt_rsc_0_6_i_qa_d(xt_rsc_0_6_i_qa_d),
      .xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_7_i_adra_d(xt_rsc_0_7_i_adra_d),
      .xt_rsc_0_7_i_da_d(xt_rsc_0_7_i_da_d),
      .xt_rsc_0_7_i_qa_d(xt_rsc_0_7_i_qa_d),
      .xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_8_i_adra_d(xt_rsc_0_8_i_adra_d),
      .xt_rsc_0_8_i_da_d(xt_rsc_0_8_i_da_d),
      .xt_rsc_0_8_i_qa_d(xt_rsc_0_8_i_qa_d),
      .xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_9_i_adra_d(xt_rsc_0_9_i_adra_d),
      .xt_rsc_0_9_i_da_d(xt_rsc_0_9_i_da_d),
      .xt_rsc_0_9_i_qa_d(xt_rsc_0_9_i_qa_d),
      .xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_10_i_adra_d(xt_rsc_0_10_i_adra_d),
      .xt_rsc_0_10_i_da_d(xt_rsc_0_10_i_da_d),
      .xt_rsc_0_10_i_qa_d(xt_rsc_0_10_i_qa_d),
      .xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_11_i_adra_d(xt_rsc_0_11_i_adra_d),
      .xt_rsc_0_11_i_da_d(xt_rsc_0_11_i_da_d),
      .xt_rsc_0_11_i_qa_d(xt_rsc_0_11_i_qa_d),
      .xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_12_i_adra_d(xt_rsc_0_12_i_adra_d),
      .xt_rsc_0_12_i_da_d(xt_rsc_0_12_i_da_d),
      .xt_rsc_0_12_i_qa_d(xt_rsc_0_12_i_qa_d),
      .xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_13_i_adra_d(xt_rsc_0_13_i_adra_d),
      .xt_rsc_0_13_i_da_d(xt_rsc_0_13_i_da_d),
      .xt_rsc_0_13_i_qa_d(xt_rsc_0_13_i_qa_d),
      .xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_14_i_adra_d(xt_rsc_0_14_i_adra_d),
      .xt_rsc_0_14_i_da_d(xt_rsc_0_14_i_da_d),
      .xt_rsc_0_14_i_qa_d(xt_rsc_0_14_i_qa_d),
      .xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_15_i_adra_d(xt_rsc_0_15_i_adra_d),
      .xt_rsc_0_15_i_da_d(xt_rsc_0_15_i_da_d),
      .xt_rsc_0_15_i_qa_d(xt_rsc_0_15_i_qa_d),
      .xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_16_i_adra_d(xt_rsc_0_16_i_adra_d),
      .xt_rsc_0_16_i_da_d(xt_rsc_0_16_i_da_d),
      .xt_rsc_0_16_i_qa_d(xt_rsc_0_16_i_qa_d),
      .xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_17_i_adra_d(xt_rsc_0_17_i_adra_d),
      .xt_rsc_0_17_i_da_d(xt_rsc_0_17_i_da_d),
      .xt_rsc_0_17_i_qa_d(xt_rsc_0_17_i_qa_d),
      .xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_18_i_adra_d(xt_rsc_0_18_i_adra_d),
      .xt_rsc_0_18_i_da_d(xt_rsc_0_18_i_da_d),
      .xt_rsc_0_18_i_qa_d(xt_rsc_0_18_i_qa_d),
      .xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_19_i_adra_d(xt_rsc_0_19_i_adra_d),
      .xt_rsc_0_19_i_da_d(xt_rsc_0_19_i_da_d),
      .xt_rsc_0_19_i_qa_d(xt_rsc_0_19_i_qa_d),
      .xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_20_i_adra_d(xt_rsc_0_20_i_adra_d),
      .xt_rsc_0_20_i_da_d(xt_rsc_0_20_i_da_d),
      .xt_rsc_0_20_i_qa_d(xt_rsc_0_20_i_qa_d),
      .xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_21_i_adra_d(xt_rsc_0_21_i_adra_d),
      .xt_rsc_0_21_i_da_d(xt_rsc_0_21_i_da_d),
      .xt_rsc_0_21_i_qa_d(xt_rsc_0_21_i_qa_d),
      .xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_22_i_adra_d(xt_rsc_0_22_i_adra_d),
      .xt_rsc_0_22_i_da_d(xt_rsc_0_22_i_da_d),
      .xt_rsc_0_22_i_qa_d(xt_rsc_0_22_i_qa_d),
      .xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_23_i_adra_d(xt_rsc_0_23_i_adra_d),
      .xt_rsc_0_23_i_da_d(xt_rsc_0_23_i_da_d),
      .xt_rsc_0_23_i_qa_d(xt_rsc_0_23_i_qa_d),
      .xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_24_i_adra_d(xt_rsc_0_24_i_adra_d),
      .xt_rsc_0_24_i_da_d(xt_rsc_0_24_i_da_d),
      .xt_rsc_0_24_i_qa_d(xt_rsc_0_24_i_qa_d),
      .xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_25_i_adra_d(xt_rsc_0_25_i_adra_d),
      .xt_rsc_0_25_i_da_d(xt_rsc_0_25_i_da_d),
      .xt_rsc_0_25_i_qa_d(xt_rsc_0_25_i_qa_d),
      .xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_26_i_adra_d(xt_rsc_0_26_i_adra_d),
      .xt_rsc_0_26_i_da_d(xt_rsc_0_26_i_da_d),
      .xt_rsc_0_26_i_qa_d(xt_rsc_0_26_i_qa_d),
      .xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_27_i_adra_d(xt_rsc_0_27_i_adra_d),
      .xt_rsc_0_27_i_da_d(xt_rsc_0_27_i_da_d),
      .xt_rsc_0_27_i_qa_d(xt_rsc_0_27_i_qa_d),
      .xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_28_i_adra_d(xt_rsc_0_28_i_adra_d),
      .xt_rsc_0_28_i_da_d(xt_rsc_0_28_i_da_d),
      .xt_rsc_0_28_i_qa_d(xt_rsc_0_28_i_qa_d),
      .xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_29_i_adra_d(xt_rsc_0_29_i_adra_d),
      .xt_rsc_0_29_i_da_d(xt_rsc_0_29_i_da_d),
      .xt_rsc_0_29_i_qa_d(xt_rsc_0_29_i_qa_d),
      .xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_30_i_adra_d(xt_rsc_0_30_i_adra_d),
      .xt_rsc_0_30_i_da_d(xt_rsc_0_30_i_da_d),
      .xt_rsc_0_30_i_qa_d(xt_rsc_0_30_i_qa_d),
      .xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .xt_rsc_0_31_i_adra_d(xt_rsc_0_31_i_adra_d),
      .xt_rsc_0_31_i_da_d(xt_rsc_0_31_i_da_d),
      .xt_rsc_0_31_i_qa_d(xt_rsc_0_31_i_qa_d),
      .xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d(xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_0_i_adra_d(twiddle_rsc_0_0_i_adra_d),
      .twiddle_rsc_0_0_i_qa_d(twiddle_rsc_0_0_i_qa_d),
      .twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_1_i_adra_d(twiddle_rsc_0_1_i_adra_d),
      .twiddle_rsc_0_1_i_qa_d(twiddle_rsc_0_1_i_qa_d),
      .twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_2_i_adra_d(twiddle_rsc_0_2_i_adra_d),
      .twiddle_rsc_0_2_i_qa_d(twiddle_rsc_0_2_i_qa_d),
      .twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_3_i_adra_d(twiddle_rsc_0_3_i_adra_d),
      .twiddle_rsc_0_3_i_qa_d(twiddle_rsc_0_3_i_qa_d),
      .twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_4_i_adra_d(twiddle_rsc_0_4_i_adra_d),
      .twiddle_rsc_0_4_i_qa_d(twiddle_rsc_0_4_i_qa_d),
      .twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_5_i_adra_d(twiddle_rsc_0_5_i_adra_d),
      .twiddle_rsc_0_5_i_qa_d(twiddle_rsc_0_5_i_qa_d),
      .twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_6_i_adra_d(twiddle_rsc_0_6_i_adra_d),
      .twiddle_rsc_0_6_i_qa_d(twiddle_rsc_0_6_i_qa_d),
      .twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_7_i_adra_d(twiddle_rsc_0_7_i_adra_d),
      .twiddle_rsc_0_7_i_qa_d(twiddle_rsc_0_7_i_qa_d),
      .twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_8_i_adra_d(twiddle_rsc_0_8_i_adra_d),
      .twiddle_rsc_0_8_i_qa_d(twiddle_rsc_0_8_i_qa_d),
      .twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_9_i_adra_d(twiddle_rsc_0_9_i_adra_d),
      .twiddle_rsc_0_9_i_qa_d(twiddle_rsc_0_9_i_qa_d),
      .twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_10_i_adra_d(twiddle_rsc_0_10_i_adra_d),
      .twiddle_rsc_0_10_i_qa_d(twiddle_rsc_0_10_i_qa_d),
      .twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_11_i_adra_d(twiddle_rsc_0_11_i_adra_d),
      .twiddle_rsc_0_11_i_qa_d(twiddle_rsc_0_11_i_qa_d),
      .twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_12_i_adra_d(twiddle_rsc_0_12_i_adra_d),
      .twiddle_rsc_0_12_i_qa_d(twiddle_rsc_0_12_i_qa_d),
      .twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_13_i_adra_d(twiddle_rsc_0_13_i_adra_d),
      .twiddle_rsc_0_13_i_qa_d(twiddle_rsc_0_13_i_qa_d),
      .twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_14_i_adra_d(twiddle_rsc_0_14_i_adra_d),
      .twiddle_rsc_0_14_i_qa_d(twiddle_rsc_0_14_i_qa_d),
      .twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_rsc_0_15_i_adra_d(twiddle_rsc_0_15_i_adra_d),
      .twiddle_rsc_0_15_i_qa_d(twiddle_rsc_0_15_i_qa_d),
      .twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_0_i_adra_d(twiddle_h_rsc_0_0_i_adra_d),
      .twiddle_h_rsc_0_0_i_qa_d(twiddle_h_rsc_0_0_i_qa_d),
      .twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_1_i_adra_d(twiddle_h_rsc_0_1_i_adra_d),
      .twiddle_h_rsc_0_1_i_qa_d(twiddle_h_rsc_0_1_i_qa_d),
      .twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_2_i_adra_d(twiddle_h_rsc_0_2_i_adra_d),
      .twiddle_h_rsc_0_2_i_qa_d(twiddle_h_rsc_0_2_i_qa_d),
      .twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_3_i_adra_d(twiddle_h_rsc_0_3_i_adra_d),
      .twiddle_h_rsc_0_3_i_qa_d(twiddle_h_rsc_0_3_i_qa_d),
      .twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_4_i_adra_d(twiddle_h_rsc_0_4_i_adra_d),
      .twiddle_h_rsc_0_4_i_qa_d(twiddle_h_rsc_0_4_i_qa_d),
      .twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_5_i_adra_d(twiddle_h_rsc_0_5_i_adra_d),
      .twiddle_h_rsc_0_5_i_qa_d(twiddle_h_rsc_0_5_i_qa_d),
      .twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_6_i_adra_d(twiddle_h_rsc_0_6_i_adra_d),
      .twiddle_h_rsc_0_6_i_qa_d(twiddle_h_rsc_0_6_i_qa_d),
      .twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_7_i_adra_d(twiddle_h_rsc_0_7_i_adra_d),
      .twiddle_h_rsc_0_7_i_qa_d(twiddle_h_rsc_0_7_i_qa_d),
      .twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_8_i_adra_d(twiddle_h_rsc_0_8_i_adra_d),
      .twiddle_h_rsc_0_8_i_qa_d(twiddle_h_rsc_0_8_i_qa_d),
      .twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_9_i_adra_d(twiddle_h_rsc_0_9_i_adra_d),
      .twiddle_h_rsc_0_9_i_qa_d(twiddle_h_rsc_0_9_i_qa_d),
      .twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_10_i_adra_d(twiddle_h_rsc_0_10_i_adra_d),
      .twiddle_h_rsc_0_10_i_qa_d(twiddle_h_rsc_0_10_i_qa_d),
      .twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_11_i_adra_d(twiddle_h_rsc_0_11_i_adra_d),
      .twiddle_h_rsc_0_11_i_qa_d(twiddle_h_rsc_0_11_i_qa_d),
      .twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_12_i_adra_d(twiddle_h_rsc_0_12_i_adra_d),
      .twiddle_h_rsc_0_12_i_qa_d(twiddle_h_rsc_0_12_i_qa_d),
      .twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_13_i_adra_d(twiddle_h_rsc_0_13_i_adra_d),
      .twiddle_h_rsc_0_13_i_qa_d(twiddle_h_rsc_0_13_i_qa_d),
      .twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_14_i_adra_d(twiddle_h_rsc_0_14_i_adra_d),
      .twiddle_h_rsc_0_14_i_qa_d(twiddle_h_rsc_0_14_i_qa_d),
      .twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .twiddle_h_rsc_0_15_i_adra_d(twiddle_h_rsc_0_15_i_adra_d),
      .twiddle_h_rsc_0_15_i_qa_d(twiddle_h_rsc_0_15_i_qa_d),
      .twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d(twiddle_h_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d),
      .yt_rsc_0_0_i_wea_d_pff(yt_rsc_0_0_i_wea_d_iff),
      .yt_rsc_0_16_i_wea_d_pff(yt_rsc_0_16_i_wea_d_iff),
      .xt_rsc_0_0_i_wea_d_pff(xt_rsc_0_0_i_wea_d_iff),
      .xt_rsc_0_16_i_wea_d_pff(xt_rsc_0_16_i_wea_d_iff)
    );
endmodule



